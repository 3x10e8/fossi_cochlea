magic
tech sky130B
magscale 1 2
timestamp 1662953364
<< metal1 >>
rect 1022 922 1457 956
rect 1423 850 1457 922
<< metal2 >>
rect 515 458 802 496
use comp_clks  comp_clks_0
timestamp 1662950490
transform 1 0 1288 0 1 544
box 0 -544 1196 640
use inv_weak_pulldown_corrected  inv_weak_pulldown_corrected_0
timestamp 1654741520
transform 1 0 276 0 1 128
box -276 -128 368 1056
use inv_weak_pulldown_corrected  inv_weak_pulldown_corrected_1
timestamp 1654741520
transform 1 0 920 0 1 128
box -276 -128 368 1056
<< end >>
