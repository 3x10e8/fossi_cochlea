VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO first_dual_core
  CLASS BLOCK ;
  FOREIGN first_dual_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 490.000 ;
  PIN cclk_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END cclk_I[0]
  PIN cclk_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END cclk_I[1]
  PIN cclk_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 45.600 400.000 46.200 ;
    END
  END cclk_Q[0]
  PIN cclk_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 259.800 400.000 260.400 ;
    END
  END cclk_Q[1]
  PIN clk_master
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END clk_master
  PIN clk_master_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 486.000 29.810 490.000 ;
    END
  END clk_master_out
  PIN clkdiv2_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END clkdiv2_I[0]
  PIN clkdiv2_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END clkdiv2_I[1]
  PIN clkdiv2_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 76.200 400.000 76.800 ;
    END
  END clkdiv2_Q[0]
  PIN clkdiv2_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 290.400 400.000 291.000 ;
    END
  END clkdiv2_Q[1]
  PIN comp_high_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END comp_high_I[0]
  PIN comp_high_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END comp_high_I[1]
  PIN comp_high_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 106.800 400.000 107.400 ;
    END
  END comp_high_Q[0]
  PIN comp_high_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 321.000 400.000 321.600 ;
    END
  END comp_high_Q[1]
  PIN cos_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END cos_out[0]
  PIN cos_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.800 4.000 413.400 ;
    END
  END cos_out[1]
  PIN cos_outb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END cos_outb[0]
  PIN cos_outb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END cos_outb[1]
  PIN div2out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 486.000 69.830 490.000 ;
    END
  END div2out
  PIN fb1_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END fb1_I[0]
  PIN fb1_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END fb1_I[1]
  PIN fb1_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 168.000 400.000 168.600 ;
    END
  END fb1_Q[0]
  PIN fb1_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 382.200 400.000 382.800 ;
    END
  END fb1_Q[1]
  PIN fb2_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END fb2_I[0]
  PIN fb2_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 486.000 370.210 490.000 ;
    END
  END fb2_I[1]
  PIN fb2_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 486.000 349.970 490.000 ;
    END
  END fb2_Q[0]
  PIN fb2_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 486.000 389.990 490.000 ;
    END
  END fb2_Q[1]
  PIN gray_clk_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 486.000 269.930 490.000 ;
    END
  END gray_clk_out[10]
  PIN gray_clk_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 486.000 90.070 490.000 ;
    END
  END gray_clk_out[1]
  PIN gray_clk_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 486.000 109.850 490.000 ;
    END
  END gray_clk_out[2]
  PIN gray_clk_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 486.000 130.090 490.000 ;
    END
  END gray_clk_out[3]
  PIN gray_clk_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 486.000 149.870 490.000 ;
    END
  END gray_clk_out[4]
  PIN gray_clk_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 486.000 170.110 490.000 ;
    END
  END gray_clk_out[5]
  PIN gray_clk_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 486.000 189.890 490.000 ;
    END
  END gray_clk_out[6]
  PIN gray_clk_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 486.000 210.130 490.000 ;
    END
  END gray_clk_out[7]
  PIN gray_clk_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 486.000 229.910 490.000 ;
    END
  END gray_clk_out[8]
  PIN gray_clk_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 486.000 250.150 490.000 ;
    END
  END gray_clk_out[9]
  PIN no_ones_below_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 486.000 290.170 490.000 ;
    END
  END no_ones_below_out[0]
  PIN no_ones_below_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 486.000 309.950 490.000 ;
    END
  END no_ones_below_out[1]
  PIN no_ones_below_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 486.000 330.190 490.000 ;
    END
  END no_ones_below_out[2]
  PIN phi1b_dig_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END phi1b_dig_I[0]
  PIN phi1b_dig_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 290.400 4.000 291.000 ;
    END
  END phi1b_dig_I[1]
  PIN phi1b_dig_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 137.400 400.000 138.000 ;
    END
  END phi1b_dig_Q[0]
  PIN phi1b_dig_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 351.600 400.000 352.200 ;
    END
  END phi1b_dig_Q[1]
  PIN read_out_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END read_out_I[0]
  PIN read_out_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END read_out_I[1]
  PIN read_out_I_top[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END read_out_I_top[0]
  PIN read_out_I_top[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.000 4.000 474.600 ;
    END
  END read_out_I_top[1]
  PIN read_out_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END read_out_Q[0]
  PIN read_out_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END read_out_Q[1]
  PIN read_out_Q_top[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 443.400 400.000 444.000 ;
    END
  END read_out_Q_top[0]
  PIN read_out_Q_top[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 474.000 400.000 474.600 ;
    END
  END read_out_Q_top[1]
  PIN rstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END rstb
  PIN rstb_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 486.000 10.030 490.000 ;
    END
  END rstb_out
  PIN sin_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 15.000 400.000 15.600 ;
    END
  END sin_out[0]
  PIN sin_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 229.200 400.000 229.800 ;
    END
  END sin_out[1]
  PIN sin_outb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 198.600 400.000 199.200 ;
    END
  END sin_outb[0]
  PIN sin_outb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 412.800 400.000 413.400 ;
    END
  END sin_outb[1]
  PIN ud_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END ud_en
  PIN ud_en_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 486.000 50.050 490.000 ;
    END
  END ud_en_out
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 478.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 478.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 478.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 478.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 478.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 394.220 478.805 ;
      LAYER met1 ;
        RECT 5.520 10.640 394.220 479.360 ;
      LAYER met2 ;
        RECT 6.990 485.720 9.470 486.610 ;
        RECT 10.310 485.720 29.250 486.610 ;
        RECT 30.090 485.720 49.490 486.610 ;
        RECT 50.330 485.720 69.270 486.610 ;
        RECT 70.110 485.720 89.510 486.610 ;
        RECT 90.350 485.720 109.290 486.610 ;
        RECT 110.130 485.720 129.530 486.610 ;
        RECT 130.370 485.720 149.310 486.610 ;
        RECT 150.150 485.720 169.550 486.610 ;
        RECT 170.390 485.720 189.330 486.610 ;
        RECT 190.170 485.720 209.570 486.610 ;
        RECT 210.410 485.720 229.350 486.610 ;
        RECT 230.190 485.720 249.590 486.610 ;
        RECT 250.430 485.720 269.370 486.610 ;
        RECT 270.210 485.720 289.610 486.610 ;
        RECT 290.450 485.720 309.390 486.610 ;
        RECT 310.230 485.720 329.630 486.610 ;
        RECT 330.470 485.720 349.410 486.610 ;
        RECT 350.250 485.720 369.650 486.610 ;
        RECT 370.490 485.720 389.430 486.610 ;
        RECT 390.270 485.720 394.130 486.610 ;
        RECT 6.990 4.280 394.130 485.720 ;
        RECT 6.990 3.670 24.650 4.280 ;
        RECT 25.490 3.670 74.330 4.280 ;
        RECT 75.170 3.670 124.470 4.280 ;
        RECT 125.310 3.670 174.610 4.280 ;
        RECT 175.450 3.670 224.750 4.280 ;
        RECT 225.590 3.670 274.430 4.280 ;
        RECT 275.270 3.670 324.570 4.280 ;
        RECT 325.410 3.670 374.710 4.280 ;
        RECT 375.550 3.670 394.130 4.280 ;
      LAYER met3 ;
        RECT 4.000 475.000 396.000 482.625 ;
        RECT 4.400 473.600 395.600 475.000 ;
        RECT 4.000 444.400 396.000 473.600 ;
        RECT 4.400 443.000 395.600 444.400 ;
        RECT 4.000 413.800 396.000 443.000 ;
        RECT 4.400 412.400 395.600 413.800 ;
        RECT 4.000 383.200 396.000 412.400 ;
        RECT 4.400 381.800 395.600 383.200 ;
        RECT 4.000 352.600 396.000 381.800 ;
        RECT 4.400 351.200 395.600 352.600 ;
        RECT 4.000 322.000 396.000 351.200 ;
        RECT 4.400 320.600 395.600 322.000 ;
        RECT 4.000 291.400 396.000 320.600 ;
        RECT 4.400 290.000 395.600 291.400 ;
        RECT 4.000 260.800 396.000 290.000 ;
        RECT 4.400 259.400 395.600 260.800 ;
        RECT 4.000 230.200 396.000 259.400 ;
        RECT 4.400 228.800 395.600 230.200 ;
        RECT 4.000 199.600 396.000 228.800 ;
        RECT 4.400 198.200 395.600 199.600 ;
        RECT 4.000 169.000 396.000 198.200 ;
        RECT 4.400 167.600 395.600 169.000 ;
        RECT 4.000 138.400 396.000 167.600 ;
        RECT 4.400 137.000 395.600 138.400 ;
        RECT 4.000 107.800 396.000 137.000 ;
        RECT 4.400 106.400 395.600 107.800 ;
        RECT 4.000 77.200 396.000 106.400 ;
        RECT 4.400 75.800 395.600 77.200 ;
        RECT 4.000 46.600 396.000 75.800 ;
        RECT 4.400 45.200 395.600 46.600 ;
        RECT 4.000 16.000 396.000 45.200 ;
        RECT 4.400 14.600 395.600 16.000 ;
        RECT 4.000 10.715 396.000 14.600 ;
      LAYER met4 ;
        RECT 47.215 479.360 380.585 482.625 ;
        RECT 47.215 177.655 97.440 479.360 ;
        RECT 99.840 177.655 174.240 479.360 ;
        RECT 176.640 177.655 251.040 479.360 ;
        RECT 253.440 177.655 327.840 479.360 ;
        RECT 330.240 177.655 380.585 479.360 ;
  END
END first_dual_core
END LIBRARY

