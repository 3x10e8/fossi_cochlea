magic
tech sky130B
magscale 1 2
timestamp 1654741520
<< metal3 >>
rect -712 2168 -390 2354
rect -712 1728 -679 2168
rect -421 2048 -390 2168
rect -44 2048 276 2354
rect -421 2046 276 2048
rect 824 2046 1144 2354
rect 1692 2048 2012 2354
rect 1692 2046 2038 2048
rect -421 2022 2038 2046
rect -421 1728 2344 2022
rect -712 1196 -390 1728
rect -68 1702 2344 1728
rect -68 1196 2036 1702
rect -712 -669 -679 1196
rect -421 1154 2036 1196
rect -421 875 2344 1154
rect -421 342 -390 875
rect -68 834 2344 875
rect -68 342 2036 834
rect -421 286 2036 342
rect -421 22 2344 286
rect -421 -380 -390 22
rect -68 -34 2344 22
rect -68 -58 2038 -34
rect -68 -380 252 -58
rect 825 -380 1145 -58
rect 1718 -380 2038 -58
rect -421 -411 2344 -380
rect 252 -669 825 -411
rect 2158 -669 2344 -411
rect -712 -702 2344 -669
<< via3 >>
rect -679 1728 -421 2168
rect -679 -411 -421 1196
rect -679 -669 252 -411
rect 825 -669 2158 -411
<< mimcap >>
rect -16 1786 1984 1994
rect -16 202 192 1786
rect 336 1066 912 1642
rect 1056 1066 1632 1642
rect 336 346 912 922
rect 1056 346 1632 922
rect 1776 202 1984 1786
rect -16 -6 1984 202
<< mimcapcontact >>
rect 192 1642 1776 1786
rect 192 1066 336 1642
rect 912 1066 1056 1642
rect 1632 1066 1776 1642
rect 192 922 1776 1066
rect 192 346 336 922
rect 912 346 1056 922
rect 1632 346 1776 922
rect 192 202 1776 346
<< metal4 >>
rect -686 2168 -414 2169
rect 36 2022 196 2354
rect 904 2022 1064 2354
rect 1772 2022 1932 2354
rect -686 1727 -414 1728
rect -44 1942 2012 2022
rect -44 1786 2344 1942
rect -686 1196 -414 1197
rect -44 202 192 1786
rect 1776 1782 2344 1786
rect 336 1066 912 1642
rect 1056 1066 1632 1642
rect 1776 1074 2012 1782
rect 336 346 912 922
rect 1056 346 1632 922
rect 1776 914 2344 1074
rect 1776 206 2012 914
rect 1776 202 2344 206
rect -44 46 2344 202
rect -44 -34 2012 46
rect 252 -676 253 -404
rect 824 -676 825 -404
rect 2158 -676 2344 -404
<< via4 >>
rect -686 1728 -679 2168
rect -679 1728 -421 2168
rect -421 1728 -414 2168
rect -686 -669 -679 1196
rect -679 -411 -421 1196
rect -421 -404 -414 1196
rect -421 -411 252 -404
rect -679 -669 252 -411
rect -686 -676 252 -669
rect 825 -411 2158 -404
rect 825 -669 2158 -411
rect 825 -676 2158 -669
<< mimcap2 >>
rect -16 1812 1984 1994
rect -16 1576 166 1812
rect 402 1576 516 1812
rect 752 1576 866 1812
rect 1102 1576 1216 1812
rect 1452 1576 1566 1812
rect 1802 1576 1984 1812
rect -16 1462 1984 1576
rect -16 1226 166 1462
rect 402 1226 866 1462
rect 1102 1226 1566 1462
rect 1802 1226 1984 1462
rect -16 1112 1984 1226
rect -16 876 166 1112
rect 402 876 516 1112
rect 752 876 866 1112
rect 1102 876 1216 1112
rect 1452 876 1566 1112
rect 1802 876 1984 1112
rect -16 762 1984 876
rect -16 526 166 762
rect 402 526 866 762
rect 1102 526 1566 762
rect 1802 526 1984 762
rect -16 412 1984 526
rect -16 176 166 412
rect 402 176 516 412
rect 752 176 866 412
rect 1102 176 1216 412
rect 1452 176 1566 412
rect 1802 176 1984 412
rect -16 -6 1984 176
<< mimcap2contact >>
rect 166 1576 402 1812
rect 516 1576 752 1812
rect 866 1576 1102 1812
rect 1216 1576 1452 1812
rect 1566 1576 1802 1812
rect 166 1226 402 1462
rect 866 1226 1102 1462
rect 1566 1226 1802 1462
rect 166 876 402 1112
rect 516 876 752 1112
rect 866 876 1102 1112
rect 1216 876 1452 1112
rect 1566 876 1802 1112
rect 166 526 402 762
rect 866 526 1102 762
rect 1566 526 1802 762
rect 166 176 402 412
rect 516 176 752 412
rect 866 176 1102 412
rect 1216 176 1452 412
rect 1566 176 1802 412
<< metal5 >>
rect -710 2168 -390 2354
rect -710 1728 -686 2168
rect -414 2048 -390 2168
rect -44 2048 276 2354
rect -414 2046 276 2048
rect 824 2046 1144 2354
rect 1692 2048 2012 2354
rect 1692 2046 2038 2048
rect -414 2022 2038 2046
rect -414 1812 2344 2022
rect -414 1728 166 1812
rect -710 1196 -390 1728
rect -68 1576 166 1728
rect 402 1576 516 1812
rect 752 1576 866 1812
rect 1102 1576 1216 1812
rect 1452 1576 1566 1812
rect 1802 1702 2344 1812
rect 1802 1576 2036 1702
rect -68 1462 2036 1576
rect -68 1226 166 1462
rect 402 1226 866 1462
rect 1102 1226 1566 1462
rect 1802 1226 2036 1462
rect -68 1196 2036 1226
rect -710 -676 -686 1196
rect -414 1154 2036 1196
rect -414 1112 2344 1154
rect -414 876 166 1112
rect 402 876 516 1112
rect 752 876 866 1112
rect 1102 876 1216 1112
rect 1452 876 1566 1112
rect 1802 876 2344 1112
rect -414 875 2344 876
rect -414 342 -390 875
rect -68 834 2344 875
rect -68 762 2036 834
rect -68 526 166 762
rect 402 526 866 762
rect 1102 526 1566 762
rect 1802 526 2036 762
rect -68 412 2036 526
rect -68 342 166 412
rect -414 176 166 342
rect 402 176 516 412
rect 752 176 866 412
rect 1102 176 1216 412
rect 1452 176 1566 412
rect 1802 286 2036 412
rect 1802 176 2344 286
rect -414 22 2344 176
rect -414 -380 -390 22
rect -68 -34 2344 22
rect -68 -58 2038 -34
rect -68 -380 252 -58
rect 825 -380 1145 -58
rect 1718 -380 2038 -58
rect -414 -404 2344 -380
rect 252 -676 825 -404
rect 2158 -676 2344 -404
rect -710 -700 2344 -676
<< end >>
