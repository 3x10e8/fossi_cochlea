magic
tech sky130B
magscale 1 2
timestamp 1654753126
<< nwell >>
rect -56 581 848 680
rect 1102 551 2007 722
<< psubdiff >>
rect 926 78 1026 127
rect 926 28 949 78
rect 1000 28 1026 78
rect 926 -11 1026 28
<< nsubdiff >>
rect 338 616 487 643
rect 338 579 396 616
rect 439 579 487 616
rect 338 563 487 579
rect 1401 620 1559 670
rect 1401 586 1462 620
rect 1496 586 1559 620
rect 1401 563 1559 586
rect 374 562 459 563
<< psubdiffcont >>
rect 949 28 1000 78
<< nsubdiffcont >>
rect 396 579 439 616
rect 1462 586 1496 620
<< locali >>
rect 378 616 455 633
rect 378 579 396 616
rect 439 579 455 616
rect 378 563 455 579
rect 1455 620 1505 637
rect 1455 586 1462 620
rect 1496 586 1505 620
rect 1455 560 1505 586
rect 949 78 1000 94
rect 949 12 1000 28
<< viali >>
rect 134 227 168 261
rect 218 228 252 262
rect 301 227 335 261
rect 747 223 781 257
rect 1353 223 1387 257
rect 1906 223 1940 257
rect 949 28 1000 78
<< metal1 >>
rect -71 262 400 272
rect -71 261 218 262
rect -71 227 134 261
rect 168 228 218 261
rect 252 261 400 262
rect 252 228 301 261
rect 168 227 301 228
rect 335 227 400 261
rect -71 214 400 227
rect 731 257 1421 267
rect 731 223 747 257
rect 781 223 1353 257
rect 1387 223 1421 257
rect 731 212 1421 223
rect 1873 257 2139 271
rect 1873 223 1906 257
rect 1940 223 2139 257
rect 1873 207 2139 223
rect 938 78 1009 97
rect 938 50 949 78
rect 802 28 949 50
rect 1000 50 1009 78
rect 1000 28 1152 50
rect 802 -46 1152 28
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 -18 0 1 2
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_1
timestamp 1644511149
transform 1 0 1140 0 1 2
box -38 -48 866 592
<< end >>
