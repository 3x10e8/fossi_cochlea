* NGSPICE file created from digital_unison.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlrtn_1 abstract view
.subckt sky130_fd_sc_hd__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_4 abstract view
.subckt sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

.subckt digital_unison cclk_I[0] cclk_I[1] cclk_Q[0] cclk_Q[1] clk_master clkdiv2_I[0]
+ clkdiv2_I[1] clkdiv2_Q[0] clkdiv2_Q[1] comp_high_I[0] comp_high_I[1] comp_high_Q[0]
+ comp_high_Q[1] cos_out[0] cos_out[1] fb1_I[0] fb1_I[1] fb1_Q[0] fb1_Q[1] phi1b_dig_I[0]
+ phi1b_dig_I[1] phi1b_dig_Q[0] phi1b_dig_Q[1] read_out_I[0] read_out_I[1] read_out_Q[0]
+ read_out_Q[1] rstb sin_out[0] sin_out[1] ud_en vccd1 vssd1
XFILLER_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1231__CLK _1357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0717__B1 _0716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1254__CLK input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1270_ _0542_/B _1270_/D _1148_/CLK vssd1 vssd1 vccd1 vccd1 _1270_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1048__31 _1052__35/A vssd1 vssd1 vccd1 vccd1 _1153_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0542__C_N _0548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0985_ _0980_/B _0984_/X _0755_/A vssd1 vssd1 vccd1 vccd1 _0986_/B sky130_fd_sc_hd__o21ai_1
XFILLER_9_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0938__B1 _0831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_TE_B _0946_/Y vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0770_ _1199_/Q _1198_/Q vssd1 vssd1 vccd1 vccd1 _0770_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_6_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1253_ _1098_/Y _1253_/D _1034_/B vssd1 vssd1 vccd1 vccd1 _1253_/Q sky130_fd_sc_hd__dfrtp_1
X_1322_ _1358_/A _1322_/D fanout46/X vssd1 vssd1 vccd1 vccd1 _1322_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1184_ _1359_/A _1184_/D fanout55/X vssd1 vssd1 vccd1 vccd1 _1184_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__0518__A _1042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0968_ _0966_/X _0967_/Y _0755_/A vssd1 vssd1 vccd1 vccd1 _0969_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__1084__A _1130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0899_ _1276_/Q _0899_/B vssd1 vssd1 vccd1 vccd1 _1276_/D sky130_fd_sc_hd__xnor2_1
XFILLER_9_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0822_ _0822_/A vssd1 vssd1 vccd1 vccd1 _0822_/Y sky130_fd_sc_hd__inv_2
X_0684_ _1332_/Q vssd1 vssd1 vccd1 vccd1 _1331_/D sky130_fd_sc_hd__inv_2
XFILLER_9_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0753_ _1013_/A _0753_/B vssd1 vssd1 vccd1 vccd1 _0754_/B sky130_fd_sc_hd__nand2_1
X_1305_ _0560_/A _1305_/D _1120__55/Y vssd1 vssd1 vccd1 vccd1 _1305_/Q sky130_fd_sc_hd__dfrtp_1
X_1236_ _0644_/D _1236_/D _1081_/Y vssd1 vssd1 vccd1 vccd1 _1236_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1098_ _1144_/A _1144_/B vssd1 vssd1 vccd1 vccd1 _1098_/Y sky130_fd_sc_hd__xnor2_2
X_1167_ _1167_/CLK _1167_/D fanout54/X vssd1 vssd1 vccd1 vccd1 _1167_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0838__C1 _0831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1021_ _1342_/Q _1341_/Q vssd1 vssd1 vccd1 vccd1 _1021_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf _1275_/Q _0952_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
X_0805_ _1222_/Q _0805_/B vssd1 vssd1 vccd1 vccd1 _1222_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__1338__CLK _1035_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0598_ _1179_/Q vssd1 vssd1 vccd1 vccd1 _1178_/D sky130_fd_sc_hd__clkinv_2
X_0667_ _1297_/Q vssd1 vssd1 vccd1 vccd1 _1298_/D sky130_fd_sc_hd__inv_2
X_0736_ _0735_/Y _0727_/B _0716_/X vssd1 vssd1 vccd1 vccd1 _0737_/B sky130_fd_sc_hd__a21o_1
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1219_ fanout34/X _1219_/D fanout58/X vssd1 vssd1 vccd1 vccd1 _1219_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0521_ _1133_/A _1133_/B vssd1 vssd1 vccd1 vccd1 _0868_/A sky130_fd_sc_hd__xor2_4
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1004_ _1324_/Q _1004_/B vssd1 vssd1 vccd1 vccd1 _1004_/X sky130_fd_sc_hd__or2_1
XANTENNA__1357__A _1357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1092__A _1097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0719_ _1185_/Q _1184_/Q _0724_/B vssd1 vssd1 vccd1 vccd1 _0719_/X sky130_fd_sc_hd__and3_1
XFILLER_26_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput20 _1365_/X vssd1 vssd1 vccd1 vccd1 cos_out[1] sky130_fd_sc_hd__buf_2
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0446__1_A _1053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1183__CLK fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1327__D _1327_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0504_ _1153_/Q vssd1 vssd1 vccd1 vccd1 _1146_/A sky130_fd_sc_hd__buf_6
XTAP_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0703__B _1180_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1087__A _1133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1127__58 _1140__64/A vssd1 vssd1 vccd1 vccd1 _1127__58/Y sky130_fd_sc_hd__inv_2
XFILLER_18_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0984_ _1318_/Q _0984_/B vssd1 vssd1 vccd1 vccd1 _0984_/X sky130_fd_sc_hd__and2b_1
XANTENNA__0804__A _1013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1370__A _1370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
+ _1186_/Q _0774_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__1221__CLK _1357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1252_ _1042_/A _1252_/D _1097_/Y vssd1 vssd1 vccd1 vccd1 _1252_/Q sky130_fd_sc_hd__dfrtp_1
X_1321_ _1358_/A _1321_/D fanout45/X vssd1 vssd1 vccd1 vccd1 _1321_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1183_ fanout31/X _1183_/D fanout52/X vssd1 vssd1 vccd1 vccd1 _1183_/Q sky130_fd_sc_hd__dfrtp_2
X_0967_ _1313_/Q _0967_/B vssd1 vssd1 vccd1 vccd1 _0967_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1365__A _1365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1084__B _1130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0898_ _0896_/X _0897_/Y _0755_/X vssd1 vssd1 vccd1 vccd1 _0899_/B sky130_fd_sc_hd__o21ai_1
XFILLER_24_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1244__CLK _1089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0821_ _1227_/Q _0821_/B vssd1 vssd1 vccd1 vccd1 _1227_/D sky130_fd_sc_hd__xnor2_1
X_0752_ _0751_/Y _0710_/C _1193_/Q vssd1 vssd1 vccd1 vccd1 _0753_/B sky130_fd_sc_hd__mux2_1
X_0683_ _1329_/Q vssd1 vssd1 vccd1 vccd1 _1330_/D sky130_fd_sc_hd__inv_2
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1304_ _0862_/A _1304_/D _1119__54/Y vssd1 vssd1 vccd1 vccd1 _1304_/Q sky130_fd_sc_hd__dfrtp_4
X_1166_ _1168_/CLK _1166_/D fanout43/X vssd1 vssd1 vccd1 vccd1 _1166_/Q sky130_fd_sc_hd__dfrtp_1
X_1235_ _0643_/Y _1235_/D _1080_/Y vssd1 vssd1 vccd1 vccd1 _1235_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1191__RESET_B fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0465__22 _0467__24/A vssd1 vssd1 vccd1 vccd1 _0465__22/Y sky130_fd_sc_hd__inv_2
XFILLER_21_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1097_ _1097_/A vssd1 vssd1 vccd1 vccd1 _1097_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1095__A _1097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout50_A fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0902__A _1277_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1020_ _1340_/Q _1339_/Q vssd1 vssd1 vccd1 vccd1 _1020_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_19_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_A _1316_/Q vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0531__B _1137_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0804_ _1013_/A _0804_/B vssd1 vssd1 vccd1 vccd1 _0805_/B sky130_fd_sc_hd__nand2_1
XANTENNA__0812__A _1224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0735_ _1188_/Q _0735_/B vssd1 vssd1 vccd1 vccd1 _0735_/Y sky130_fd_sc_hd__nand2_1
X_0597_ _1176_/Q vssd1 vssd1 vccd1 vccd1 _1177_/D sky130_fd_sc_hd__inv_2
X_0666_ _1298_/Q vssd1 vssd1 vccd1 vccd1 _1297_/D sky130_fd_sc_hd__inv_2
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1149_ _1149_/CLK _1149_/D fanout44/X vssd1 vssd1 vccd1 vccd1 _1149_/Q sky130_fd_sc_hd__dfrtp_1
X_1218_ _1357_/A _1218_/D fanout56/X vssd1 vssd1 vccd1 vccd1 _1218_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0520_ _1166_/Q vssd1 vssd1 vccd1 vccd1 _1133_/B sky130_fd_sc_hd__buf_6
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1003_ _1326_/Q _1352_/D vssd1 vssd1 vccd1 vccd1 _1004_/B sky130_fd_sc_hd__or2_1
XFILLER_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1305__CLK _0560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0542__A _0548_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0718_ _1182_/Q _0718_/B vssd1 vssd1 vccd1 vccd1 _1182_/D sky130_fd_sc_hd__xnor2_1
X_0649_ _1266_/Q _0650_/B vssd1 vssd1 vccd1 vccd1 _1265_/D sky130_fd_sc_hd__xnor2_2
XANTENNA__1373__A _1373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput21 _1366_/X vssd1 vssd1 vccd1 vccd1 fb1_I[0] sky130_fd_sc_hd__buf_2
XFILLER_1_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1223__RESET_B fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0503_ _1151_/Q vssd1 vssd1 vccd1 vccd1 _1151_/D sky130_fd_sc_hd__inv_2
XTAP_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0537__A _0560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1148_/CLK fanout41/X vssd1 vssd1 vccd1 vccd1 _1368_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__1087__B _1133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0447__A _1053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0983_ _1319_/Q _0983_/B vssd1 vssd1 vccd1 vccd1 _0984_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1098__A _1144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1054__36 _1058__40/A vssd1 vssd1 vccd1 vccd1 _1163_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0730__A _1185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf _1283_/Q _0944_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1320_ _1356_/A _1320_/D fanout46/X vssd1 vssd1 vccd1 vccd1 _1320_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1251_ _1096_/Y _1251_/D _0470_/Y vssd1 vssd1 vccd1 vccd1 _1251_/Q sky130_fd_sc_hd__dfrtp_1
X_1182_ _1359_/A _1182_/D fanout52/X vssd1 vssd1 vccd1 vccd1 _1182_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0550__A _1142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0966_ _1314_/Q _1313_/Q _0970_/B vssd1 vssd1 vccd1 vccd1 _0966_/X sky130_fd_sc_hd__and3_1
X_0897_ _1277_/Q _0897_/B vssd1 vssd1 vccd1 vccd1 _0897_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1326__RESET_B fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0820_ _0816_/B _0819_/Y _0755_/X vssd1 vssd1 vccd1 vccd1 _0821_/B sky130_fd_sc_hd__o21ai_1
X_0751_ _0751_/A vssd1 vssd1 vccd1 vccd1 _0751_/Y sky130_fd_sc_hd__inv_2
X_0682_ _1330_/Q vssd1 vssd1 vccd1 vccd1 _1329_/D sky130_fd_sc_hd__inv_2
X_1303_ _1118_/X _1303_/D _0461__18/Y vssd1 vssd1 vccd1 vccd1 _1303_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1165_ _1165_/CLK _1165_/D fanout50/X vssd1 vssd1 vccd1 vccd1 _1165_/Q sky130_fd_sc_hd__dfrtp_1
X_1096_ _1142_/A _1142_/B vssd1 vssd1 vccd1 vccd1 _1096_/Y sky130_fd_sc_hd__xnor2_2
X_1234_ _1078_/X _1234_/D _0478_/Y vssd1 vssd1 vccd1 vccd1 _1234_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0545__A _1042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0949_ _1302_/Q _1301_/Q vssd1 vssd1 vccd1 vccd1 _0949_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout43_A fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1211__CLK _1035_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1143__3_A _1053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output24_A _1369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0665_ _1295_/Q vssd1 vssd1 vccd1 vccd1 _1296_/D sky130_fd_sc_hd__inv_2
X_0734_ _1186_/Q _0734_/B vssd1 vssd1 vccd1 vccd1 _1186_/D sky130_fd_sc_hd__xnor2_1
X_0803_ _1224_/Q _1223_/Q _0806_/B _0800_/B vssd1 vssd1 vccd1 vccd1 _0804_/B sky130_fd_sc_hd__a31o_1
XANTENNA__0756__B1 _0755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0596_ _1177_/Q vssd1 vssd1 vccd1 vccd1 _1176_/D sky130_fd_sc_hd__inv_2
XFILLER_26_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1217_ _0546_/A _1217_/D _0479_/Y vssd1 vssd1 vccd1 vccd1 _1217_/Q sky130_fd_sc_hd__dfrtp_1
X_1079_ _1079_/A vssd1 vssd1 vccd1 vccd1 _1097_/A sky130_fd_sc_hd__buf_4
X_1148_ _1148_/CLK _1148_/D fanout42/X vssd1 vssd1 vccd1 vccd1 _1148_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1234__CLK _1078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0706__C _1188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__0311_ clkbuf_0__0311_/X vssd1 vssd1 vccd1 vccd1 _1049__32/A sky130_fd_sc_hd__clkbuf_16
XFILLER_12_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1257__CLK input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1002_ _1326_/Q _1352_/D _1324_/Q vssd1 vssd1 vccd1 vccd1 _1002_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__0542__B _0542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0977__B1 _0974_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1099_/A fanout58/X vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__dlrtn_1
X_0648_ _0644_/C _0585_/B _0870_/A vssd1 vssd1 vccd1 vccd1 _0650_/B sky130_fd_sc_hd__mux2_1
X_0717_ _0708_/X _0713_/Y _0716_/X vssd1 vssd1 vccd1 vccd1 _0718_/B sky130_fd_sc_hd__a21o_1
XANTENNA__0729__B1 _0998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0579_ _1170_/Q vssd1 vssd1 vccd1 vccd1 _1130_/B sky130_fd_sc_hd__buf_4
XANTENNA__0901__B1 _0831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0733__A _1013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0968__B1 _0755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput22 _1367_/X vssd1 vssd1 vccd1 vccd1 fb1_I[1] sky130_fd_sc_hd__buf_2
Xoutput11 _1356_/X vssd1 vssd1 vccd1 vccd1 cclk_I[0] sky130_fd_sc_hd__clkbuf_1
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0908__A _0998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0643__A _0643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0974__A_N _1315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0502_ _1150_/Q vssd1 vssd1 vccd1 vccd1 _1150_/D sky130_fd_sc_hd__clkinv_2
XFILLER_8_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0537__B _0560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0553__A _0560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1168_/CLK fanout42/X vssd1 vssd1 vccd1 vccd1 _1366_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_27_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf _1325_/Q _1023_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_1_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0982_ _1316_/Q _0982_/B vssd1 vssd1 vccd1 vccd1 _1316_/D sky130_fd_sc_hd__xnor2_1
XFILLER_9_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1098__B _1144_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0458__A _1122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1181_ _1066_/Y _1181_/D _0490__25/Y vssd1 vssd1 vccd1 vccd1 _1181_/Q sky130_fd_sc_hd__dfrtp_1
X_1250_ _0518_/Y _1250_/D _1095_/Y vssd1 vssd1 vccd1 vccd1 _1250_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0965_ _1311_/Q _0965_/B vssd1 vssd1 vccd1 vccd1 _1311_/D sky130_fd_sc_hd__xnor2_1
X_0896_ _1278_/Q _1277_/Q _0900_/B vssd1 vssd1 vccd1 vccd1 _0896_/X sky130_fd_sc_hd__and3_1
XANTENNA__0831__A _0831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_A _1279_/Q vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1259__D _1259_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0741__A _1188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1120__55 _1120__55/A vssd1 vssd1 vccd1 vccd1 _1120__55/Y sky130_fd_sc_hd__inv_2
XFILLER_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1169__D _1169_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0681_ _1327_/Q vssd1 vssd1 vccd1 vccd1 _1328_/D sky130_fd_sc_hd__inv_2
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0750_ _1191_/Q _0750_/B vssd1 vssd1 vccd1 vccd1 _1191_/D sky130_fd_sc_hd__xnor2_1
X_1302_ _1035_/B _1302_/D _1117__53/Y vssd1 vssd1 vccd1 vccd1 _1302_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_2_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1233_ fanout34/X _1233_/D fanout55/X vssd1 vssd1 vccd1 vccd1 _1233_/Q sky130_fd_sc_hd__dfrtp_2
X_1164_ _1360_/A _1164_/D fanout45/X vssd1 vssd1 vccd1 vccd1 _1164_/Q sky130_fd_sc_hd__dfrtp_1
X_1095_ _1097_/A vssd1 vssd1 vccd1 vccd1 _1095_/Y sky130_fd_sc_hd__inv_2
X_0948_ _1300_/Q _1299_/Q vssd1 vssd1 vccd1 vccd1 _0948_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_20_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0545__B _0560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0879_ _0879_/A _0879_/B vssd1 vssd1 vccd1 vccd1 _1365_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0471__A _0479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0646__A _1264_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0802_ _1221_/Q _0802_/B vssd1 vssd1 vccd1 vccd1 _1221_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__1186__CLK fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0664_ _1296_/Q vssd1 vssd1 vccd1 vccd1 _1295_/D sky130_fd_sc_hd__inv_2
XFILLER_6_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0733_ _1013_/A _0733_/B vssd1 vssd1 vccd1 vccd1 _0734_/B sky130_fd_sc_hd__nand2_1
XFILLER_7_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0595_ _1174_/Q vssd1 vssd1 vccd1 vccd1 _1175_/D sky130_fd_sc_hd__inv_2
X_1216_ _1042_/A _1216_/D _1077_/Y vssd1 vssd1 vccd1 vccd1 _1216_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_26_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0556__A _1139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1078_ _1263_/Q _1264_/Q vssd1 vssd1 vccd1 vccd1 _1078_/X sky130_fd_sc_hd__xor2_2
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
+ _1221_/Q _0846_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__0913__B _0913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1001_ _1322_/Q _1001_/B vssd1 vssd1 vccd1 vccd1 _1322_/D sky130_fd_sc_hd__xnor2_1
X_0578_ _1171_/Q vssd1 vssd1 vccd1 vccd1 _1130_/A sky130_fd_sc_hd__buf_4
X_0647_ _1266_/Q _1265_/Q vssd1 vssd1 vccd1 vccd1 _0870_/A sky130_fd_sc_hd__xnor2_1
X_0716_ _0831_/A vssd1 vssd1 vccd1 vccd1 _0716_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1351__CLK input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1079_/A fanout57/X vssd1 vssd1 vccd1 vccd1 _1367_/A sky130_fd_sc_hd__dlrtn_1
Xoutput12 _1357_/X vssd1 vssd1 vccd1 vccd1 cclk_I[1] sky130_fd_sc_hd__buf_2
XFILLER_21_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput23 _1368_/X vssd1 vssd1 vccd1 vccd1 fb1_Q[0] sky130_fd_sc_hd__buf_2
XFILLER_5_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1224__CLK _1357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0501_ _1105_/A _0548_/B vssd1 vssd1 vccd1 vccd1 _1149_/D sky130_fd_sc_hd__xnor2_1
XTAP_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0553__B _0862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0834__A _1259_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input8_A phi1b_dig_Q[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1247__CLK _1035_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0919__A _1282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0981_ _0980_/Y _0973_/B _0831_/A vssd1 vssd1 vccd1 vccd1 _0982_/B sky130_fd_sc_hd__a21o_1
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0801__B1 _0755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0829__A _1259_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0548__B _0548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0564__A _0873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0474__A _0479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1036__B1 _0548_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1180_ _1035_/A _1180_/D _1065__45/Y vssd1 vssd1 vccd1 vccd1 _1180_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_13_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0964_ _0958_/X _0963_/Y _0831_/X vssd1 vssd1 vccd1 vccd1 _0965_/B sky130_fd_sc_hd__a21o_1
X_0895_ _1275_/Q _0895_/B vssd1 vssd1 vccd1 vccd1 _1275_/D sky130_fd_sc_hd__xnor2_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_GATE_N
+ _1099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0469__A _1363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0932__A _1290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0680_ _1328_/Q vssd1 vssd1 vccd1 vccd1 _1327_/D sky130_fd_sc_hd__inv_2
XFILLER_10_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1301_ _1116_/X _1301_/D _0462__19/Y vssd1 vssd1 vccd1 vccd1 _1301_/Q sky130_fd_sc_hd__dfrtp_2
X_1232_ _1357_/A _1232_/D fanout57/X vssd1 vssd1 vccd1 vccd1 _1232_/Q sky130_fd_sc_hd__dfstp_1
X_1163_ _1163_/CLK _1163_/D fanout50/X vssd1 vssd1 vccd1 vccd1 _1163_/Q sky130_fd_sc_hd__dfrtp_1
X_1094_ _1097_/A vssd1 vssd1 vccd1 vccd1 _1094_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0947_ _1298_/Q _1297_/Q vssd1 vssd1 vccd1 vccd1 _0947_/Y sky130_fd_sc_hd__xnor2_2
X_0878_ _1045_/A _0865_/X _0877_/X vssd1 vssd1 vccd1 vccd1 _0879_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0456__14 _0448__6/A vssd1 vssd1 vccd1 vccd1 _0456__14/Y sky130_fd_sc_hd__inv_2
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0646__B _0646_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0662__A _1294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0801_ _0796_/B _0800_/X _0755_/X vssd1 vssd1 vccd1 vccd1 _0802_/B sky130_fd_sc_hd__o21ai_1
X_0663_ _1293_/Q vssd1 vssd1 vccd1 vccd1 _1294_/D sky130_fd_sc_hd__inv_2
X_0594_ _1175_/Q vssd1 vssd1 vccd1 vccd1 _1174_/D sky130_fd_sc_hd__inv_2
X_0732_ _1188_/Q _1187_/Q _0735_/B _0728_/B vssd1 vssd1 vccd1 vccd1 _0733_/B sky130_fd_sc_hd__a31o_1
XFILLER_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1146_ _1146_/A _1146_/B vssd1 vssd1 vccd1 vccd1 _1146_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__0556__B _0557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1215_ _1042_/B _1215_/D _0481_/Y vssd1 vssd1 vccd1 vccd1 _1215_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__0837__A _1259_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf _1318_/Q _1015_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
X_1077_ _1077_/A vssd1 vssd1 vccd1 vccd1 _1077_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1350__RESET_B fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0482__A _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1000_ _0960_/C _0996_/Y _0755_/A vssd1 vssd1 vccd1 vccd1 _1001_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0977__A2 _1316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0715_ _0755_/A vssd1 vssd1 vccd1 vccd1 _0831_/A sky130_fd_sc_hd__inv_4
X_0577_ _1132_/A _0577_/B vssd1 vssd1 vccd1 vccd1 _1169_/D sky130_fd_sc_hd__xor2_4
X_0646_ _1264_/Q _0646_/B vssd1 vssd1 vccd1 vccd1 _1264_/D sky130_fd_sc_hd__xor2_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0567__A _1135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput24 _1369_/X vssd1 vssd1 vccd1 vccd1 fb1_Q[1] sky130_fd_sc_hd__buf_2
Xoutput13 _1358_/X vssd1 vssd1 vccd1 vccd1 cclk_Q[0] sky130_fd_sc_hd__clkbuf_1
XANTENNA__1176__CLK _1035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0477__A _0479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0940__A _1290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0500_ _1105_/B _0548_/B vssd1 vssd1 vccd1 vccd1 _1148_/D sky130_fd_sc_hd__xnor2_1
XTAP_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0537__D _0873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0629_ _1240_/Q vssd1 vssd1 vccd1 vccd1 _1241_/D sky130_fd_sc_hd__clkinv_2
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0877__A1 _0546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0980_ _1317_/Q _0980_/B vssd1 vssd1 vccd1 vccd1 _0980_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__1341__CLK _0560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0548__C _0548_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1141__65 _1141__65/A vssd1 vssd1 vccd1 vccd1 _1141__65/Y sky130_fd_sc_hd__inv_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0580__A _1130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
+ _1183_/Q _0777_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout59_A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1214__CLK _0560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0755__A _0755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1036__A1 _0546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0492__26 _1049__32/A vssd1 vssd1 vccd1 vccd1 _0492__26/Y sky130_fd_sc_hd__inv_2
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0894_ _0888_/X _0893_/Y _0831_/X vssd1 vssd1 vccd1 vccd1 _0895_/B sky130_fd_sc_hd__a21o_1
X_0963_ _1314_/Q _1313_/Q _1312_/Q _0970_/B vssd1 vssd1 vccd1 vccd1 _0963_/Y sky130_fd_sc_hd__nand4_1
XFILLER_9_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0575__A _1045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_TE_B _0947_/Y vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0485__A _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0932__B _1348_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1300_ _0868_/B _1300_/D _1115__52/Y vssd1 vssd1 vccd1 vccd1 _1300_/Q sky130_fd_sc_hd__dfrtp_2
X_1162_ _1360_/A _1162_/D fanout44/X vssd1 vssd1 vccd1 vccd1 _1162_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1231_ _1357_/A _1231_/D fanout56/X vssd1 vssd1 vccd1 vccd1 _1231_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1093_ _1139_/A _1139_/B vssd1 vssd1 vccd1 vccd1 _1093_/X sky130_fd_sc_hd__xor2_2
XANTENNA__1003__B _1352_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0877_ _0546_/A _0872_/X _0874_/X _0876_/X _0868_/A vssd1 vssd1 vccd1 vccd1 _0877_/X
+ sky130_fd_sc_hd__o311a_1
X_0946_ _1296_/Q _1295_/Q vssd1 vssd1 vccd1 vccd1 _0946_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1104__A _1105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0943__A _1013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0800_ _1222_/Q _0800_/B vssd1 vssd1 vccd1 vccd1 _0800_/X sky130_fd_sc_hd__and2b_1
XFILLER_6_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0731_ _0755_/A vssd1 vssd1 vccd1 vccd1 _1013_/A sky130_fd_sc_hd__buf_4
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0662_ _1294_/Q vssd1 vssd1 vccd1 vccd1 _1293_/D sky130_fd_sc_hd__inv_2
X_0593_ _0593_/A vssd1 vssd1 vccd1 vccd1 _1355_/D sky130_fd_sc_hd__inv_2
X_1214_ _0560_/A _1214_/D _1076_/Y vssd1 vssd1 vccd1 vccd1 _1214_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1076_ _1077_/A vssd1 vssd1 vccd1 vccd1 _1076_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0929_ _1285_/Q _0929_/B vssd1 vssd1 vccd1 vccd1 _1285_/D sky130_fd_sc_hd__xnor2_1
XFILLER_1_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output22_A _1367_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0714_ _0714_/A vssd1 vssd1 vccd1 vccd1 _0755_/A sky130_fd_sc_hd__buf_4
X_0645_ _1263_/Q _0646_/B vssd1 vssd1 vccd1 vccd1 _1263_/D sky130_fd_sc_hd__xor2_1
X_0576_ _1132_/B _0577_/B vssd1 vssd1 vccd1 vccd1 _1168_/D sky130_fd_sc_hd__xor2_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0583__A _0590_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1128_ _1128_/A _1128_/B vssd1 vssd1 vccd1 vccd1 _1128_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_22_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput25 _1370_/X vssd1 vssd1 vccd1 vccd1 read_out_I[0] sky130_fd_sc_hd__buf_2
Xoutput14 _1359_/X vssd1 vssd1 vccd1 vccd1 cclk_Q[1] sky130_fd_sc_hd__buf_2
XFILLER_1_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0940__B _1275_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1270__CLK _0542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0628_ _1241_/Q vssd1 vssd1 vccd1 vccd1 _1240_/D sky130_fd_sc_hd__inv_2
XFILLER_8_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0559_ _0568_/B _1042_/C vssd1 vssd1 vccd1 vccd1 _0865_/C sky130_fd_sc_hd__nand2_1
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1293__CLK _0581_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0488__A _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1099_/A fanout58/X vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__1112__A _1133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1039__C1 _1035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf _1280_/Q _0947_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_9_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1163__RESET_B fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0580__B _1130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0861__A _1034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1107__A _1128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1189__CLK fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0681__A _1327_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0893_ _1278_/Q _1277_/Q _1276_/Q _0900_/B vssd1 vssd1 vccd1 vccd1 _0893_/Y sky130_fd_sc_hd__nand4_1
X_0962_ _1317_/Q _1316_/Q _1315_/Q _0980_/B vssd1 vssd1 vccd1 vccd1 _0970_/B sky130_fd_sc_hd__and4_2
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1168_/CLK fanout42/X vssd1 vssd1 vccd1 vccd1 _1366_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_9_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1017__A _1334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0538__A1 _1045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0575__B _0590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0591__A _1128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1331__CLK _0590_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1161_ _1161_/CLK _1161_/D fanout44/X vssd1 vssd1 vccd1 vccd1 _1161_/Q sky130_fd_sc_hd__dfrtp_1
X_1092_ _1097_/A vssd1 vssd1 vccd1 vccd1 _1092_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1230_ _1357_/A _1230_/D fanout56/X vssd1 vssd1 vccd1 vccd1 _1230_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1204__CLK _0590_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0945_ _1294_/Q _1293_/Q vssd1 vssd1 vccd1 vccd1 _0945_/Y sky130_fd_sc_hd__xnor2_2
X_0876_ _1042_/B _0873_/B _0862_/Y _0875_/X vssd1 vssd1 vccd1 vccd1 _0876_/X sky130_fd_sc_hd__a31o_1
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1354__CLK input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1102__47 _1117__53/A vssd1 vssd1 vccd1 vccd1 _1266_/CLK sky130_fd_sc_hd__inv_2
X_1359_ _1359_/A vssd1 vssd1 vccd1 vccd1 _1359_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_TE_B
+ _0771_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1266__RESET_B fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0462__19 _0467__24/A vssd1 vssd1 vccd1 vccd1 _0462__19/Y sky130_fd_sc_hd__inv_2
XANTENNA__0943__B _1290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f__0308_ clkbuf_0__0308_/X vssd1 vssd1 vccd1 vccd1 _0467__24/A sky130_fd_sc_hd__clkbuf_16
X_0661_ _1291_/Q vssd1 vssd1 vccd1 vccd1 _1292_/D sky130_fd_sc_hd__inv_2
XFILLER_11_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0730_ _1185_/Q _0730_/B vssd1 vssd1 vccd1 vccd1 _1185_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__1227__CLK _1357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1213_ _0862_/A _1213_/D _1075_/Y vssd1 vssd1 vccd1 vccd1 _1213_/Q sky130_fd_sc_hd__dfrtp_1
X_0592_ _1128_/A _0592_/B vssd1 vssd1 vccd1 vccd1 _1173_/D sky130_fd_sc_hd__xnor2_1
XFILLER_3_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1014__B _1327_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1144_ _1144_/A _1144_/B vssd1 vssd1 vccd1 vccd1 _1144_/Y sky130_fd_sc_hd__xnor2_1
X_1075_ _1077_/A vssd1 vssd1 vccd1 vccd1 _1075_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0859_ _0859_/A _0859_/B vssd1 vssd1 vccd1 vccd1 _0860_/A sky130_fd_sc_hd__or2_1
XFILLER_20_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0928_ _0998_/A _0928_/B vssd1 vssd1 vccd1 vccd1 _0929_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0644_ _0879_/A _0644_/B _0644_/C _0644_/D vssd1 vssd1 vccd1 vccd1 _0646_/B sky130_fd_sc_hd__and4_4
X_0713_ _1185_/Q _1184_/Q _1183_/Q _0724_/B vssd1 vssd1 vccd1 vccd1 _0713_/Y sky130_fd_sc_hd__nand4_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0575_ _1045_/A _0590_/B vssd1 vssd1 vccd1 vccd1 _0577_/B sky130_fd_sc_hd__nor2_2
XANTENNA__0898__B1 _0755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1188__RESET_B fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0583__B _0644_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput15 _1360_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_I[0] sky130_fd_sc_hd__clkbuf_1
Xoutput26 _1371_/X vssd1 vssd1 vccd1 vccd1 read_out_I[1] sky130_fd_sc_hd__buf_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0684__A _1332_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0558_ _0873_/A _0874_/D vssd1 vssd1 vccd1 vccd1 _1042_/C sky130_fd_sc_hd__nand2_1
X_0627_ _1238_/Q vssd1 vssd1 vccd1 vccd1 _1239_/D sky130_fd_sc_hd__inv_2
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0594__A _1175_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0489_ _0593_/A vssd1 vssd1 vccd1 vccd1 _0489_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1112__B _1133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1099_/A fanout58/X vssd1 vssd1 vccd1 vccd1 _1367_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1__f_w0.cclk_I clkbuf_0_w0.cclk_I/X vssd1 vssd1 vccd1 vccd1 _1356_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input6_A phi1b_dig_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1117__53 _1117__53/A vssd1 vssd1 vccd1 vccd1 _1117__53/Y sky130_fd_sc_hd__inv_2
XFILLER_15_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1260__CLK input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1107__B _1128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1123__56 _1140__64/A vssd1 vssd1 vccd1 vccd1 _1123__56/Y sky130_fd_sc_hd__inv_2
X_0961_ _1320_/Q _1319_/Q _1318_/Q _0990_/B vssd1 vssd1 vccd1 vccd1 _0980_/B sky130_fd_sc_hd__and4_1
X_0892_ _1281_/Q _1280_/Q _1279_/Q _0910_/B vssd1 vssd1 vccd1 vccd1 _0900_/B sky130_fd_sc_hd__and4_1
XFILLER_9_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1017__B _1333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0538__A2 _0590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1375_ _1375_/A vssd1 vssd1 vccd1 vccd1 _1375_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0591__B _0592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1050__33 _1052__35/A vssd1 vssd1 vccd1 vccd1 _1157_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout50 fanout51/X vssd1 vssd1 vccd1 vccd1 fanout50/X sky130_fd_sc_hd__clkbuf_4
XFILLER_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1118__A _1139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0957__A _1316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1160_ _1360_/A _1160_/D fanout44/X vssd1 vssd1 vccd1 vccd1 _1160_/Q sky130_fd_sc_hd__dfrtp_1
X_1091_ _1137_/A _1137_/B vssd1 vssd1 vccd1 vccd1 _1091_/X sky130_fd_sc_hd__xor2_1
XANTENNA__0692__A _1340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0944_ _1292_/Q _1291_/Q vssd1 vssd1 vccd1 vccd1 _0944_/Y sky130_fd_sc_hd__xnor2_2
X_0875_ _0560_/A _0532_/Y _0868_/B _1042_/A vssd1 vssd1 vccd1 vccd1 _0875_/X sky130_fd_sc_hd__a31o_1
X_1358_ _1358_/A vssd1 vssd1 vccd1 vccd1 _1358_/X sky130_fd_sc_hd__buf_2
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1289_ _1325_/CLK _1289_/D fanout48/X vssd1 vssd1 vccd1 vccd1 _1289_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_24_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__0307_ clkbuf_0__0307_/X vssd1 vssd1 vccd1 vccd1 _0451__9/A sky130_fd_sc_hd__clkbuf_16
X_0660_ _1292_/Q vssd1 vssd1 vccd1 vccd1 _1291_/D sky130_fd_sc_hd__inv_2
X_0591_ _1128_/B _0592_/B vssd1 vssd1 vccd1 vccd1 _1172_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0687__A _1333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1212_ _0873_/A _1212_/D _0482_/Y vssd1 vssd1 vccd1 vccd1 _1212_/Q sky130_fd_sc_hd__dfrtp_1
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
+ _1218_/Q _0849_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_19_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1074_ _1077_/A vssd1 vssd1 vccd1 vccd1 _1074_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0927_ _0926_/Y _0890_/C _1286_/Q vssd1 vssd1 vccd1 vccd1 _0928_/B sky130_fd_sc_hd__mux2_1
X_0858_ _1260_/D _1261_/Q vssd1 vssd1 vccd1 vccd1 _0859_/B sky130_fd_sc_hd__and2b_1
XANTENNA__0597__A _1176_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0789_ _1221_/Q _1220_/Q _1219_/Q _0796_/B vssd1 vssd1 vccd1 vccd1 _0789_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_1__f_clk_master clkbuf_0_clk_master/X vssd1 vssd1 vccd1 vccd1 _1168_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0954__B _1352_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0574_ _0879_/A vssd1 vssd1 vccd1 vccd1 _0590_/C sky130_fd_sc_hd__inv_2
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0712_ _1188_/Q _1187_/Q _1186_/Q _0735_/B vssd1 vssd1 vccd1 vccd1 _0724_/B sky130_fd_sc_hd__and4_1
X_0643_ _0643_/A vssd1 vssd1 vccd1 vccd1 _0643_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1126_ _1146_/A _1146_/B vssd1 vssd1 vccd1 vccd1 _1126_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput16 _1361_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_I[1] sky130_fd_sc_hd__buf_2
Xoutput27 _1372_/X vssd1 vssd1 vccd1 vccd1 read_out_Q[0] sky130_fd_sc_hd__buf_2
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1217__CLK _0546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0949__B _1301_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0626_ _1239_/Q vssd1 vssd1 vccd1 vccd1 _1238_/D sky130_fd_sc_hd__inv_2
X_0557_ _1139_/B _0557_/B vssd1 vssd1 vccd1 vccd1 _1161_/D sky130_fd_sc_hd__xnor2_1
XFILLER_26_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1109_ _1130_/A _1130_/B vssd1 vssd1 vccd1 vccd1 _1109_/Y sky130_fd_sc_hd__xnor2_1
X_0488_ _0593_/A vssd1 vssd1 vccd1 vccd1 _0488_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0740__B1 _0998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1057__39 _1058__40/A vssd1 vssd1 vccd1 vccd1 _1169_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0769__B _1013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0785__A _1259_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0722__B1 _0998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0609_ _1204_/Q vssd1 vssd1 vccd1 vccd1 _1205_/D sky130_fd_sc_hd__inv_2
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0962__B _1316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0960_ _1322_/Q _1321_/Q _0960_/C vssd1 vssd1 vccd1 vccd1 _0990_/B sky130_fd_sc_hd__and3_1
X_0891_ _1284_/Q _1283_/Q _1282_/Q _0920_/B vssd1 vssd1 vccd1 vccd1 _0910_/B sky130_fd_sc_hd__and4_1
X_1374_ _1374_/A vssd1 vssd1 vccd1 vccd1 _1374_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1353__RESET_B fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout51 input9/X vssd1 vssd1 vccd1 vccd1 fanout51/X sky130_fd_sc_hd__clkbuf_4
Xfanout40 _1363_/A vssd1 vssd1 vccd1 vccd1 _1099_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1118__B _1139_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0957__B _1315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0973__A _1316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1090_ _1097_/A vssd1 vssd1 vccd1 vccd1 _1090_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0874_ _1035_/C _0871_/Y _0874_/C _0874_/D vssd1 vssd1 vccd1 vccd1 _0874_/X sky130_fd_sc_hd__and4bb_1
XFILLER_9_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0943_ _1013_/A _1290_/Q vssd1 vssd1 vccd1 vccd1 _1290_/D sky130_fd_sc_hd__xor2_1
X_1357_ _1357_/A vssd1 vssd1 vccd1 vccd1 _1357_/X sky130_fd_sc_hd__clkbuf_1
X_1145__4 _1053_/A vssd1 vssd1 vccd1 vccd1 _1145__4/Y sky130_fd_sc_hd__inv_2
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1362_/A fanout42/X vssd1 vssd1 vccd1 vccd1 _1368_/A sky130_fd_sc_hd__dlrtn_1
X_1288_ _1326_/CLK _1288_/D fanout48/X vssd1 vssd1 vccd1 vccd1 _1288_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf _1315_/Q _1018_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__0306_ clkbuf_0__0306_/X vssd1 vssd1 vccd1 vccd1 _1122_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0590_ _0868_/A _0590_/B _0590_/C _0644_/B vssd1 vssd1 vccd1 vccd1 _0592_/B sky130_fd_sc_hd__or4_4
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1142_ _1142_/A _1142_/B vssd1 vssd1 vccd1 vccd1 _1142_/Y sky130_fd_sc_hd__xnor2_1
X_1211_ _1035_/B _1211_/D _1074_/Y vssd1 vssd1 vccd1 vccd1 _1211_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1073_ _1077_/A vssd1 vssd1 vccd1 vccd1 _1073_/Y sky130_fd_sc_hd__inv_2
X_0857_ _0857_/A vssd1 vssd1 vccd1 vccd1 _0859_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0926_ _0926_/A vssd1 vssd1 vccd1 vccd1 _0926_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1011__C1 _0831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0788_ _1224_/Q _1223_/Q _1222_/Q _0806_/B vssd1 vssd1 vccd1 vccd1 _0796_/B sky130_fd_sc_hd__and4_1
XFILLER_25_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0452__10 _0451__9/A vssd1 vssd1 vccd1 vccd1 _0452__10/Y sky130_fd_sc_hd__inv_2
XFILLER_8_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0788__A _1224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0970__B _0970_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0711_ _1191_/Q _1190_/Q _1189_/Q _0745_/B vssd1 vssd1 vccd1 vccd1 _0735_/B sky130_fd_sc_hd__and4_1
X_0573_ _1132_/A _1132_/B vssd1 vssd1 vccd1 vccd1 _0879_/A sky130_fd_sc_hd__xnor2_4
X_0642_ _1263_/Q _1264_/Q vssd1 vssd1 vccd1 vccd1 _0643_/A sky130_fd_sc_hd__xor2_4
XFILLER_3_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1041__B _1041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0909_ _1279_/Q _0909_/B vssd1 vssd1 vccd1 vccd1 _1279_/D sky130_fd_sc_hd__xnor2_1
Xoutput17 _1362_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_Q[0] sky130_fd_sc_hd__clkbuf_1
Xoutput28 _1373_/X vssd1 vssd1 vccd1 vccd1 read_out_Q[1] sky130_fd_sc_hd__buf_2
Xclkbuf_0__0308_ _0458_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0308_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1138__63 _1141__65/A vssd1 vssd1 vccd1 vccd1 _1138__63/Y sky130_fd_sc_hd__inv_2
XANTENNA__1142__A _1142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0625_ _1236_/Q vssd1 vssd1 vccd1 vccd1 _1237_/D sky130_fd_sc_hd__clkinv_2
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0487_ _0593_/A vssd1 vssd1 vccd1 vccd1 _0487_/Y sky130_fd_sc_hd__inv_2
X_0556_ _1139_/A _0557_/B vssd1 vssd1 vccd1 vccd1 _1160_/D sky130_fd_sc_hd__xnor2_1
XFILLER_27_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1039_ _0865_/A _0874_/D _1035_/C _1038_/Y _1035_/A vssd1 vssd1 vccd1 vccd1 _1040_/B
+ sky130_fd_sc_hd__o311a_1
XANTENNA__0891__A _1284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1334__CLK _1045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1039__A2 _0874_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1207__CLK _1045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0608_ _1205_/Q vssd1 vssd1 vccd1 vccd1 _1204_/D sky130_fd_sc_hd__clkinv_2
XFILLER_27_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0539_ _1041_/A _0590_/B _0538_/Y vssd1 vssd1 vccd1 vccd1 _0541_/B sky130_fd_sc_hd__o21ai_1
XFILLER_27_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
+ _1226_/Q _0841_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[0\].w1.ro_block_Q.ro_pol.tribuf.t_buf _0855_/X _0700_/Y vssd1
+ vssd1 vccd1 vccd1 _1372_/A sky130_fd_sc_hd__ebufn_4
XFILLER_14_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0962__C _1315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0890_ _1286_/Q _1285_/Q _0890_/C vssd1 vssd1 vccd1 vccd1 _0920_/B sky130_fd_sc_hd__and3_1
XFILLER_5_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1373_ _1373_/A vssd1 vssd1 vccd1 vccd1 _1373_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1079_/A fanout57/X vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__dlrtn_1
X_0459__16 _0490__25/A vssd1 vssd1 vccd1 vccd1 _0459__16/Y sky130_fd_sc_hd__inv_2
XANTENNA__0555__S _0560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout52 fanout53/X vssd1 vssd1 vccd1 vccd1 fanout52/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout41 fanout42/X vssd1 vssd1 vccd1 vccd1 fanout41/X sky130_fd_sc_hd__buf_2
XANTENNA__0782__C _1224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0973__B _0973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0873_ _0873_/A _0873_/B vssd1 vssd1 vccd1 vccd1 _0874_/C sky130_fd_sc_hd__nand2_1
X_0942_ _1289_/Q _0942_/B vssd1 vssd1 vccd1 vccd1 _1289_/D sky130_fd_sc_hd__xnor2_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1356_ _1356_/A vssd1 vssd1 vccd1 vccd1 _1356_/X sky130_fd_sc_hd__buf_2
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1287_ _1358_/A _1287_/D fanout47/X vssd1 vssd1 vccd1 vccd1 _1287_/Q sky130_fd_sc_hd__dfrtp_1
X_1110__50 _1117__53/A vssd1 vssd1 vccd1 vccd1 _1110__50/Y sky130_fd_sc_hd__inv_2
XFILLER_3_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1168_/CLK fanout42/X vssd1 vssd1 vccd1 vccd1 _1366_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_8_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__0305_ clkbuf_0__0305_/X vssd1 vssd1 vccd1 vccd1 _1140__64/A sky130_fd_sc_hd__clkbuf_16
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1072_ _1077_/A vssd1 vssd1 vccd1 vccd1 _1072_/Y sky130_fd_sc_hd__inv_2
X_1210_ _0874_/D _1210_/D _0483_/Y vssd1 vssd1 vccd1 vccd1 _1210_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0856_ _1261_/Q _1260_/D vssd1 vssd1 vccd1 vccd1 _0857_/A sky130_fd_sc_hd__and2b_1
X_0787_ _1227_/Q _1226_/Q _1225_/Q _0816_/B vssd1 vssd1 vccd1 vccd1 _0806_/B sky130_fd_sc_hd__and4_1
X_0925_ _1284_/Q _0925_/B vssd1 vssd1 vccd1 vccd1 _1284_/D sky130_fd_sc_hd__xnor2_1
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1339_ _1139_/X _1339_/D _0450__8/Y vssd1 vssd1 vccd1 vccd1 _1339_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0641_ _1252_/Q vssd1 vssd1 vccd1 vccd1 _1253_/D sky130_fd_sc_hd__inv_2
XANTENNA__0979__A _1315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0710_ _1193_/Q _1192_/Q _0710_/C vssd1 vssd1 vccd1 vccd1 _0745_/B sky130_fd_sc_hd__and3_1
XANTENNA__1240__CLK _0590_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0572_ _1168_/Q vssd1 vssd1 vccd1 vccd1 _1132_/B sky130_fd_sc_hd__buf_6
X_1124_ _1144_/A _1144_/B vssd1 vssd1 vccd1 vccd1 _1124_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0807__B1 _0716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0908_ _0998_/A _0908_/B vssd1 vssd1 vccd1 vccd1 _0909_/B sky130_fd_sc_hd__nand2_1
X_0839_ _1232_/Q _0839_/B vssd1 vssd1 vccd1 vccd1 _1232_/D sky130_fd_sc_hd__xnor2_1
Xoutput18 _1363_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_Q[1] sky130_fd_sc_hd__buf_2
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput29 _1374_/X vssd1 vssd1 vccd1 vccd1 sin_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0889__A _1290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0__0307_ _0447_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0307_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_5_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout32_A _1357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1142__B _1142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[0\].w1.ro_block_Q.ro_pol.tribuf.t_buf_TE_B _0700_/Y vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0624_ _1237_/Q vssd1 vssd1 vccd1 vccd1 _1236_/D sky130_fd_sc_hd__inv_2
X_0486_ _0593_/A vssd1 vssd1 vccd1 vccd1 _0486_/Y sky130_fd_sc_hd__inv_2
X_0555_ _0554_/Y _0862_/A _0560_/B vssd1 vssd1 vccd1 vccd1 _0557_/B sky130_fd_sc_hd__mux2_2
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf _1277_/Q _0950_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_26_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1107_ _1128_/A _1128_/B vssd1 vssd1 vccd1 vccd1 _1107_/Y sky130_fd_sc_hd__xnor2_1
X_1038_ _1042_/A _0874_/D _0547_/X _0873_/A vssd1 vssd1 vccd1 vccd1 _1038_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_22_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1347__RESET_B fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1039__A3 _1035_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1137__B _1137_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0992__A _1319_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_A _1280_/Q vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1047__30 _1049__32/A vssd1 vssd1 vccd1 vccd1 _1150_/CLK sky130_fd_sc_hd__inv_2
X_0607_ _1202_/Q vssd1 vssd1 vccd1 vccd1 _1203_/D sky130_fd_sc_hd__inv_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0538_ _1045_/A _0590_/B _1041_/A vssd1 vssd1 vccd1 vccd1 _0538_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__0886__B _1282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0469_ _1363_/A vssd1 vssd1 vccd1 vccd1 _0479_/A sky130_fd_sc_hd__buf_4
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1301__CLK _1116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1372_ _1372_/A vssd1 vssd1 vccd1 vccd1 _1372_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1031__A_N _1353_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A comp_high_Q[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0897__A _1277_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1099_/A fanout58/X vssd1 vssd1 vccd1 vccd1 _1367_/A sky130_fd_sc_hd__dlrtn_1
Xfanout53 fanout54/X vssd1 vssd1 vccd1 vccd1 fanout53/X sky130_fd_sc_hd__buf_4
XFILLER_13_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout42 fanout51/X vssd1 vssd1 vccd1 vccd1 fanout42/X sky130_fd_sc_hd__buf_2
XFILLER_11_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout31 fanout34/X vssd1 vssd1 vccd1 vccd1 fanout31/X sky130_fd_sc_hd__buf_2
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0957__D _0973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0941_ _0888_/X _0893_/Y _0940_/X _0831_/A vssd1 vssd1 vccd1 vccd1 _0942_/B sky130_fd_sc_hd__a211o_1
X_0872_ _0862_/Y _0871_/Y _0560_/A vssd1 vssd1 vccd1 vccd1 _0872_/X sky130_fd_sc_hd__o21a_1
X_1355_ _1355_/CLK _1355_/D fanout53/X vssd1 vssd1 vccd1 vccd1 _1363_/A sky130_fd_sc_hd__dfrtp_4
X_1286_ _1358_/A _1286_/D fanout47/X vssd1 vssd1 vccd1 vccd1 _1286_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0907__A2 _1280_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f__0304_ clkbuf_0__0304_/X vssd1 vssd1 vccd1 vccd1 _1120__55/A sky130_fd_sc_hd__clkbuf_16
XFILLER_7_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0914__A_N _1282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1071_ _1077_/A vssd1 vssd1 vccd1 vccd1 _1071_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
+ _1188_/Q _0772_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_0924_ _0920_/B _0923_/Y _0755_/X vssd1 vssd1 vccd1 vccd1 _0925_/B sky130_fd_sc_hd__o21ai_1
X_0855_ _0855_/A vssd1 vssd1 vccd1 vccd1 _0855_/X sky130_fd_sc_hd__clkbuf_1
X_0786_ _1229_/Q _1228_/Q _0786_/C vssd1 vssd1 vccd1 vccd1 _0816_/B sky130_fd_sc_hd__and3_1
X_1338_ _1035_/B _1338_/D _1138__63/Y vssd1 vssd1 vccd1 vccd1 _1338_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1071__A _1077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1269_ _1103_/Y _1269_/D _1148_/CLK vssd1 vssd1 vccd1 vccd1 _1269_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_10_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0761__B1 _0716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1192__CLK fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0571_ _1169_/Q vssd1 vssd1 vccd1 vccd1 _1132_/A sky130_fd_sc_hd__buf_6
X_0640_ _1253_/Q vssd1 vssd1 vccd1 vccd1 _1252_/D sky130_fd_sc_hd__inv_2
XFILLER_11_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0907_ _1281_/Q _1280_/Q _0910_/B _0904_/B vssd1 vssd1 vccd1 vccd1 _0908_/B sky130_fd_sc_hd__a31o_1
Xoutput19 _1364_/X vssd1 vssd1 vccd1 vccd1 cos_out[0] sky130_fd_sc_hd__buf_2
Xclkbuf_0__0306_ _0445_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0306_/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__0991__B1 _0831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0838_ _0784_/X _0789_/Y _0837_/X _0831_/A vssd1 vssd1 vccd1 vccd1 _0839_/B sky130_fd_sc_hd__a211o_1
XANTENNA__0889__B _1348_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0769_ _1197_/Q _1013_/A vssd1 vssd1 vccd1 vccd1 _1197_/D sky130_fd_sc_hd__xor2_1
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0554_ _1035_/C _0866_/B vssd1 vssd1 vccd1 vccd1 _0554_/Y sky130_fd_sc_hd__nor2_1
X_0623_ _1234_/Q vssd1 vssd1 vccd1 vccd1 _1235_/D sky130_fd_sc_hd__inv_2
XANTENNA__0725__B1 _0716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0485_ _0593_/A vssd1 vssd1 vccd1 vccd1 _0485_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1037_ _0871_/Y _1035_/X _1036_/X _0873_/B vssd1 vssd1 vccd1 vccd1 _1040_/A sky130_fd_sc_hd__o22a_1
XANTENNA__0891__C _1282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0964__B1 _0831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1316__RESET_B fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1230__CLK _1357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0513__A _1144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0606_ _1203_/Q vssd1 vssd1 vccd1 vccd1 _1202_/D sky130_fd_sc_hd__clkinv_2
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0537_ _0560_/A _0560_/B _0568_/B _0873_/B vssd1 vssd1 vccd1 vccd1 _0590_/B sky130_fd_sc_hd__or4_4
XFILLER_26_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1253__CLK _1098_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0468_ _1099_/A vssd1 vssd1 vccd1 vccd1 _1034_/B sky130_fd_sc_hd__inv_2
XFILLER_23_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1131__60 _1141__65/A vssd1 vssd1 vccd1 vccd1 _1131__60/Y sky130_fd_sc_hd__inv_2
XFILLER_17_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1371_ _1371_/A vssd1 vssd1 vccd1 vccd1 _1371_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0508__A _0542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1074__A _1077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout54 input9/X vssd1 vssd1 vccd1 vccd1 fanout54/X sky130_fd_sc_hd__buf_4
Xfanout43 fanout51/X vssd1 vssd1 vccd1 vccd1 fanout43/X sky130_fd_sc_hd__clkbuf_4
Xfanout32 _1357_/A vssd1 vssd1 vccd1 vccd1 _1359_/A sky130_fd_sc_hd__buf_2
XFILLER_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_A
+ _1185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0940_ _1290_/Q _1275_/Q vssd1 vssd1 vccd1 vccd1 _0940_/X sky130_fd_sc_hd__xor2_1
X_0871_ _0873_/A _0873_/B vssd1 vssd1 vccd1 vccd1 _0871_/Y sky130_fd_sc_hd__nor2_2
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0998__A _0998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1354_ input5/X _1354_/D fanout53/X vssd1 vssd1 vccd1 vccd1 _1354_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1285_ _1358_/A _1285_/D fanout47/X vssd1 vssd1 vccd1 vccd1 _1285_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0464__21 _0467__24/A vssd1 vssd1 vccd1 vccd1 _0464__21/Y sky130_fd_sc_hd__inv_2
XFILLER_20_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1069__A _1077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout55_A fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1253__RESET_B _1034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1070_ _1077_/A vssd1 vssd1 vccd1 vccd1 _1070_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_TE_B
+ _0772_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0923_ _1286_/Q _1285_/Q _0926_/A vssd1 vssd1 vccd1 vccd1 _0923_/Y sky130_fd_sc_hd__nor3_1
X_0854_ _0854_/A _0854_/B vssd1 vssd1 vccd1 vccd1 _0855_/A sky130_fd_sc_hd__or2_1
XANTENNA__0521__A _1133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0785_ _1259_/D _1233_/Q _1231_/Q _1230_/Q vssd1 vssd1 vccd1 vccd1 _0786_/C sky130_fd_sc_hd__and4_1
X_1337_ _1137_/X _1337_/D _0451__9/Y vssd1 vssd1 vccd1 vccd1 _1337_/Q sky130_fd_sc_hd__dfrtp_4
X_1268_ _0542_/B _1268_/D _1148_/CLK vssd1 vssd1 vccd1 vccd1 _1268_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1199_ _0643_/Y _1199_/D _1068_/Y vssd1 vssd1 vccd1 vccd1 _1199_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1362_/A fanout41/X vssd1 vssd1 vccd1 vccd1 _1368_/A sky130_fd_sc_hd__dlrtn_1
X_0570_ _1133_/A _0570_/B vssd1 vssd1 vccd1 vccd1 _1167_/D sky130_fd_sc_hd__xnor2_1
XFILLER_3_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1122_ _1122_/A vssd1 vssd1 vccd1 vccd1 _1122_/X sky130_fd_sc_hd__buf_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1053_ _1053_/A vssd1 vssd1 vccd1 vccd1 _1053_/X sky130_fd_sc_hd__buf_1
X_0837_ _1259_/D _1218_/Q vssd1 vssd1 vccd1 vccd1 _0837_/X sky130_fd_sc_hd__xor2_1
X_0906_ _1278_/Q _0906_/B vssd1 vssd1 vccd1 vccd1 _1278_/D sky130_fd_sc_hd__xnor2_1
Xclkbuf_0__0305_ _1122_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0305_/X sky130_fd_sc_hd__clkbuf_16
X_0699_ _1345_/Q vssd1 vssd1 vccd1 vccd1 _1346_/D sky130_fd_sc_hd__inv_2
X_0768_ _1196_/Q _0768_/B vssd1 vssd1 vccd1 vccd1 _1196_/D sky130_fd_sc_hd__xnor2_1
XFILLER_25_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1082__A _1128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf_A _1275_/Q vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0904__A_N _1279_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0553_ _0560_/A _0862_/A vssd1 vssd1 vccd1 vccd1 _0866_/B sky130_fd_sc_hd__nor2_1
X_0484_ _0593_/A vssd1 vssd1 vccd1 vccd1 _0484_/Y sky130_fd_sc_hd__inv_2
X_0622_ _1235_/Q vssd1 vssd1 vccd1 vccd1 _1234_/D sky130_fd_sc_hd__clkinv_2
XFILLER_3_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1105_ _1105_/A _1105_/B vssd1 vssd1 vccd1 vccd1 _1105_/Y sky130_fd_sc_hd__xnor2_1
X_1036_ _0546_/A _0568_/B _0548_/C vssd1 vssd1 vccd1 vccd1 _1036_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1077__A _1077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0513__B _1144_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0536_ _1135_/A _1135_/B vssd1 vssd1 vccd1 vccd1 _0873_/B sky130_fd_sc_hd__xor2_4
X_0605_ _1200_/Q vssd1 vssd1 vccd1 vccd1 _1201_/D sky130_fd_sc_hd__inv_2
XANTENNA__0886__D _0913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1019_ _1338_/Q _1337_/Q vssd1 vssd1 vccd1 vccd1 _1019_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_23_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1190__RESET_B fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1370_ _1370_/A vssd1 vssd1 vccd1 vccd1 _1370_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0508__B _0548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0524__A _0542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1220__CLK fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0519_ _1167_/Q vssd1 vssd1 vccd1 vccd1 _1133_/A sky130_fd_sc_hd__buf_6
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1090__A _1097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout44 fanout45/X vssd1 vssd1 vccd1 vccd1 fanout44/X sky130_fd_sc_hd__clkbuf_4
XFILLER_15_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout33 fanout34/X vssd1 vssd1 vccd1 vccd1 _1357_/A sky130_fd_sc_hd__clkbuf_4
Xfanout55 fanout59/X vssd1 vssd1 vccd1 vccd1 fanout55/X sky130_fd_sc_hd__clkbuf_4
XFILLER_23_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0870_ _0870_/A _0870_/B vssd1 vssd1 vccd1 vccd1 _1375_/A sky130_fd_sc_hd__xor2_1
XFILLER_14_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf _1312_/Q _1021_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XANTENNA__1243__CLK _1045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1353_ input5/X _1353_/D fanout54/X vssd1 vssd1 vccd1 vccd1 _1354_/D sky130_fd_sc_hd__dfrtp_1
X_1284_ _1326_/CLK _1284_/D fanout48/X vssd1 vssd1 vccd1 vccd1 _1284_/Q sky130_fd_sc_hd__dfrtp_2
X_0999_ _1321_/Q _0999_/B vssd1 vssd1 vccd1 vccd1 _1321_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__0701__B _1176_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1085__A _1097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout48_A fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1005__B1 _0831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout38/X fanout56/X vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0922_ _1283_/Q _0922_/B vssd1 vssd1 vccd1 vccd1 _1283_/D sky130_fd_sc_hd__xnor2_1
X_0853_ _1256_/D _1257_/Q vssd1 vssd1 vccd1 vccd1 _0854_/B sky130_fd_sc_hd__and2b_1
XANTENNA__1222__RESET_B fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0521__B _1133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0784_ _1220_/Q _1219_/Q _0793_/B vssd1 vssd1 vccd1 vccd1 _0784_/X sky130_fd_sc_hd__or3_1
Xinput1 comp_high_I[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
X_1336_ _0868_/B _1336_/D _1136__62/Y vssd1 vssd1 vccd1 vccd1 _1336_/Q sky130_fd_sc_hd__dfrtp_2
X_1198_ _0643_/A _1198_/D _0489_/Y vssd1 vssd1 vccd1 vccd1 _1198_/Q sky130_fd_sc_hd__dfrtp_1
X_1267_ _0548_/A _1267_/D _1362_/A vssd1 vssd1 vccd1 vccd1 _1267_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_90 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0712__A _1188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1121_ _1142_/A _1142_/B vssd1 vssd1 vccd1 vccd1 _1121_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_22_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_GATE_N
+ _1099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0767_ _0708_/X _0713_/Y _0766_/X _0831_/A vssd1 vssd1 vccd1 vccd1 _0768_/B sky130_fd_sc_hd__a211o_1
X_0905_ _0900_/B _0904_/X _0755_/X vssd1 vssd1 vccd1 vccd1 _0906_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__0532__A _0874_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0836_ _1231_/Q _0836_/B vssd1 vssd1 vccd1 vccd1 _1231_/D sky130_fd_sc_hd__xnor2_1
X_0698_ _1346_/Q vssd1 vssd1 vccd1 vccd1 _1345_/D sky130_fd_sc_hd__clkinv_2
Xclkbuf_0__0304_ _1100_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0304_/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__1363__A _1363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1082__B _1128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1319_ _1356_/A _1319_/D fanout46/X vssd1 vssd1 vccd1 vccd1 _1319_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__0707__A _1187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0874__B_N _0871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1304__CLK _0862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1059__41 _1065__45/A vssd1 vssd1 vccd1 vccd1 _1173_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0621_ _1216_/Q vssd1 vssd1 vccd1 vccd1 _1217_/D sky130_fd_sc_hd__inv_2
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0552_ _1042_/B _0873_/A vssd1 vssd1 vccd1 vccd1 _1035_/C sky130_fd_sc_hd__nor2_2
X_0483_ _0593_/A vssd1 vssd1 vccd1 vccd1 _0483_/Y sky130_fd_sc_hd__inv_2
X_1035_ _1035_/A _1035_/B _1035_/C _1035_/D vssd1 vssd1 vccd1 vccd1 _1035_/X sky130_fd_sc_hd__or4_1
X_1104_ _1105_/A _1105_/B vssd1 vssd1 vccd1 vccd1 _1104_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__0527__A _1139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1327__CLK _0644_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0819_ _1229_/Q _1228_/Q _0822_/A vssd1 vssd1 vccd1 vccd1 _0819_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__1093__A _1139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
+ _1223_/Q _0844_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__0900__A _1278_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0604_ _1201_/Q vssd1 vssd1 vccd1 vccd1 _1200_/D sky130_fd_sc_hd__inv_2
XFILLER_8_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0535_ _1164_/Q vssd1 vssd1 vccd1 vccd1 _1135_/B sky130_fd_sc_hd__buf_4
XFILLER_23_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1018_ _1336_/Q _1335_/Q vssd1 vssd1 vccd1 vccd1 _1018_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1088__A _1097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0864__A1 _0546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0524__B _1035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0518_ _1042_/B vssd1 vssd1 vccd1 vccd1 _0518_/Y sky130_fd_sc_hd__inv_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1371__A _1371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1113__51 _1120__55/A vssd1 vssd1 vccd1 vccd1 _1113__51/Y sky130_fd_sc_hd__inv_2
Xfanout45 fanout51/X vssd1 vssd1 vccd1 vccd1 fanout45/X sky130_fd_sc_hd__buf_2
XFILLER_10_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout34 _0861_/Y vssd1 vssd1 vccd1 vccd1 fanout34/X sky130_fd_sc_hd__buf_2
XANTENNA__0715__A _0755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout56 fanout57/X vssd1 vssd1 vccd1 vccd1 fanout56/X sky130_fd_sc_hd__buf_2
XFILLER_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1195__CLK fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input10_A ud_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1352_ input5/X _1352_/D fanout54/X vssd1 vssd1 vccd1 vccd1 _1353_/D sky130_fd_sc_hd__dfrtp_1
X_1283_ _1326_/CLK _1283_/D fanout48/X vssd1 vssd1 vccd1 vccd1 _1283_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1169__RESET_B fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0998_ _0998_/A _0998_/B vssd1 vssd1 vccd1 vccd1 _0999_/B sky130_fd_sc_hd__nand2_1
XANTENNA_input2_A comp_high_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__0301_ clkbuf_0__0301_/X vssd1 vssd1 vccd1 vccd1 _1058__40/A sky130_fd_sc_hd__clkbuf_16
XFILLER_11_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0764__B1 _0716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1210__CLK _0874_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0921_ _0920_/Y _0913_/B _0831_/X vssd1 vssd1 vccd1 vccd1 _0922_/B sky130_fd_sc_hd__a21o_1
XANTENNA__1262__RESET_B fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0783_ _1223_/Q _1222_/Q _1221_/Q _0799_/B vssd1 vssd1 vccd1 vccd1 _0793_/B sky130_fd_sc_hd__or4_1
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout38/X fanout56/X vssd1 vssd1 vccd1 vccd1 _1367_/A sky130_fd_sc_hd__dlrtn_1
X_0852_ _0852_/A vssd1 vssd1 vccd1 vccd1 _0854_/A sky130_fd_sc_hd__clkbuf_1
X_1335_ _1135_/X _1335_/D _0452__10/Y vssd1 vssd1 vccd1 vccd1 _1335_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput2 comp_high_I[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1266_ _1266_/CLK _1266_/D fanout53/X vssd1 vssd1 vccd1 vccd1 _1266_/Q sky130_fd_sc_hd__dfrtp_2
X_1197_ _1359_/A _1197_/D fanout52/X vssd1 vssd1 vccd1 vccd1 _1197_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_91 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1096__A _1142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0994__B1 _0755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0746__B1 _0716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0712__B _1187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1233__CLK fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0903__A _1280_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0985__B1 _0755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0904_ _1279_/Q _0904_/B vssd1 vssd1 vccd1 vccd1 _0904_/X sky130_fd_sc_hd__and2b_1
X_0697_ _1343_/Q vssd1 vssd1 vccd1 vccd1 _1344_/D sky130_fd_sc_hd__inv_2
X_0766_ _1255_/D _1182_/Q vssd1 vssd1 vccd1 vccd1 _0766_/X sky130_fd_sc_hd__xor2_1
X_0835_ _0834_/Y _0830_/B _0831_/X vssd1 vssd1 vccd1 vccd1 _0836_/B sky130_fd_sc_hd__a21o_1
X_1318_ _1356_/A _1318_/D fanout46/X vssd1 vssd1 vccd1 vccd1 _1318_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__1256__CLK input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1249_ _0862_/A _1249_/D _1094_/Y vssd1 vssd1 vccd1 vccd1 _1249_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0723__A _1183_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf _1289_/Q _0953_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0551_ _1142_/B _0551_/B vssd1 vssd1 vccd1 vccd1 _1159_/D sky130_fd_sc_hd__xnor2_1
X_0620_ _1217_/Q vssd1 vssd1 vccd1 vccd1 _1216_/D sky130_fd_sc_hd__inv_2
XFILLER_8_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0482_ _0593_/A vssd1 vssd1 vccd1 vccd1 _0482_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1034_ _1034_/A _1034_/B vssd1 vssd1 vccd1 vccd1 _1034_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__0527__B _1139_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1103_ _1105_/A _1105_/B vssd1 vssd1 vccd1 vccd1 _1103_/Y sky130_fd_sc_hd__xnor2_1
X_1065__45 _1065__45/A vssd1 vssd1 vccd1 vccd1 _1065__45/Y sky130_fd_sc_hd__inv_2
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0543__A _1144_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1093__B _1139_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0749_ _0745_/B _0748_/Y _0998_/A vssd1 vssd1 vccd1 vccd1 _0750_/B sky130_fd_sc_hd__o21ai_1
X_0818_ _1226_/Q _0818_/B vssd1 vssd1 vccd1 vccd1 _1226_/D sky130_fd_sc_hd__xnor2_1
XFILLER_26_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0534_ _1165_/Q vssd1 vssd1 vccd1 vccd1 _1135_/A sky130_fd_sc_hd__buf_4
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0603_ _1198_/Q vssd1 vssd1 vccd1 vccd1 _1199_/D sky130_fd_sc_hd__inv_2
XFILLER_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0867__C1 _0874_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1017_ _1334_/Q _1333_/Q vssd1 vssd1 vccd1 vccd1 _1017_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_23_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1108__49 _1117__53/A vssd1 vssd1 vccd1 vccd1 _1108__49/Y sky130_fd_sc_hd__inv_2
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1254__D input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0561__A1 _1035_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1164__D _1164_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0864__A2 _1035_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0524__C _1042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0517_ _1142_/A _1142_/B vssd1 vssd1 vccd1 vccd1 _1042_/B sky130_fd_sc_hd__xnor2_4
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1099__A _1099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout35 _0532_/Y vssd1 vssd1 vccd1 vccd1 _1035_/B sky130_fd_sc_hd__buf_2
Xfanout46 fanout47/X vssd1 vssd1 vccd1 vccd1 fanout46/X sky130_fd_sc_hd__clkbuf_4
XFILLER_13_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout57 fanout58/X vssd1 vssd1 vccd1 vccd1 fanout57/X sky130_fd_sc_hd__buf_2
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0731__A _0755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0906__A _1278_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1351_ input5/X input1/X fanout49/X vssd1 vssd1 vccd1 vccd1 _1352_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_6_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2__f_w0.cclk_I clkbuf_0_w0.cclk_I/X vssd1 vssd1 vccd1 vccd1 _1326_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_23_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1282_ _1325_/CLK _1282_/D fanout46/X vssd1 vssd1 vccd1 vccd1 _1282_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0551__A _1142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0997_ _0996_/Y _0960_/C _1322_/Q vssd1 vssd1 vccd1 vccd1 _0998_/B sky130_fd_sc_hd__mux2_1
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
+ _1185_/Q _0775_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0455__13 _0448__6/A vssd1 vssd1 vccd1 vccd1 _0455__13/Y sky130_fd_sc_hd__inv_2
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0920_ _1284_/Q _0920_/B vssd1 vssd1 vccd1 vccd1 _0920_/Y sky130_fd_sc_hd__nand2_1
X_0782_ _1226_/Q _1225_/Q _1224_/Q _0809_/B vssd1 vssd1 vccd1 vccd1 _0799_/B sky130_fd_sc_hd__or4_1
X_0851_ _1257_/Q _1256_/D vssd1 vssd1 vccd1 vccd1 _0852_/A sky130_fd_sc_hd__and2b_1
XFILLER_6_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1352__D _1352_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1334_ _1045_/A _1334_/D _1134__61/Y vssd1 vssd1 vccd1 vccd1 _1334_/Q sky130_fd_sc_hd__dfrtp_2
X_1265_ _1360_/A _1265_/D fanout45/X vssd1 vssd1 vccd1 vccd1 _1265_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0546__A _0546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1196_ _1359_/A _1196_/D fanout55/X vssd1 vssd1 vccd1 vccd1 _1196_/Q sky130_fd_sc_hd__dfstp_1
XTAP_81 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 comp_high_Q[0] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XTAP_70 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_92 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1096__B _1142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout53_A fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0903_ _1280_/Q _0903_/B vssd1 vssd1 vccd1 vccd1 _0904_/B sky130_fd_sc_hd__nor2_1
X_0834_ _1259_/D _1233_/Q vssd1 vssd1 vccd1 vccd1 _0834_/Y sky130_fd_sc_hd__nand2_1
X_0696_ _1344_/Q vssd1 vssd1 vccd1 vccd1 _1343_/D sky130_fd_sc_hd__inv_2
X_0765_ _1195_/Q _0765_/B vssd1 vssd1 vccd1 vccd1 _1195_/D sky130_fd_sc_hd__xnor2_1
X_1317_ _1356_/A _1317_/D fanout46/X vssd1 vssd1 vccd1 vccd1 _1317_/Q sky130_fd_sc_hd__dfrtp_2
X_1248_ _1093_/X _1248_/D _0471_/Y vssd1 vssd1 vccd1 vccd1 _1248_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1179_ _1064_/Y _1179_/D _0492__26/Y vssd1 vssd1 vccd1 vccd1 _1179_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__0707__C _1185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1200__CLK _0644_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0550_ _1142_/A _0551_/B vssd1 vssd1 vccd1 vccd1 _1158_/D sky130_fd_sc_hd__xnor2_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0481_ _0593_/A vssd1 vssd1 vccd1 vccd1 _0481_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0894__B1 _0831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1033_ _1033_/A vssd1 vssd1 vccd1 vccd1 _1033_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0824__A _1013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0817_ _0816_/Y _0809_/B _0716_/X vssd1 vssd1 vccd1 vccd1 _0818_/B sky130_fd_sc_hd__a21o_1
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0679_ _1309_/Q vssd1 vssd1 vccd1 vccd1 _1310_/D sky130_fd_sc_hd__inv_2
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1362_/A fanout41/X vssd1 vssd1 vccd1 vccd1 _1368_/A sky130_fd_sc_hd__dlrtn_1
X_0748_ _1193_/Q _1192_/Q _0751_/A vssd1 vssd1 vccd1 vccd1 _0748_/Y sky130_fd_sc_hd__nor3_1
XFILLER_25_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0448__6 _0448__6/A vssd1 vssd1 vccd1 vccd1 _0448__6/Y sky130_fd_sc_hd__inv_2
XANTENNA__0909__A _1279_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1134__61 _1141__65/A vssd1 vssd1 vccd1 vccd1 _1134__61/Y sky130_fd_sc_hd__inv_2
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0533_ _0862_/A _1035_/B vssd1 vssd1 vccd1 vccd1 _0568_/B sky130_fd_sc_hd__nand2_1
X_0602_ _1199_/Q vssd1 vssd1 vccd1 vccd1 _1198_/D sky130_fd_sc_hd__clkinv_2
XFILLER_26_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0554__A _1035_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1016_ _1332_/Q _1331_/Q vssd1 vssd1 vccd1 vccd1 _1016_/Y sky130_fd_sc_hd__xnor2_2
X_1140__64 _1140__64/A vssd1 vssd1 vccd1 vccd1 _1140__64/Y sky130_fd_sc_hd__inv_2
XFILLER_27_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1180__D _1180_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1256__RESET_B fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f__0308_ clkbuf_0__0308_/X vssd1 vssd1 vccd1 vccd1 _0490__25/A sky130_fd_sc_hd__clkbuf_16
XFILLER_8_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0447_ _1053_/A vssd1 vssd1 vccd1 vccd1 _0447_/X sky130_fd_sc_hd__buf_1
X_0516_ _1158_/Q vssd1 vssd1 vccd1 vccd1 _1142_/B sky130_fd_sc_hd__buf_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout36 _0518_/Y vssd1 vssd1 vccd1 vccd1 _0560_/A sky130_fd_sc_hd__clkbuf_4
Xfanout47 fanout49/X vssd1 vssd1 vccd1 vccd1 fanout47/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout58 fanout59/X vssd1 vssd1 vccd1 vccd1 fanout58/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1265__D _1265_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1008__B1 _0831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0767__C1 _0831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1175__D _1175_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf _1282_/Q _0945_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
X_1281_ _1326_/CLK _1281_/D fanout48/X vssd1 vssd1 vccd1 vccd1 _1281_/Q sky130_fd_sc_hd__dfrtp_2
X_1350_ input7/X _1350_/D fanout50/X vssd1 vssd1 vccd1 vccd1 _1350_/Q sky130_fd_sc_hd__dfrtp_1
X_0996_ _0996_/A vssd1 vssd1 vccd1 vccd1 _0996_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1307__CLK _0514_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0850_ _1253_/Q _1252_/Q vssd1 vssd1 vccd1 vccd1 _0850_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_14_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0781_ _1229_/Q _1228_/Q _1227_/Q _0822_/A vssd1 vssd1 vccd1 vccd1 _0809_/B sky130_fd_sc_hd__or4_1
X_1333_ _1133_/X _1333_/D _0453__11/Y vssd1 vssd1 vccd1 vccd1 _1333_/Q sky130_fd_sc_hd__dfrtp_2
X_1264_ _1264_/CLK _1264_/D fanout59/X vssd1 vssd1 vccd1 vccd1 _1264_/Q sky130_fd_sc_hd__dfrtp_4
Xinput4 comp_high_Q[1] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0546__B _1042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_82 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_93 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_60 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1195_ fanout31/X _1195_/D fanout52/X vssd1 vssd1 vccd1 vccd1 _1195_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0979_ _1315_/Q _0979_/B vssd1 vssd1 vccd1 vccd1 _1315_/D sky130_fd_sc_hd__xnor2_1
XFILLER_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0737__A _1187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_w0.ro_block_I.ro_pol_eve.tribuf.t_buf_TE_B _0883_/Y vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0472__A _0479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0902_ _1277_/Q _0902_/B vssd1 vssd1 vccd1 vccd1 _1277_/D sky130_fd_sc_hd__xnor2_1
X_0833_ _1230_/Q _0833_/B vssd1 vssd1 vccd1 vccd1 _1230_/D sky130_fd_sc_hd__xnor2_1
Xclkbuf_0__0301_ _1053_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0301_/X sky130_fd_sc_hd__clkbuf_16
X_0695_ _1341_/Q vssd1 vssd1 vccd1 vccd1 _1342_/D sky130_fd_sc_hd__inv_2
XFILLER_6_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0764_ _0763_/Y _0760_/B _0716_/X vssd1 vssd1 vccd1 vccd1 _0765_/B sky130_fd_sc_hd__a21o_1
X_1178_ _1035_/A _1178_/D _1063__44/Y vssd1 vssd1 vccd1 vccd1 _1178_/Q sky130_fd_sc_hd__dfrtp_4
X_1316_ _1356_/A _1316_/D fanout49/X vssd1 vssd1 vccd1 vccd1 _1316_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__0557__A _1139_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1247_ _1035_/B _1247_/D _1092_/Y vssd1 vssd1 vccd1 vccd1 _1247_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout38/X fanout56/X vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1193__RESET_B fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0480_ _1099_/A vssd1 vssd1 vccd1 vccd1 _0593_/A sky130_fd_sc_hd__buf_6
XFILLER_7_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1032_ _1032_/A _1032_/B vssd1 vssd1 vccd1 vccd1 _1033_/A sky130_fd_sc_hd__or2_1
X_1129__59 _1140__64/A vssd1 vssd1 vccd1 vccd1 _1129__59/Y sky130_fd_sc_hd__inv_2
XANTENNA__1175__CLK _0548_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0840__A _1013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0816_ _1227_/Q _0816_/B vssd1 vssd1 vccd1 vccd1 _0816_/Y sky130_fd_sc_hd__nand2_1
X_0747_ _1190_/Q _0747_/B vssd1 vssd1 vccd1 vccd1 _1190_/D sky130_fd_sc_hd__xnor2_1
X_0678_ _1310_/Q vssd1 vssd1 vccd1 vccd1 _1309_/D sky130_fd_sc_hd__inv_2
XFILLER_26_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.ro_block_I.ro_pol.tribuf.t_buf _1033_/X _0882_/Y vssd1 vssd1 vccd1 vccd1 _1370_/A
+ sky130_fd_sc_hd__ebufn_2
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1168_/CLK fanout43/X vssd1 vssd1 vccd1 vccd1 _1366_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1198__CLK _0643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0876__A1 _1042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0925__A _1284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0601_ _1180_/Q vssd1 vssd1 vccd1 vccd1 _1181_/D sky130_fd_sc_hd__inv_2
XANTENNA__0660__A _1292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0532_ _0874_/D vssd1 vssd1 vccd1 vccd1 _0532_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0867__A1 _0546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1015_ _1330_/Q _1329_/Q vssd1 vssd1 vccd1 vccd1 _1015_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_22_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1044__A1 _0873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1340__CLK _0862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0570__A _1133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0480__A _1099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0794__B1 _0755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0450__8 _0451__9/A vssd1 vssd1 vccd1 vccd1 _0450__8/Y sky130_fd_sc_hd__inv_2
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1213__CLK _0862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__0307_ clkbuf_0__0307_/X vssd1 vssd1 vccd1 vccd1 _0448__6/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__1225__RESET_B fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0515_ _1159_/Q vssd1 vssd1 vccd1 vccd1 _1142_/A sky130_fd_sc_hd__buf_4
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout37 _0514_/Y vssd1 vssd1 vccd1 vccd1 _1042_/A sky130_fd_sc_hd__buf_4
XANTENNA_w0.ro_block_I.ro_pol.tribuf.t_buf_TE_B _0882_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout59 input9/X vssd1 vssd1 vccd1 vccd1 fanout59/X sky130_fd_sc_hd__buf_2
Xfanout48 fanout49/X vssd1 vssd1 vccd1 vccd1 fanout48/X sky130_fd_sc_hd__clkbuf_4
XFILLER_13_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0475__A _0479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1236__CLK _0644_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1280_ _1358_/A _1280_/D fanout46/X vssd1 vssd1 vccd1 vccd1 _1280_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0995_ _1320_/Q _0995_/B vssd1 vssd1 vccd1 vccd1 _1320_/D sky130_fd_sc_hd__xnor2_1
XFILLER_9_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1259__CLK input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0930__B1 _0755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1101__46 _1120__55/A vssd1 vssd1 vccd1 vccd1 _1264_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0749__B1 _0998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1276__D _1276_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0921__B1 _0831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0461__18 _0467__24/A vssd1 vssd1 vccd1 vccd1 _0461__18/Y sky130_fd_sc_hd__inv_2
XANTENNA__0933__A _1290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0780_ _1259_/D _1233_/Q _1231_/Q _1230_/Q vssd1 vssd1 vccd1 vccd1 _0822_/A sky130_fd_sc_hd__or4_2
XFILLER_6_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 phi1b_dig_I[0] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
X_1332_ _1132_/Y _1332_/D _0454__12/Y vssd1 vssd1 vccd1 vccd1 _1332_/Q sky130_fd_sc_hd__dfrtp_4
X_1263_ _1362_/A _1263_/D fanout45/X vssd1 vssd1 vccd1 vccd1 _1263_/Q sky130_fd_sc_hd__dfrtp_4
X_1194_ fanout34/X _1194_/D fanout52/X vssd1 vssd1 vccd1 vccd1 _1194_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_83 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0978_ _0998_/A _0978_/B vssd1 vssd1 vccd1 vccd1 _0979_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout39_A _1099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0753__A _1013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0647__B _1265_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0928__A _0998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0663__A _1293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0901_ _0900_/Y _0897_/B _0831_/X vssd1 vssd1 vccd1 vccd1 _0902_/B sky130_fd_sc_hd__a21o_1
X_0832_ _0828_/Y _0830_/X _0831_/X vssd1 vssd1 vccd1 vccd1 _0833_/B sky130_fd_sc_hd__a21o_1
X_0763_ _1255_/D _1197_/Q vssd1 vssd1 vccd1 vccd1 _0763_/Y sky130_fd_sc_hd__nand2_1
X_0694_ _1342_/Q vssd1 vssd1 vccd1 vccd1 _1341_/D sky130_fd_sc_hd__inv_2
X_1315_ _1356_/A _1315_/D fanout49/X vssd1 vssd1 vccd1 vccd1 _1315_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1177_ _1062_/Y _1177_/D _0493__27/Y vssd1 vssd1 vccd1 vccd1 _1177_/Q sky130_fd_sc_hd__dfrtp_2
X_1246_ _1091_/X _1246_/D _0472_/Y vssd1 vssd1 vccd1 vccd1 _1246_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__0557__B _0557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0573__A _1132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0483__A _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1079_/A fanout56/X vssd1 vssd1 vccd1 vccd1 _1367_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_11_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1031_ _1353_/D _1354_/Q vssd1 vssd1 vccd1 vccd1 _1032_/B sky130_fd_sc_hd__and2b_1
X_1100_ _1122_/A vssd1 vssd1 vccd1 vccd1 _1100_/X sky130_fd_sc_hd__buf_1
XFILLER_19_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
+ _1220_/Q _0847_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_7_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0815_ _1225_/Q _0815_/B vssd1 vssd1 vccd1 vccd1 _1225_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0746_ _0745_/Y _0738_/B _0716_/X vssd1 vssd1 vccd1 vccd1 _0747_/B sky130_fd_sc_hd__a21o_1
X_0677_ _1307_/Q vssd1 vssd1 vccd1 vccd1 _1308_/D sky130_fd_sc_hd__clkinv_2
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_A _1313_/Q vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1229_ fanout34/X _1229_/D fanout55/X vssd1 vssd1 vccd1 vccd1 _1229_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_3__f_clk_master clkbuf_0_clk_master/X vssd1 vssd1 vccd1 vccd1 _1360_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0876__A2 _0873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0478__A _0479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0644__C _0644_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1038__C1 _0873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0600_ _1181_/Q vssd1 vssd1 vccd1 vccd1 _1180_/D sky130_fd_sc_hd__inv_2
X_0531_ _1137_/A _1137_/B vssd1 vssd1 vccd1 vccd1 _0874_/D sky130_fd_sc_hd__xor2_4
XFILLER_8_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1014_ _1328_/Q _1327_/Q vssd1 vssd1 vccd1 vccd1 _1014_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__0570__B _0570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0555__A1 _0862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0729_ _0724_/B _0728_/X _0998_/A vssd1 vssd1 vccd1 vccd1 _0730_/B sky130_fd_sc_hd__o21ai_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0446__2_A _1053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0671__A _1301_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__0306_ clkbuf_0__0306_/X vssd1 vssd1 vccd1 vccd1 _1053_/A sky130_fd_sc_hd__clkbuf_16
X_0514_ _0546_/A vssd1 vssd1 vccd1 vccd1 _0514_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0445_ _1360_/A vssd1 vssd1 vccd1 vccd1 _0445_/X sky130_fd_sc_hd__buf_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0467__24 _0467__24/A vssd1 vssd1 vccd1 vccd1 _0467__24/Y sky130_fd_sc_hd__inv_2
XANTENNA__0565__B _0873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout49 fanout51/X vssd1 vssd1 vccd1 vccd1 fanout49/X sky130_fd_sc_hd__clkbuf_4
Xfanout38 _1079_/A vssd1 vssd1 vccd1 vccd1 fanout38/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1188__CLK fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0491__A _1053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0994_ _0990_/B _0993_/Y _0755_/A vssd1 vssd1 vccd1 vccd1 _0995_/B sky130_fd_sc_hd__o21ai_1
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0576__A _1132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1353__CLK input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0486__A _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0933__B _1348_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1331_ _0590_/C _1331_/D _1131__60/Y vssd1 vssd1 vccd1 vccd1 _1331_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 phi1b_dig_I[1] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
X_1262_ _1099_/Y _1262_/D fanout59/X vssd1 vssd1 vccd1 vccd1 _1262_/Q sky130_fd_sc_hd__dfrtp_1
X_1193_ fanout31/X _1193_/D fanout54/X vssd1 vssd1 vccd1 vccd1 _1193_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1020__A _1340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_84 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0977_ _1317_/Q _1316_/Q _0980_/B _0974_/B vssd1 vssd1 vccd1 vccd1 _0978_/B sky130_fd_sc_hd__a31o_1
XFILLER_9_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1105__A _1105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0944__A _1292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0900_ _1278_/Q _0900_/B vssd1 vssd1 vccd1 vccd1 _0900_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__1249__CLK _0862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0693_ _1339_/Q vssd1 vssd1 vccd1 vccd1 _1340_/D sky130_fd_sc_hd__inv_2
X_0831_ _0831_/A vssd1 vssd1 vccd1 vccd1 _0831_/X sky130_fd_sc_hd__buf_4
X_0762_ _1194_/Q _0762_/B vssd1 vssd1 vccd1 vccd1 _1194_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1314_ _1325_/CLK _1314_/D fanout49/X vssd1 vssd1 vccd1 vccd1 _1314_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1015__A _1330_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1176_ _1035_/A _1176_/D _1061__43/Y vssd1 vssd1 vccd1 vccd1 _1176_/Q sky130_fd_sc_hd__dfrtp_2
X_1245_ _0868_/B _1245_/D _1090_/Y vssd1 vssd1 vccd1 vccd1 _1245_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0573__B _1132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout51_A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf _1317_/Q _1016_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_12_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1030_ _1030_/A vssd1 vssd1 vccd1 vccd1 _1032_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_19_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0814_ _1013_/A _0814_/B vssd1 vssd1 vccd1 vccd1 _0815_/B sky130_fd_sc_hd__nand2_1
X_0676_ _1308_/Q vssd1 vssd1 vccd1 vccd1 _1307_/D sky130_fd_sc_hd__inv_2
XFILLER_6_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0745_ _1191_/Q _0745_/B vssd1 vssd1 vccd1 vccd1 _0745_/Y sky130_fd_sc_hd__nand2_1
X_1228_ _1357_/A _1228_/D fanout55/X vssd1 vssd1 vccd1 vccd1 _1228_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_GATE_N
+ _1099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1056__38 _1058__40/A vssd1 vssd1 vccd1 vccd1 _1167_/CLK sky130_fd_sc_hd__inv_2
X_1159_ _1159_/CLK _1159_/D fanout44/X vssd1 vssd1 vccd1 vccd1 _1159_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__0584__A _1130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1312__RESET_B fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0644__D _0644_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0530_ _1162_/Q vssd1 vssd1 vccd1 vccd1 _1137_/B sky130_fd_sc_hd__clkbuf_4
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1013_ _1013_/A _1326_/Q vssd1 vssd1 vccd1 vccd1 _1326_/D sky130_fd_sc_hd__xor2_1
XFILLER_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0659_ _1273_/Q vssd1 vssd1 vccd1 vccd1 _1274_/D sky130_fd_sc_hd__inv_2
X_0728_ _1186_/Q _0728_/B vssd1 vssd1 vccd1 vccd1 _0728_/X sky130_fd_sc_hd__and2b_1
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0489__A _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1148_/CLK fanout41/X vssd1 vssd1 vccd1 vccd1 _1368_/A sky130_fd_sc_hd__dlrtn_1
Xclkbuf_1_0__f__0305_ clkbuf_0__0305_/X vssd1 vssd1 vccd1 vccd1 _1141__65/A sky130_fd_sc_hd__clkbuf_16
X_0513_ _1144_/A _1144_/B vssd1 vssd1 vccd1 vccd1 _0546_/A sky130_fd_sc_hd__xnor2_4
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0565__C _1035_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1007__B _1352_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0862__A _0862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout39 _1099_/A vssd1 vssd1 vccd1 vccd1 _1079_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
+ _1182_/Q _0778_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_10_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0682__A _1330_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0993_ _1322_/Q _1321_/Q _0996_/A vssd1 vssd1 vccd1 vccd1 _0993_/Y sky130_fd_sc_hd__nor3_1
XFILLER_8_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0592__A _1128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0921__A2 _0913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1261_ input6/X _1261_/D fanout53/X vssd1 vssd1 vccd1 vccd1 _1261_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1178__CLK _1035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1330_ _1130_/Y _1330_/D _0455__13/Y vssd1 vssd1 vccd1 vccd1 _1330_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_85 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 phi1b_dig_Q[0] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
XTAP_63 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1192_ fanout31/X _1192_/D fanout50/X vssd1 vssd1 vccd1 vccd1 _1192_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1020__B _1339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0976_ _1314_/Q _0976_/B vssd1 vssd1 vccd1 vccd1 _1314_/D sky130_fd_sc_hd__xnor2_1
XTAP_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_A _1276_/Q vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0497__A _1105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1121__A _1142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0830_ _1231_/Q _0830_/B vssd1 vssd1 vccd1 vccd1 _0830_/X sky130_fd_sc_hd__or2_1
X_0692_ _1340_/Q vssd1 vssd1 vccd1 vccd1 _1339_/D sky130_fd_sc_hd__inv_2
X_0761_ _0758_/Y _0760_/X _0716_/X vssd1 vssd1 vccd1 vccd1 _0762_/B sky130_fd_sc_hd__a21o_1
XANTENNA__1015__B _1329_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1313_ _1356_/A _1313_/D fanout45/X vssd1 vssd1 vccd1 vccd1 _1313_/Q sky130_fd_sc_hd__dfrtp_4
X_1244_ _1089_/X _1244_/D _0473_/Y vssd1 vssd1 vccd1 vccd1 _1244_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1175_ _0548_/C _1175_/D _0494__28/Y vssd1 vssd1 vccd1 vccd1 _1175_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__1343__CLK _1042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0959_ _1326_/Q _1352_/D _1324_/Q _1323_/Q vssd1 vssd1 vccd1 vccd1 _0960_/C sky130_fd_sc_hd__and4_1
XFILLER_24_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0780__A _1259_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1171__RESET_B fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1216__CLK _1042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1259__RESET_B fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0690__A _1338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput10 ud_en vssd1 vssd1 vccd1 vccd1 _0714_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__0803__A1 _1224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0813_ _1227_/Q _1226_/Q _0816_/B _0810_/B vssd1 vssd1 vccd1 vccd1 _0814_/B sky130_fd_sc_hd__a31o_1
X_0675_ _1305_/Q vssd1 vssd1 vccd1 vccd1 _1306_/D sky130_fd_sc_hd__inv_2
X_0744_ _1189_/Q _0744_/B vssd1 vssd1 vccd1 vccd1 _1189_/D sky130_fd_sc_hd__xnor2_1
XFILLER_26_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1143__3 _1053_/A vssd1 vssd1 vccd1 vccd1 _1143__3/Y sky130_fd_sc_hd__inv_2
XANTENNA__0584__B _0585_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1158_ _1360_/A _1158_/D fanout44/X vssd1 vssd1 vccd1 vccd1 _1158_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__0568__C _0868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1227_ _1357_/A _1227_/D fanout55/X vssd1 vssd1 vccd1 vccd1 _1227_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1089_ _1135_/A _1135_/B vssd1 vssd1 vccd1 vccd1 _1089_/X sky130_fd_sc_hd__xor2_2
XFILLER_16_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1352__RESET_B fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0797__B1 _0716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1038__A1 _1042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0549__A0 _1042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0685__A _1331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1012_ _1325_/Q _1012_/B vssd1 vssd1 vccd1 vccd1 _1325_/D sky130_fd_sc_hd__xnor2_1
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout38/X fanout56/X vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0727_ _1187_/Q _0727_/B vssd1 vssd1 vccd1 vccd1 _0728_/B sky130_fd_sc_hd__nor2_1
X_0658_ _1274_/Q vssd1 vssd1 vccd1 vccd1 _1273_/D sky130_fd_sc_hd__clkinv_2
X_0589_ _0589_/A vssd1 vssd1 vccd1 vccd1 _0644_/D sky130_fd_sc_hd__clkinv_2
XFILLER_26_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__0304_ clkbuf_0__0304_/X vssd1 vssd1 vccd1 vccd1 _1117__53/A sky130_fd_sc_hd__clkbuf_16
XFILLER_8_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0512_ _1156_/Q vssd1 vssd1 vccd1 vccd1 _1144_/B sky130_fd_sc_hd__buf_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1168_/CLK fanout42/X vssd1 vssd1 vccd1 vccd1 _1366_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_22_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0862__B _1035_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf _1279_/Q _0948_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_2_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0924__B1 _0755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1124__A _1144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0992_ _1319_/Q _0992_/B vssd1 vssd1 vccd1 vccd1 _1319_/D sky130_fd_sc_hd__xnor2_1
XFILLER_12_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0915__B1 _0755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0592__B _0592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0873__A _0873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1260_ input6/X _1260_/D fanout53/X vssd1 vssd1 vccd1 vccd1 _1261_/D sky130_fd_sc_hd__dfrtp_1
XANTENNA__0958__A _1313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 phi1b_dig_Q[1] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_2
X_1191_ fanout31/X _1191_/D fanout54/X vssd1 vssd1 vccd1 vccd1 _1191_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__0693__A _1339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_86 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0975_ _0970_/B _0974_/X _0755_/A vssd1 vssd1 vccd1 vccd1 _0976_/B sky130_fd_sc_hd__o21ai_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1272__CLK _0542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1121__B _1142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0760_ _1195_/Q _0760_/B vssd1 vssd1 vccd1 vccd1 _0760_/X sky130_fd_sc_hd__or2_1
X_0691_ _1337_/Q vssd1 vssd1 vccd1 vccd1 _1338_/D sky130_fd_sc_hd__inv_2
XANTENNA__1295__CLK _0590_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1174_ _1035_/A _1174_/D _1060__42/Y vssd1 vssd1 vccd1 vccd1 _1174_/Q sky130_fd_sc_hd__dfrtp_1
X_1312_ _1325_/CLK _1312_/D fanout49/X vssd1 vssd1 vccd1 vccd1 _1312_/Q sky130_fd_sc_hd__dfrtp_2
X_1243_ _1045_/A _1243_/D _1088_/Y vssd1 vssd1 vccd1 vccd1 _1243_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0958_ _1313_/Q _1312_/Q _0967_/B vssd1 vssd1 vccd1 vccd1 _0958_/X sky130_fd_sc_hd__or3_1
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0889_ _1290_/Q _1348_/D _1288_/Q _1287_/Q vssd1 vssd1 vccd1 vccd1 _0890_/C sky130_fd_sc_hd__and4_1
XANTENNA__0598__A _1179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout37_A _0514_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1116__B _1137_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1132__A _1132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0812_ _1224_/Q _0812_/B vssd1 vssd1 vccd1 vccd1 _1224_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0743_ _1013_/A _0743_/B vssd1 vssd1 vccd1 vccd1 _0744_/B sky130_fd_sc_hd__nand2_1
X_0674_ _1306_/Q vssd1 vssd1 vccd1 vccd1 _1305_/D sky130_fd_sc_hd__inv_2
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
+ _1190_/Q _0770_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_26_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1042__A _1042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1157_ _1157_/CLK _1157_/D fanout44/X vssd1 vssd1 vccd1 vccd1 _1157_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__0865__B _0873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1226_ _1359_/A _1226_/D fanout55/X vssd1 vssd1 vccd1 vccd1 _1226_/Q sky130_fd_sc_hd__dfrtp_2
X_1088_ _1097_/A vssd1 vssd1 vccd1 vccd1 _1088_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1038__A2 _0874_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_GATE_N
+ _1099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1011_ _0958_/X _0963_/Y _1010_/X _0831_/A vssd1 vssd1 vccd1 vccd1 _1012_/B sky130_fd_sc_hd__a211o_1
XFILLER_23_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1061__43 _1065__45/A vssd1 vssd1 vccd1 vccd1 _1061__43/Y sky130_fd_sc_hd__inv_2
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout38/X fanout57/X vssd1 vssd1 vccd1 vccd1 _1367_/A sky130_fd_sc_hd__dlrtn_1
X_0726_ _1184_/Q _0726_/B vssd1 vssd1 vccd1 vccd1 _1184_/D sky130_fd_sc_hd__xnor2_1
XFILLER_8_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0588_ _1128_/A _1128_/B vssd1 vssd1 vccd1 vccd1 _0589_/A sky130_fd_sc_hd__xnor2_1
X_0657_ _1271_/Q vssd1 vssd1 vccd1 vccd1 _1272_/D sky130_fd_sc_hd__inv_2
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1209_ _0868_/B _1209_/D _1073_/Y vssd1 vssd1 vccd1 vccd1 _1209_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0511_ _1157_/Q vssd1 vssd1 vccd1 vccd1 _1144_/A sky130_fd_sc_hd__buf_4
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1229__CLK fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0709_ _1255_/D _1197_/Q _1195_/Q _1194_/Q vssd1 vssd1 vccd1 vccd1 _0710_/C sky130_fd_sc_hd__and4_1
XANTENNA_input9_A rstb vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1124__B _1144_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0963__B _1313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0991_ _0990_/Y _0983_/B _0831_/A vssd1 vssd1 vccd1 vccd1 _0992_/B sky130_fd_sc_hd__a21o_1
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1034__B _1034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0873__B _0873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1165__RESET_B fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_TE_B _0950_/Y vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 rstb vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1135__A _1135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1190_ fanout31/X _1190_/D fanout50/X vssd1 vssd1 vccd1 vccd1 _1190_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_18_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_87 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0974_ _1315_/Q _0974_/B vssd1 vssd1 vccd1 vccd1 _0974_/X sky130_fd_sc_hd__and2b_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1029__B _1353_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1045__A _1045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0868__B _0868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0884__A _1290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0690_ _1338_/Q vssd1 vssd1 vccd1 vccd1 _1337_/D sky130_fd_sc_hd__inv_2
XFILLER_10_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1311_ _1325_/CLK _1311_/D fanout48/X vssd1 vssd1 vccd1 vccd1 _1311_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_2_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1173_ _1173_/CLK _1173_/D fanout51/X vssd1 vssd1 vccd1 vccd1 _1173_/Q sky130_fd_sc_hd__dfrtp_1
X_1242_ _1087_/X _1242_/D _0474_/Y vssd1 vssd1 vccd1 vccd1 _1242_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0957_ _1316_/Q _1315_/Q _1314_/Q _0973_/B vssd1 vssd1 vccd1 vccd1 _0967_/B sky130_fd_sc_hd__or4_1
X_0888_ _1277_/Q _1276_/Q _0897_/B vssd1 vssd1 vccd1 vccd1 _0888_/X sky130_fd_sc_hd__or3_1
XFILLER_9_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
+ _1232_/Q _0850_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1132__B _1132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0673_ _1303_/Q vssd1 vssd1 vccd1 vccd1 _1304_/D sky130_fd_sc_hd__inv_2
XFILLER_7_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_0__f_clk_master clkbuf_0_clk_master/X vssd1 vssd1 vccd1 vccd1 _1148_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_0811_ _0806_/B _0810_/X _0755_/X vssd1 vssd1 vccd1 vccd1 _0812_/B sky130_fd_sc_hd__o21ai_1
XFILLER_6_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0742_ _1191_/Q _1190_/Q _0745_/B _0739_/B vssd1 vssd1 vccd1 vccd1 _0743_/B sky130_fd_sc_hd__a31o_1
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1042__B _1042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1087_ _1133_/A _1133_/B vssd1 vssd1 vccd1 vccd1 _1087_/X sky130_fd_sc_hd__xor2_1
X_1156_ _1168_/CLK _1156_/D fanout43/X vssd1 vssd1 vccd1 vccd1 _1156_/Q sky130_fd_sc_hd__dfrtp_1
X_1225_ _1359_/A _1225_/D fanout53/X vssd1 vssd1 vccd1 vccd1 _1225_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0966__B _1313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0494__28 _1049__32/A vssd1 vssd1 vccd1 vccd1 _0494__28/Y sky130_fd_sc_hd__inv_2
XANTENNA__0982__A _1316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1010_ _1326_/Q _1311_/Q vssd1 vssd1 vccd1 vccd1 _1010_/X sky130_fd_sc_hd__xor2_1
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0656_ _1272_/Q vssd1 vssd1 vccd1 vccd1 _1271_/D sky130_fd_sc_hd__inv_2
X_0725_ _0724_/Y _0720_/B _0716_/X vssd1 vssd1 vccd1 vccd1 _0726_/B sky130_fd_sc_hd__a21o_1
XFILLER_7_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1208_ _0873_/B _1208_/D _0484_/Y vssd1 vssd1 vccd1 vccd1 _1208_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1053__A _1053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0587_ _1172_/Q vssd1 vssd1 vccd1 vccd1 _1128_/B sky130_fd_sc_hd__buf_4
XFILLER_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1139_ _1139_/A _1139_/B vssd1 vssd1 vccd1 vccd1 _1139_/X sky130_fd_sc_hd__xor2_1
XFILLER_22_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1300__CLK _0868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0510_ _1146_/A _0510_/B vssd1 vssd1 vccd1 vccd1 _1153_/D sky130_fd_sc_hd__xnor2_1
XFILLER_8_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0639_ _1250_/Q vssd1 vssd1 vccd1 vccd1 _1251_/D sky130_fd_sc_hd__clkinv_2
X_0708_ _1184_/Q _1183_/Q _0720_/B vssd1 vssd1 vccd1 vccd1 _0708_/X sky130_fd_sc_hd__or3_1
XANTENNA__0887__A _1280_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0924__A2 _0923_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0990_ _1320_/Q _0990_/B vssd1 vssd1 vccd1 vccd1 _0990_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0463__20 _0490__25/A vssd1 vssd1 vccd1 vccd1 _0463__20/Y sky130_fd_sc_hd__inv_2
XANTENNA__1346__CLK _1146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1362_/A fanout41/X vssd1 vssd1 vccd1 vccd1 _1368_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1135__B _1135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0974__B _0974_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1219__CLK fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0446__1 _1053_/A vssd1 vssd1 vccd1 vccd1 _0446__1/Y sky130_fd_sc_hd__inv_2
XFILLER_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_88 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0973_ _1316_/Q _0973_/B vssd1 vssd1 vccd1 vccd1 _0974_/B sky130_fd_sc_hd__nor2_1
XANTENNA__1045__B _1045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0884__B _1348_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1315__RESET_B fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_3__f_w0.cclk_I clkbuf_0_w0.cclk_I/X vssd1 vssd1 vccd1 vccd1 _1325_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1310_ _1126_/Y _1310_/D _0457__15/Y vssd1 vssd1 vccd1 vccd1 _1310_/Q sky130_fd_sc_hd__dfrtp_2
X_1241_ _1086_/Y _1241_/D _0475_/Y vssd1 vssd1 vccd1 vccd1 _1241_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf _1314_/Q _1019_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
X_1172_ _1360_/A _1172_/D fanout41/X vssd1 vssd1 vccd1 vccd1 _1172_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1191__CLK fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0956_ _1319_/Q _1318_/Q _1317_/Q _0983_/B vssd1 vssd1 vccd1 vccd1 _0973_/B sky130_fd_sc_hd__or4_2
X_0887_ _1280_/Q _1279_/Q _1278_/Q _0903_/B vssd1 vssd1 vccd1 vccd1 _0897_/B sky130_fd_sc_hd__or4_1
XANTENNA__0895__A _1275_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0981__B1 _0831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0810_ _1225_/Q _0810_/B vssd1 vssd1 vccd1 vccd1 _0810_/X sky130_fd_sc_hd__and2b_1
X_0672_ _1304_/Q vssd1 vssd1 vccd1 vccd1 _1303_/D sky130_fd_sc_hd__inv_2
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0741_ _1188_/Q _0741_/B vssd1 vssd1 vccd1 vccd1 _1188_/D sky130_fd_sc_hd__xnor2_1
X_1224_ _1357_/A _1224_/D fanout55/X vssd1 vssd1 vccd1 vccd1 _1224_/Q sky130_fd_sc_hd__dfrtp_4
X_1086_ _1132_/A _1132_/B vssd1 vssd1 vccd1 vccd1 _1086_/Y sky130_fd_sc_hd__xnor2_1
X_1155_ _1155_/CLK _1155_/D fanout44/X vssd1 vssd1 vccd1 vccd1 _1155_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0939_ _1288_/Q _0939_/B vssd1 vssd1 vccd1 vccd1 _1288_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1119__54 _1120__55/A vssd1 vssd1 vccd1 vccd1 _1119__54/Y sky130_fd_sc_hd__inv_2
XFILLER_24_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout42_A fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_A _1319_/Q vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0966__C _0970_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1125__57 _1141__65/A vssd1 vssd1 vccd1 vccd1 _1125__57/Y sky130_fd_sc_hd__inv_2
XFILLER_22_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0586_ _1173_/Q vssd1 vssd1 vccd1 vccd1 _1128_/A sky130_fd_sc_hd__buf_4
X_0655_ _1269_/Q vssd1 vssd1 vccd1 vccd1 _1270_/D sky130_fd_sc_hd__inv_2
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0724_ _1185_/Q _0724_/B vssd1 vssd1 vccd1 vccd1 _0724_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1207_ _1045_/A _1207_/D _1072_/Y vssd1 vssd1 vccd1 vccd1 _1207_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1069_ _1077_/A vssd1 vssd1 vccd1 vccd1 _1069_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0892__B _1280_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1252__CLK _1042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__0301_ clkbuf_0__0301_/X vssd1 vssd1 vccd1 vccd1 _1065__45/A sky130_fd_sc_hd__clkbuf_16
XFILLER_12_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0707_ _1187_/Q _1186_/Q _1185_/Q _0727_/B vssd1 vssd1 vccd1 vccd1 _0720_/B sky130_fd_sc_hd__or4_1
X_0569_ _1133_/B _0570_/B vssd1 vssd1 vccd1 vccd1 _1166_/D sky130_fd_sc_hd__xnor2_1
X_0638_ _1251_/Q vssd1 vssd1 vccd1 vccd1 _1250_/D sky130_fd_sc_hd__inv_2
XANTENNA__0887__B _1279_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout38/X fanout56/X vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_1_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0963__D _0970_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1298__CLK _1045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
+ _1225_/Q _0842_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_9_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0500__B _0548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0988__A _0998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1168_/CLK fanout43/X vssd1 vssd1 vccd1 vccd1 _1366_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_10_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0601__A _1180_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0446__2 _1053_/A vssd1 vssd1 vccd1 vccd1 _1034_/A sky130_fd_sc_hd__inv_2
XTAP_67 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0972_ _1313_/Q _0972_/B vssd1 vssd1 vccd1 vccd1 _1313_/D sky130_fd_sc_hd__xnor2_1
XTAP_89 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1355__RESET_B fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1336__CLK _0868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1171_ _1171_/CLK _1171_/D fanout54/X vssd1 vssd1 vccd1 vccd1 _1171_/Q sky130_fd_sc_hd__dfrtp_1
X_1240_ _0590_/C _1240_/D _1085_/Y vssd1 vssd1 vccd1 vccd1 _1240_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0955_ _1322_/Q _1321_/Q _1320_/Q _0996_/A vssd1 vssd1 vccd1 vccd1 _0983_/B sky130_fd_sc_hd__or4_1
X_0886_ _1283_/Q _1282_/Q _1281_/Q _0913_/B vssd1 vssd1 vccd1 vccd1 _0903_/B sky130_fd_sc_hd__or4_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1072__A _1077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1369_ _1369_/A vssd1 vssd1 vccd1 vccd1 _1369_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1209__CLK _0868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_0_clk_master_A clk_master vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1058__40 _1058__40/A vssd1 vssd1 vccd1 vccd1 _1171_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0740_ _0735_/B _0739_/X _0998_/A vssd1 vssd1 vccd1 vccd1 _0741_/B sky130_fd_sc_hd__o21ai_1
X_0671_ _1301_/Q vssd1 vssd1 vccd1 vccd1 _1302_/D sky130_fd_sc_hd__inv_2
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1154_ _1360_/A _1154_/D fanout43/X vssd1 vssd1 vccd1 vccd1 _1154_/Q sky130_fd_sc_hd__dfrtp_1
X_1223_ _1359_/A _1223_/D fanout53/X vssd1 vssd1 vccd1 vccd1 _1223_/Q sky130_fd_sc_hd__dfrtp_2
X_1085_ _1097_/A vssd1 vssd1 vccd1 vccd1 _1085_/Y sky130_fd_sc_hd__inv_2
X_0869_ _0873_/B _0864_/X _0865_/X _1045_/A _0868_/X vssd1 vssd1 vccd1 vccd1 _0870_/B
+ sky130_fd_sc_hd__o221a_1
X_0938_ _0937_/Y _0934_/B _0831_/X vssd1 vssd1 vccd1 vccd1 _0939_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1181__CLK _1066_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0723_ _1183_/Q _0723_/B vssd1 vssd1 vccd1 vccd1 _1183_/D sky130_fd_sc_hd__xnor2_1
X_0585_ _1130_/A _0585_/B vssd1 vssd1 vccd1 vccd1 _1171_/D sky130_fd_sc_hd__xnor2_1
X_0654_ _1270_/Q vssd1 vssd1 vccd1 vccd1 _1269_/D sky130_fd_sc_hd__clkinv_2
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1137_ _1137_/A _1137_/B vssd1 vssd1 vccd1 vccd1 _1137_/X sky130_fd_sc_hd__xor2_1
X_1206_ _0868_/A _1206_/D _0485_/Y vssd1 vssd1 vccd1 vccd1 _1206_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__0892__C _1279_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1068_ _1077_/A vssd1 vssd1 vccd1 vccd1 _1068_/Y sky130_fd_sc_hd__inv_2
X_1052__35 _1052__35/A vssd1 vssd1 vccd1 vccd1 _1161_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0872__B1 _0560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf _1276_/Q _0951_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0863__B1 _1042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0514__A _0546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0706_ _1190_/Q _1189_/Q _1188_/Q _0738_/B vssd1 vssd1 vccd1 vccd1 _0727_/B sky130_fd_sc_hd__or4_2
X_0568_ _0568_/A _0568_/B _0868_/B vssd1 vssd1 vccd1 vccd1 _0570_/B sky130_fd_sc_hd__or3_4
X_0499_ _1150_/Q _1151_/Q vssd1 vssd1 vccd1 vccd1 _0548_/B sky130_fd_sc_hd__xor2_4
X_0637_ _1248_/Q vssd1 vssd1 vccd1 vccd1 _1249_/D sky130_fd_sc_hd__inv_2
XANTENNA__0887__C _1278_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_A
+ _1224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1080__A _1097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout38/X fanout57/X vssd1 vssd1 vccd1 vccd1 _1367_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA_wrapper_cell_loop\[0\].w1.ro_block_I.ro_pol.tribuf.t_buf_TE_B _0702_/Y vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1075__A _1077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input7_A phi1b_dig_Q[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_79 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0971_ _0970_/Y _0967_/B _0831_/X vssd1 vssd1 vccd1 vccd1 _0972_/B sky130_fd_sc_hd__a21o_1
XFILLER_4_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[0\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf _0854_/A _0701_/Y vssd1
+ vssd1 vccd1 vccd1 _1373_/A sky130_fd_sc_hd__ebufn_4
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0702__A _1179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1170_ _1360_/A _1170_/D fanout51/X vssd1 vssd1 vccd1 vccd1 _1170_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_A _1282_/Q vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0954_ _1326_/Q _1352_/D _1324_/Q _1323_/Q vssd1 vssd1 vccd1 vccd1 _0996_/A sky130_fd_sc_hd__or4_2
X_0885_ _1286_/Q _1285_/Q _1284_/Q _0926_/A vssd1 vssd1 vccd1 vccd1 _0913_/B sky130_fd_sc_hd__or4_2
X_1299_ _1114_/X _1299_/D _0463__20/Y vssd1 vssd1 vccd1 vccd1 _1299_/Q sky130_fd_sc_hd__dfrtp_2
X_1368_ _1368_/A vssd1 vssd1 vccd1 vccd1 _1368_/X sky130_fd_sc_hd__clkbuf_1
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
+ _1187_/Q _0773_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0981__A2 _0973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1303__CLK _1118_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0670_ _1302_/Q vssd1 vssd1 vccd1 vccd1 _1301_/D sky130_fd_sc_hd__clkinv_2
XFILLER_11_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1084_ _1130_/A _1130_/B vssd1 vssd1 vccd1 vccd1 _1084_/Y sky130_fd_sc_hd__xnor2_1
X_1153_ _1153_/CLK _1153_/D fanout44/X vssd1 vssd1 vccd1 vccd1 _1153_/Q sky130_fd_sc_hd__dfrtp_1
X_1222_ _1359_/A _1222_/D fanout53/X vssd1 vssd1 vccd1 vccd1 _1222_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0517__A _1142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0868_ _0868_/A _0868_/B _0868_/C vssd1 vssd1 vccd1 vccd1 _0868_/X sky130_fd_sc_hd__or3_1
X_0799_ _1223_/Q _0799_/B vssd1 vssd1 vccd1 vccd1 _0800_/B sky130_fd_sc_hd__nor2_1
X_0937_ _1290_/Q _1348_/D vssd1 vssd1 vccd1 vccd1 _0937_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__1083__A _1097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0722_ _0719_/X _0720_/Y _0998_/A vssd1 vssd1 vccd1 vccd1 _0723_/B sky130_fd_sc_hd__o21ai_1
XFILLER_8_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0653_ _1267_/Q vssd1 vssd1 vccd1 vccd1 _1268_/D sky130_fd_sc_hd__inv_2
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0584_ _1130_/B _0585_/B vssd1 vssd1 vccd1 vccd1 _1170_/D sky130_fd_sc_hd__xnor2_1
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1205_ _0879_/A _1205_/D _0486_/Y vssd1 vssd1 vccd1 vccd1 _1205_/Q sky130_fd_sc_hd__dfrtp_1
X_1067_ _1079_/A vssd1 vssd1 vccd1 vccd1 _1077_/A sky130_fd_sc_hd__buf_6
XFILLER_21_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0863__A1 _0560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0636_ _1249_/Q vssd1 vssd1 vccd1 vccd1 _1248_/D sky130_fd_sc_hd__inv_2
X_0705_ _1193_/Q _1192_/Q _1191_/Q _0751_/A vssd1 vssd1 vccd1 vccd1 _0738_/B sky130_fd_sc_hd__or4_1
XFILLER_26_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1361__A _1363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0567_ _1135_/A _0567_/B vssd1 vssd1 vccd1 vccd1 _1165_/D sky130_fd_sc_hd__xnor2_1
X_0498_ _0548_/A vssd1 vssd1 vccd1 vccd1 _0542_/B sky130_fd_sc_hd__inv_2
XANTENNA__1261__RESET_B fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0790__B1 _0716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1349__RESET_B fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1194__CLK fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0619_ _1214_/Q vssd1 vssd1 vccd1 vccd1 _1215_/D sky130_fd_sc_hd__clkinv_2
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0454__12 _0448__6/A vssd1 vssd1 vccd1 vccd1 _0454__12/Y sky130_fd_sc_hd__inv_2
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_69 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0970_ _1314_/Q _0970_/B vssd1 vssd1 vccd1 vccd1 _0970_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1086__A _1132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0702__B _1178_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout58_A fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0736__B1 _0716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1232__CLK _1357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1325__SET_B fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1148_/CLK fanout41/X vssd1 vssd1 vccd1 vccd1 _1368_/A sky130_fd_sc_hd__dlrtn_1
X_0953_ _1310_/Q _1309_/Q vssd1 vssd1 vccd1 vccd1 _0953_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__0975__B1 _0755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0884_ _1290_/Q _1348_/D _1288_/Q _1287_/Q vssd1 vssd1 vccd1 vccd1 _0926_/A sky130_fd_sc_hd__or4_1
X_1367_ _1367_/A vssd1 vssd1 vccd1 vccd1 _1367_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1298_ _1045_/A _1298_/D _1113__51/Y vssd1 vssd1 vccd1 vccd1 _1298_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0713__A _1185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1255__CLK input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1221_ _1357_/A _1221_/D fanout55/X vssd1 vssd1 vccd1 vccd1 _1221_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1152_ _1168_/CLK _1152_/D fanout43/X vssd1 vssd1 vccd1 vccd1 _1152_/Q sky130_fd_sc_hd__dfrtp_1
X_1083_ _1097_/A vssd1 vssd1 vccd1 vccd1 _1083_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0517__B _1142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0533__A _0862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0936_ _1287_/Q _0936_/B vssd1 vssd1 vccd1 vccd1 _1287_/D sky130_fd_sc_hd__xnor2_1
X_0867_ _0546_/A _0554_/Y _1035_/D _0874_/D vssd1 vssd1 vccd1 vccd1 _0868_/C sky130_fd_sc_hd__o211a_1
X_0798_ _1220_/Q _0798_/B vssd1 vssd1 vccd1 vccd1 _1220_/D sky130_fd_sc_hd__xnor2_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_A
+ _1187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0583_ _0590_/C _0644_/C vssd1 vssd1 vccd1 vccd1 _0585_/B sky130_fd_sc_hd__nand2_4
X_0721_ _0755_/A vssd1 vssd1 vccd1 vccd1 _0998_/A sky130_fd_sc_hd__buf_4
X_0652_ _1268_/Q vssd1 vssd1 vccd1 vccd1 _1267_/D sky130_fd_sc_hd__clkinv_2
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1204_ _0590_/C _1204_/D _1071_/Y vssd1 vssd1 vccd1 vccd1 _1204_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_26_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0528__A _0873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1066_ _1146_/A _1146_/B vssd1 vssd1 vccd1 vccd1 _1066_/Y sky130_fd_sc_hd__xnor2_4
X_1135_ _1135_/A _1135_/B vssd1 vssd1 vccd1 vccd1 _1135_/X sky130_fd_sc_hd__xor2_1
XFILLER_22_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0919_ _1282_/Q _0919_/B vssd1 vssd1 vccd1 vccd1 _1282_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__1078__B _1264_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1094__A _1097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout40_A _1363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0872__A2 _0871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0863__A2 _1035_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0566_ _1135_/B _0567_/B vssd1 vssd1 vccd1 vccd1 _1164_/D sky130_fd_sc_hd__xnor2_1
X_0635_ _1246_/Q vssd1 vssd1 vccd1 vccd1 _1247_/D sky130_fd_sc_hd__clkinv_2
X_0704_ _1255_/D _1197_/Q _1195_/Q _1194_/Q vssd1 vssd1 vccd1 vccd1 _0751_/A sky130_fd_sc_hd__or4_1
XFILLER_7_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0497_ _1105_/A _1105_/B vssd1 vssd1 vccd1 vccd1 _0548_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__1089__A _1135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1118_ _1139_/A _1139_/B vssd1 vssd1 vccd1 vccd1 _1118_/X sky130_fd_sc_hd__xor2_2
XFILLER_22_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0721__A _0755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0806__A _1224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0549_ _1042_/B _0547_/X _0549_/S vssd1 vssd1 vccd1 vccd1 _0551_/B sky130_fd_sc_hd__mux2_1
X_0618_ _1215_/Q vssd1 vssd1 vccd1 vccd1 _1214_/D sky130_fd_sc_hd__inv_2
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_A _1277_/Q vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1372__A _1372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1091__B _1137_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0716__A _0831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_59 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout38/X fanout56/X vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0536__A _1135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1086__B _1132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf _1311_/Q _1022_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0952_ _1308_/Q _1307_/Q vssd1 vssd1 vccd1 vccd1 _0952_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0975__A1 _0970_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0883_ _1274_/Q _1273_/Q vssd1 vssd1 vccd1 vccd1 _0883_/Y sky130_fd_sc_hd__xnor2_4
X_1366_ _1366_/A vssd1 vssd1 vccd1 vccd1 _1366_/X sky130_fd_sc_hd__clkbuf_1
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1168_/CLK fanout43/X vssd1 vssd1 vccd1 vccd1 _1366_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_23_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1297_ _1112_/X _1297_/D _0464__21/Y vssd1 vssd1 vccd1 vccd1 _1297_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1097__A _1097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1151_ _1168_/CLK _1151_/D fanout43/X vssd1 vssd1 vccd1 vccd1 _1151_/Q sky130_fd_sc_hd__dfrtp_4
X_1220_ fanout34/X _1220_/D fanout57/X vssd1 vssd1 vccd1 vccd1 _1220_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_2_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1049__32 _1049__32/A vssd1 vssd1 vccd1 vccd1 _1155_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1082_ _1128_/A _1128_/B vssd1 vssd1 vccd1 vccd1 _1082_/Y sky130_fd_sc_hd__xnor2_1
X_0866_ _1042_/A _0866_/B vssd1 vssd1 vccd1 vccd1 _1035_/D sky130_fd_sc_hd__or2_1
XFILLER_9_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0814__A _1013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0935_ _0932_/Y _0934_/X _0831_/X vssd1 vssd1 vccd1 vccd1 _0936_/B sky130_fd_sc_hd__a21o_1
XANTENNA__0533__B _1035_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0797_ _0796_/Y _0793_/B _0716_/X vssd1 vssd1 vccd1 vccd1 _0798_/B sky130_fd_sc_hd__a21o_1
XANTENNA__0708__B _1183_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1255__RESET_B fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1349_ input7/X _1349_/D fanout50/X vssd1 vssd1 vccd1 vccd1 _1350_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_25_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0724__A _1185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0875__B1 _1042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0720_ _1184_/Q _0720_/B vssd1 vssd1 vccd1 vccd1 _0720_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0651_ _1262_/Q vssd1 vssd1 vccd1 vccd1 _1262_/D sky130_fd_sc_hd__inv_2
X_0582_ _0868_/A _0590_/B vssd1 vssd1 vccd1 vccd1 _0644_/C sky130_fd_sc_hd__nor2_2
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1203_ _0644_/B _1203_/D _0487_/Y vssd1 vssd1 vccd1 vccd1 _1203_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0544__A _1144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1043__B1 _0868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0849_ _1251_/Q _1250_/Q vssd1 vssd1 vccd1 vccd1 _0849_/Y sky130_fd_sc_hd__xnor2_2
X_0918_ _0998_/A _0918_/B vssd1 vssd1 vccd1 vccd1 _0919_/B sky130_fd_sc_hd__nand2_1
XANTENNA__1245__CLK _0868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[0\].w1.ro_block_I.ro_pol_eve.tribuf.t_buf _0859_/A _0703_/Y vssd1
+ vssd1 vccd1 vccd1 _1371_/A sky130_fd_sc_hd__ebufn_2
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0719__A _1185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout33_A fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1268__CLK _0542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0490__25 _0490__25/A vssd1 vssd1 vccd1 vccd1 _0490__25/Y sky130_fd_sc_hd__inv_2
X_0703_ _1181_/Q _1180_/Q vssd1 vssd1 vccd1 vccd1 _0703_/Y sky130_fd_sc_hd__xnor2_1
X_0565_ _0568_/A _0873_/A _1035_/B vssd1 vssd1 vccd1 vccd1 _0567_/B sky130_fd_sc_hd__or3_2
X_0634_ _1247_/Q vssd1 vssd1 vccd1 vccd1 _1246_/D sky130_fd_sc_hd__inv_2
X_0496_ _1148_/Q vssd1 vssd1 vccd1 vccd1 _1105_/B sky130_fd_sc_hd__buf_2
XFILLER_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
+ _1222_/Q _0845_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_22_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1089__B _1135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0912__A _1280_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_GATE_N
+ _1099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0617_ _1212_/Q vssd1 vssd1 vccd1 vccd1 _1213_/D sky130_fd_sc_hd__clkinv_2
X_0548_ _0548_/A _0548_/B _0548_/C vssd1 vssd1 vccd1 vccd1 _0549_/S sky130_fd_sc_hd__and3_1
X_0479_ _0479_/A vssd1 vssd1 vccd1 vccd1 _0479_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1306__CLK _1121_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0460__17 _0490__25/A vssd1 vssd1 vccd1 vccd1 _0460__17/Y sky130_fd_sc_hd__inv_2
XANTENNA__1192__RESET_B fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0536__B _1135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0552__A _1042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout38/X fanout57/X vssd1 vssd1 vccd1 vccd1 _1367_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input5_A phi1b_dig_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0727__A _1187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1329__CLK _0581_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.ro_block_Q.ro_pol_eve.tribuf.t_buf _1027_/A _0881_/Y vssd1 vssd1 vccd1 vccd1 _1373_/A
+ sky130_fd_sc_hd__ebufn_4
X_0951_ _1306_/Q _1305_/Q vssd1 vssd1 vccd1 vccd1 _0951_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0882_ _1272_/Q _1271_/Q vssd1 vssd1 vccd1 vccd1 _0882_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__1353__D _1353_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1365_ _1365_/A vssd1 vssd1 vccd1 vccd1 _1365_/X sky130_fd_sc_hd__clkbuf_1
X_1296_ _1111_/Y _1296_/D _0465__22/Y vssd1 vssd1 vccd1 vccd1 _1296_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0713__C _1183_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1147__5_A _1122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0920__A _1284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1150_ _1150_/CLK _1150_/D fanout44/X vssd1 vssd1 vccd1 vccd1 _1150_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1081_ _1097_/A vssd1 vssd1 vccd1 vccd1 _1081_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0865_ _0865_/A _0873_/B _0865_/C vssd1 vssd1 vccd1 vccd1 _0865_/X sky130_fd_sc_hd__and3_1
XANTENNA__1348__D _1348_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0934_ _1288_/Q _0934_/B vssd1 vssd1 vccd1 vccd1 _0934_/X sky130_fd_sc_hd__or2_1
X_0796_ _1221_/Q _0796_/B vssd1 vssd1 vccd1 vccd1 _0796_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1174__CLK _1035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1279_ _1356_/A _1279_/D fanout46/X vssd1 vssd1 vccd1 vccd1 _1279_/Q sky130_fd_sc_hd__dfrtp_4
X_1348_ input7/X _1348_/D fanout50/X vssd1 vssd1 vccd1 vccd1 _1349_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_25_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0875__A1 _0560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0650__A _1265_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0581_ _0644_/B vssd1 vssd1 vccd1 vccd1 _0581_/Y sky130_fd_sc_hd__clkinv_2
X_0650_ _1265_/Q _0650_/B vssd1 vssd1 vccd1 vccd1 _1266_/D sky130_fd_sc_hd__xnor2_1
XFILLER_3_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1202_ _0581_/Y _1202_/D _1070_/Y vssd1 vssd1 vccd1 vccd1 _1202_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1064_ _1146_/A _1146_/B vssd1 vssd1 vccd1 vccd1 _1064_/Y sky130_fd_sc_hd__xnor2_1
X_1133_ _1133_/A _1133_/B vssd1 vssd1 vccd1 vccd1 _1133_/X sky130_fd_sc_hd__xor2_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0560__A _0560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0779_ _1217_/Q _1216_/Q vssd1 vssd1 vccd1 vccd1 _0779_/Y sky130_fd_sc_hd__xnor2_2
X_0848_ _1249_/Q _1248_/Q vssd1 vssd1 vccd1 vccd1 _0848_/Y sky130_fd_sc_hd__xnor2_2
X_0917_ _1284_/Q _1283_/Q _0920_/B _0914_/B vssd1 vssd1 vccd1 vccd1 _0918_/B sky130_fd_sc_hd__a31o_1
XFILLER_1_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0735__A _1188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0470__A _0479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf _1319_/Q _1014_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_15_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0702_ _1179_/Q _1178_/Q vssd1 vssd1 vccd1 vccd1 _0702_/Y sky130_fd_sc_hd__xnor2_2
X_0633_ _1244_/Q vssd1 vssd1 vccd1 vccd1 _1245_/D sky130_fd_sc_hd__clkinv_2
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0495_ _1149_/Q vssd1 vssd1 vccd1 vccd1 _1105_/A sky130_fd_sc_hd__clkbuf_4
X_0564_ _0873_/B vssd1 vssd1 vccd1 vccd1 _0868_/B sky130_fd_sc_hd__inv_2
X_0466__23 _0490__25/A vssd1 vssd1 vccd1 vccd1 _0466__23/Y sky130_fd_sc_hd__inv_2
XANTENNA__1212__CLK _0873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1116_ _1137_/A _1137_/B vssd1 vssd1 vccd1 vccd1 _1116_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0616_ _1213_/Q vssd1 vssd1 vccd1 vccd1 _1212_/D sky130_fd_sc_hd__inv_2
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0547_ _0865_/A _0547_/B vssd1 vssd1 vccd1 vccd1 _0547_/X sky130_fd_sc_hd__or2_1
X_0478_ _0479_/A vssd1 vssd1 vccd1 vccd1 _0478_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1258__CLK input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0642__B _1264_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0911__B1 _0831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0552__B _0873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_0__0306__A _0445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0743__A _1013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0918__A _0998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
+ _1184_/Q _0776_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_0950_ _1304_/Q _1303_/Q vssd1 vssd1 vccd1 vccd1 _0950_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0881_ _1270_/Q _1269_/Q vssd1 vssd1 vccd1 vccd1 _0881_/Y sky130_fd_sc_hd__xnor2_2
X_1364_ _1364_/A vssd1 vssd1 vccd1 vccd1 _1364_/X sky130_fd_sc_hd__clkbuf_1
X_1295_ _0590_/C _1295_/D _1110__50/Y vssd1 vssd1 vccd1 vccd1 _1295_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__0828__A _1259_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0563__A _1137_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0473__A _0479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1080_ _1097_/A vssd1 vssd1 vccd1 vccd1 _1080_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0864_ _0546_/A _1035_/C _0862_/Y _0863_/X vssd1 vssd1 vccd1 vccd1 _0864_/X sky130_fd_sc_hd__o31a_1
XFILLER_13_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0795_ _1219_/Q _0795_/B vssd1 vssd1 vccd1 vccd1 _1219_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0933_ _1290_/Q _1348_/D vssd1 vssd1 vccd1 vccd1 _0934_/B sky130_fd_sc_hd__or2_1
XANTENNA__0558__A _0873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1347_ input7/X input3/X fanout50/X vssd1 vssd1 vccd1 vccd1 _1348_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1278_ _1326_/CLK _1278_/D fanout48/X vssd1 vssd1 vccd1 vccd1 _1278_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1055__37 _1058__40/A vssd1 vssd1 vccd1 vccd1 _1165_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__1264__RESET_B fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1168_/CLK fanout41/X vssd1 vssd1 vccd1 vccd1 _1368_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0468__A _1099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0580_ _1130_/A _1130_/B vssd1 vssd1 vccd1 vccd1 _0644_/B sky130_fd_sc_hd__xnor2_2
X_1201_ _0589_/A _1201_/D _0488_/Y vssd1 vssd1 vccd1 vccd1 _1201_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1132_ _1132_/A _1132_/B vssd1 vssd1 vccd1 vccd1 _1132_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0916_ _1281_/Q _0916_/B vssd1 vssd1 vccd1 vccd1 _1281_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__0560__B _0560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0778_ _1215_/Q _1214_/Q vssd1 vssd1 vccd1 vccd1 _0778_/Y sky130_fd_sc_hd__xnor2_2
X_0847_ _1247_/Q _1246_/Q vssd1 vssd1 vccd1 vccd1 _0847_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1291__CLK _0644_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1115__52 _1117__53/A vssd1 vssd1 vccd1 vccd1 _1115__52/Y sky130_fd_sc_hd__inv_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0449__7 _0451__9/A vssd1 vssd1 vccd1 vccd1 _0449__7/Y sky130_fd_sc_hd__inv_2
XFILLER_16_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0645__B _0646_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0563_ _1137_/B _0563_/B vssd1 vssd1 vccd1 vccd1 _1163_/D sky130_fd_sc_hd__xnor2_1
X_0701_ _1177_/Q _1176_/Q vssd1 vssd1 vccd1 vccd1 _0701_/Y sky130_fd_sc_hd__xnor2_2
X_0632_ _1245_/Q vssd1 vssd1 vccd1 vccd1 _1244_/D sky130_fd_sc_hd__inv_2
XFILLER_11_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0481__A _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1187__CLK fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0546_ _0546_/A _1042_/B vssd1 vssd1 vccd1 vccd1 _0547_/B sky130_fd_sc_hd__nor2_1
X_0615_ _1210_/Q vssd1 vssd1 vccd1 vccd1 _1211_/D sky130_fd_sc_hd__clkinv_2
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0566__A _1135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0477_ _0479_/A vssd1 vssd1 vccd1 vccd1 _0477_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1029_ _1354_/Q _1353_/D vssd1 vssd1 vccd1 vccd1 _1030_/A sky130_fd_sc_hd__and2b_1
XFILLER_22_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0476__A _0479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1100__A _1122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1202__CLK _0581_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1352__CLK input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0529_ _1163_/Q vssd1 vssd1 vccd1 vccd1 _1137_/A sky130_fd_sc_hd__buf_4
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf _1281_/Q _0946_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0880_ _1268_/Q _1267_/Q vssd1 vssd1 vccd1 vccd1 _0880_/Y sky130_fd_sc_hd__xnor2_2
X_1363_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1363_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1294_ _1109_/Y _1294_/D _0466__23/Y vssd1 vssd1 vccd1 vccd1 _1294_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__0648__A0 _0644_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1248__CLK _1093_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0820__B1 _0755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout49_A fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0811__B1 _0755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0932_ _1290_/Q _1348_/D _1288_/Q vssd1 vssd1 vccd1 vccd1 _0932_/Y sky130_fd_sc_hd__nand3_1
X_0863_ _0560_/A _1035_/B _1042_/A vssd1 vssd1 vccd1 vccd1 _0863_/X sky130_fd_sc_hd__a21o_1
X_0794_ _0792_/X _0793_/Y _0755_/X vssd1 vssd1 vccd1 vccd1 _0795_/B sky130_fd_sc_hd__o21ai_1
XFILLER_9_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0869__B1 _0865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0558__B _0874_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1346_ _1146_/Y _1346_/D _0446__1/Y vssd1 vssd1 vccd1 vccd1 _1346_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1277_ _1325_/CLK _1277_/D fanout48/X vssd1 vssd1 vccd1 vccd1 _1277_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0875__A3 _0868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0484__A _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1168_/CLK fanout43/X vssd1 vssd1 vccd1 vccd1 _1366_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1200_ _0644_/D _1200_/D _1069_/Y vssd1 vssd1 vccd1 vccd1 _1200_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1062_ _1146_/A _1146_/B vssd1 vssd1 vccd1 vccd1 _1062_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0915_ _0910_/B _0914_/X _0755_/X vssd1 vssd1 vccd1 vccd1 _0916_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__1002__B _1352_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0777_ _1213_/Q _1212_/Q vssd1 vssd1 vccd1 vccd1 _0777_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__0569__A _1133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0846_ _1245_/Q _1244_/Q vssd1 vssd1 vccd1 vccd1 _0846_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1329_ _0581_/Y _1329_/D _1129__59/Y vssd1 vssd1 vccd1 vccd1 _1329_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0479__A _0479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1103__A _1105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1309__CLK _1035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0700_ _1175_/Q _1174_/Q vssd1 vssd1 vccd1 vccd1 _0700_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_16_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.ro_block_I.ro_pol_eve.tribuf.t_buf _1032_/A _0883_/Y vssd1 vssd1 vccd1 vccd1 _1371_/A
+ sky130_fd_sc_hd__ebufn_2
X_0562_ _1137_/A _0563_/B vssd1 vssd1 vccd1 vccd1 _1162_/D sky130_fd_sc_hd__xnor2_1
X_0631_ _1242_/Q vssd1 vssd1 vccd1 vccd1 _1243_/D sky130_fd_sc_hd__inv_2
XFILLER_7_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1114_ _1135_/A _1135_/B vssd1 vssd1 vccd1 vccd1 _1114_/X sky130_fd_sc_hd__xor2_1
XANTENNA__0941__C1 _0831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1045_ _1045_/A _1045_/B vssd1 vssd1 vccd1 vccd1 _1364_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__1013__A _1013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0829_ _1259_/D _1233_/Q vssd1 vssd1 vccd1 vccd1 _0830_/B sky130_fd_sc_hd__or2_1
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[0\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf_TE_B _0701_/Y
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout31_A fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0451__9 _0451__9/A vssd1 vssd1 vccd1 vccd1 _0451__9/Y sky130_fd_sc_hd__inv_2
XFILLER_5_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0937__A _1290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0476_ _0479_/A vssd1 vssd1 vccd1 vccd1 _0476_/Y sky130_fd_sc_hd__inv_2
X_0545_ _1042_/A _0560_/A vssd1 vssd1 vccd1 vccd1 _0865_/A sky130_fd_sc_hd__nor2_1
X_0614_ _1211_/Q vssd1 vssd1 vccd1 vccd1 _1210_/D sky130_fd_sc_hd__clkinv_2
XFILLER_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1028_ _1028_/A vssd1 vssd1 vccd1 vccd1 _1028_/X sky130_fd_sc_hd__clkbuf_1
Xwrapper_cell_loop\[0\].w1.ro_block_I.ro_pol.tribuf.t_buf _0860_/X _0702_/Y vssd1
+ vssd1 vccd1 vccd1 _1370_/A sky130_fd_sc_hd__ebufn_2
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0987__A2 _1319_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1170__RESET_B fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1258__RESET_B fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0577__A _1132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0528_ _0873_/A vssd1 vssd1 vccd1 vccd1 _0862_/A sky130_fd_sc_hd__inv_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0487__A _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1111__A _1132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1293_ _0581_/Y _1293_/D _1108__49/Y vssd1 vssd1 vccd1 vccd1 _1293_/Q sky130_fd_sc_hd__dfrtp_2
X_1362_ _1362_/A vssd1 vssd1 vccd1 vccd1 _1362_/X sky130_fd_sc_hd__buf_2
XANTENNA__1351__RESET_B fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0648__A1 _0585_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1021__A _1342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input3_A comp_high_Q[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__0311_ clkbuf_0__0311_/X vssd1 vssd1 vccd1 vccd1 _1052__35/A sky130_fd_sc_hd__clkbuf_16
XFILLER_10_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0878__A1 _1045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0945__A _1294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1136__62 _1141__65/A vssd1 vssd1 vccd1 vccd1 _1136__62/Y sky130_fd_sc_hd__inv_2
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1079_/A fanout57/X vssd1 vssd1 vccd1 vccd1 _1367_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0862_ _0862_/A _1035_/B vssd1 vssd1 vccd1 vccd1 _0862_/Y sky130_fd_sc_hd__nor2_1
X_0931_ _1286_/Q _0931_/B vssd1 vssd1 vccd1 vccd1 _1286_/D sky130_fd_sc_hd__xnor2_1
X_0793_ _1220_/Q _0793_/B vssd1 vssd1 vccd1 vccd1 _0793_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__0869__A1 _0873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0869__B2 _1045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1016__A _1332_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1345_ _1035_/A _1345_/D _1145__4/Y vssd1 vssd1 vccd1 vccd1 _1345_/Q sky130_fd_sc_hd__dfrtp_1
X_1276_ _1325_/CLK _1276_/D fanout48/X vssd1 vssd1 vccd1 vccd1 _1276_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__1215__CLK _1042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1037__A1 _0871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1037__B2 _0873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1238__CLK _0581_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1130_ _1130_/A _1130_/B vssd1 vssd1 vccd1 vccd1 _1130_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_19_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0845_ _1243_/Q _1242_/Q vssd1 vssd1 vccd1 vccd1 _0845_/Y sky130_fd_sc_hd__xnor2_2
X_0914_ _1282_/Q _0914_/B vssd1 vssd1 vccd1 vccd1 _0914_/X sky130_fd_sc_hd__and2b_1
X_1060__42 _1065__45/A vssd1 vssd1 vccd1 vccd1 _1060__42/Y sky130_fd_sc_hd__inv_2
X_0776_ _1211_/Q _1210_/Q vssd1 vssd1 vccd1 vccd1 _0776_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__0569__B _0570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1259_ input6/X _1259_/D fanout53/X vssd1 vssd1 vccd1 vccd1 _1260_/D sky130_fd_sc_hd__dfrtp_1
XANTENNA__0585__A _1130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1328_ _1128_/Y _1328_/D _0456__14/Y vssd1 vssd1 vccd1 vccd1 _1328_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
+ _1219_/Q _0848_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_4_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0561_ _0865_/C _1035_/B _0568_/A vssd1 vssd1 vccd1 vccd1 _0563_/B sky130_fd_sc_hd__mux2_1
X_0630_ _1243_/Q vssd1 vssd1 vccd1 vccd1 _1242_/D sky130_fd_sc_hd__clkinv_2
XFILLER_19_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1044_ _0873_/B _1035_/X _1040_/B _1043_/X vssd1 vssd1 vccd1 vccd1 _1045_/B sky130_fd_sc_hd__o22a_2
XFILLER_0_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_2__f_clk_master clkbuf_0_clk_master/X vssd1 vssd1 vccd1 vccd1 _1362_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_21_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0828_ _1259_/D _1233_/Q _1231_/Q vssd1 vssd1 vccd1 vccd1 _0828_/Y sky130_fd_sc_hd__nand3_1
X_0759_ _1255_/D _1197_/Q vssd1 vssd1 vccd1 vccd1 _0760_/B sky130_fd_sc_hd__or2_1
X_0457__15 _0448__6/A vssd1 vssd1 vccd1 vccd1 _0457__15/Y sky130_fd_sc_hd__inv_2
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1114__A _1135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0937__B _1348_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0953__A _1310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0613_ _1208_/Q vssd1 vssd1 vccd1 vccd1 _1209_/D sky130_fd_sc_hd__clkinv_2
XFILLER_8_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0544_ _1144_/A _0544_/B vssd1 vssd1 vccd1 vccd1 _1157_/D sky130_fd_sc_hd__xnor2_1
X_0475_ _0479_/A vssd1 vssd1 vccd1 vccd1 _0475_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1027_ _1027_/A _1027_/B vssd1 vssd1 vccd1 vccd1 _1028_/A sky130_fd_sc_hd__or2_1
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0582__B _0590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0905__B1 _0755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1109__A _1130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0683__A _1329_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1019__A _1338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_A _1315_/Q vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0458_ _1122_/A vssd1 vssd1 vccd1 vccd1 _0458_/X sky130_fd_sc_hd__buf_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0527_ _1139_/A _1139_/B vssd1 vssd1 vccd1 vccd1 _0873_/A sky130_fd_sc_hd__xor2_4
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0593__A _0593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1111__B _1132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf_TE_B _0952_/Y vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0678__A _1310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1292_ _1107_/Y _1292_/D _0467__24/Y vssd1 vssd1 vccd1 vccd1 _1292_/Q sky130_fd_sc_hd__dfrtp_2
X_1361_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1361_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0588__A _1128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0878__A2 _0865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1122__A _1122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0945__B _1293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0861_ _1034_/B _1262_/D vssd1 vssd1 vccd1 vccd1 _0861_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0792_ _1221_/Q _1220_/Q _0796_/B vssd1 vssd1 vccd1 vccd1 _0792_/X sky130_fd_sc_hd__and3_1
XFILLER_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0930_ _0890_/C _0926_/Y _0755_/A vssd1 vssd1 vccd1 vccd1 _0931_/B sky130_fd_sc_hd__o21ai_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1016__B _1331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1344_ _1144_/Y _1344_/D _0448__6/Y vssd1 vssd1 vccd1 vccd1 _1344_/Q sky130_fd_sc_hd__dfrtp_2
X_1275_ _1325_/CLK _1275_/D fanout46/X vssd1 vssd1 vccd1 vccd1 _1275_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0871__A _0873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0590__B _0590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout54_A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1046__29 _1049__32/A vssd1 vssd1 vccd1 vccd1 _1149_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0956__A _1319_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0691__A _1337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0493__27 _1049__32/A vssd1 vssd1 vccd1 vccd1 _0493__27/Y sky130_fd_sc_hd__inv_2
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0775_ _1209_/Q _1208_/Q vssd1 vssd1 vccd1 vccd1 _0775_/Y sky130_fd_sc_hd__xnor2_2
X_0844_ _1241_/Q _1240_/Q vssd1 vssd1 vccd1 vccd1 _0844_/Y sky130_fd_sc_hd__xnor2_2
X_0913_ _1283_/Q _0913_/B vssd1 vssd1 vccd1 vccd1 _0914_/B sky130_fd_sc_hd__nor2_1
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf _1316_/Q _1017_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
X_1258_ input6/X input2/X fanout59/X vssd1 vssd1 vccd1 vccd1 _1259_/D sky130_fd_sc_hd__dfrtp_4
XANTENNA__0585__B _0585_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1327_ _0644_/D _1327_/D _1127__58/Y vssd1 vssd1 vccd1 vccd1 _1327_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__0866__A _1042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1189_ fanout31/X _1189_/D fanout50/X vssd1 vssd1 vccd1 vccd1 _1189_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_4_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0491_ _1053_/A vssd1 vssd1 vccd1 vccd1 _0491_/X sky130_fd_sc_hd__buf_1
X_0560_ _0560_/A _0560_/B vssd1 vssd1 vccd1 vccd1 _0568_/A sky130_fd_sc_hd__or2_1
XFILLER_3_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0686__A _1334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1112_ _1133_/A _1133_/B vssd1 vssd1 vccd1 vccd1 _1112_/X sky130_fd_sc_hd__xor2_1
X_1043_ _1036_/X _1042_/X _0868_/B vssd1 vssd1 vccd1 vccd1 _1043_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1362_/A fanout41/X vssd1 vssd1 vccd1 vccd1 _1368_/A sky130_fd_sc_hd__dlrtn_1
X_0827_ _1229_/Q _0827_/B vssd1 vssd1 vccd1 vccd1 _1229_/D sky130_fd_sc_hd__xnor2_1
X_0758_ _1255_/D _1197_/Q _1195_/Q vssd1 vssd1 vccd1 vccd1 _0758_/Y sky130_fd_sc_hd__nand3_1
X_0689_ _1335_/Q vssd1 vssd1 vccd1 vccd1 _1336_/D sky130_fd_sc_hd__inv_2
XFILLER_25_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1228__CLK _1357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1114__B _1135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1130__A _1130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0612_ _1209_/Q vssd1 vssd1 vccd1 vccd1 _1208_/D sky130_fd_sc_hd__clkinv_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0543_ _1144_/B _0544_/B vssd1 vssd1 vccd1 vccd1 _1156_/D sky130_fd_sc_hd__xnor2_1
X_0474_ _0479_/A vssd1 vssd1 vccd1 vccd1 _0474_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1026_ _1349_/D _1350_/Q vssd1 vssd1 vccd1 vccd1 _1027_/B sky130_fd_sc_hd__and2b_1
XFILLER_2_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1109__B _1130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.ro_block_Q.ro_pol.tribuf.t_buf _1028_/X _0880_/Y vssd1 vssd1 vccd1 vccd1 _1372_/A
+ sky130_fd_sc_hd__ebufn_4
XFILLER_5_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0832__B1 _0831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1019__B _1337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0526_ _1160_/Q vssd1 vssd1 vccd1 vccd1 _1139_/B sky130_fd_sc_hd__buf_4
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
+ _1196_/Q _0779_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1035__A _1035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1009_ _1324_/Q _1009_/B vssd1 vssd1 vccd1 vccd1 _1324_/D sky130_fd_sc_hd__xnor2_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1000__B1 _0755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1360_ _1360_/A vssd1 vssd1 vccd1 vccd1 _1360_/X sky130_fd_sc_hd__buf_2
XANTENNA__0694__A _1342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1291_ _0644_/D _1291_/D _1106__48/Y vssd1 vssd1 vccd1 vccd1 _1291_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0509_ _1146_/B _0510_/B vssd1 vssd1 vccd1 vccd1 _1152_/D sky130_fd_sc_hd__xnor2_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_A
+ _1188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0588__B _1128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0961__B _1319_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1189__RESET_B fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0860_ _0860_/A vssd1 vssd1 vccd1 vccd1 _0860_/X sky130_fd_sc_hd__clkbuf_1
X_0791_ _1218_/Q _0791_/B vssd1 vssd1 vccd1 vccd1 _1218_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1343_ _1042_/A _1343_/D _1143__3/Y vssd1 vssd1 vccd1 vccd1 _1343_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1274_ _0542_/B _1274_/D _1148_/CLK vssd1 vssd1 vccd1 vccd1 _1274_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__0590__C _0590_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0871__B _0873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1261__CLK input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0599__A _1178_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0989_ _1318_/Q _0989_/B vssd1 vssd1 vccd1 vccd1 _1318_/D sky130_fd_sc_hd__xnor2_1
XFILLER_27_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout47_A fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1133__A _1133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0972__A _1313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0912_ _1280_/Q _0912_/B vssd1 vssd1 vccd1 vccd1 _1280_/D sky130_fd_sc_hd__xnor2_1
X_0843_ _1239_/Q _1238_/Q vssd1 vssd1 vccd1 vccd1 _0843_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__0539__A2 _0590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0774_ _1207_/Q _1206_/Q vssd1 vssd1 vccd1 vccd1 _0774_/Y sky130_fd_sc_hd__xnor2_2
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1099_/A fanout55/X vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_25_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__0311_ _0491_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0311_/X sky130_fd_sc_hd__clkbuf_16
X_1326_ _1326_/CLK _1326_/D fanout49/X vssd1 vssd1 vccd1 vccd1 _1326_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1257_ input8/X _1257_/D fanout52/X vssd1 vssd1 vccd1 vccd1 _1257_/Q sky130_fd_sc_hd__dfrtp_1
X_1188_ fanout31/X _1188_/D fanout54/X vssd1 vssd1 vccd1 vccd1 _1188_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1128__A _1128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0967__A _1313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1111_ _1132_/A _1132_/B vssd1 vssd1 vccd1 vccd1 _1111_/Y sky130_fd_sc_hd__xnor2_1
X_1042_ _1042_/A _1042_/B _1042_/C vssd1 vssd1 vccd1 vccd1 _1042_/X sky130_fd_sc_hd__or3_1
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0688_ _1336_/Q vssd1 vssd1 vccd1 vccd1 _1335_/D sky130_fd_sc_hd__inv_2
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0757_ _1193_/Q _0757_/B vssd1 vssd1 vccd1 vccd1 _1193_/D sky130_fd_sc_hd__xnor2_1
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_A _1278_/Q vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0826_ _0786_/C _0822_/Y _0755_/X vssd1 vssd1 vccd1 vccd1 _0827_/B sky130_fd_sc_hd__o21ai_1
X_1309_ _1035_/A _1309_/D _1125__57/Y vssd1 vssd1 vccd1 vccd1 _1309_/Q sky130_fd_sc_hd__dfrtp_2
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1168_/CLK fanout42/X vssd1 vssd1 vccd1 vccd1 _1366_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_25_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0874__A_N _1035_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1130__B _1130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0542_ _0548_/C _0542_/B _0548_/B vssd1 vssd1 vccd1 vccd1 _0544_/B sky130_fd_sc_hd__or3b_1
X_0611_ _1206_/Q vssd1 vssd1 vccd1 vccd1 _1207_/D sky130_fd_sc_hd__inv_2
XFILLER_4_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0473_ _0479_/A vssd1 vssd1 vccd1 vccd1 _0473_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1314__RESET_B fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1025_ _1025_/A vssd1 vssd1 vccd1 vccd1 _1027_/A sky130_fd_sc_hd__clkbuf_1
X_0809_ _1226_/Q _0809_/B vssd1 vssd1 vccd1 vccd1 _0810_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1345__CLK _1035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf _1278_/Q _0949_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0525_ _1161_/Q vssd1 vssd1 vccd1 vccd1 _1139_/A sky130_fd_sc_hd__buf_4
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1145__4_A _1053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1035__B _1035_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1218__CLK _1357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1008_ _1007_/Y _1004_/B _0831_/A vssd1 vssd1 vccd1 vccd1 _1009_/B sky130_fd_sc_hd__a21o_1
XFILLER_2_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0524__D_N _0548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0959__B _1352_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1290_ _1326_/CLK _1290_/D fanout48/X vssd1 vssd1 vccd1 vccd1 _1290_/Q sky130_fd_sc_hd__dfrtp_4
X_0508_ _0542_/B _0548_/B vssd1 vssd1 vccd1 vccd1 _0510_/B sky130_fd_sc_hd__nand2_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1190__CLK fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk_master clk_master vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk_master/X sky130_fd_sc_hd__clkbuf_16
XFILLER_23_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0790_ _0784_/X _0789_/Y _0716_/X vssd1 vssd1 vccd1 vccd1 _0791_/B sky130_fd_sc_hd__a21o_1
XFILLER_9_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1342_ _1142_/Y _1342_/D _0449__7/Y vssd1 vssd1 vccd1 vccd1 _1342_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__0971__B1 _0831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1273_ _1105_/Y _1273_/D _1362_/A vssd1 vssd1 vccd1 vccd1 _1273_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_1_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0988_ _0998_/A _0988_/B vssd1 vssd1 vccd1 vccd1 _0989_/B sky130_fd_sc_hd__nand2_1
XANTENNA_input1_A comp_high_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1133__B _1133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0842_ _1237_/Q _1236_/Q vssd1 vssd1 vccd1 vccd1 _0842_/Y sky130_fd_sc_hd__xnor2_2
X_0911_ _0910_/Y _0903_/B _0831_/X vssd1 vssd1 vccd1 vccd1 _0912_/B sky130_fd_sc_hd__a21o_1
X_0773_ _1205_/Q _1204_/Q vssd1 vssd1 vccd1 vccd1 _0773_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1325_ _1325_/CLK _1325_/D fanout49/X vssd1 vssd1 vccd1 vccd1 _1325_/Q sky130_fd_sc_hd__dfstp_1
X_1256_ input8/X _1256_/D fanout54/X vssd1 vssd1 vccd1 vccd1 _1257_/D sky130_fd_sc_hd__dfrtp_1
X_1187_ fanout31/X _1187_/D fanout52/X vssd1 vssd1 vccd1 vccd1 _1187_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1051__34 _1052__35/A vssd1 vssd1 vccd1 vccd1 _1159_/CLK sky130_fd_sc_hd__inv_2
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout38/X fanout57/X vssd1 vssd1 vccd1 vccd1 _1367_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__0549__S _0549_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0935__B1 _0831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
+ _1189_/Q _0771_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_15_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1128__B _1128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1144__A _1144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1173__RESET_B fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1041_ _1041_/A _1041_/B vssd1 vssd1 vccd1 vccd1 _1374_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__0983__A _1319_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1251__CLK _1096_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0825_ _1228_/Q _0825_/B vssd1 vssd1 vccd1 vccd1 _1228_/D sky130_fd_sc_hd__xnor2_1
X_0687_ _1333_/Q vssd1 vssd1 vccd1 vccd1 _1334_/D sky130_fd_sc_hd__inv_2
X_0756_ _0710_/C _0751_/Y _0755_/X vssd1 vssd1 vccd1 vccd1 _0757_/B sky130_fd_sc_hd__o21ai_1
XFILLER_6_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1308_ _1124_/Y _1308_/D _0459__16/Y vssd1 vssd1 vccd1 vccd1 _1308_/Q sky130_fd_sc_hd__dfrtp_2
X_1239_ _1084_/Y _1239_/D _0476_/Y vssd1 vssd1 vccd1 vccd1 _1239_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__0893__A _1278_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1274__CLK _0542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1139__A _1139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0978__A _0998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0541_ _1154_/Q _0541_/B vssd1 vssd1 vccd1 vccd1 _1155_/D sky130_fd_sc_hd__xnor2_1
X_0610_ _1207_/Q vssd1 vssd1 vccd1 vccd1 _1206_/D sky130_fd_sc_hd__clkinv_2
X_0472_ _0479_/A vssd1 vssd1 vccd1 vccd1 _0472_/Y sky130_fd_sc_hd__inv_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1354__RESET_B fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1024_ _1350_/Q _1349_/D vssd1 vssd1 vccd1 vccd1 _1025_/A sky130_fd_sc_hd__and2b_1
XFILLER_22_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0888__A _1277_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0808_ _1223_/Q _0808_/B vssd1 vssd1 vccd1 vccd1 _1223_/D sky130_fd_sc_hd__xnor2_1
X_0739_ _1189_/Q _0739_/B vssd1 vssd1 vccd1 vccd1 _0739_/X sky130_fd_sc_hd__and2b_1
XFILLER_26_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_A
+ _1183_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1035__C _1035_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0501__A _1105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0524_ _0542_/B _1035_/A _1042_/A _0548_/B vssd1 vssd1 vccd1 vccd1 _0560_/B sky130_fd_sc_hd__or4b_2
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1007_ _1326_/Q _1352_/D vssd1 vssd1 vccd1 vccd1 _1007_/Y sky130_fd_sc_hd__nand2_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_GATE_N
+ _1099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1147__5 _1122_/A vssd1 vssd1 vccd1 vccd1 _1355_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0507_ _0548_/C vssd1 vssd1 vccd1 vccd1 _1035_/A sky130_fd_sc_hd__inv_2
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0732__A1 _1188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1208__CLK _0873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1341_ _0560_/A _1341_/D _1141__65/Y vssd1 vssd1 vccd1 vccd1 _1341_/Q sky130_fd_sc_hd__dfrtp_2
X_1272_ _0542_/B _1272_/D _1148_/CLK vssd1 vssd1 vccd1 vccd1 _1272_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_1_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0987_ _1320_/Q _1319_/Q _0990_/B _0984_/B vssd1 vssd1 vccd1 vccd1 _0988_/B sky130_fd_sc_hd__a31o_1
XANTENNA__0896__A _1278_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1180__CLK _1035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0772_ _1203_/Q _1202_/Q vssd1 vssd1 vccd1 vccd1 _0772_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_15_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0910_ _1281_/Q _0910_/B vssd1 vssd1 vccd1 vccd1 _0910_/Y sky130_fd_sc_hd__nand2_1
X_0841_ _1235_/Q _1234_/Q vssd1 vssd1 vccd1 vccd1 _0841_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1186_ fanout31/X _1186_/D fanout52/X vssd1 vssd1 vccd1 vccd1 _1186_/Q sky130_fd_sc_hd__dfrtp_1
X_1255_ input8/X _1255_/D fanout54/X vssd1 vssd1 vccd1 vccd1 _1256_/D sky130_fd_sc_hd__dfrtp_1
X_1324_ _1326_/CLK _1324_/D fanout47/X vssd1 vssd1 vccd1 vccd1 _1324_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout52_A fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1144__B _1144_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1040_ _1040_/A _1040_/B vssd1 vssd1 vccd1 vccd1 _1041_/B sky130_fd_sc_hd__or2_2
XANTENNA__1310__D _1310_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0755_ _0755_/A vssd1 vssd1 vccd1 vccd1 _0755_/X sky130_fd_sc_hd__clkbuf_4
X_0824_ _1013_/A _0824_/B vssd1 vssd1 vccd1 vccd1 _0825_/B sky130_fd_sc_hd__nand2_1
XANTENNA__0917__A1 _1284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0686_ _1334_/Q vssd1 vssd1 vccd1 vccd1 _1333_/D sky130_fd_sc_hd__inv_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1070__A _1077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1307_ _0514_/Y _1307_/D _1123__56/Y vssd1 vssd1 vccd1 vccd1 _1307_/Q sky130_fd_sc_hd__dfrtp_4
X_1169_ _1169_/CLK _1169_/D fanout50/X vssd1 vssd1 vccd1 vccd1 _1169_/Q sky130_fd_sc_hd__dfrtp_1
X_1238_ _0581_/Y _1238_/D _1083_/Y vssd1 vssd1 vccd1 vccd1 _1238_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__0893__B _1277_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1139__B _1139_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0540_ _1155_/Q _0541_/B vssd1 vssd1 vccd1 vccd1 _1154_/D sky130_fd_sc_hd__xnor2_1
X_0471_ _0479_/A vssd1 vssd1 vccd1 vccd1 _0471_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1023_ _1346_/Q _1345_/Q vssd1 vssd1 vccd1 vccd1 _1023_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_15_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0835__B1 _0831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0807_ _0806_/Y _0799_/B _0716_/X vssd1 vssd1 vccd1 vccd1 _0808_/B sky130_fd_sc_hd__a21o_1
XANTENNA__0888__B _1276_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0738_ _1190_/Q _0738_/B vssd1 vssd1 vccd1 vccd1 _0739_/B sky130_fd_sc_hd__nor2_1
X_0669_ _1299_/Q vssd1 vssd1 vccd1 vccd1 _1300_/D sky130_fd_sc_hd__inv_2
XFILLER_25_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0826__B1 _0755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0453__11 _0448__6/A vssd1 vssd1 vccd1 vccd1 _0453__11/Y sky130_fd_sc_hd__inv_2
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1148_/CLK fanout41/X vssd1 vssd1 vccd1 vccd1 _1368_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_17_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0817__B1 _0716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0523_ _1155_/Q _1154_/Q vssd1 vssd1 vccd1 vccd1 _1041_/A sky130_fd_sc_hd__xnor2_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0501__B _0548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0874__D _0874_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1006_ _1323_/Q _1006_/B vssd1 vssd1 vccd1 vccd1 _1323_/D sky130_fd_sc_hd__xnor2_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0899__A _1276_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0506_ _1146_/A _1146_/B vssd1 vssd1 vccd1 vccd1 _0548_/C sky130_fd_sc_hd__xnor2_4
XFILLER_8_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0885__C _1284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0732__A2 _1187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1340_ _0862_/A _1340_/D _1140__64/Y vssd1 vssd1 vccd1 vccd1 _1340_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1167__RESET_B fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1313__D _1313_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1271_ _1104_/Y _1271_/D _1168_/CLK vssd1 vssd1 vccd1 vccd1 _1271_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0507__A _0548_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1063__44 _1065__45/A vssd1 vssd1 vccd1 vccd1 _1063__44/Y sky130_fd_sc_hd__inv_2
XANTENNA__1302__CLK _1035_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0986_ _1317_/Q _0986_/B vssd1 vssd1 vccd1 vccd1 _1317_/D sky130_fd_sc_hd__xnor2_1
XFILLER_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1073__A _1077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0896__B _1277_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf _1313_/Q _1020_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_11_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1260__RESET_B fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0771_ _1201_/Q _1200_/Q vssd1 vssd1 vccd1 vccd1 _0771_/Y sky130_fd_sc_hd__xnor2_4
X_0840_ _1013_/A _1233_/Q vssd1 vssd1 vccd1 vccd1 _1233_/D sky130_fd_sc_hd__xor2_1
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1323_ _1326_/CLK _1323_/D fanout46/X vssd1 vssd1 vccd1 vccd1 _1323_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1348__RESET_B fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1185_ _1359_/A _1185_/D fanout52/X vssd1 vssd1 vccd1 vccd1 _1185_/Q sky130_fd_sc_hd__dfrtp_4
X_1254_ input8/X input4/X fanout52/X vssd1 vssd1 vccd1 vccd1 _1255_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_21_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0969_ _1312_/Q _0969_/B vssd1 vssd1 vccd1 vccd1 _1312_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__1068__A _1077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0700__A _1175_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout45_A fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1106__48 _1117__53/A vssd1 vssd1 vccd1 vccd1 _1106__48/Y sky130_fd_sc_hd__inv_2
XFILLER_12_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0685_ _1331_/Q vssd1 vssd1 vccd1 vccd1 _1332_/D sky130_fd_sc_hd__inv_2
XFILLER_7_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0823_ _0822_/Y _0786_/C _1229_/Q vssd1 vssd1 vccd1 vccd1 _0824_/B sky130_fd_sc_hd__mux2_1
X_0754_ _1192_/Q _0754_/B vssd1 vssd1 vccd1 vccd1 _1192_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1306_ _1121_/Y _1306_/D _0460__17/Y vssd1 vssd1 vccd1 vccd1 _1306_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1099_ _1099_/A vssd1 vssd1 vccd1 vccd1 _1099_/Y sky130_fd_sc_hd__clkinv_2
X_1168_ _1168_/CLK _1168_/D fanout43/X vssd1 vssd1 vccd1 vccd1 _1168_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0893__C _1276_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1237_ _1082_/Y _1237_/D _0477_/Y vssd1 vssd1 vccd1 vccd1 _1237_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1099_/A fanout58/X vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_24_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0470_ _0479_/A vssd1 vssd1 vccd1 vccd1 _0470_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1022_ _1344_/Q _1343_/Q vssd1 vssd1 vccd1 vccd1 _1022_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_22_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0668_ _1300_/Q vssd1 vssd1 vccd1 vccd1 _1299_/D sky130_fd_sc_hd__inv_2
XFILLER_7_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0806_ _1224_/Q _0806_/B vssd1 vssd1 vccd1 vccd1 _0806_/Y sky130_fd_sc_hd__nand2_1
X_0737_ _1187_/Q _0737_/B vssd1 vssd1 vccd1 vccd1 _1187_/D sky130_fd_sc_hd__xnor2_1
X_0599_ _1178_/Q vssd1 vssd1 vccd1 vccd1 _1179_/D sky130_fd_sc_hd__inv_2
XANTENNA__1193__CLK fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1081__A _1097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0_w0.cclk_I _1034_/Y vssd1 vssd1 vccd1 vccd1 clkbuf_0_w0.cclk_I/X sky130_fd_sc_hd__clkbuf_16
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _1148_/CLK fanout42/X vssd1 vssd1 vccd1 vccd1 _1366_/A sky130_fd_sc_hd__dlrtn_1
X_0522_ _0868_/A vssd1 vssd1 vccd1 vccd1 _1045_/A sky130_fd_sc_hd__inv_6
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1005_ _1002_/Y _1004_/X _0831_/A vssd1 vssd1 vccd1 vccd1 _1006_/B sky130_fd_sc_hd__a21o_1
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
+ _1224_/Q _0843_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__1076__A _1077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_0__f_w0.cclk_I clkbuf_0_w0.cclk_I/X vssd1 vssd1 vccd1 vccd1 _1358_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput30 _1375_/X vssd1 vssd1 vccd1 vccd1 sin_out[1] sky130_fd_sc_hd__buf_2
XFILLER_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0505_ _1152_/Q vssd1 vssd1 vccd1 vccd1 _1146_/B sky130_fd_sc_hd__clkbuf_8
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

