magic
tech sky130A
timestamp 1654156409
use cap_10_10_x2  cap_10_10_x2_0
array 0 7 1098 0 3 1098
timestamp 1654156239
transform 1 0 61 0 1 48
box -57 -52 1041 1046
<< labels >>
flabel space 4 -4 8788 4388 0 FreeSans 4000 0 0 0 12.8pF
<< end >>
