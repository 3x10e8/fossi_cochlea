magic
tech sky130A
timestamp 1645590992
<< nwell >>
rect 7602 78 8019 162
rect 11733 100 12150 184
rect 1599 -44 2016 40
<< nmos >>
rect 7679 -4 7694 38
rect 7959 -4 7974 38
rect 11810 18 11825 60
rect 12090 18 12105 60
rect 1676 -126 1691 -84
rect 1956 -126 1971 -84
<< pmos >>
rect 7679 96 7694 138
rect 7959 96 7974 138
rect 11810 118 11825 160
rect 12090 118 12105 160
rect 1676 -26 1691 16
rect 1956 -26 1971 16
<< ndiff >>
rect 11781 48 11810 60
rect 7650 26 7679 38
rect 7650 9 7656 26
rect 7673 9 7679 26
rect 7650 -4 7679 9
rect 7694 26 7721 38
rect 7694 9 7700 26
rect 7717 9 7721 26
rect 7694 -4 7721 9
rect 7929 26 7959 38
rect 7929 9 7936 26
rect 7953 9 7959 26
rect 7929 -4 7959 9
rect 7974 26 8001 38
rect 7974 9 7980 26
rect 7997 9 8001 26
rect 11781 31 11787 48
rect 11804 31 11810 48
rect 11781 18 11810 31
rect 11825 48 11852 60
rect 11825 31 11831 48
rect 11848 31 11852 48
rect 11825 18 11852 31
rect 12060 48 12090 60
rect 12060 31 12067 48
rect 12084 31 12090 48
rect 12060 18 12090 31
rect 12105 48 12132 60
rect 12105 31 12111 48
rect 12128 31 12132 48
rect 12105 18 12132 31
rect 7974 -4 8001 9
rect 1646 -96 1676 -84
rect 1646 -113 1653 -96
rect 1670 -113 1676 -96
rect 1646 -126 1676 -113
rect 1691 -96 1718 -84
rect 1691 -113 1697 -96
rect 1714 -113 1718 -96
rect 1691 -126 1718 -113
rect 1926 -96 1956 -84
rect 1926 -113 1933 -96
rect 1950 -113 1956 -96
rect 1926 -126 1956 -113
rect 1971 -96 1998 -84
rect 1971 -113 1977 -96
rect 1994 -113 1998 -96
rect 1971 -126 1998 -113
<< pdiff >>
rect 11780 148 11810 160
rect 7649 126 7679 138
rect 7649 109 7656 126
rect 7673 109 7679 126
rect 7649 96 7679 109
rect 7694 126 7721 138
rect 7694 109 7700 126
rect 7717 109 7721 126
rect 7694 96 7721 109
rect 7929 126 7959 138
rect 7929 109 7936 126
rect 7953 109 7959 126
rect 7929 96 7959 109
rect 7974 126 8001 138
rect 7974 109 7980 126
rect 7997 109 8001 126
rect 11780 131 11787 148
rect 11804 131 11810 148
rect 11780 118 11810 131
rect 11825 148 11852 160
rect 11825 131 11831 148
rect 11848 131 11852 148
rect 11825 118 11852 131
rect 12060 148 12090 160
rect 12060 131 12067 148
rect 12084 131 12090 148
rect 12060 118 12090 131
rect 12105 148 12132 160
rect 12105 131 12111 148
rect 12128 131 12132 148
rect 12105 118 12132 131
rect 7974 96 8001 109
rect 1646 4 1676 16
rect 1646 -13 1653 4
rect 1670 -13 1676 4
rect 1646 -26 1676 -13
rect 1691 4 1718 16
rect 1691 -13 1697 4
rect 1714 -13 1718 4
rect 1691 -26 1718 -13
rect 1926 4 1956 16
rect 1926 -13 1933 4
rect 1950 -13 1956 4
rect 1926 -26 1956 -13
rect 1971 4 1998 16
rect 1971 -13 1977 4
rect 1994 -13 1998 4
rect 1971 -26 1998 -13
<< ndiffc >>
rect 7656 9 7673 26
rect 7700 9 7717 26
rect 7936 9 7953 26
rect 7980 9 7997 26
rect 11787 31 11804 48
rect 11831 31 11848 48
rect 12067 31 12084 48
rect 12111 31 12128 48
rect 1653 -113 1670 -96
rect 1697 -113 1714 -96
rect 1933 -113 1950 -96
rect 1977 -113 1994 -96
<< pdiffc >>
rect 7656 109 7673 126
rect 7700 109 7717 126
rect 7936 109 7953 126
rect 7980 109 7997 126
rect 11787 131 11804 148
rect 11831 131 11848 148
rect 12067 131 12084 148
rect 12111 131 12128 148
rect 1653 -13 1670 4
rect 1697 -13 1714 4
rect 1933 -13 1950 4
rect 1977 -13 1994 4
<< psubdiff >>
rect 5850 145 5986 211
rect 5850 55 5869 145
rect 5968 55 5986 145
rect 5850 7 5986 55
<< nsubdiff >>
rect 11751 147 11780 160
rect 7620 125 7649 138
rect 7620 108 7622 125
rect 7639 108 7649 125
rect 7620 96 7649 108
rect 11751 130 11753 147
rect 11770 130 11780 147
rect 11751 118 11780 130
<< psubdiffcont >>
rect 5869 55 5968 145
<< nsubdiffcont >>
rect 7622 108 7639 125
rect 11753 130 11770 147
<< poly >>
rect 11808 202 11835 210
rect 7677 180 7704 188
rect 7677 163 7682 180
rect 7699 163 7704 180
rect 7677 155 7704 163
rect 7957 180 7984 188
rect 7957 163 7962 180
rect 7979 163 7984 180
rect 11808 185 11813 202
rect 11830 185 11835 202
rect 11808 177 11835 185
rect 12088 202 12115 210
rect 12088 185 12093 202
rect 12110 185 12115 202
rect 12088 177 12115 185
rect 7957 155 7984 163
rect 11810 160 11825 177
rect 12090 160 12105 177
rect 1674 58 1701 66
rect 1674 41 1679 58
rect 1696 41 1701 58
rect 1674 33 1701 41
rect 1954 58 1981 66
rect 1954 41 1959 58
rect 1976 41 1981 58
rect 1954 33 1981 41
rect 7679 138 7694 155
rect 7959 138 7974 155
rect 11810 105 11825 118
rect 12090 105 12105 118
rect 7679 83 7694 96
rect 7959 83 7974 96
rect 11810 60 11825 73
rect 12090 60 12105 73
rect 1676 16 1691 33
rect 1956 16 1971 33
rect 7679 38 7694 51
rect 7959 38 7974 51
rect 11810 1 11825 18
rect 12090 1 12105 18
rect 7679 -21 7694 -4
rect 7959 -21 7974 -4
rect 11810 -7 11837 1
rect 1676 -39 1691 -26
rect 1956 -39 1971 -26
rect 7679 -29 7706 -21
rect 7679 -46 7684 -29
rect 7701 -46 7706 -29
rect 7679 -54 7706 -46
rect 7949 -29 7976 -21
rect 7949 -46 7954 -29
rect 7971 -46 7976 -29
rect 11810 -24 11815 -7
rect 11832 -24 11837 -7
rect 11810 -32 11837 -24
rect 12080 -7 12107 1
rect 12080 -24 12085 -7
rect 12102 -24 12107 -7
rect 12080 -32 12107 -24
rect 7949 -54 7976 -46
rect 1676 -84 1691 -71
rect 1956 -84 1971 -71
rect 1676 -143 1691 -126
rect 1956 -143 1971 -126
rect 1676 -151 1703 -143
rect 1676 -168 1681 -151
rect 1698 -168 1703 -151
rect 1676 -176 1703 -168
rect 1946 -151 1973 -143
rect 1946 -168 1951 -151
rect 1968 -168 1973 -151
rect 1946 -176 1973 -168
<< polycont >>
rect 7682 163 7699 180
rect 7962 163 7979 180
rect 11813 185 11830 202
rect 12093 185 12110 202
rect 1679 41 1696 58
rect 1959 41 1976 58
rect 7684 -46 7701 -29
rect 7954 -46 7971 -29
rect 11815 -24 11832 -7
rect 12085 -24 12102 -7
rect 1681 -168 1698 -151
rect 1951 -168 1968 -151
<< locali >>
rect 5850 146 5986 211
rect 11808 202 11835 210
rect 7677 180 7704 188
rect 7677 163 7682 180
rect 7699 163 7704 180
rect 7677 155 7704 163
rect 7957 180 7984 188
rect 7957 163 7962 180
rect 7979 163 7984 180
rect 11808 185 11813 202
rect 11830 185 11835 202
rect 11808 177 11835 185
rect 12088 202 12115 210
rect 12088 185 12093 202
rect 12110 185 12115 202
rect 12088 177 12115 185
rect 7957 155 7984 163
rect 1674 58 1701 66
rect 1674 41 1679 58
rect 1696 41 1701 58
rect 1674 33 1701 41
rect 1954 58 1981 66
rect 1954 41 1959 58
rect 1976 41 1981 58
rect 1954 33 1981 41
rect 5850 53 5867 146
rect 5969 53 5986 146
rect 11751 148 11808 160
rect 11751 147 11787 148
rect 7620 126 7677 138
rect 7620 125 7656 126
rect 7620 108 7622 125
rect 7639 109 7656 125
rect 7673 109 7677 126
rect 7639 108 7677 109
rect 7620 96 7677 108
rect 7696 126 7721 138
rect 7696 109 7700 126
rect 7717 109 7721 126
rect 7696 96 7721 109
rect 7929 126 7957 138
rect 7929 109 7936 126
rect 7953 109 7957 126
rect 7929 96 7957 109
rect 7976 126 8001 138
rect 7976 109 7980 126
rect 7997 109 8001 126
rect 11751 130 11753 147
rect 11770 131 11787 147
rect 11804 131 11808 148
rect 11770 130 11808 131
rect 11751 118 11808 130
rect 11827 148 11852 160
rect 11827 131 11831 148
rect 11848 131 11852 148
rect 11827 118 11852 131
rect 12060 148 12088 160
rect 12060 131 12067 148
rect 12084 131 12088 148
rect 12060 118 12088 131
rect 12107 148 12132 160
rect 12107 131 12111 148
rect 12128 131 12132 148
rect 12107 118 12132 131
rect 7976 96 8001 109
rect 1646 4 1674 16
rect 1646 -13 1653 4
rect 1670 -13 1674 4
rect 1646 -26 1674 -13
rect 1693 4 1718 16
rect 1693 -13 1697 4
rect 1714 -13 1718 4
rect 1693 -26 1718 -13
rect 1926 4 1954 16
rect 1926 -13 1933 4
rect 1950 -13 1954 4
rect 1926 -26 1954 -13
rect 1973 4 1998 16
rect 5850 7 5986 53
rect 7653 38 7670 96
rect 7703 72 7721 96
rect 7789 72 7847 79
rect 7933 72 7950 96
rect 7703 63 7950 72
rect 7703 55 7801 63
rect 7703 38 7721 55
rect 7650 26 7677 38
rect 7650 14 7656 26
rect 7630 9 7656 14
rect 7673 9 7677 26
rect 1973 -13 1977 4
rect 1994 -13 1998 4
rect 1973 -26 1998 -13
rect 7630 -4 7677 9
rect 7696 26 7721 38
rect 7696 9 7700 26
rect 7717 9 7721 26
rect 7789 31 7801 55
rect 7833 55 7950 63
rect 7833 31 7847 55
rect 7933 38 7950 55
rect 7983 61 8001 96
rect 7983 38 8611 61
rect 11784 60 11801 118
rect 11834 94 11852 118
rect 11920 94 11978 101
rect 12064 94 12081 118
rect 11834 85 12081 94
rect 11834 77 11932 85
rect 11834 60 11852 77
rect 7789 21 7847 31
rect 7929 26 7957 38
rect 7696 -4 7721 9
rect 7929 9 7936 26
rect 7953 9 7957 26
rect 7929 -4 7957 9
rect 7976 26 8001 38
rect 7976 9 7980 26
rect 7997 9 8001 26
rect 7976 -4 8001 9
rect 1650 -84 1667 -26
rect 1700 -50 1718 -26
rect 1786 -50 1844 -43
rect 1930 -50 1947 -26
rect 1700 -59 1947 -50
rect 1700 -67 1798 -59
rect 1700 -84 1718 -67
rect 1646 -96 1674 -84
rect 1646 -113 1653 -96
rect 1670 -113 1674 -96
rect 1646 -126 1674 -113
rect 1693 -96 1718 -84
rect 1693 -113 1697 -96
rect 1714 -113 1718 -96
rect 1786 -91 1798 -67
rect 1830 -67 1947 -59
rect 1830 -91 1844 -67
rect 1930 -84 1947 -67
rect 1980 -61 1998 -26
rect 3001 -61 3257 -16
rect 1980 -68 3257 -61
rect 1980 -84 3057 -68
rect 1786 -101 1844 -91
rect 1926 -96 1954 -84
rect 1693 -126 1718 -113
rect 1926 -113 1933 -96
rect 1950 -113 1954 -96
rect 1926 -126 1954 -113
rect 1973 -96 1998 -84
rect 1973 -113 1977 -96
rect 1994 -113 1998 -96
rect 1973 -126 1998 -113
rect 1676 -151 1703 -143
rect 1676 -168 1681 -151
rect 1698 -168 1703 -151
rect 1676 -176 1703 -168
rect 1946 -151 1973 -143
rect 1946 -168 1951 -151
rect 1968 -168 1973 -151
rect 1946 -176 1973 -168
rect 3001 -192 3057 -84
rect 3208 -108 3257 -68
rect 7630 -108 7662 -4
rect 7679 -29 7706 -21
rect 7679 -46 7684 -29
rect 7701 -46 7706 -29
rect 7679 -54 7706 -46
rect 7949 -29 7976 -21
rect 7949 -46 7954 -29
rect 7971 -46 7976 -29
rect 7949 -54 7976 -46
rect 8592 -78 8611 38
rect 11781 48 11808 60
rect 11781 37 11787 48
rect 11748 31 11787 37
rect 11804 31 11808 48
rect 11748 18 11808 31
rect 11827 48 11852 60
rect 11827 31 11831 48
rect 11848 31 11852 48
rect 11920 53 11932 77
rect 11964 77 12081 85
rect 11964 53 11978 77
rect 12064 60 12081 77
rect 12114 83 12132 118
rect 12250 91 12299 101
rect 12250 83 12260 91
rect 12114 61 12260 83
rect 12289 61 12299 91
rect 12114 60 12299 61
rect 11920 43 11978 53
rect 12060 48 12088 60
rect 11827 18 11852 31
rect 12060 31 12067 48
rect 12084 31 12088 48
rect 12060 18 12088 31
rect 12107 48 12132 60
rect 12250 54 12299 60
rect 12107 31 12111 48
rect 12128 31 12132 48
rect 12107 18 12132 31
rect 11748 14 11790 18
rect 8747 -78 9003 -33
rect 8592 -85 9003 -78
rect 8592 -101 8803 -85
rect 3208 -190 7662 -108
rect 3208 -192 3257 -190
rect 3001 -249 3257 -192
rect 8747 -209 8803 -101
rect 8954 -95 9003 -85
rect 11748 -95 11777 14
rect 11810 -7 11837 1
rect 11810 -24 11815 -7
rect 11832 -24 11837 -7
rect 11810 -32 11837 -24
rect 12080 -7 12107 1
rect 12080 -24 12085 -7
rect 12102 -24 12107 -7
rect 12080 -32 12107 -24
rect 8954 -133 11777 -95
rect 8954 -209 9003 -133
rect 11748 -134 11777 -133
rect 8747 -266 9003 -209
<< viali >>
rect 5867 145 5969 146
rect 5867 55 5869 145
rect 5869 55 5968 145
rect 5968 55 5969 145
rect 5867 53 5969 55
rect 7801 31 7833 63
rect 1798 -91 1830 -59
rect 3057 -192 3208 -68
rect 11932 53 11964 85
rect 12260 61 12289 91
rect 8803 -209 8954 -85
<< metal1 >>
rect 5849 146 5986 402
rect 5849 53 5867 146
rect 5969 53 5986 146
rect 11920 85 11978 101
rect 5849 7 5986 53
rect 7789 63 7847 79
rect 7789 31 7801 63
rect 7833 31 7847 63
rect 11920 53 11932 85
rect 11964 53 11978 85
rect 12250 91 12299 101
rect 12250 61 12260 91
rect 12289 61 12299 91
rect 12250 54 12299 61
rect 11920 43 11978 53
rect 7789 21 7847 31
rect 1786 -59 1844 -43
rect 1786 -91 1798 -59
rect 1830 -91 1844 -59
rect 1786 -101 1844 -91
rect 3000 -68 3256 -17
rect 3000 -192 3057 -68
rect 3208 -192 3256 -68
rect 3000 -251 3256 -192
rect 8746 -85 9002 -34
rect 8746 -209 8803 -85
rect 8954 -209 9002 -85
rect 8746 -268 9002 -209
<< via1 >>
rect 5867 53 5969 146
rect 7801 31 7833 63
rect 11932 53 11964 85
rect 12260 61 12289 91
rect 1798 -91 1830 -59
rect 3057 -192 3208 -68
rect 8803 -209 8954 -85
<< metal2 >>
rect 5849 146 5986 402
rect 5849 53 5867 146
rect 5969 53 5986 146
rect 11920 85 11978 101
rect 5849 7 5986 53
rect 7789 63 7847 79
rect 7789 31 7801 63
rect 7833 31 7847 63
rect 11920 53 11932 85
rect 11964 53 11978 85
rect 12250 91 12299 101
rect 12250 61 12260 91
rect 12289 61 12299 91
rect 12250 54 12299 61
rect 11920 43 11978 53
rect 7789 21 7847 31
rect 1786 -59 1844 -43
rect 1786 -91 1798 -59
rect 1830 -91 1844 -59
rect 1786 -101 1844 -91
rect 3000 -68 3256 -17
rect 3000 -192 3057 -68
rect 3208 -192 3256 -68
rect 3000 -251 3256 -192
rect 8746 -85 9002 -34
rect 8746 -209 8803 -85
rect 8954 -209 9002 -85
rect 8746 -268 9002 -209
<< via2 >>
rect 5867 53 5969 146
rect 7801 31 7833 63
rect 11932 53 11964 85
rect 12260 61 12289 91
rect 1798 -91 1830 -59
rect 3057 -192 3208 -68
rect 8803 -209 8954 -85
<< metal3 >>
rect -303 316 5811 6428
rect 563 -43 1291 260
rect 2883 -16 3384 316
rect 6038 276 10964 2704
rect 11255 292 14033 3070
rect 5849 146 5986 245
rect 5849 53 5867 146
rect 5969 53 5986 146
rect 5849 7 5986 53
rect 7158 79 7575 195
rect 7158 63 7847 79
rect 7158 40 7801 63
rect 7158 21 7620 40
rect 7650 31 7801 40
rect 7833 31 7847 63
rect 7650 21 7847 31
rect 563 -59 1844 -43
rect 563 -91 1798 -59
rect 1830 -91 1844 -59
rect 563 -101 1844 -91
rect 563 -468 1291 -101
rect 2883 -249 3001 -16
rect 3254 -249 3384 -16
rect 7158 -222 7575 21
rect 8629 -33 9130 276
rect 11402 101 11660 220
rect 11402 85 11978 101
rect 11402 63 11932 85
rect 11402 43 11744 63
rect 11781 53 11932 63
rect 11964 53 11978 85
rect 11781 43 11978 53
rect 12241 91 12305 292
rect 12241 61 12260 91
rect 12289 61 12305 91
rect 12241 46 12305 61
rect 11402 -28 11660 43
rect 2883 -381 3384 -249
rect 8629 -266 8747 -33
rect 9000 -266 9130 -33
rect 8629 -398 9130 -266
<< via3 >>
rect 5867 53 5969 146
rect 3001 -68 3254 -16
rect 3001 -192 3057 -68
rect 3057 -192 3208 -68
rect 3208 -192 3254 -68
rect 3001 -249 3254 -192
rect 8747 -85 9000 -33
rect 8747 -209 8803 -85
rect 8803 -209 8954 -85
rect 8954 -209 9000 -85
rect 8747 -266 9000 -209
<< mimcap >>
rect -289 6254 2711 6414
rect -289 6136 2071 6254
rect 2189 6136 2711 6254
rect -289 5941 2711 6136
rect -289 5823 -180 5941
rect -62 5823 2711 5941
rect -289 3983 2711 5823
rect -289 3865 -156 3983
rect -38 3865 2711 3983
rect -289 3414 2711 3865
rect 2795 6276 5797 6414
rect 2795 6158 3259 6276
rect 3377 6158 5797 6276
rect 2795 5930 5797 6158
rect 2795 5812 5538 5930
rect 5656 5812 5797 5930
rect 2795 3947 5797 5812
rect 2795 3829 5542 3947
rect 5660 3829 5797 3947
rect 2795 3414 5797 3829
rect -289 2886 2711 3330
rect -289 2768 -180 2886
rect -62 2768 2711 2886
rect -289 863 2711 2768
rect -289 745 -199 863
rect -81 745 2711 863
rect -289 530 2711 745
rect -289 412 2075 530
rect 2193 412 2711 530
rect -289 330 2711 412
rect 2795 2913 5797 3330
rect 2795 2795 5558 2913
rect 5676 2795 5797 2913
rect 2795 536 5797 2795
rect 2795 418 3249 536
rect 3367 418 5211 536
rect 5329 418 5797 536
rect 2795 330 5797 418
rect 6052 2609 8452 2690
rect 6052 2491 6368 2609
rect 6486 2584 8452 2609
rect 6486 2491 7939 2584
rect 6052 2466 7939 2491
rect 8057 2466 8452 2584
rect 6052 473 8452 2466
rect 6052 456 7959 473
rect 6052 338 6360 456
rect 6478 355 7959 456
rect 8077 355 8452 473
rect 6478 338 8452 355
rect 6052 290 8452 338
rect 8550 2565 10950 2690
rect 8550 2447 8929 2565
rect 9047 2548 10950 2565
rect 9047 2447 10489 2548
rect 8550 2430 10489 2447
rect 10607 2430 10950 2548
rect 8550 473 10950 2430
rect 8550 471 10483 473
rect 8550 353 8915 471
rect 9033 355 10483 471
rect 10601 355 10950 473
rect 9033 353 10950 355
rect 8550 290 10950 353
rect 11269 463 14019 3056
rect 11269 363 11470 463
rect 11570 363 14019 463
rect 11269 306 14019 363
rect 577 201 1277 246
rect 577 113 1137 201
rect 1229 113 1277 201
rect 577 -454 1277 113
rect 7172 145 7561 181
rect 7172 27 7398 145
rect 7516 27 7561 145
rect 7172 -208 7561 27
rect 11416 152 11646 206
rect 11416 52 11474 152
rect 11574 52 11646 152
rect 11416 -14 11646 52
<< mimcapcontact >>
rect 2071 6136 2189 6254
rect -180 5823 -62 5941
rect -156 3865 -38 3983
rect 3259 6158 3377 6276
rect 5538 5812 5656 5930
rect 5542 3829 5660 3947
rect -180 2768 -62 2886
rect -199 745 -81 863
rect 2075 412 2193 530
rect 5558 2795 5676 2913
rect 3249 418 3367 536
rect 5211 418 5329 536
rect 6368 2491 6486 2609
rect 7939 2466 8057 2584
rect 6360 338 6478 456
rect 7959 355 8077 473
rect 8929 2447 9047 2565
rect 10489 2430 10607 2548
rect 8915 353 9033 471
rect 10483 355 10601 473
rect 11470 363 11570 463
rect 1137 113 1229 201
rect 7398 27 7516 145
rect 11474 52 11574 152
<< metal4 >>
rect -303 6276 5811 6428
rect -303 6254 3259 6276
rect -303 6136 2071 6254
rect 2189 6158 3259 6254
rect 3377 6158 5811 6276
rect 2189 6136 5811 6158
rect -303 5941 5811 6136
rect -303 5823 -180 5941
rect -62 5930 5811 5941
rect -62 5823 5538 5930
rect -303 5812 5538 5823
rect 5656 5812 5811 5930
rect -303 3983 5811 5812
rect -303 3865 -156 3983
rect -38 3947 5811 3983
rect -38 3865 5542 3947
rect -303 3829 5542 3865
rect 5660 3829 5811 3947
rect -303 2913 5811 3829
rect -303 2886 5558 2913
rect -303 2768 -180 2886
rect -62 2795 5558 2886
rect 5676 2795 5811 2913
rect -62 2768 5811 2795
rect -303 2704 5811 2768
rect -303 2609 10964 2704
rect -303 2491 6368 2609
rect 6486 2584 10964 2609
rect 6486 2491 7939 2584
rect -303 2466 7939 2491
rect 8057 2565 10964 2584
rect 8057 2466 8929 2565
rect -303 2447 8929 2466
rect 9047 2548 10964 2565
rect 9047 2447 10489 2548
rect -303 2430 10489 2447
rect 10607 2430 10964 2548
rect -303 863 10964 2430
rect -303 745 -199 863
rect -81 745 10964 863
rect -303 536 10964 745
rect -303 530 3249 536
rect -303 412 2075 530
rect 2193 418 3249 530
rect 3367 418 5211 536
rect 5329 485 10964 536
rect 11459 485 11582 506
rect 5329 473 11582 485
rect 5329 456 7959 473
rect 5329 418 6360 456
rect 2193 412 6360 418
rect -303 338 6360 412
rect 6478 355 7959 456
rect 8077 471 10483 473
rect 8077 355 8915 471
rect 6478 353 8915 355
rect 9033 355 10483 471
rect 10601 463 11582 473
rect 10601 365 11470 463
rect 10601 355 10964 365
rect 9033 353 10964 355
rect 6478 338 10964 353
rect -303 316 10964 338
rect 1125 201 1245 316
rect 5848 245 5985 316
rect 6038 276 10964 316
rect 11459 363 11470 365
rect 11570 363 11582 463
rect 5848 226 5986 245
rect 1125 113 1137 201
rect 1229 113 1245 201
rect 1125 93 1245 113
rect 5849 146 5986 226
rect 5849 53 5867 146
rect 5969 53 5986 146
rect 2970 -16 3284 11
rect 5849 7 5986 53
rect 7385 145 7534 276
rect 7385 27 7398 145
rect 7516 27 7534 145
rect 11459 152 11582 363
rect 11459 52 11474 152
rect 11574 52 11582 152
rect 11459 30 11582 52
rect 7385 8 7534 27
rect 2970 -249 3001 -16
rect 3254 -249 3284 -16
rect 2970 -278 3284 -249
rect 8716 -33 9030 -6
rect 8716 -266 8747 -33
rect 9000 -266 9030 -33
rect 8716 -295 9030 -266
<< via4 >>
rect 3001 -249 3254 -16
rect 8747 -266 9000 -33
<< mimcap2 >>
rect -289 6272 2711 6414
rect -289 6154 -182 6272
rect -64 6262 2711 6272
rect -64 6154 2435 6262
rect -289 6144 2435 6154
rect 2553 6144 2711 6262
rect -289 3647 2711 6144
rect -289 3642 2440 3647
rect -289 3524 -164 3642
rect -46 3529 2440 3642
rect 2558 3529 2711 3647
rect -46 3524 2711 3529
rect -289 3414 2711 3524
rect 2795 6277 5797 6414
rect 2795 6159 2925 6277
rect 3043 6267 5797 6277
rect 3043 6159 5548 6267
rect 2795 6149 5548 6159
rect 5666 6149 5797 6267
rect 2795 3663 5797 6149
rect 2795 3545 2923 3663
rect 3041 3658 5797 3663
rect 3041 3545 5540 3658
rect 2795 3540 5540 3545
rect 5658 3540 5797 3658
rect 2795 3414 5797 3540
rect -289 3214 2711 3330
rect -289 3096 -174 3214
rect -56 3199 2711 3214
rect -56 3096 2453 3199
rect -289 3081 2453 3096
rect 2571 3081 2711 3199
rect -289 529 2711 3081
rect -289 516 2411 529
rect -289 398 -216 516
rect -98 411 2411 516
rect 2529 411 2711 529
rect -98 398 2711 411
rect -289 330 2711 398
rect 2795 3201 5797 3330
rect 2795 3196 5558 3201
rect 2795 3078 2917 3196
rect 3035 3083 5558 3196
rect 5676 3083 5797 3201
rect 3035 3078 5797 3083
rect 2795 553 5797 3078
rect 2795 532 5574 553
rect 2795 414 2915 532
rect 3033 435 5574 532
rect 5694 435 5797 553
rect 3033 414 5797 435
rect 2795 330 5797 414
rect 6052 2612 8452 2690
rect 6052 2494 6101 2612
rect 6219 2576 8452 2612
rect 6219 2494 8182 2576
rect 6052 2458 8182 2494
rect 8300 2458 8452 2576
rect 6052 472 8452 2458
rect 6052 455 8181 472
rect 6052 337 6102 455
rect 6220 354 8181 455
rect 8299 354 8452 472
rect 6220 337 8452 354
rect 6052 290 8452 337
rect 8550 2562 10950 2690
rect 8550 2444 8657 2562
rect 8775 2548 10950 2562
rect 8775 2444 10731 2548
rect 8550 2430 10731 2444
rect 10849 2430 10950 2548
rect 8550 475 10950 2430
rect 8550 464 10704 475
rect 8550 346 8650 464
rect 8768 357 10704 464
rect 10822 357 10950 475
rect 8768 346 10950 357
rect 8550 290 10950 346
<< mimcap2contact >>
rect -182 6154 -64 6272
rect 2435 6144 2553 6262
rect -164 3524 -46 3642
rect 2440 3529 2558 3647
rect 2925 6159 3043 6277
rect 5548 6149 5666 6267
rect 2923 3545 3041 3663
rect 5540 3540 5658 3658
rect -174 3096 -56 3214
rect 2453 3081 2571 3199
rect -216 398 -98 516
rect 2411 411 2529 529
rect 2917 3078 3035 3196
rect 5558 3083 5676 3201
rect 2915 414 3033 532
rect 5574 435 5694 553
rect 6101 2494 6219 2612
rect 8182 2458 8300 2576
rect 6102 337 6220 455
rect 8181 354 8299 472
rect 8657 2444 8775 2562
rect 10731 2430 10849 2548
rect 8650 346 8768 464
rect 10704 357 10822 475
<< metal5 >>
rect -226 6314 5746 6316
rect -238 6277 5746 6314
rect -238 6272 2925 6277
rect -238 6154 -182 6272
rect -64 6262 2925 6272
rect -64 6154 2435 6262
rect -238 6144 2435 6154
rect 2553 6159 2925 6262
rect 3043 6267 5746 6277
rect 3043 6159 5548 6267
rect 2553 6149 5548 6159
rect 5666 6149 5746 6267
rect 2553 6144 5746 6149
rect -238 6116 5746 6144
rect -238 3719 -14 6116
rect 5518 3719 5746 6116
rect -243 3663 5748 3719
rect -243 3647 2923 3663
rect -243 3642 2440 3647
rect -243 3524 -164 3642
rect -46 3529 2440 3642
rect 2558 3545 2923 3647
rect 3041 3658 5748 3663
rect 3041 3545 5540 3658
rect 2558 3540 5540 3545
rect 5658 3540 5748 3658
rect 2558 3529 5748 3540
rect -46 3524 5748 3529
rect -243 3470 5748 3524
rect -238 3244 -14 3470
rect 5518 3244 5746 3470
rect -240 3214 5751 3244
rect -240 3096 -174 3214
rect -56 3201 5751 3214
rect -56 3199 5558 3201
rect -56 3096 2453 3199
rect -240 3081 2453 3096
rect 2571 3196 5558 3199
rect 2571 3081 2917 3196
rect -240 3078 2917 3081
rect 3035 3083 5558 3196
rect 5676 3083 5751 3201
rect 3035 3078 5751 3083
rect -240 2995 5751 3078
rect -238 603 -14 2995
rect 5518 603 5746 2995
rect -238 553 5746 603
rect -238 532 5574 553
rect -238 529 2915 532
rect -238 516 2411 529
rect -238 398 -216 516
rect -98 411 2411 516
rect 2529 414 2915 529
rect 3033 435 5574 532
rect 5694 435 5746 553
rect 3033 414 5746 435
rect 2529 411 5746 414
rect -98 398 5746 411
rect -238 366 5746 398
rect 2883 -16 3384 366
rect 5518 357 5746 366
rect 6079 2612 6244 2646
rect 6079 2494 6101 2612
rect 6219 2611 6244 2612
rect 10664 2611 10883 2662
rect 6219 2576 10891 2611
rect 6219 2494 8182 2576
rect 6079 2458 8182 2494
rect 8300 2562 10891 2576
rect 8300 2458 8657 2562
rect 6079 2444 8657 2458
rect 8775 2548 10891 2562
rect 8775 2444 10731 2548
rect 6079 2430 10731 2444
rect 10849 2430 10891 2548
rect 6079 2417 10891 2430
rect 6079 524 6244 2417
rect 10664 524 10883 2417
rect 6079 475 10883 524
rect 6079 472 10704 475
rect 6079 455 8181 472
rect 6079 337 6102 455
rect 6220 354 8181 455
rect 8299 464 10704 472
rect 8299 354 8650 464
rect 6220 346 8650 354
rect 8768 357 10704 464
rect 10822 357 10883 475
rect 8768 346 10883 357
rect 6220 337 10883 346
rect 6079 317 10883 337
rect 2883 -249 3001 -16
rect 3254 -249 3384 -16
rect 2883 -381 3384 -249
rect 8629 -33 9130 317
rect 8629 -266 8747 -33
rect 9000 -266 9130 -33
rect 8629 -398 9130 -266
<< labels >>
rlabel metal4 1245 279 1245 279 3 gnd
rlabel locali 1650 -62 1650 -62 7 in
rlabel locali 1690 -176 1690 -176 5 phi1
rlabel locali 1689 66 1689 66 1 phi1b
rlabel locali 1969 66 1969 66 1 phi2b
rlabel locali 1959 -176 1959 -176 1 phi2
rlabel metal3 1375 -101 1375 -101 5 cs1top
rlabel locali 7693 -54 7693 -54 5 phi1
rlabel locali 7692 188 7692 188 1 phi1b
rlabel locali 7972 188 7972 188 1 phi2b
rlabel locali 7962 -54 7962 -54 1 phi2
rlabel locali 11824 -32 11824 -32 5 phi1
rlabel locali 11823 210 11823 210 1 phi1b
rlabel locali 12103 210 12103 210 1 phi2b
rlabel locali 12093 -32 12093 -32 1 phi2
rlabel metal3 12288 292 12288 292 5 out3
rlabel locali 2123 -84 2123 -84 5 out1
rlabel metal3 7592 21 7592 21 5 mimsmall2
rlabel metal3 11688 43 11688 43 5 mimsmall3
rlabel locali 9657 -133 9657 -133 5 out2
<< end >>
