magic
tech sky130A
timestamp 1654307754
use cap_10_10_center_x2  cap_10_10_center_x2_0
array 0 0 -1052 0 5 1742
timestamp 1654307754
transform 0 1 374 -1 0 1018
box -34 -374 1018 1368
use cap_10_10_side2_x2  cap_10_10_side2_x2_0
timestamp 1654307754
transform 0 -1 -374 1 0 34
box -34 -374 1018 1023
use cap_10_10_side2_x2  cap_10_10_side2_x2_1
timestamp 1654307754
transform 0 1 10826 -1 0 1018
box -34 -374 1018 1023
<< end >>
