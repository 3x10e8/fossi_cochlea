magic
tech sky130A
timestamp 1654156743
use cap_10_10_x2  cap_10_10_x2_0
array 0 7 1098 0 0 1098
timestamp 1654156239
transform 1 0 50 0 1 54
box -57 -52 1041 1046
<< labels >>
flabel space -7 2 8777 1100 0 FreeSans 4000 0 0 0 3.2pF
<< end >>
