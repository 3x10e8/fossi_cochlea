magic
tech sky130A
magscale 1 2
timestamp 1654737118
<< obsli1 >>
rect 1104 2159 78844 57681
<< obsm1 >>
rect 1104 2128 79382 59288
<< metal2 >>
rect 2226 59200 2282 60000
rect 6642 59200 6698 60000
rect 11058 59200 11114 60000
rect 15566 59200 15622 60000
rect 19982 59200 20038 60000
rect 24398 59200 24454 60000
rect 28906 59200 28962 60000
rect 33322 59200 33378 60000
rect 37738 59200 37794 60000
rect 42246 59200 42302 60000
rect 46662 59200 46718 60000
rect 51078 59200 51134 60000
rect 55586 59200 55642 60000
rect 60002 59200 60058 60000
rect 64418 59200 64474 60000
rect 68926 59200 68982 60000
rect 73342 59200 73398 60000
rect 77758 59200 77814 60000
rect 4434 0 4490 800
rect 13266 0 13322 800
rect 22190 0 22246 800
rect 31114 0 31170 800
rect 39946 0 40002 800
rect 48870 0 48926 800
rect 57794 0 57850 800
rect 66626 0 66682 800
rect 75550 0 75606 800
<< obsm2 >>
rect 1398 59144 2170 59809
rect 2338 59144 6586 59809
rect 6754 59144 11002 59809
rect 11170 59144 15510 59809
rect 15678 59144 19926 59809
rect 20094 59144 24342 59809
rect 24510 59144 28850 59809
rect 29018 59144 33266 59809
rect 33434 59144 37682 59809
rect 37850 59144 42190 59809
rect 42358 59144 46606 59809
rect 46774 59144 51022 59809
rect 51190 59144 55530 59809
rect 55698 59144 59946 59809
rect 60114 59144 64362 59809
rect 64530 59144 68870 59809
rect 69038 59144 73286 59809
rect 73454 59144 77702 59809
rect 77870 59144 79376 59809
rect 1398 856 79376 59144
rect 1398 800 4378 856
rect 4546 800 13210 856
rect 13378 800 22134 856
rect 22302 800 31058 856
rect 31226 800 39890 856
rect 40058 800 48814 856
rect 48982 800 57738 856
rect 57906 800 66570 856
rect 66738 800 75494 856
rect 75662 800 79376 856
<< metal3 >>
rect 0 57944 800 58064
rect 79200 58080 80000 58200
rect 79200 54544 80000 54664
rect 0 54136 800 54256
rect 79200 51008 80000 51128
rect 0 50464 800 50584
rect 79200 47472 80000 47592
rect 0 46656 800 46776
rect 79200 43936 80000 44056
rect 0 42984 800 43104
rect 79200 40400 80000 40520
rect 0 39176 800 39296
rect 79200 36864 80000 36984
rect 0 35504 800 35624
rect 79200 33328 80000 33448
rect 0 31696 800 31816
rect 79200 29792 80000 29912
rect 0 27888 800 28008
rect 79200 26256 80000 26376
rect 0 24216 800 24336
rect 79200 22720 80000 22840
rect 0 20408 800 20528
rect 79200 19184 80000 19304
rect 0 16736 800 16856
rect 79200 15648 80000 15768
rect 0 12928 800 13048
rect 79200 12112 80000 12232
rect 0 9256 800 9376
rect 79200 8576 80000 8696
rect 0 5448 800 5568
rect 79200 5040 80000 5160
rect 0 1776 800 1896
rect 79200 1640 80000 1760
<< obsm3 >>
rect 800 58280 79200 59940
rect 800 58144 79120 58280
rect 880 58000 79120 58144
rect 880 57864 79200 58000
rect 800 54744 79200 57864
rect 800 54464 79120 54744
rect 800 54336 79200 54464
rect 880 54056 79200 54336
rect 800 51208 79200 54056
rect 800 50928 79120 51208
rect 800 50664 79200 50928
rect 880 50384 79200 50664
rect 800 47672 79200 50384
rect 800 47392 79120 47672
rect 800 46856 79200 47392
rect 880 46576 79200 46856
rect 800 44136 79200 46576
rect 800 43856 79120 44136
rect 800 43184 79200 43856
rect 880 42904 79200 43184
rect 800 40600 79200 42904
rect 800 40320 79120 40600
rect 800 39376 79200 40320
rect 880 39096 79200 39376
rect 800 37064 79200 39096
rect 800 36784 79120 37064
rect 800 35704 79200 36784
rect 880 35424 79200 35704
rect 800 33528 79200 35424
rect 800 33248 79120 33528
rect 800 31896 79200 33248
rect 880 31616 79200 31896
rect 800 29992 79200 31616
rect 800 29712 79120 29992
rect 800 28088 79200 29712
rect 880 27808 79200 28088
rect 800 26456 79200 27808
rect 800 26176 79120 26456
rect 800 24416 79200 26176
rect 880 24136 79200 24416
rect 800 22920 79200 24136
rect 800 22640 79120 22920
rect 800 20608 79200 22640
rect 880 20328 79200 20608
rect 800 19384 79200 20328
rect 800 19104 79120 19384
rect 800 16936 79200 19104
rect 880 16656 79200 16936
rect 800 15848 79200 16656
rect 800 15568 79120 15848
rect 800 13128 79200 15568
rect 880 12848 79200 13128
rect 800 12312 79200 12848
rect 800 12032 79120 12312
rect 800 9456 79200 12032
rect 880 9176 79200 9456
rect 800 8776 79200 9176
rect 800 8496 79120 8776
rect 800 5648 79200 8496
rect 880 5368 79200 5648
rect 800 5240 79200 5368
rect 800 4960 79120 5240
rect 800 1976 79200 4960
rect 880 1840 79200 1976
rect 880 1696 79120 1840
rect 800 1667 79120 1696
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
rect 65648 2128 65968 57712
<< obsm4 >>
rect 8155 57792 76485 59941
rect 8155 2048 19488 57792
rect 19968 2048 34848 57792
rect 35328 2048 50208 57792
rect 50688 2048 65568 57792
rect 66048 2048 76485 57792
rect 8155 1939 76485 2048
<< labels >>
rlabel metal3 s 0 20408 800 20528 6 cclk_I[0]
port 1 nsew signal output
rlabel metal3 s 0 46656 800 46776 6 cclk_I[1]
port 2 nsew signal output
rlabel metal3 s 79200 5040 80000 5160 6 cclk_Q[0]
port 3 nsew signal output
rlabel metal3 s 79200 29792 80000 29912 6 cclk_Q[1]
port 4 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 clk_master
port 5 nsew signal input
rlabel metal2 s 6642 59200 6698 60000 6 clk_master_out
port 6 nsew signal output
rlabel metal3 s 0 16736 800 16856 6 clkdiv2_I[0]
port 7 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 clkdiv2_I[1]
port 8 nsew signal output
rlabel metal3 s 79200 8576 80000 8696 6 clkdiv2_Q[0]
port 9 nsew signal output
rlabel metal3 s 79200 33328 80000 33448 6 clkdiv2_Q[1]
port 10 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 comp_high_I[0]
port 11 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 comp_high_I[1]
port 12 nsew signal input
rlabel metal3 s 79200 12112 80000 12232 6 comp_high_Q[0]
port 13 nsew signal input
rlabel metal3 s 79200 36864 80000 36984 6 comp_high_Q[1]
port 14 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 cos_out[0]
port 15 nsew signal output
rlabel metal3 s 0 50464 800 50584 6 cos_out[1]
port 16 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 cos_outb[0]
port 17 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 cos_outb[1]
port 18 nsew signal output
rlabel metal2 s 15566 59200 15622 60000 6 div2out
port 19 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 fb1_I[0]
port 20 nsew signal output
rlabel metal3 s 0 31696 800 31816 6 fb1_I[1]
port 21 nsew signal output
rlabel metal3 s 79200 19184 80000 19304 6 fb1_Q[0]
port 22 nsew signal output
rlabel metal3 s 79200 43936 80000 44056 6 fb1_Q[1]
port 23 nsew signal output
rlabel metal3 s 79200 58080 80000 58200 6 fb2_I[0]
port 24 nsew signal output
rlabel metal2 s 66626 0 66682 800 6 fb2_I[1]
port 25 nsew signal output
rlabel metal2 s 77758 59200 77814 60000 6 fb2_Q[0]
port 26 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 fb2_Q[1]
port 27 nsew signal output
rlabel metal2 s 60002 59200 60058 60000 6 gray_clk_out[10]
port 28 nsew signal output
rlabel metal2 s 19982 59200 20038 60000 6 gray_clk_out[1]
port 29 nsew signal output
rlabel metal2 s 24398 59200 24454 60000 6 gray_clk_out[2]
port 30 nsew signal output
rlabel metal2 s 28906 59200 28962 60000 6 gray_clk_out[3]
port 31 nsew signal output
rlabel metal2 s 33322 59200 33378 60000 6 gray_clk_out[4]
port 32 nsew signal output
rlabel metal2 s 37738 59200 37794 60000 6 gray_clk_out[5]
port 33 nsew signal output
rlabel metal2 s 42246 59200 42302 60000 6 gray_clk_out[6]
port 34 nsew signal output
rlabel metal2 s 46662 59200 46718 60000 6 gray_clk_out[7]
port 35 nsew signal output
rlabel metal2 s 51078 59200 51134 60000 6 gray_clk_out[8]
port 36 nsew signal output
rlabel metal2 s 55586 59200 55642 60000 6 gray_clk_out[9]
port 37 nsew signal output
rlabel metal2 s 64418 59200 64474 60000 6 no_ones_below_out[0]
port 38 nsew signal output
rlabel metal2 s 68926 59200 68982 60000 6 no_ones_below_out[1]
port 39 nsew signal output
rlabel metal2 s 73342 59200 73398 60000 6 no_ones_below_out[2]
port 40 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 phi1b_dig_I[0]
port 41 nsew signal input
rlabel metal3 s 0 35504 800 35624 6 phi1b_dig_I[1]
port 42 nsew signal input
rlabel metal3 s 79200 15648 80000 15768 6 phi1b_dig_Q[0]
port 43 nsew signal input
rlabel metal3 s 79200 40400 80000 40520 6 phi1b_dig_Q[1]
port 44 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 read_out_I[0]
port 45 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 read_out_I[1]
port 46 nsew signal output
rlabel metal3 s 0 54136 800 54256 6 read_out_I_top[0]
port 47 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 read_out_I_top[1]
port 48 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 read_out_Q[0]
port 49 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 read_out_Q[1]
port 50 nsew signal output
rlabel metal3 s 79200 51008 80000 51128 6 read_out_Q_top[0]
port 51 nsew signal output
rlabel metal3 s 79200 54544 80000 54664 6 read_out_Q_top[1]
port 52 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 rstb
port 53 nsew signal input
rlabel metal2 s 2226 59200 2282 60000 6 rstb_out
port 54 nsew signal output
rlabel metal3 s 79200 1640 80000 1760 6 sin_out[0]
port 55 nsew signal output
rlabel metal3 s 79200 26256 80000 26376 6 sin_out[1]
port 56 nsew signal output
rlabel metal3 s 79200 22720 80000 22840 6 sin_outb[0]
port 57 nsew signal output
rlabel metal3 s 79200 47472 80000 47592 6 sin_outb[1]
port 58 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 ud_en
port 59 nsew signal input
rlabel metal2 s 11058 59200 11114 60000 6 ud_en_out
port 60 nsew signal output
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 61 nsew power input
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 61 nsew power input
rlabel metal4 s 65648 2128 65968 57712 6 vccd1
port 61 nsew power input
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 62 nsew ground input
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 62 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 80000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7786664
string GDS_FILE /Volumes/export/isn/abhinav/fossi_cochlea/openlane/first_dual_core/runs/first_dual_core/results/finishing/first_dual_core.magic.gds
string GDS_START 424876
<< end >>

