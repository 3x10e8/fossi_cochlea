VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO first_dual_core
  CLASS BLOCK ;
  FOREIGN first_dual_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 300.000 ;
  PIN cclk_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END cclk_I[0]
  PIN cclk_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END cclk_I[1]
  PIN cclk_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 25.200 400.000 25.800 ;
    END
  END cclk_Q[0]
  PIN cclk_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 148.960 400.000 149.560 ;
    END
  END cclk_Q[1]
  PIN clk_master
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END clk_master
  PIN clk_master_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 296.000 33.490 300.000 ;
    END
  END clk_master_out
  PIN clkdiv2_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END clkdiv2_I[0]
  PIN clkdiv2_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END clkdiv2_I[1]
  PIN clkdiv2_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 42.880 400.000 43.480 ;
    END
  END clkdiv2_Q[0]
  PIN clkdiv2_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 166.640 400.000 167.240 ;
    END
  END clkdiv2_Q[1]
  PIN comp_high_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END comp_high_I[0]
  PIN comp_high_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END comp_high_I[1]
  PIN comp_high_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 60.560 400.000 61.160 ;
    END
  END comp_high_Q[0]
  PIN comp_high_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 184.320 400.000 184.920 ;
    END
  END comp_high_Q[1]
  PIN cos_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END cos_out[0]
  PIN cos_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.320 4.000 252.920 ;
    END
  END cos_out[1]
  PIN cos_outb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END cos_outb[0]
  PIN cos_outb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END cos_outb[1]
  PIN div2out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 296.000 78.110 300.000 ;
    END
  END div2out
  PIN fb1_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END fb1_I[0]
  PIN fb1_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END fb1_I[1]
  PIN fb1_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 95.920 400.000 96.520 ;
    END
  END fb1_Q[0]
  PIN fb1_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 219.680 400.000 220.280 ;
    END
  END fb1_Q[1]
  PIN fb2_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 290.400 400.000 291.000 ;
    END
  END fb2_I[0]
  PIN fb2_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END fb2_I[1]
  PIN fb2_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 296.000 389.070 300.000 ;
    END
  END fb2_Q[0]
  PIN fb2_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END fb2_Q[1]
  PIN gray_clk_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 296.000 300.290 300.000 ;
    END
  END gray_clk_out[10]
  PIN gray_clk_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 296.000 100.190 300.000 ;
    END
  END gray_clk_out[1]
  PIN gray_clk_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 296.000 122.270 300.000 ;
    END
  END gray_clk_out[2]
  PIN gray_clk_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 296.000 144.810 300.000 ;
    END
  END gray_clk_out[3]
  PIN gray_clk_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 296.000 166.890 300.000 ;
    END
  END gray_clk_out[4]
  PIN gray_clk_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 296.000 188.970 300.000 ;
    END
  END gray_clk_out[5]
  PIN gray_clk_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 296.000 211.510 300.000 ;
    END
  END gray_clk_out[6]
  PIN gray_clk_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 296.000 233.590 300.000 ;
    END
  END gray_clk_out[7]
  PIN gray_clk_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 296.000 255.670 300.000 ;
    END
  END gray_clk_out[8]
  PIN gray_clk_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 296.000 278.210 300.000 ;
    END
  END gray_clk_out[9]
  PIN no_ones_below_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 296.000 322.370 300.000 ;
    END
  END no_ones_below_out[0]
  PIN no_ones_below_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 296.000 344.910 300.000 ;
    END
  END no_ones_below_out[1]
  PIN no_ones_below_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 296.000 366.990 300.000 ;
    END
  END no_ones_below_out[2]
  PIN phi1b_dig_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END phi1b_dig_I[0]
  PIN phi1b_dig_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.520 4.000 178.120 ;
    END
  END phi1b_dig_I[1]
  PIN phi1b_dig_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 78.240 400.000 78.840 ;
    END
  END phi1b_dig_Q[0]
  PIN phi1b_dig_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 202.000 400.000 202.600 ;
    END
  END phi1b_dig_Q[1]
  PIN read_out_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END read_out_I[0]
  PIN read_out_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END read_out_I[1]
  PIN read_out_I_top[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END read_out_I_top[0]
  PIN read_out_I_top[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END read_out_I_top[1]
  PIN read_out_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END read_out_Q[0]
  PIN read_out_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END read_out_Q[1]
  PIN read_out_Q_top[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 255.040 400.000 255.640 ;
    END
  END read_out_Q_top[0]
  PIN read_out_Q_top[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 272.720 400.000 273.320 ;
    END
  END read_out_Q_top[1]
  PIN rstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END rstb
  PIN rstb_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 296.000 11.410 300.000 ;
    END
  END rstb_out
  PIN sin_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 8.200 400.000 8.800 ;
    END
  END sin_out[0]
  PIN sin_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 131.280 400.000 131.880 ;
    END
  END sin_out[1]
  PIN sin_outb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 113.600 400.000 114.200 ;
    END
  END sin_outb[0]
  PIN sin_outb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 237.360 400.000 237.960 ;
    END
  END sin_outb[1]
  PIN ud_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END ud_en
  PIN ud_en_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 296.000 55.570 300.000 ;
    END
  END ud_en_out
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 394.220 288.405 ;
      LAYER met1 ;
        RECT 5.520 10.640 396.910 296.440 ;
      LAYER met2 ;
        RECT 6.990 295.720 10.850 299.045 ;
        RECT 11.690 295.720 32.930 299.045 ;
        RECT 33.770 295.720 55.010 299.045 ;
        RECT 55.850 295.720 77.550 299.045 ;
        RECT 78.390 295.720 99.630 299.045 ;
        RECT 100.470 295.720 121.710 299.045 ;
        RECT 122.550 295.720 144.250 299.045 ;
        RECT 145.090 295.720 166.330 299.045 ;
        RECT 167.170 295.720 188.410 299.045 ;
        RECT 189.250 295.720 210.950 299.045 ;
        RECT 211.790 295.720 233.030 299.045 ;
        RECT 233.870 295.720 255.110 299.045 ;
        RECT 255.950 295.720 277.650 299.045 ;
        RECT 278.490 295.720 299.730 299.045 ;
        RECT 300.570 295.720 321.810 299.045 ;
        RECT 322.650 295.720 344.350 299.045 ;
        RECT 345.190 295.720 366.430 299.045 ;
        RECT 367.270 295.720 388.510 299.045 ;
        RECT 389.350 295.720 396.880 299.045 ;
        RECT 6.990 4.280 396.880 295.720 ;
        RECT 6.990 4.000 21.890 4.280 ;
        RECT 22.730 4.000 66.050 4.280 ;
        RECT 66.890 4.000 110.670 4.280 ;
        RECT 111.510 4.000 155.290 4.280 ;
        RECT 156.130 4.000 199.450 4.280 ;
        RECT 200.290 4.000 244.070 4.280 ;
        RECT 244.910 4.000 288.690 4.280 ;
        RECT 289.530 4.000 332.850 4.280 ;
        RECT 333.690 4.000 377.470 4.280 ;
        RECT 378.310 4.000 396.880 4.280 ;
      LAYER met3 ;
        RECT 4.000 291.400 396.000 299.700 ;
        RECT 4.000 290.720 395.600 291.400 ;
        RECT 4.400 290.000 395.600 290.720 ;
        RECT 4.400 289.320 396.000 290.000 ;
        RECT 4.000 273.720 396.000 289.320 ;
        RECT 4.000 272.320 395.600 273.720 ;
        RECT 4.000 271.680 396.000 272.320 ;
        RECT 4.400 270.280 396.000 271.680 ;
        RECT 4.000 256.040 396.000 270.280 ;
        RECT 4.000 254.640 395.600 256.040 ;
        RECT 4.000 253.320 396.000 254.640 ;
        RECT 4.400 251.920 396.000 253.320 ;
        RECT 4.000 238.360 396.000 251.920 ;
        RECT 4.000 236.960 395.600 238.360 ;
        RECT 4.000 234.280 396.000 236.960 ;
        RECT 4.400 232.880 396.000 234.280 ;
        RECT 4.000 220.680 396.000 232.880 ;
        RECT 4.000 219.280 395.600 220.680 ;
        RECT 4.000 215.920 396.000 219.280 ;
        RECT 4.400 214.520 396.000 215.920 ;
        RECT 4.000 203.000 396.000 214.520 ;
        RECT 4.000 201.600 395.600 203.000 ;
        RECT 4.000 196.880 396.000 201.600 ;
        RECT 4.400 195.480 396.000 196.880 ;
        RECT 4.000 185.320 396.000 195.480 ;
        RECT 4.000 183.920 395.600 185.320 ;
        RECT 4.000 178.520 396.000 183.920 ;
        RECT 4.400 177.120 396.000 178.520 ;
        RECT 4.000 167.640 396.000 177.120 ;
        RECT 4.000 166.240 395.600 167.640 ;
        RECT 4.000 159.480 396.000 166.240 ;
        RECT 4.400 158.080 396.000 159.480 ;
        RECT 4.000 149.960 396.000 158.080 ;
        RECT 4.000 148.560 395.600 149.960 ;
        RECT 4.000 140.440 396.000 148.560 ;
        RECT 4.400 139.040 396.000 140.440 ;
        RECT 4.000 132.280 396.000 139.040 ;
        RECT 4.000 130.880 395.600 132.280 ;
        RECT 4.000 122.080 396.000 130.880 ;
        RECT 4.400 120.680 396.000 122.080 ;
        RECT 4.000 114.600 396.000 120.680 ;
        RECT 4.000 113.200 395.600 114.600 ;
        RECT 4.000 103.040 396.000 113.200 ;
        RECT 4.400 101.640 396.000 103.040 ;
        RECT 4.000 96.920 396.000 101.640 ;
        RECT 4.000 95.520 395.600 96.920 ;
        RECT 4.000 84.680 396.000 95.520 ;
        RECT 4.400 83.280 396.000 84.680 ;
        RECT 4.000 79.240 396.000 83.280 ;
        RECT 4.000 77.840 395.600 79.240 ;
        RECT 4.000 65.640 396.000 77.840 ;
        RECT 4.400 64.240 396.000 65.640 ;
        RECT 4.000 61.560 396.000 64.240 ;
        RECT 4.000 60.160 395.600 61.560 ;
        RECT 4.000 47.280 396.000 60.160 ;
        RECT 4.400 45.880 396.000 47.280 ;
        RECT 4.000 43.880 396.000 45.880 ;
        RECT 4.000 42.480 395.600 43.880 ;
        RECT 4.000 28.240 396.000 42.480 ;
        RECT 4.400 26.840 396.000 28.240 ;
        RECT 4.000 26.200 396.000 26.840 ;
        RECT 4.000 24.800 395.600 26.200 ;
        RECT 4.000 9.880 396.000 24.800 ;
        RECT 4.400 9.200 396.000 9.880 ;
        RECT 4.400 8.480 395.600 9.200 ;
        RECT 4.000 8.335 395.600 8.480 ;
      LAYER met4 ;
        RECT 40.775 288.960 382.425 299.705 ;
        RECT 40.775 10.240 97.440 288.960 ;
        RECT 99.840 10.240 174.240 288.960 ;
        RECT 176.640 10.240 251.040 288.960 ;
        RECT 253.440 10.240 327.840 288.960 ;
        RECT 330.240 10.240 382.425 288.960 ;
        RECT 40.775 9.695 382.425 10.240 ;
  END
END first_dual_core
END LIBRARY

