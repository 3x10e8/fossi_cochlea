magic
tech sky130B
magscale 1 2
timestamp 1663962710
<< metal1 >>
rect 406166 23488 406172 23588
rect 406272 23488 407704 23588
rect 406466 19488 406472 19588
rect 406572 19488 407704 19588
rect 406766 15488 406772 15588
rect 406872 15488 407704 15588
rect 407066 11488 407072 11588
rect 407172 11488 407704 11588
rect 407366 7488 407372 7588
rect 407472 7488 407704 7588
rect 406462 3595 406575 3601
rect 406462 3494 406468 3595
rect 406569 3494 407704 3595
rect 406462 3488 406575 3494
rect 406162 -384 406274 -378
rect 406162 -484 406168 -384
rect 406268 -484 407704 -384
rect 406162 -490 406274 -484
<< via1 >>
rect 406172 23488 406272 23588
rect 406472 19488 406572 19588
rect 406772 15488 406872 15588
rect 407072 11488 407172 11588
rect 407372 7488 407472 7588
rect 406468 3494 406569 3595
rect 406168 -484 406268 -384
<< metal2 >>
rect 406172 23588 406272 23594
rect 406172 7292 406272 23488
rect 406472 19588 406572 19594
rect 406168 7287 406276 7292
rect 406168 7197 406177 7287
rect 406267 7197 406276 7287
rect 406168 7188 406276 7197
rect 406472 7096 406572 19488
rect 406472 7006 406477 7096
rect 406567 7006 406572 7096
rect 406472 7001 406572 7006
rect 406772 15588 406872 15594
rect 406477 6997 406567 7001
rect 406772 6159 406872 15488
rect 406772 6069 406777 6159
rect 406867 6069 406872 6159
rect 406772 6064 406872 6069
rect 407072 11588 407172 11594
rect 406777 6060 406867 6064
rect 407072 5959 407172 11488
rect 407072 5869 407077 5959
rect 407167 5869 407172 5959
rect 407072 5864 407172 5869
rect 407372 7588 407472 7594
rect 407077 5860 407167 5864
rect 407372 5759 407472 7488
rect 407372 5669 407377 5759
rect 407467 5669 407472 5759
rect 407372 5664 407472 5669
rect 407377 5660 407467 5664
rect 406473 5210 406563 5214
rect 406468 5205 406568 5210
rect 406468 5115 406473 5205
rect 406563 5115 406568 5205
rect 406173 5010 406263 5014
rect 406168 5005 406268 5010
rect 406168 4915 406173 5005
rect 406263 4915 406268 5005
rect 5078 -490 5134 1110
rect 13542 -490 13598 1110
rect 22006 -490 22062 1110
rect 30470 -490 30526 1110
rect 38934 -490 38990 1110
rect 47398 -490 47454 1110
rect 55862 -490 55918 1110
rect 64326 -490 64382 1110
rect 72790 -490 72846 1110
rect 81254 -490 81310 1110
rect 89718 -490 89774 1110
rect 98182 -490 98238 1110
rect 106646 -490 106702 1110
rect 115110 -490 115166 1110
rect 123574 -490 123630 1110
rect 132038 -490 132094 1110
rect 140502 -490 140558 1110
rect 148966 -490 149022 1110
rect 157430 -490 157486 1110
rect 165894 -490 165950 1110
rect 174358 -490 174414 1110
rect 182822 -490 182878 1110
rect 191286 -490 191342 1110
rect 199750 -490 199806 1110
rect 208214 -490 208270 1110
rect 216678 -490 216734 1110
rect 225142 -490 225198 1110
rect 233606 -490 233662 1110
rect 242070 -490 242126 1110
rect 250534 -490 250590 1110
rect 258998 -490 259054 1110
rect 267462 -490 267518 1110
rect 275926 -490 275982 1110
rect 284390 -490 284446 1110
rect 292854 -490 292910 1110
rect 301318 -490 301374 1110
rect 309782 -490 309838 1110
rect 318246 -490 318302 1110
rect 326710 -490 326766 1110
rect 335174 -490 335230 1110
rect 343638 -490 343694 1110
rect 352102 -490 352158 1110
rect 360566 -490 360622 1110
rect 369030 -490 369086 1110
rect 377494 -490 377550 1110
rect 385958 -490 386014 1110
rect 394422 -490 394478 1110
rect 402886 -490 402942 1110
rect 406168 -378 406268 4915
rect 406468 4478 406568 5115
rect 406468 3601 406569 4478
rect 406462 3595 406575 3601
rect 406462 3494 406468 3595
rect 406569 3494 406575 3595
rect 406462 3488 406575 3494
rect 406162 -384 406274 -378
rect 406162 -484 406168 -384
rect 406268 -484 406274 -384
rect 406162 -490 406274 -484
<< via2 >>
rect 406177 7197 406267 7287
rect 406477 7006 406567 7096
rect 406777 6069 406867 6159
rect 407077 5869 407167 5959
rect 407377 5669 407467 5759
rect 406473 5115 406563 5205
rect 406173 4915 406263 5005
<< metal3 >>
rect 406172 7287 406272 7292
rect 406172 7197 406177 7287
rect 406267 7197 406272 7287
rect 406172 7192 406272 7197
rect 406154 7096 406572 7101
rect 406154 7006 406477 7096
rect 406567 7006 406572 7096
rect 406154 7001 406572 7006
rect 406168 6159 406872 6164
rect 406168 6069 406777 6159
rect 406867 6069 406872 6159
rect 406168 6064 406872 6069
rect 406172 5959 407172 5964
rect 406172 5869 407077 5959
rect 407167 5869 407172 5959
rect 406172 5864 407172 5869
rect 406172 5759 407472 5764
rect 406172 5669 407377 5759
rect 407467 5669 407472 5759
rect 406172 5664 407472 5669
rect 406170 5205 406568 5210
rect 406170 5115 406473 5205
rect 406563 5115 406568 5205
rect 406170 5110 406568 5115
rect 406168 5005 406268 5010
rect 406168 4915 406173 5005
rect 406263 4915 406268 5005
rect 406168 4910 406268 4915
use filter_p_m  filter_p_m_0
array 0 7 50784 0 0 13945
timestamp 1663891137
transform 1 0 26 0 -1 36650
box -26 -328 50758 37140
<< labels >>
flabel metal2 5078 -490 5134 -490 1 FreeSans 1600 0 0 0 fb1[0]
port 1 s default input
flabel metal2 55862 -490 55918 -490 5 FreeSans 1600 0 0 0 fb1[1]
port 2 n default input
flabel metal2 106646 -490 106702 -490 5 FreeSans 1600 0 0 0 fb1[2]
port 3 n default input
flabel metal2 157430 -490 157486 -490 5 FreeSans 1600 0 0 0 fb1[3]
port 4 n default input
flabel metal2 208214 -490 208270 -490 5 FreeSans 1600 0 0 0 fb1[4]
port 5 n default input
flabel metal2 258998 -490 259054 -490 5 FreeSans 1600 0 0 0 fb1[5]
port 6 n default input
flabel metal2 309782 -490 309838 -490 5 FreeSans 1600 0 0 0 fb1[6]
port 7 n default input
flabel metal2 360566 -490 360622 -490 5 FreeSans 1600 0 0 0 fb1[7]
port 8 n default input
flabel metal2 13542 -490 13598 -490 5 FreeSans 1600 0 0 0 cclk[0]
port 9 n default input
flabel metal2 64326 -490 64382 -490 5 FreeSans 1600 0 0 0 cclk[1]
port 10 n default input
flabel metal2 115110 -490 115166 -490 5 FreeSans 1600 0 0 0 cclk[2]
port 11 n default input
flabel metal2 165894 -490 165950 -490 5 FreeSans 1600 0 0 0 cclk[3]
port 12 n default input
flabel metal2 216678 -490 216734 -490 5 FreeSans 1600 0 0 0 cclk[4]
port 13 n default input
flabel metal2 267462 -490 267518 -490 5 FreeSans 1600 0 0 0 cclk[5]
port 14 n default input
flabel metal2 318246 -490 318302 -490 5 FreeSans 1600 0 0 0 cclk[6]
port 15 n default input
flabel metal2 369030 -490 369086 -490 5 FreeSans 1600 0 0 0 cclk[7]
port 16 n default input
flabel metal2 22006 -490 22062 -490 5 FreeSans 1600 0 0 0 div2[0]
port 17 n default input
flabel metal2 72790 -490 72846 -490 5 FreeSans 1600 0 0 0 div2[1]
port 18 n default input
flabel metal2 123574 -490 123630 -490 5 FreeSans 1600 0 0 0 div2[2]
port 19 n default input
flabel metal2 174358 -490 174414 -490 5 FreeSans 1600 0 0 0 div2[3]
port 20 n default input
flabel metal2 225142 -490 225198 -490 5 FreeSans 1600 0 0 0 div2[4]
port 21 n default input
flabel metal2 275926 -490 275982 -490 5 FreeSans 1600 0 0 0 div2[5]
port 22 n default input
flabel metal2 326710 -490 326766 -490 5 FreeSans 1600 0 0 0 div2[6]
port 23 n default input
flabel metal2 377494 -490 377550 -490 5 FreeSans 1600 0 0 0 div2[7]
port 24 n default input
flabel metal2 30470 -490 30526 -490 5 FreeSans 1600 0 0 0 high_buf[0]
port 25 n default output
flabel metal2 81254 -490 81310 -490 5 FreeSans 1600 0 0 0 high_buf[1]
port 26 n default output
flabel metal2 132038 -490 132094 -490 5 FreeSans 1600 0 0 0 high_buf[2]
port 27 n default output
flabel metal2 182822 -490 182878 -490 5 FreeSans 1600 0 0 0 high_buf[3]
port 28 n default output
flabel metal2 233606 -490 233662 -490 5 FreeSans 1600 0 0 0 high_buf[4]
port 29 n default output
flabel metal2 284390 -490 284446 -490 5 FreeSans 1600 0 0 0 high_buf[5]
port 30 n default output
flabel metal2 335174 -490 335230 -490 5 FreeSans 1600 0 0 0 high_buf[6]
port 31 n default output
flabel metal2 385958 -490 386014 -490 5 FreeSans 1600 0 0 0 high_buf[7]
port 32 n default output
flabel metal2 38934 -490 38990 -490 5 FreeSans 1600 0 0 0 phi1b_dig[0]
port 33 n default output
flabel metal2 89718 -490 89774 -490 5 FreeSans 1600 0 0 0 phi1b_dig[1]
port 34 n default output
flabel metal2 140502 -490 140558 -490 5 FreeSans 1600 0 0 0 phi1b_dig[2]
port 35 n default output
flabel metal2 191286 -490 191342 -490 5 FreeSans 1600 0 0 0 phi1b_dig[3]
port 36 n default output
flabel metal2 242070 -490 242126 -490 5 FreeSans 1600 0 0 0 phi1b_dig[4]
port 37 n default output
flabel metal2 292854 -490 292910 -490 5 FreeSans 1600 0 0 0 phi1b_dig[5]
port 38 n default output
flabel metal2 343638 -490 343694 -490 5 FreeSans 1600 0 0 0 phi1b_dig[6]
port 39 n default output
flabel metal2 394422 -490 394478 -490 5 FreeSans 1600 0 0 0 phi1b_dig[7]
port 40 n default output
flabel metal2 47398 -490 47454 -490 5 FreeSans 1600 0 0 0 lo[0]
port 41 n default input
flabel metal2 98182 -490 98238 -490 5 FreeSans 1600 0 0 0 lo[1]
port 42 n default input
flabel metal2 148966 -490 149022 -490 5 FreeSans 1600 0 0 0 lo[2]
port 43 n default input
flabel metal2 199750 -490 199806 -490 5 FreeSans 1600 0 0 0 lo[3]
port 44 n default input
flabel metal2 250534 -490 250590 -490 5 FreeSans 1600 0 0 0 lo[4]
port 45 n default input
flabel metal2 301318 -490 301374 -490 5 FreeSans 1600 0 0 0 lo[5]
port 46 n default input
flabel metal2 352102 -490 352158 -490 5 FreeSans 1600 0 0 0 lo[6]
port 47 n default input
flabel metal2 402886 -490 402942 -490 5 FreeSans 1600 0 0 0 lo[7]
port 48 n default input
flabel metal1 407704 -484 407704 -384 5 FreeSans 1600 0 0 0 vnb
port 49 n default bidirectional
flabel metal1 407704 3494 407704 3595 5 FreeSans 1600 0 0 0 vpb
port 50 n default bidirectional
flabel metal1 407704 7488 407704 7588 5 FreeSans 1600 0 0 0 vccd1
port 51 n power bidirectional
flabel metal1 407704 11488 407704 11588 5 FreeSans 1600 0 0 0 th1
port 52 n default bidirectional
flabel metal1 407704 15488 407704 15588 5 FreeSans 1600 0 0 0 th2
port 53 n default bidirectional
flabel metal1 407704 19488 407704 19588 5 FreeSans 1600 0 0 0 vssd1
port 54 n ground bidirectional
flabel metal1 407704 23488 407704 23588 5 FreeSans 1600 0 0 0 vdda1
port 55 n power bidirectional
<< end >>
