** sch_path: /local_disk/fossi_cochlea/xschem/tryandtest/for_lvs.sch
.subckt for_lvs inp inm vdda vccd fb1 vssd div2 cclk phi1b_dig high_buf th1 th2 vpb vnb lo
*.PININFO inp:I inm:I vdda:B vccd:B fb1:I vssd:B div2:I cclk:I phi1b_dig:O high_buf:O th1:B th2:B
*+ vpb:B vnb:B lo:I
x1 cclk phi2b phi2 phi1b phi1 cclkb_ana cclk_ana vpb vnb vdda vssd vccd div2
+ filter_clkgen_balanced_clks
XC7 net1 vssd sky130_fd_pr__cap_mim_m3_1 W=6.7 L=6 MF=1 m=1
XC8 net5 vssd sky130_fd_pr__cap_mim_m3_1 W=3.4 L=3 MF=1 m=1
XC9 net3 vssd sky130_fd_pr__cap_mim_m3_1 W=4 L=5 MF=1 m=1
XC10 net4 vssd sky130_fd_pr__cap_mim_m3_1 W=3.4 L=3 MF=1 m=1
x2 th2 th1 cclk_ana cclkb_ana net6 vssd vdda analogMux
XC17 net7 vssd sky130_fd_pr__cap_mim_m3_1 W=6.7 L=6 MF=1 m=1
XC18 net11 vssd sky130_fd_pr__cap_mim_m3_1 W=3.4 L=3 MF=1 m=1
XC19 net9 vssd sky130_fd_pr__cap_mim_m3_1 W=4 L=5 MF=1 m=1
XC20 net10 vssd sky130_fd_pr__cap_mim_m3_1 W=3.4 L=3 MF=1 m=1
x4 th1 th2 cclk_ana cclkb_ana net12 vssd vdda analogMux
x5 inm inp ctrl ctrl_ net13 vssd vdda analogMux
x6 inp inm ctrl ctrl_ net20 vssd vdda analogMux
x7 inm inp ctrl ctrl_ net21 vssd vdda analogMux
x8 inp inm ctrl ctrl_ net14 vssd vdda analogMux
x13 fb_inv net5 phi1b phi1 vdda vssd switch Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
x9 net2 vssd mim_cap_stacked_12pF
x10 net8 vssd mim_cap_stacked_12pF
x11 net16 vssd mim_cap_stacked_6pF
x12 high net6 mim_cap_stacked_3pF
x29 net17 vssd mim_cap_stacked_6pF
x30 low net12 mim_cap_stacked_3pF
x33 vdda net19 fb_inv fb vssd net18 level_up_shifter_no_inv
X34 fb1 net18 net19 vccd vssd comp_clks_1stage Wpmos=1.26 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x35 high low high_buf phi1_dig phi1b_dig net15 vccd vssd comparator_single_tail Wplus=0.42
+ Lplus=0.42 Wminus=0.42 Lminus=0.15
x3 vdda vccd phi1 phi1_dig vssd level_down_shifter
x31 vdda vccd phi1b phi1b_dig vssd level_down_shifter
x14 net5 net2 phi2b phi2 vdda vssd switch Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
x15 net13 net1 phi1b phi1 vdda vssd switch Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
x16 net1 net2 phi2b phi2 vdda vssd switch Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
x17 net2 net3 phi1b phi1 vdda vssd switch Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
x18 net3 net16 phi2b phi2 vdda vssd switch Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
x19 net16 net4 phi1b phi1 vdda vssd switch Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
x20 net4 high phi2b phi2 vdda vssd switch Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
x21 fb net11 phi1b phi1 vdda vssd switch Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
x22 net11 net8 phi2b phi2 vdda vssd switch Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
x23 net14 net7 phi1b phi1 vdda vssd switch Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
x24 net7 net8 phi2b phi2 vdda vssd switch Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
x25 net8 net9 phi1b phi1 vdda vssd switch Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
x26 net9 net17 phi2b phi2 vdda vssd switch Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
x27 net17 net10 phi1b phi1 vdda vssd switch Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
x28 net10 low phi2b phi2 vdda vssd switch Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
x32 vdda net23 ctrl_ ctrl vssd net22 level_up_shifter_no_inv
X36 lo net22 net23 vccd vssd comp_clks_1stage Wpmos=1.26 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
**** begin user architecture code
 .lib /local_disk/fossi_cochlea/dependencies/pdks/sky130B/libs.tech/ngspice/sky130.lib.spice tt
.include /local_disk/fossi_cochlea/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
.ends

* expanding   symbol:  clkgen/filter_clkgen_balanced_clks.sym # of pins=13
** sym_path: /local_disk/fossi_cochlea/xschem/clkgen/filter_clkgen_balanced_clks.sym
** sch_path: /local_disk/fossi_cochlea/xschem/clkgen/filter_clkgen_balanced_clks.sch
.subckt filter_clkgen_balanced_clks cclk phi2b phi2 phi1b phi1 cclkb_ana cclk_ana vpb vnb vdda vssd
+ vccd div2
*.PININFO div2:I phi2:O phi2b:O phi1:O phi1b:O cclk_ana:O cclkb_ana:O vpb:I vnb:I cclk:I vdda:B
*+ vccd:B vssd:B
X4 phi2dd phi2 phi2b vdda vssd comp_clks Wpmos=1.26 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
X7 phi1dd phi1 phi1b vdda vssd comp_clks Wpmos=1.26 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
X10 div2dd cclk_ana cclkb_ana vdda vssd comp_clks Wpmos=1.26 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
X2 net1 phi2d vnb vdda vssd inv_weak_pulldown Wpmos=1.26 Lpmos= Wnmos= Lnmos=0.54
X5 net2 phi1d vnb vdda vssd inv_weak_pulldown Wpmos=1.26 Lpmos= Wnmos= Lnmos=0.54
X8 net3 div2d vnb vdda vssd inv_weak_pulldown Wpmos=1.26 Lpmos= Wnmos= Lnmos=0.54
X9 div2d div2dd vnb vdda vssd inv_weak_pulldown Wpmos=1.26 Lpmos= Wnmos= Lnmos=0.54
X3 phi2d phi2dd vpb vdda vssd inv_weak_pullup Wpmos=1.26 Lpmos=0.54 Wnmos= Lnmos=
X6 phi1d phi1dd vpb vdda vssd inv_weak_pullup Wpmos=1.26 Lpmos=0.54 Wnmos= Lnmos=
x12 vdda vccd vssd div2 net2 net1 level_up_shifter_d_a
x1 vdda vccd vssd cclk net4 net3 level_up_shifter_d_a
.ends


* expanding   symbol:  mux/analogMux.sym # of pins=7
** sym_path: /local_disk/fossi_cochlea/xschem/mux/analogMux.sym
** sch_path: /local_disk/fossi_cochlea/xschem/mux/analogMux.sch
.subckt analogMux vref2 vref1 c cbar out vssa vdda
*.PININFO vref1:I out:O vref2:I c:I cbar:I vssa:I vdda:I
XM2 vref1 c out vssa sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 vref1 cbar out vdda sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 out cbar vref2 vssa sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 out c vref2 vdda sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  transmission_gate/switch.sym # of pins=6
** sym_path: /local_disk/fossi_cochlea/xschem/transmission_gate/switch.sym
** sch_path: /local_disk/fossi_cochlea/xschem/transmission_gate/switch.sch
.subckt switch in out ctrl_ ctrl vdd vss   Wpmos=Wpmos Lpmos=Lpmos Wnmos=Wnmos Lnmos=Lnmos
*.PININFO in:B out:B ctrl_:I ctrl:I vdd:B vss:B
XM1 out ctrl in vss sky130_fd_pr__nfet_01v8 L=Lnmos W=Wnmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out ctrl_ in vdd sky130_fd_pr__pfet_01v8 L=Lpmos W=Wpmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  Switched_Caps/mim_cap_stacked_12pF.sym # of pins=2
** sym_path: /local_disk/fossi_cochlea/xschem/Switched_Caps/mim_cap_stacked_12pF.sym
** sch_path: /local_disk/fossi_cochlea/xschem/Switched_Caps/mim_cap_stacked_12pF.sch
.subckt mim_cap_stacked_12pF sig vss
*.PININFO sig:B vss:B
XC1 sig vss sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=32 m=32
XC2 vss sig sky130_fd_pr__cap_mim_m3_2 W=10 L=10 VM=32 m=32
.ends


* expanding   symbol:  Switched_Caps/mim_cap_stacked_6pF.sym # of pins=2
** sym_path: /local_disk/fossi_cochlea/xschem/Switched_Caps/mim_cap_stacked_6pF.sym
** sch_path: /local_disk/fossi_cochlea/xschem/Switched_Caps/mim_cap_stacked_6pF.sch
.subckt mim_cap_stacked_6pF sig vss
*.PININFO sig:B vss:B
XC1 sig vss sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=16 m=16
XC2 vss sig sky130_fd_pr__cap_mim_m3_2 W=10 L=10 VM=16 m=16
.ends


* expanding   symbol:  Switched_Caps/mim_cap_stacked_3pF.sym # of pins=2
** sym_path: /local_disk/fossi_cochlea/xschem/Switched_Caps/mim_cap_stacked_3pF.sym
** sch_path: /local_disk/fossi_cochlea/xschem/Switched_Caps/mim_cap_stacked_3pF.sch
.subckt mim_cap_stacked_3pF sig ref
*.PININFO sig:B ref:B
XC1 sig ref sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=8 m=8
XC2 ref sig sky130_fd_pr__cap_mim_m3_2 W=10 L=10 VM=8 m=8
.ends


* expanding   symbol:  level_shifter/level_up_shifter_no_inv.sym # of pins=6
** sym_path: /local_disk/fossi_cochlea/xschem/level_shifter/level_up_shifter_no_inv.sym
** sch_path: /local_disk/fossi_cochlea/xschem/level_shifter/level_up_shifter_no_inv.sch
.subckt level_up_shifter_no_inv vdd in outb out vss inb
*.PININFO in:I vdd:B out:O outb:O inb:I vss:B
XM7 outb out vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 out outb vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 outb inb vdd vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM3 outb in vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM4 vss in outb vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM5 out inb vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM6 vss inb out vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM9 vdd in out vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM10 out in vdd vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM11 vdd inb outb vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
.ends


* expanding   symbol:  clkgen/comp_clks_1stage.sym # of pins=5
** sym_path: /local_disk/fossi_cochlea/xschem/clkgen/comp_clks_1stage.sym
** sch_path: /local_disk/fossi_cochlea/xschem/clkgen/comp_clks_1stage.sch
.subckt comp_clks_1stage clk clka clkb vdd vss   Wpmos=1.26 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
*.PININFO clk:I clka:O clkb:O vdd:B vss:B
X1 clk clka vdd vss inv Wpmos=Wpmos Lpmos=Lpmos Wnmos=Wnmos Lnmos=Lnmos
x2 clk clkb vss vdd vdd vss tg
.ends


* expanding   symbol:  xschem/comparator_latest/comparator_single_tail.sym # of pins=8
** sym_path: /local_disk/fossi_cochlea/xschem/comparator_latest/comparator_single_tail.sym
** sch_path: /local_disk/fossi_cochlea/xschem/comparator_latest/comparator_single_tail.sch
.subckt comparator_single_tail inp inm high_buf phi1 phi1b low_buf vccd vssd   Wplus=0.42 Lplus=0.15
+ Wminus=0.42 Lminus=0.15
*.PININFO phi1:I phi1b:I inp:I inm:I low_buf:O vccd:B vssd:B high_buf:O
XM12 FP inp tail vssd sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM13 FN inm tail vssd sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM14 pfetw low vccd vccd sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 high FP pfetw vccd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 pfete FN low vccd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 vccd high pfete vccd sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 low high vssd vssd sky130_fd_pr__nfet_01v8_lvt L=2 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 high low vssd vssd sky130_fd_pr__nfet_01v8_lvt L=2 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 tail phi1 vssd vssd sky130_fd_pr__nfet_01v8_lvt L=2 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 vccd phi1 FP vccd sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 FN phi1 vccd vccd sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
X1 high net1 vccd vssd inv Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
X2 net1 net2 vccd vssd inv Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
X3 net2 net3 vccd vssd inv Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
X4 net3 high_buf vccd vssd inv Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
X5 low net4 vccd vssd inv Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
X6 net4 net5 vccd vssd inv Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
X7 net5 net6 vccd vssd inv Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
X8 net6 low_buf vccd vssd inv Wpmos=0.42 Lpmos=0.15 Wnmos=0.42 Lnmos=0.15
XM4 high phi1b vssd vssd sky130_fd_pr__nfet_01v8_lvt L=2 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 low phi1b vssd vssd sky130_fd_pr__nfet_01v8_lvt L=2 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  xschem/level_shifter/level_down_shifter.sym # of pins=5
** sym_path: /local_disk/fossi_cochlea/xschem/level_shifter/level_down_shifter.sym
** sch_path: /local_disk/fossi_cochlea/xschem/level_shifter/level_down_shifter.sch
.subckt level_down_shifter vdda vccd in out vssd
*.PININFO in:I vssd:B vdda:B out:O vccd:B
x1 in vssd vssd vdda vdda net1 sky130_fd_sc_hd__inv_8
x2 net1 vssd vssd vccd vccd out sky130_fd_sc_hd__inv_8
.ends


* expanding   symbol:  clkgen/comp_clks.sym # of pins=5
** sym_path: /local_disk/fossi_cochlea/xschem/clkgen/comp_clks.sym
** sch_path: /local_disk/fossi_cochlea/xschem/clkgen/comp_clks.sch
.subckt comp_clks clk clka clkb vdd vss   Wpmos=Wpmos Lpmos=Lpmos Wnmos=Wnmos Lnmos=Lnmos
*.PININFO clk:I clka:O clkb:O vdd:B vss:B
X1 clk clki vdd vss inv Wpmos=Wpmos Lpmos=Lpmos Wnmos=Wnmos Lnmos=Lnmos
X2 clki clka vdd vss inv Wpmos=Wpmos Lpmos=Lpmos Wnmos=Wnmos Lnmos=Lnmos
X4 clkt clkb vdd vss inv Wpmos=Wpmos Lpmos=Lpmos Wnmos=Wnmos Lnmos=Lnmos
x3 clk clkt vss vdd vdd vss tg
.ends


* expanding   symbol:  inv/inv_weak_pulldown.sym # of pins=5
** sym_path: /local_disk/fossi_cochlea/xschem/inv/inv_weak_pulldown.sym
** sch_path: /local_disk/fossi_cochlea/xschem/inv/inv_weak_pulldown.sch
.subckt inv_weak_pulldown in out Vnb vdda vssa   Wpmos=1.26 Lmin=0.18 Wmin=0.42 Lnmos=0.54
*.PININFO in:I out:B Vnb:I vdda:I vssa:I
XM1 net1 in vssa vssa sky130_fd_pr__nfet_01v8 L=Lmin W=Wmin nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 out Vnb net1 vssa sky130_fd_pr__nfet_01v8 L=Lnmos W=Wmin nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 out in vdda vdda sky130_fd_pr__pfet_01v8 L=Lmin W=Wpmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  inv/inv_weak_pullup.sym # of pins=5
** sym_path: /local_disk/fossi_cochlea/xschem/inv/inv_weak_pullup.sym
** sch_path: /local_disk/fossi_cochlea/xschem/inv/inv_weak_pullup.sch
.subckt inv_weak_pullup in out Vpb vdda vssa   Wpmos=1.26 Lpmos=0.54 Wmin=0.42 Lmin=0.18
*.PININFO in:I out:B Vpb:I vdda:I vssa:I
XM1 out in vssa vssa sky130_fd_pr__nfet_01v8 L=Lmin W=Wmin nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 out Vpb net1 vdda sky130_fd_pr__pfet_01v8 L=Lpmos W=Wpmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net1 in vdda vdda sky130_fd_pr__pfet_01v8 L=Lmin W=Wpmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  xschem/level_shifter/level_up_shifter_d_a.sym # of pins=6
** sym_path: /local_disk/fossi_cochlea/xschem/level_shifter/level_up_shifter_d_a.sym
** sch_path: /local_disk/fossi_cochlea/xschem/level_shifter/level_up_shifter_d_a.sch
.subckt level_up_shifter_d_a vdda vccd vssd clk outb out
*.PININFO clk:I outb:O out:O vdda:B vccd:B vssd:B
X1 clk net1 net2 vccd vssd comp_clks_1stage Wpmos=1.26 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x15 vdda net1 outb out vssd net2 level_up_shifter_no_inv
.ends


* expanding   symbol:  inv/inv.sym # of pins=4
** sym_path: /local_disk/fossi_cochlea/xschem/inv/inv.sym
** sch_path: /local_disk/fossi_cochlea/xschem/inv/inv.sch
.subckt inv in out vdd vss   Wpmos=Wpmos Lpmos=Lpmos Wnmos=Wnmos Lnmos=Lnmos
*.PININFO in:I out:B vdd:B vss:B
XM1 vss in out vss sky130_fd_pr__nfet_01v8 L=Lnmos W=Wnmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 vdd in out vdd sky130_fd_pr__pfet_01v8 L=Lpmos W=Wpmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  xschem/transmission_gate/tg.sym # of pins=6
** sym_path: /local_disk/fossi_cochlea/xschem/transmission_gate/tg.sym
** sch_path: /local_disk/fossi_cochlea/xschem/transmission_gate/tg.sch
.subckt tg in out ctrl_ ctrl vdd vss
*.PININFO in:B out:B ctrl_:I ctrl:I vdd:B vss:B
XM1 out ctrl in vss sky130_fd_pr__nfet_01v8 L=0.18 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out ctrl_ in vdd sky130_fd_pr__pfet_01v8 L=0.18 W=0.63 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
.ends

.end
