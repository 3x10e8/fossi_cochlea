magic
tech sky130B
magscale 1 2
timestamp 1661198472
<< error_p >>
rect -35473 138898 -35064 139218
rect 13209 138898 13618 139218
rect -35483 138003 -35074 138323
rect 13199 138003 13608 138323
rect -35491 136881 -35039 137201
rect -14891 136881 -14439 137201
rect 13191 136881 13643 137201
rect 33791 136881 34243 137201
rect -35470 135450 -35061 135770
rect -14869 135450 -14460 135770
rect 13212 135450 13621 135770
rect 33813 135450 34222 135770
rect -25008 133789 -24931 133795
rect 23674 133789 23751 133795
rect -24998 133725 -24942 133731
rect -24937 133725 -24931 133789
rect 23684 133725 23740 133731
rect 23745 133725 23751 133789
rect -25008 133716 -24931 133725
rect 23674 133716 23751 133725
rect -24998 133703 -24942 133716
rect 23684 133703 23740 133716
rect -48509 133244 -48503 133250
rect -48463 133244 -48457 133250
rect -48515 133238 -48451 133244
rect -48509 133198 -48457 133238
rect -48252 133206 -48218 133240
rect -48072 133206 -48038 133256
rect -47815 133239 -47809 133245
rect -47769 133239 -47763 133245
rect -47821 133233 -47757 133239
rect -25734 133236 -25657 133242
rect -24282 133237 -24205 133242
rect -2167 133239 -2161 133245
rect -2121 133239 -2115 133245
rect -48515 133192 -48451 133198
rect -47815 133193 -47763 133233
rect -48509 133186 -48503 133192
rect -48463 133186 -48457 133192
rect -47821 133187 -47757 133193
rect -47815 133181 -47809 133187
rect -47769 133181 -47763 133187
rect -25664 133172 -25657 133236
rect -25734 133166 -25657 133172
rect -24211 133171 -24205 133237
rect -2173 133233 -2109 133239
rect -2167 133193 -2115 133233
rect -1892 133206 -1858 133256
rect -1473 133244 -1467 133250
rect -1427 133244 -1421 133250
rect 173 133244 179 133250
rect 219 133244 225 133250
rect -1712 133206 -1678 133240
rect -1479 133238 -1415 133244
rect 167 133238 231 133244
rect -1473 133198 -1421 133238
rect 173 133198 225 133238
rect 430 133206 464 133240
rect 610 133206 644 133256
rect 867 133239 873 133245
rect 913 133239 919 133245
rect 861 133233 925 133239
rect 22948 133236 23025 133242
rect 24400 133237 24477 133242
rect 46515 133239 46521 133245
rect 46561 133239 46567 133245
rect -2173 133187 -2109 133193
rect -1479 133192 -1415 133198
rect 167 133192 231 133198
rect 867 133193 919 133233
rect -2167 133181 -2161 133187
rect -2121 133181 -2115 133187
rect -1473 133186 -1467 133192
rect -1427 133186 -1421 133192
rect 173 133186 179 133192
rect 219 133186 225 133192
rect 861 133187 925 133193
rect 867 133181 873 133187
rect 913 133181 919 133187
rect 23018 133172 23025 133236
rect -24282 133166 -24205 133171
rect 22948 133166 23025 133172
rect 24471 133171 24477 133237
rect 46509 133233 46573 133239
rect 46515 133193 46567 133233
rect 46790 133206 46824 133256
rect 47209 133244 47215 133250
rect 47255 133244 47261 133250
rect 46970 133206 47004 133240
rect 47203 133238 47267 133244
rect 47209 133198 47261 133238
rect 46509 133187 46573 133193
rect 47203 133192 47267 133198
rect 46515 133181 46521 133187
rect 46561 133181 46567 133187
rect 47209 133186 47215 133192
rect 47255 133186 47261 133192
rect 24400 133166 24477 133171
rect -24997 133102 -24991 133108
rect -24951 133102 -24945 133108
rect 23685 133102 23691 133108
rect 23731 133102 23737 133108
rect -25003 133096 -24939 133102
rect 23679 133096 23743 133102
rect -24997 133056 -24945 133096
rect 23685 133056 23737 133096
rect -25003 133050 -24939 133056
rect 23679 133050 23743 133056
rect -24997 133044 -24991 133050
rect -24951 133044 -24945 133050
rect 23685 133044 23691 133050
rect 23731 133044 23737 133050
rect -26788 131091 -26747 131125
rect -23167 131091 -23129 131142
rect 21894 131091 21935 131125
rect 25515 131091 25553 131142
rect -27873 130420 -27867 130426
rect -27827 130420 -27821 130426
rect -22109 130420 -22103 130426
rect -22063 130420 -22057 130426
rect 20809 130420 20815 130426
rect 20855 130420 20861 130426
rect 26573 130420 26579 130426
rect 26619 130420 26625 130426
rect -27879 130414 -27815 130420
rect -22115 130414 -22051 130420
rect 20803 130414 20867 130420
rect 26567 130414 26631 130420
rect -27873 130374 -27821 130414
rect -22109 130374 -22057 130414
rect 20809 130374 20861 130414
rect 26573 130374 26625 130414
rect -27879 130368 -27815 130374
rect -22115 130368 -22051 130374
rect 20803 130368 20867 130374
rect 26567 130368 26631 130374
rect -27873 130362 -27867 130368
rect -27827 130362 -27821 130368
rect -22109 130362 -22103 130368
rect -22063 130362 -22057 130368
rect 20809 130362 20815 130368
rect 20855 130362 20861 130368
rect 26573 130362 26579 130368
rect 26619 130362 26625 130368
rect -26542 127532 -26536 127538
rect -26496 127532 -26490 127538
rect 22140 127532 22146 127538
rect 22186 127532 22192 127538
rect -26548 127526 -26484 127532
rect 22134 127526 22198 127532
rect -26542 127486 -26490 127526
rect 22140 127486 22192 127526
rect -26548 127480 -26484 127486
rect 22134 127480 22198 127486
rect -26542 127474 -26536 127480
rect -26496 127474 -26490 127480
rect 22140 127474 22146 127480
rect 22186 127474 22192 127480
rect -27187 127224 -27181 127230
rect -27141 127224 -27135 127230
rect 21495 127224 21501 127230
rect 21541 127224 21547 127230
rect -27193 127218 -27129 127224
rect 21489 127218 21553 127224
rect -27187 127178 -27135 127218
rect 21495 127178 21547 127218
rect -27193 127172 -27129 127178
rect 21489 127172 21553 127178
rect -27187 127166 -27181 127172
rect -27141 127166 -27135 127172
rect 21495 127166 21501 127172
rect 21541 127166 21547 127172
rect -26238 126937 -26187 126987
rect 22444 126937 22495 126987
rect -27186 126750 -27180 126756
rect -27140 126750 -27134 126756
rect 21496 126750 21502 126756
rect 21542 126750 21548 126756
rect -27192 126744 -27128 126750
rect 21490 126744 21554 126750
rect -27186 126704 -27134 126744
rect 21496 126704 21548 126744
rect -27192 126698 -27128 126704
rect 21490 126698 21554 126704
rect -27186 126692 -27180 126698
rect -27140 126692 -27134 126698
rect 21496 126692 21502 126698
rect 21542 126692 21548 126698
rect -26651 126386 -26547 126450
rect 22031 126386 22135 126450
rect -26547 126302 -26483 126386
rect 22135 126302 22199 126386
rect -3708 43434 -3702 43440
rect -3606 43434 -3600 43440
rect -3714 43428 -3708 43434
rect -3600 43428 -3594 43434
rect -3714 42866 -3708 42872
rect -3600 42866 -3594 42872
rect -3708 42860 -3702 42866
rect -3606 42860 -3600 42866
rect 25235 38680 25299 38764
rect 25299 38616 25403 38680
rect 25886 38368 25892 38374
rect 25932 38368 25938 38374
rect 25880 38362 25944 38368
rect 25886 38322 25938 38362
rect 25880 38316 25944 38322
rect 25886 38310 25892 38316
rect 25932 38310 25938 38316
rect 24939 38079 24990 38129
rect 25887 37894 25893 37900
rect 25933 37894 25939 37900
rect 25881 37888 25945 37894
rect 25887 37848 25939 37888
rect 25881 37842 25945 37848
rect 25887 37836 25893 37842
rect 25933 37836 25939 37842
rect 25242 37586 25248 37592
rect 25288 37586 25294 37592
rect 25236 37580 25300 37586
rect 25242 37540 25294 37580
rect 25236 37534 25300 37540
rect 25242 37528 25248 37534
rect 25288 37528 25294 37534
rect 20809 34698 20815 34704
rect 20855 34698 20861 34704
rect 26573 34698 26579 34704
rect 26619 34698 26625 34704
rect 20803 34692 20867 34698
rect 26567 34692 26631 34698
rect 20809 34652 20861 34692
rect 26573 34652 26625 34692
rect 20803 34646 20867 34652
rect 26567 34646 26631 34652
rect 20809 34640 20815 34646
rect 20855 34640 20861 34646
rect 26573 34640 26579 34646
rect 26619 34640 26625 34646
rect 21881 33924 21919 33975
rect 25499 33941 25540 33975
rect 23697 32016 23703 32022
rect 23743 32016 23749 32022
rect 23691 32010 23755 32016
rect 23697 31970 23749 32010
rect 23691 31964 23755 31970
rect 23697 31958 23703 31964
rect 23743 31958 23749 31964
rect -48509 31874 -48503 31880
rect -48463 31874 -48457 31880
rect -47815 31879 -47809 31885
rect -47769 31879 -47763 31885
rect -48515 31868 -48451 31874
rect -47821 31873 -47757 31879
rect -48509 31828 -48457 31868
rect -48515 31822 -48451 31828
rect -48252 31826 -48218 31860
rect -48509 31816 -48503 31822
rect -48463 31816 -48457 31822
rect -48072 31810 -48038 31860
rect -47815 31833 -47763 31873
rect -47821 31827 -47757 31833
rect 22957 31895 23034 31900
rect -2167 31879 -2161 31885
rect -2121 31879 -2115 31885
rect -2173 31873 -2109 31879
rect -1473 31874 -1467 31880
rect -1427 31874 -1421 31880
rect 173 31874 179 31880
rect 219 31874 225 31880
rect 867 31879 873 31885
rect 913 31879 919 31885
rect -2167 31833 -2115 31873
rect -1479 31868 -1415 31874
rect 167 31868 231 31874
rect 861 31873 925 31879
rect -47815 31821 -47809 31827
rect -47769 31821 -47763 31827
rect -2173 31827 -2109 31833
rect -2167 31821 -2161 31827
rect -2121 31821 -2115 31827
rect -1892 31810 -1858 31860
rect -1712 31826 -1678 31860
rect -1473 31828 -1421 31868
rect 173 31828 225 31868
rect -1479 31822 -1415 31828
rect 167 31822 231 31828
rect 430 31826 464 31860
rect -1473 31816 -1467 31822
rect -1427 31816 -1421 31822
rect 173 31816 179 31822
rect 219 31816 225 31822
rect 610 31810 644 31860
rect 867 31833 919 31873
rect 861 31827 925 31833
rect 22957 31829 22963 31895
rect 24409 31894 24486 31900
rect 24409 31830 24416 31894
rect 46515 31879 46521 31885
rect 46561 31879 46567 31885
rect 46509 31873 46573 31879
rect 47209 31874 47215 31880
rect 47255 31874 47261 31880
rect 46515 31833 46567 31873
rect 47203 31868 47267 31874
rect 867 31821 873 31827
rect 913 31821 919 31827
rect 22957 31824 23034 31829
rect 24409 31824 24486 31830
rect 46509 31827 46573 31833
rect 46515 31821 46521 31827
rect 46561 31821 46567 31827
rect 46790 31810 46824 31860
rect 46970 31826 47004 31860
rect 47209 31828 47261 31868
rect 47203 31822 47267 31828
rect 47209 31816 47215 31822
rect 47255 31816 47261 31822
rect 23694 31350 23750 31363
rect 23683 31341 23760 31350
rect 23683 31277 23689 31341
rect 23694 31335 23750 31341
rect 23683 31271 23760 31277
rect -35470 29296 -35061 29616
rect -14869 29296 -14460 29616
rect 13212 29296 13621 29616
rect 33813 29296 34222 29616
rect -35491 27865 -35039 28185
rect -14891 27865 -14439 28185
rect 13191 27865 13643 28185
rect 33791 27865 34243 28185
rect -14856 26743 -14447 27063
rect 33826 26743 34235 27063
rect -14866 25848 -14457 26168
rect 33816 25848 34225 26168
<< error_s >>
rect -26513 41980 -26507 41986
rect -26461 41980 -26455 41986
rect -26519 41974 -26449 41980
rect -26513 41930 -26455 41974
rect -26519 41924 -26449 41930
rect -26513 41918 -26507 41924
rect -26461 41918 -26455 41924
rect -26049 40896 -26043 40902
rect -25995 40896 -25989 40902
rect -26055 40890 -26049 40896
rect -25989 40890 -25983 40896
rect -26055 40838 -26049 40844
rect -25989 40838 -25983 40844
rect -26049 40832 -26043 40838
rect -25995 40832 -25989 40838
rect -23447 38680 -23383 38784
rect -23383 38616 -23279 38680
rect -22796 38368 -22790 38374
rect -22750 38368 -22744 38374
rect -22802 38362 -22738 38368
rect -22796 38322 -22744 38362
rect -22802 38316 -22738 38322
rect -22796 38310 -22790 38316
rect -22750 38310 -22744 38316
rect -23743 38079 -23692 38129
rect -22795 37894 -22789 37900
rect -22749 37894 -22743 37900
rect -22801 37888 -22737 37894
rect -22795 37848 -22743 37888
rect -22801 37842 -22737 37848
rect -22795 37836 -22789 37842
rect -22749 37836 -22743 37842
rect -23440 37586 -23434 37592
rect -23394 37586 -23388 37592
rect -23446 37580 -23382 37586
rect -23440 37540 -23388 37580
rect -23446 37534 -23382 37540
rect -23440 37528 -23434 37534
rect -23394 37528 -23388 37534
rect -27873 34698 -27867 34704
rect -27827 34698 -27821 34704
rect -22109 34698 -22103 34704
rect -22063 34698 -22057 34704
rect -27879 34692 -27815 34698
rect -22115 34692 -22051 34698
rect -27873 34652 -27821 34692
rect -22109 34652 -22057 34692
rect -27879 34646 -27815 34652
rect -22115 34646 -22051 34652
rect -27873 34640 -27867 34646
rect -27827 34640 -27821 34646
rect -22109 34640 -22103 34646
rect -22063 34640 -22057 34646
rect -26801 33924 -26763 33975
rect -23183 33941 -23142 33975
rect -24985 32016 -24979 32022
rect -24939 32016 -24933 32022
rect -24991 32010 -24927 32016
rect -24985 31970 -24933 32010
rect -24991 31964 -24927 31970
rect -24985 31958 -24979 31964
rect -24939 31958 -24933 31964
rect -25725 31895 -25648 31900
rect -25725 31829 -25719 31895
rect -24273 31894 -24196 31900
rect -24273 31830 -24266 31894
rect -25725 31824 -25648 31829
rect -24273 31824 -24196 31830
rect -24988 31350 -24932 31363
rect -24999 31341 -24922 31350
rect -24999 31277 -24993 31341
rect -24988 31335 -24932 31341
rect -24999 31271 -24922 31277
<< viali >>
rect -9808 42802 -9634 43538
<< metal1 >>
rect -9846 43538 -9590 43598
rect -9846 42802 -9808 43538
rect -9634 42802 -9590 43538
rect -9846 42746 -9590 42802
rect -9733 37898 -9671 42746
rect -22638 37836 -9671 37898
rect -19438 34012 -6846 34030
rect -19438 33954 -19418 34012
rect -19366 33954 -6846 34012
rect -19438 33938 -6846 33954
rect -19010 32590 -18874 32596
rect -19010 32546 -19004 32590
rect -26706 32540 -19004 32546
rect -26710 32470 -19004 32540
rect -18882 32524 -18874 32590
rect -18882 32470 -18872 32524
rect -26710 32422 -18872 32470
rect -26710 31910 -26674 32422
rect -6956 31274 -6864 33938
<< via1 >>
rect -9808 42802 -9634 43538
rect -19418 33954 -19366 34012
rect -19004 32470 -18882 32590
<< metal2 >>
rect -9846 43538 -9590 43598
rect -16028 43328 -15818 43354
rect -16028 42794 -15982 43328
rect -15842 42794 -15818 43328
rect -16028 42780 -15818 42794
rect -9846 42802 -9808 43538
rect -9634 42802 -9590 43538
rect -15987 42731 -15861 42780
rect -9846 42746 -9590 42802
rect -19008 42605 -15861 42731
rect -26160 42242 -26108 42272
rect -35742 42190 -26108 42242
rect -35742 36712 -35690 42190
rect -26160 41392 -26108 42190
rect -26856 41224 -26778 41234
rect -26856 41216 -26848 41224
rect -27750 41166 -26848 41216
rect -26788 41166 -26778 41224
rect -26856 41160 -26778 41166
rect -26818 40948 -26638 41000
rect -26818 40378 -26774 40948
rect -26818 40334 -19370 40378
rect -30362 38244 -30272 38254
rect -30362 38182 -30352 38244
rect -30282 38182 -30272 38244
rect -30362 38172 -30272 38182
rect -30360 37638 -30278 37648
rect -30360 37578 -30350 37638
rect -30288 37578 -30278 37638
rect -30360 37568 -30278 37578
rect -43040 36660 -35690 36712
rect -43040 36376 -42988 36660
rect -43040 31302 -42986 36376
rect -19414 34022 -19370 40334
rect -19424 34012 -19360 34022
rect -19424 33954 -19418 34012
rect -19366 33954 -19360 34012
rect -19424 33944 -19360 33954
rect -19008 32596 -18882 42605
rect -19010 32590 -18874 32596
rect -19010 32470 -19004 32590
rect -18882 32470 -18874 32590
rect -19010 32464 -18874 32470
<< via2 >>
rect -15982 42794 -15842 43328
rect -9808 42802 -9634 43538
rect -26848 41166 -26788 41224
rect -30352 38182 -30282 38244
rect -30350 37578 -30288 37638
<< metal3 >>
rect -28384 43127 -28044 43602
rect -9846 43538 -9590 43598
rect -31098 42941 -28044 43127
rect -31098 41582 -30912 42941
rect -28384 42788 -28044 42941
rect -22424 42535 -21460 43508
rect -16028 43328 -15818 43354
rect -16028 42794 -15982 43328
rect -15842 42794 -15818 43328
rect -16028 42780 -15818 42794
rect -9846 42802 -9808 43538
rect -9634 42802 -9590 43538
rect -9846 42746 -9590 42802
rect -30758 42456 -21460 42535
rect -30758 42436 -21927 42456
rect -31098 37650 -30916 41582
rect -30758 38252 -30659 42436
rect -22081 42408 -21927 42436
rect -26876 41234 -26770 41268
rect -26876 41160 -26856 41234
rect -26778 41160 -26770 41234
rect -26876 41136 -26770 41160
rect -30366 38252 -30272 38254
rect -30758 38244 -30272 38252
rect -30758 38182 -30352 38244
rect -30282 38182 -30272 38244
rect -30758 38172 -30272 38182
rect -30758 38170 -30274 38172
rect -30366 38168 -30274 38170
rect -31098 37638 -30278 37650
rect -31098 37578 -30350 37638
rect -30288 37578 -30278 37638
rect -31098 37568 -30278 37578
<< via3 >>
rect -3708 42866 -3600 43434
rect -26856 41224 -26778 41234
rect -26856 41166 -26848 41224
rect -26848 41166 -26788 41224
rect -26788 41166 -26778 41224
rect -26856 41160 -26778 41166
<< metal4 >>
rect -3730 43434 -3554 43600
rect -3730 42866 -3708 43434
rect -3600 42866 -3554 43434
rect -26876 41234 -26770 41268
rect -26876 41160 -26856 41234
rect -26778 41232 -26770 41234
rect -3730 41232 -3554 42866
rect -26778 41160 -3507 41232
rect -26876 41150 -3507 41160
rect -26876 41136 -26770 41150
rect -3730 41134 -3554 41150
use filter_p_m  filter_p_m_0
array 0 1 -48682 0 0 34550
timestamp 1661198472
transform 1 0 -321 0 1 5258
box -26 0 48102 37136
use filter_p_m  filter_p_m_1
array 0 1 -48682 0 0 34550
timestamp 1661198472
transform -1 0 -927 0 -1 159808
box -26 0 48102 37136
use first_dual_core  first_dual_core_0 ./mag/final_designs/digital/
timestamp 1661193354
transform 0 -1 48362 1 0 42794
box 0 0 80000 98000
<< end >>
