magic
tech sky130A
magscale 1 2
timestamp 1647917973
<< error_s >>
rect 8141 15958 8147 15964
rect 10933 15958 10939 15964
rect 3130 15949 3150 15955
rect 5522 15949 5542 15955
rect 8173 15934 8177 15954
rect 10903 15934 10907 15954
rect 3675 15923 3684 15933
rect 6067 15923 6076 15933
rect 6887 15931 6900 15933
rect 6934 15931 6953 15933
rect 6934 15923 6935 15931
rect 3108 15901 3109 15913
rect 5500 15901 5501 15913
rect 3641 15889 3650 15899
rect 6033 15889 6042 15899
rect 6853 15897 6866 15899
rect 6968 15897 6987 15899
rect 6968 15889 6969 15897
rect 3079 15871 3091 15883
rect 5471 15871 5483 15883
rect 3347 15850 3359 15859
rect 5739 15850 5751 15859
rect 8215 15846 8219 15866
rect 10861 15846 10865 15866
rect 8171 15824 8177 15830
rect 10903 15824 10909 15830
rect 3385 15812 3397 15821
rect 5777 15812 5789 15821
rect 2523 15797 2540 15803
rect 4915 15797 4932 15803
rect 1885 15468 1891 15474
rect 2779 15468 2796 15469
rect 1917 15444 1921 15464
rect 2813 15434 2830 15435
rect 1959 15356 1963 15376
rect 7797 15369 7813 15371
rect 9429 15369 9442 15371
rect 9544 15369 9563 15371
rect 1915 15334 1921 15340
rect 7763 15335 7779 15337
rect 9463 15335 9476 15337
rect 9510 15335 9529 15337
rect 2747 14843 2760 14845
rect 2794 14843 2813 14845
rect 5783 14843 5796 14845
rect 5830 14843 5849 14845
rect 7159 14843 7178 14845
rect 7212 14843 7225 14845
rect 8723 14843 8742 14845
rect 8776 14843 8789 14845
rect 10707 14843 10723 14845
rect 2794 14835 2795 14843
rect 2713 14809 2726 14811
rect 2828 14809 2847 14811
rect 5749 14809 5762 14811
rect 5864 14809 5883 14811
rect 7125 14809 7144 14811
rect 7246 14809 7259 14811
rect 8689 14809 8708 14811
rect 8810 14809 8823 14811
rect 10741 14809 10757 14811
rect 2828 14801 2829 14809
rect 11117 14380 11123 14386
rect 2426 14359 2427 14365
rect 11087 14356 11091 14376
rect 2460 14325 2461 14331
rect 7051 14283 7052 14291
rect 2345 14281 2358 14283
rect 2460 14281 2479 14283
rect 3841 14281 3857 14283
rect 5289 14281 5302 14283
rect 5404 14281 5423 14283
rect 7033 14281 7052 14283
rect 7154 14281 7167 14283
rect 7679 14281 7695 14283
rect 9705 14281 9718 14283
rect 9820 14281 9839 14283
rect 10347 14281 10363 14283
rect 11045 14268 11049 14288
rect 7085 14249 7086 14257
rect 2379 14247 2392 14249
rect 2426 14247 2445 14249
rect 3807 14247 3823 14249
rect 5323 14247 5336 14249
rect 5370 14247 5389 14249
rect 7067 14247 7086 14249
rect 7120 14247 7133 14249
rect 7713 14247 7729 14249
rect 9739 14247 9752 14249
rect 9786 14247 9805 14249
rect 10381 14247 10397 14249
rect 11087 14246 11093 14252
rect 3099 13954 3108 13960
rect 3071 13926 3080 13932
rect 1885 13782 1891 13788
rect 1917 13758 1921 13778
rect 4863 13755 4876 13757
rect 4910 13755 4929 13757
rect 4829 13721 4842 13723
rect 4944 13721 4963 13723
rect 1959 13670 1963 13690
rect 1915 13648 1921 13654
rect 10522 13327 10539 13333
rect 9703 13271 9715 13280
rect 10051 13251 10063 13263
rect 9741 13233 9753 13242
rect 10021 13209 10022 13221
rect 2461 13193 2477 13195
rect 4459 13193 4475 13195
rect 5745 13193 5764 13195
rect 5866 13193 5879 13195
rect 9992 13179 10012 13185
rect 2427 13159 2443 13161
rect 4493 13159 4509 13161
rect 5779 13159 5798 13161
rect 5832 13159 5845 13161
rect 10268 12866 10276 12872
rect 10296 12838 10304 12844
rect 2498 12685 2518 12691
rect 1964 12659 1973 12669
rect 6567 12667 6583 12669
rect 7211 12667 7227 12669
rect 8267 12667 8280 12669
rect 8314 12667 8333 12669
rect 9827 12667 9846 12669
rect 9880 12667 9893 12669
rect 2539 12637 2540 12649
rect 1998 12625 2007 12635
rect 6601 12633 6617 12635
rect 7245 12633 7261 12635
rect 8233 12633 8246 12635
rect 8348 12633 8367 12635
rect 9793 12633 9812 12635
rect 9914 12633 9927 12635
rect 2557 12607 2569 12619
rect 2289 12586 2301 12595
rect 2251 12548 2263 12557
rect 3108 12533 3125 12539
rect 3205 12239 3222 12245
rect 8774 12239 8791 12245
rect 1885 12204 1891 12210
rect 5505 12204 5511 12210
rect 10013 12204 10019 12210
rect 10993 12204 10999 12210
rect 1917 12180 1921 12200
rect 4029 12183 4041 12192
rect 5475 12180 5479 12200
rect 7955 12183 7967 12192
rect 9983 12180 9987 12200
rect 11025 12180 11029 12200
rect 3681 12163 3693 12175
rect 8303 12163 8315 12175
rect 3991 12145 4003 12154
rect 7993 12145 8005 12154
rect 3722 12121 3723 12133
rect 8273 12121 8274 12133
rect 1959 12092 1963 12112
rect 4285 12105 4294 12115
rect 3732 12091 3752 12097
rect 5433 12092 5437 12112
rect 7702 12105 7711 12115
rect 8244 12091 8264 12097
rect 9941 12092 9945 12112
rect 11067 12092 11071 12112
rect 1915 12070 1921 12076
rect 4319 12071 4328 12081
rect 5475 12070 5481 12076
rect 7668 12071 7677 12081
rect 9983 12070 9989 12076
rect 11023 12070 11029 12076
rect 5614 11597 5634 11603
rect 10582 11597 10602 11603
rect 6159 11571 6168 11581
rect 8173 11579 8189 11581
rect 11127 11571 11136 11581
rect 5592 11549 5593 11561
rect 10560 11549 10561 11561
rect 6125 11537 6134 11547
rect 8139 11545 8155 11547
rect 11093 11537 11102 11547
rect 5563 11519 5575 11531
rect 10531 11519 10543 11531
rect 5831 11498 5843 11507
rect 10799 11498 10811 11507
rect 2910 11481 2927 11482
rect 5869 11460 5881 11469
rect 10837 11460 10849 11469
rect 2944 11447 2961 11448
rect 5007 11445 5024 11451
rect 9975 11445 9992 11451
<< nwell >>
rect 2242 16212 2564 16281
rect 14580 11851 14755 12005
rect 2654 11088 2854 11097
rect 2654 11031 2854 11039
rect 2617 10618 2940 10807
<< pwell >>
rect 2405 11057 2561 11242
rect 2404 11031 2534 11045
<< ndiff >>
rect 2404 11031 2534 11045
<< pdiff >>
rect 2654 11031 2854 11039
<< psubdiff >>
rect 2372 11209 2518 11214
rect 2372 11174 2427 11209
rect 2462 11174 2518 11209
rect 2372 11165 2518 11174
<< nsubdiff >>
rect 2654 11093 2854 11097
rect 2654 11059 2730 11093
rect 2764 11059 2854 11093
rect 2654 11039 2854 11059
<< psubdiffcont >>
rect 2427 11174 2462 11209
<< nsubdiffcont >>
rect 2730 11059 2764 11093
<< locali >>
rect 14927 11592 14959 11593
rect 14927 11462 14961 11592
rect 2340 11214 2374 11268
rect 2340 11209 2518 11214
rect 2340 11174 2427 11209
rect 2462 11174 2518 11209
rect 2340 11165 2518 11174
rect 2340 11096 2374 11165
rect 2656 11093 2885 11099
rect 2656 11059 2730 11093
rect 2764 11059 2885 11093
rect 2656 11031 2885 11059
<< viali >>
rect 2399 17319 2433 17353
rect 2577 16831 2612 16865
rect 2396 16456 2431 16491
rect 2575 16375 2609 16410
rect 14926 11764 14961 11800
rect 15036 11721 15070 11755
rect 14926 11677 14960 11711
rect 14547 11543 14583 11579
rect 15037 11384 15071 11418
rect 14927 11340 14961 11374
rect 14927 11252 14961 11286
rect 14549 11206 14583 11240
rect 2572 10985 2606 11019
rect 2737 10904 2773 10940
rect 2559 10619 2593 10653
rect 2737 10131 2771 10165
<< metal1 >>
rect 2389 17363 2444 17369
rect 2389 17303 2444 17311
rect 2566 16879 2623 16882
rect 2566 16876 2625 16879
rect 2623 16821 2625 16876
rect 2566 16815 2625 16821
rect 2383 16499 2443 16505
rect 2383 16441 2443 16447
rect 2561 16419 2624 16425
rect 2561 16366 2567 16419
rect 2619 16366 2624 16419
rect 2561 16358 2624 16366
rect 2233 16222 2329 16299
rect 16975 13103 17027 13109
rect 16568 13061 16975 13095
rect 16975 13045 17027 13051
rect 17185 12728 17237 12734
rect 16544 12681 17185 12715
rect 17185 12665 17237 12671
rect 17115 12474 17167 12480
rect 15002 12421 15008 12473
rect 15060 12421 15066 12473
rect 16544 12429 17115 12463
rect 17115 12409 17167 12415
rect 14533 12103 14595 12110
rect 16906 12093 16958 12099
rect 16575 12049 16906 12083
rect 14533 12028 14595 12035
rect 16906 12033 16958 12039
rect 14898 11752 14908 11812
rect 14973 11752 14986 11812
rect 14913 11711 14975 11719
rect 15020 11711 15027 11765
rect 15079 11711 15086 11765
rect 14913 11677 14926 11711
rect 14960 11682 14975 11711
rect 17044 11698 17096 11704
rect 14960 11677 17044 11682
rect 14913 11654 17044 11677
rect 17044 11631 17096 11637
rect 14531 11533 14540 11595
rect 14592 11533 14598 11595
rect 14934 11483 15143 11484
rect 14930 11468 15143 11483
rect 17255 11483 17308 11489
rect 14930 11456 17255 11468
rect 14930 11440 14993 11456
rect 15115 11440 17255 11456
rect 14930 11381 14962 11440
rect 14915 11374 14973 11381
rect 15021 11374 15027 11428
rect 15080 11374 15087 11428
rect 17255 11418 17308 11424
rect 14915 11340 14927 11374
rect 14961 11340 14973 11374
rect 14915 11330 14973 11340
rect 2340 11241 2374 11268
rect 2309 11081 2405 11241
rect 14533 11196 14540 11256
rect 14592 11196 14599 11256
rect 14903 11240 14915 11298
rect 14976 11240 14988 11298
rect 2561 11032 2619 11038
rect 2561 10967 2619 10973
rect 2726 10956 2783 10962
rect 2726 10883 2783 10889
rect 2553 10662 2608 10669
rect 2605 10610 2608 10662
rect 2553 10603 2608 10610
rect 2727 10174 2781 10181
rect 2727 10115 2781 10122
<< via1 >>
rect 2389 17353 2444 17363
rect 2389 17319 2399 17353
rect 2399 17319 2433 17353
rect 2433 17319 2444 17353
rect 2389 17311 2444 17319
rect 2566 16865 2623 16876
rect 2566 16831 2577 16865
rect 2577 16831 2612 16865
rect 2612 16831 2623 16865
rect 2566 16821 2623 16831
rect 2383 16491 2443 16499
rect 2383 16456 2396 16491
rect 2396 16456 2431 16491
rect 2431 16456 2443 16491
rect 2383 16447 2443 16456
rect 2567 16410 2619 16419
rect 2567 16375 2575 16410
rect 2575 16375 2609 16410
rect 2609 16375 2619 16410
rect 2567 16366 2619 16375
rect 2793 16337 2846 16396
rect 2784 15599 2851 15669
rect 16975 13051 17027 13103
rect 17185 12671 17237 12728
rect 15008 12421 15060 12473
rect 17115 12415 17167 12474
rect 14533 12035 14595 12103
rect 16906 12039 16958 12093
rect 2851 11801 2904 11859
rect 14908 11800 14973 11812
rect 14908 11764 14926 11800
rect 14926 11764 14961 11800
rect 14961 11764 14973 11800
rect 14908 11752 14973 11764
rect 15027 11755 15079 11765
rect 15027 11721 15036 11755
rect 15036 11721 15070 11755
rect 15070 11721 15079 11755
rect 15027 11711 15079 11721
rect 17044 11637 17096 11698
rect 14540 11579 14592 11595
rect 14540 11543 14547 11579
rect 14547 11543 14583 11579
rect 14583 11543 14592 11579
rect 14540 11533 14592 11543
rect 15027 11418 15080 11428
rect 15027 11384 15037 11418
rect 15037 11384 15071 11418
rect 15071 11384 15080 11418
rect 15027 11374 15080 11384
rect 17255 11424 17308 11483
rect 14540 11240 14592 11256
rect 14540 11206 14549 11240
rect 14549 11206 14583 11240
rect 14583 11206 14592 11240
rect 14540 11196 14592 11206
rect 14915 11286 14976 11298
rect 14915 11252 14927 11286
rect 14927 11252 14961 11286
rect 14961 11252 14976 11286
rect 14915 11240 14976 11252
rect 2561 11019 2619 11032
rect 2561 10985 2572 11019
rect 2572 10985 2606 11019
rect 2606 10985 2619 11019
rect 2561 10973 2619 10985
rect 2726 10940 2783 10956
rect 2726 10904 2737 10940
rect 2737 10904 2773 10940
rect 2773 10904 2783 10940
rect 2874 10931 2926 10984
rect 2726 10889 2783 10904
rect 2553 10653 2605 10662
rect 2553 10619 2559 10653
rect 2559 10619 2593 10653
rect 2593 10619 2605 10653
rect 2553 10610 2605 10619
rect 2727 10165 2781 10174
rect 2727 10131 2737 10165
rect 2737 10131 2771 10165
rect 2771 10131 2781 10165
rect 2727 10122 2781 10131
<< metal2 >>
rect 10657 19424 10723 19433
rect 10657 19364 10662 19424
rect 10718 19364 10723 19424
rect 10657 19359 10723 19364
rect 7989 19274 8055 19283
rect 7989 19214 7994 19274
rect 8050 19214 8055 19274
rect 7989 19208 8055 19214
rect 5229 18520 5295 18529
rect 5229 18464 5234 18520
rect 5290 18464 5295 18520
rect 5229 18453 5295 18464
rect 2389 17363 2444 17369
rect 2389 17303 2444 17311
rect 2391 16505 2439 17303
rect 2566 16876 2623 16882
rect 2566 16647 2623 16821
rect 2383 16499 2443 16505
rect 5234 16471 5290 18453
rect 7994 16825 8050 19208
rect 10662 16715 10718 19359
rect 11977 18224 12045 18233
rect 11977 18164 11982 18224
rect 12038 18164 12045 18224
rect 11977 18158 12045 18164
rect 2383 16441 2443 16447
rect 2793 16396 2846 16402
rect 2793 16331 2846 16337
rect 2796 15675 2842 16331
rect 2784 15669 2851 15675
rect 2784 15593 2851 15599
rect 11982 13151 12038 18158
rect 11982 13086 12038 13095
rect 15002 12421 15008 12473
rect 15060 12421 15066 12473
rect 14533 12103 14595 12110
rect 14533 12028 14595 12035
rect 2847 11859 2909 11871
rect 2847 11801 2851 11859
rect 2904 11801 2909 11859
rect 2847 11785 2909 11801
rect 2556 11032 2623 11047
rect 2556 10973 2561 11032
rect 2619 10973 2623 11032
rect 2556 10967 2623 10973
rect 2874 10990 2903 11785
rect 14548 11595 14582 12028
rect 14900 11752 14908 11812
rect 14973 11752 14986 11812
rect 15020 11765 15063 12421
rect 14531 11533 14540 11595
rect 14592 11533 14598 11595
rect 14549 11256 14582 11533
rect 14926 11298 14964 11752
rect 15020 11711 15027 11765
rect 15079 11711 15086 11765
rect 15037 11428 15070 11711
rect 15021 11374 15027 11428
rect 15080 11374 15087 11428
rect 14533 11196 14540 11256
rect 14592 11196 14599 11256
rect 14903 11240 14915 11298
rect 14976 11240 14988 11298
rect 2874 10984 2926 10990
rect 2567 10669 2610 10967
rect 2726 10956 2783 10962
rect 2874 10924 2926 10931
rect 2726 10883 2783 10889
rect 2553 10662 2610 10669
rect 2605 10617 2610 10662
rect 2553 10604 2605 10610
rect 2737 10181 2772 10883
rect 2727 10174 2781 10181
rect 2727 10115 2781 10122
rect 16846 9072 16876 21510
rect 16916 12099 16946 21515
rect 16986 13109 17016 21515
rect 16975 13103 17027 13109
rect 16975 13045 17027 13051
rect 16906 12093 16958 12099
rect 16906 12033 16958 12039
rect 16916 9077 16946 12033
rect 16986 9077 17016 13045
rect 17056 11704 17086 21514
rect 17126 12480 17156 21513
rect 17196 12734 17226 21509
rect 17185 12728 17237 12734
rect 17185 12665 17237 12671
rect 17115 12474 17167 12480
rect 17115 12409 17167 12415
rect 17044 11698 17096 11704
rect 17044 11631 17096 11637
rect 17056 9076 17086 11631
rect 17126 9075 17156 12409
rect 17196 9071 17226 12665
rect 17266 11489 17296 21514
rect 17255 11483 17308 11489
rect 17255 11418 17308 11424
rect 17266 9076 17296 11418
<< via2 >>
rect 10662 19364 10718 19424
rect 7994 19214 8050 19274
rect 5234 18464 5290 18520
rect 11982 18164 12038 18224
rect 11982 13095 12038 13151
<< metal3 >>
rect 1037 20714 34034 20774
rect 1037 20564 34034 20624
rect 1037 20414 34034 20474
rect 1037 20264 34034 20324
rect 1037 20114 34034 20174
rect 1037 19964 34034 20024
rect 1037 19814 34034 19874
rect 1037 19664 34034 19724
rect 1037 19514 34034 19574
rect 10657 19424 10723 19433
rect 1037 19364 10662 19424
rect 10718 19364 34034 19424
rect 10657 19359 10723 19364
rect 7989 19274 8055 19283
rect 1037 19214 7994 19274
rect 8050 19214 34034 19274
rect 7989 19208 8055 19214
rect 1037 19064 34034 19124
rect 1037 18914 34034 18974
rect 1037 18764 34034 18824
rect 1037 18614 34034 18674
rect 5229 18524 5295 18529
rect 1037 18520 34034 18524
rect 1037 18464 5234 18520
rect 5290 18464 34034 18520
rect 5229 18453 5295 18464
rect 1037 18314 34034 18374
rect 11977 18224 12045 18233
rect 1037 18164 11982 18224
rect 12038 18164 34034 18224
rect 11977 18158 12045 18164
use filter_p_m_fin  filter_p_m_fin_0
timestamp 1647909829
transform 1 0 5620 0 1 2680
box -5284 -10468 28186 6398
use multiplier  multiplier_1 ~/cochlea_latest/fossi_cochlea/mag/Switched_Caps
timestamp 1647558825
transform -1 0 2517 0 -1 17227
box -426 -152 472 480
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1 ~/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1647912899
transform 0 -1 2825 1 0 16295
box -38 -48 314 592
use mux  mux_1
timestamp 1647510647
transform 0 -1 14945 1 0 11300
box -118 -152 220 422
use mux  mux_0
timestamp 1647510647
transform 0 -1 14944 1 0 11637
box -118 -152 220 422
use filter_clkgen  filter_clkgen_0 ~/cochlea_latest/fossi_cochlea/mag/clkgen
timestamp 1647878126
transform 1 0 15039 0 1 11191
box -1895 666 1540 2096
use lo_gen  lo_gen_0
timestamp 1647915447
transform 1 0 1260 0 1 9106
box 0 1500 10882 7765
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1647912899
transform 0 1 2357 -1 0 11099
box -38 -48 314 592
use multiplier  multiplier_0
timestamp 1647558825
transform 1 0 2653 0 1 10257
box -426 -152 472 480
use filter_p_m_fin  filter_p_m_fin_1
timestamp 1647909829
transform 1 0 5620 0 -1 26676
box -5284 -10468 28186 6398
<< labels >>
rlabel metal2 17283 9078 17283 9078 1 thresh_m
rlabel metal2 17071 9078 17071 9078 3 thresh_p
rlabel metal2 16862 9078 16862 9078 1 VDD
rlabel metal2 16930 9078 16930 9078 1 phi1
rlabel metal2 17001 9078 17001 9078 1 phi2
rlabel metal2 17139 9078 17139 9078 1 phi1b
rlabel metal2 17211 9078 17211 9078 1 phi2b
rlabel metal1 16579 13078 16579 13078 3 phi2
rlabel metal1 16557 12699 16557 12699 3 phi2b
rlabel metal1 16557 12447 16557 12447 3 phi1b
rlabel metal1 16579 12066 16579 12066 3 phi1
<< end >>
