** sch_path: /local_disk/fossi_cochlea/xschem/Switched_Caps/mim_cap_stacked_3pF.sch
.subckt mim_cap_stacked_3pF sig ref
*.PININFO sig:B ref:B
XC1 sig ref sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=8 m=8
XC2 ref sig sky130_fd_pr__cap_mim_m3_2 W=10 L=10 VM=8 m=8
.ends
.end
