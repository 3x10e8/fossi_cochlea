VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO analog_core_I
  CLASS BLOCK ;
  FOREIGN analog_core_I ;
  ORIGIN 0.000 2.450 ;
  SIZE 2038.520 BY 187.340 ;
  PIN fb1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.390 -2.455 25.670 -2.445 ;
    END
  END fb1[0]
  PIN fb1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 279.310 -2.455 279.590 -2.445 ;
    END
  END fb1[1]
  PIN fb1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 533.230 -2.455 533.510 -2.445 ;
    END
  END fb1[2]
  PIN fb1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.150 -2.455 787.430 -2.445 ;
    END
  END fb1[3]
  PIN fb1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1041.070 -2.455 1041.350 -2.445 ;
    END
  END fb1[4]
  PIN fb1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1294.990 -2.455 1295.270 -2.445 ;
    END
  END fb1[5]
  PIN fb1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1548.910 -2.455 1549.190 -2.445 ;
    END
  END fb1[6]
  PIN fb1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1802.830 -2.455 1803.110 -2.445 ;
    END
  END fb1[7]
  PIN cclk[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.710 -2.455 67.990 -2.445 ;
    END
  END cclk[0]
  PIN cclk[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 321.630 -2.455 321.910 -2.445 ;
    END
  END cclk[1]
  PIN cclk[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 575.550 -2.455 575.830 -2.445 ;
    END
  END cclk[2]
  PIN cclk[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.470 -2.455 829.750 -2.445 ;
    END
  END cclk[3]
  PIN cclk[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1083.390 -2.455 1083.670 -2.445 ;
    END
  END cclk[4]
  PIN cclk[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1337.310 -2.455 1337.590 -2.445 ;
    END
  END cclk[5]
  PIN cclk[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1591.230 -2.455 1591.510 -2.445 ;
    END
  END cclk[6]
  PIN cclk[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.150 -2.455 1845.430 -2.445 ;
    END
  END cclk[7]
  PIN div2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.030 -2.455 110.310 -2.445 ;
    END
  END div2[0]
  PIN div2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 363.950 -2.455 364.230 -2.445 ;
    END
  END div2[1]
  PIN div2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 617.870 -2.455 618.150 -2.445 ;
    END
  END div2[2]
  PIN div2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 871.790 -2.455 872.070 -2.445 ;
    END
  END div2[3]
  PIN div2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1125.710 -2.455 1125.990 -2.445 ;
    END
  END div2[4]
  PIN div2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1379.630 -2.455 1379.910 -2.445 ;
    END
  END div2[5]
  PIN div2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1633.550 -2.455 1633.830 -2.445 ;
    END
  END div2[6]
  PIN div2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1887.470 -2.455 1887.750 -2.445 ;
    END
  END div2[7]
  PIN high_buf[0]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 152.350 -2.455 152.630 -2.445 ;
    END
  END high_buf[0]
  PIN high_buf[1]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 406.270 -2.455 406.550 -2.445 ;
    END
  END high_buf[1]
  PIN high_buf[2]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 660.190 -2.455 660.470 -2.445 ;
    END
  END high_buf[2]
  PIN high_buf[3]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 914.110 -2.455 914.390 -2.445 ;
    END
  END high_buf[3]
  PIN high_buf[4]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.030 -2.455 1168.310 -2.445 ;
    END
  END high_buf[4]
  PIN high_buf[5]
    DIRECTION OUTPUT ;
    PORT