magic
tech sky130A
magscale 1 2
timestamp 1654741520
<< metal3 >>
rect -710 2224 -388 2354
rect -710 -180 -677 2224
rect -419 1808 -388 2224
rect -44 2048 276 2354
rect -68 2046 276 2048
rect 824 2046 1144 2354
rect 1692 2048 2012 2354
rect 2356 2224 2678 2354
rect 1692 2046 2036 2048
rect -68 1808 2036 2046
rect 2356 1808 2387 2224
rect -419 1485 2387 1808
rect -419 461 -388 1485
rect -68 461 2036 1485
rect 2356 461 2387 1485
rect -419 138 2387 461
rect -419 -180 -388 138
rect -68 -58 2036 138
rect -68 -60 276 -58
rect -710 -366 -388 -180
rect -44 -366 276 -60
rect 824 -366 1144 -58
rect 1692 -60 2036 -58
rect 1692 -366 2012 -60
rect 2356 -180 2387 138
rect 2645 -180 2678 2224
rect 2356 -366 2678 -180
<< via3 >>
rect -677 -180 -419 2224
rect 2387 -180 2645 2224
<< mimcap >>
rect -16 1786 1984 1994
rect -16 202 192 1786
rect 336 1066 912 1642
rect 1056 1066 1632 1642
rect 336 346 912 922
rect 1056 346 1632 922
rect 1776 202 1984 1786
rect -16 -6 1984 202
<< mimcapcontact >>
rect 192 1642 1776 1786
rect 192 1066 336 1642
rect 912 1066 1056 1642
rect 1632 1066 1776 1642
rect 192 922 1776 1066
rect 192 346 336 922
rect 912 346 1056 922
rect 1632 346 1776 922
rect 192 202 1776 346
<< metal4 >>
rect -685 2224 -412 2354
rect -685 2168 -684 2224
rect 36 2022 196 2354
rect 904 2022 1064 2354
rect 1772 2022 1932 2354
rect 2379 2224 2652 2354
rect 2379 2168 2380 2224
rect -44 1786 2012 2022
rect -44 202 192 1786
rect 336 1066 912 1642
rect 1056 1066 1632 1642
rect 336 346 912 922
rect 1056 346 1632 922
rect 1776 202 2012 1786
rect -44 -34 2012 202
rect -684 -366 -411 -180
rect 36 -366 196 -34
rect 904 -366 1064 -34
rect 1772 -366 1932 -34
rect 2380 -366 2653 -180
<< via4 >>
rect -684 -180 -677 2224
rect -677 -180 -419 2224
rect -419 -180 -412 2224
rect 2380 -180 2387 2224
rect 2387 -180 2645 2224
rect 2645 -180 2652 2224
<< mimcap2 >>
rect -16 1812 1984 1994
rect -16 1576 166 1812
rect 402 1576 516 1812
rect 752 1576 866 1812
rect 1102 1576 1216 1812
rect 1452 1576 1566 1812
rect 1802 1576 1984 1812
rect -16 1462 1984 1576
rect -16 1226 166 1462
rect 402 1226 866 1462
rect 1102 1226 1566 1462
rect 1802 1226 1984 1462
rect -16 1112 1984 1226
rect -16 876 166 1112
rect 402 876 516 1112
rect 752 876 866 1112
rect 1102 876 1216 1112
rect 1452 876 1566 1112
rect 1802 876 1984 1112
rect -16 762 1984 876
rect -16 526 166 762
rect 402 526 866 762
rect 1102 526 1566 762
rect 1802 526 1984 762
rect -16 412 1984 526
rect -16 176 166 412
rect 402 176 516 412
rect 752 176 866 412
rect 1102 176 1216 412
rect 1452 176 1566 412
rect 1802 176 1984 412
rect -16 -6 1984 176
<< mimcap2contact >>
rect 166 1576 402 1812
rect 516 1576 752 1812
rect 866 1576 1102 1812
rect 1216 1576 1452 1812
rect 1566 1576 1802 1812
rect 166 1226 402 1462
rect 866 1226 1102 1462
rect 1566 1226 1802 1462
rect 166 876 402 1112
rect 516 876 752 1112
rect 866 876 1102 1112
rect 1216 876 1452 1112
rect 1566 876 1802 1112
rect 166 526 402 762
rect 866 526 1102 762
rect 1566 526 1802 762
rect 166 176 402 412
rect 516 176 752 412
rect 866 176 1102 412
rect 1216 176 1452 412
rect 1566 176 1802 412
<< metal5 >>
rect -708 2224 -388 2354
rect -708 -180 -684 2224
rect -412 1808 -388 2224
rect -44 2048 276 2354
rect -68 2046 276 2048
rect 824 2046 1144 2354
rect 1692 2048 2012 2354
rect 2356 2224 2676 2354
rect 1692 2046 2036 2048
rect -68 1812 2036 2046
rect -68 1808 166 1812
rect -412 1576 166 1808
rect 402 1576 516 1812
rect 752 1576 866 1812
rect 1102 1576 1216 1812
rect 1452 1576 1566 1812
rect 1802 1808 2036 1812
rect 2356 1808 2380 2224
rect 1802 1576 2380 1808
rect -412 1485 2380 1576
rect -412 461 -388 1485
rect -68 1462 2036 1485
rect -68 1226 166 1462
rect 402 1226 866 1462
rect 1102 1226 1566 1462
rect 1802 1226 2036 1462
rect -68 1112 2036 1226
rect -68 876 166 1112
rect 402 876 516 1112
rect 752 876 866 1112
rect 1102 876 1216 1112
rect 1452 876 1566 1112
rect 1802 876 2036 1112
rect -68 762 2036 876
rect -68 526 166 762
rect 402 526 866 762
rect 1102 526 1566 762
rect 1802 526 2036 762
rect -68 461 2036 526
rect 2356 461 2380 1485
rect -412 412 2380 461
rect -412 176 166 412
rect 402 176 516 412
rect 752 176 866 412
rect 1102 176 1216 412
rect 1452 176 1566 412
rect 1802 176 2380 412
rect -412 138 2380 176
rect -412 -180 -388 138
rect -68 -58 2036 138
rect -68 -60 276 -58
rect -708 -366 -388 -180
rect -44 -366 276 -60
rect 824 -366 1144 -58
rect 1692 -60 2036 -58
rect 1692 -366 2012 -60
rect 2356 -180 2380 138
rect 2652 -180 2676 2224
rect 2356 -366 2676 -180
<< end >>
