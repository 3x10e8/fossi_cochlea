magic
tech sky130A
magscale 1 2
timestamp 1647899285
<< error_p >>
rect 16880 40500 16898 40520
rect 24755 40161 24761 40167
rect 24803 40161 24809 40167
rect 24749 40155 24815 40161
rect 24755 40115 24809 40155
rect 24749 40109 24815 40115
rect 24755 40103 24761 40109
rect 24803 40103 24809 40109
rect 24755 39703 24761 39709
rect 24803 39703 24809 39709
rect 24749 39697 24815 39703
rect 24755 39657 24809 39697
rect 24749 39651 24815 39657
rect 24755 39645 24761 39651
rect 24803 39645 24809 39651
rect 16880 39352 16958 39372
use filter_i_q  filter_i_q_0
array 0 7 33844 0 5 40080
timestamp 1647899285
transform 1 0 -336 0 1 7788
box 336 -7788 33806 31944
<< end >>
