magic
tech sky130A
magscale 1 2
timestamp 1647898595
<< nwell >>
rect 14580 11851 14755 12005
<< locali >>
rect 14927 11592 14959 11593
rect 14927 11462 14961 11592
<< viali >>
rect 14926 11764 14961 11800
rect 15036 11721 15070 11755
rect 14926 11677 14960 11711
rect 14547 11543 14583 11579
rect 15037 11384 15071 11418
rect 14927 11340 14961 11374
rect 14927 11252 14961 11286
rect 14549 11206 14583 11240
<< metal1 >>
rect 16975 13103 17027 13109
rect 16568 13061 16975 13095
rect 16975 13045 17027 13051
rect 17185 12728 17237 12734
rect 16544 12681 17185 12715
rect 17185 12665 17237 12671
rect 17115 12474 17167 12480
rect 15002 12421 15008 12473
rect 15060 12421 15066 12473
rect 16544 12429 17115 12463
rect 17115 12409 17167 12415
rect 14533 12103 14595 12110
rect 16906 12093 16958 12099
rect 16575 12049 16906 12083
rect 14533 12028 14595 12035
rect 16906 12033 16958 12039
rect 14898 11752 14908 11812
rect 14973 11752 14986 11812
rect 14913 11711 14975 11719
rect 15020 11711 15027 11765
rect 15079 11711 15086 11765
rect 14913 11677 14926 11711
rect 14960 11682 14975 11711
rect 17044 11698 17096 11704
rect 14960 11677 17044 11682
rect 14913 11654 17044 11677
rect 17044 11631 17096 11637
rect 14531 11533 14540 11595
rect 14592 11533 14598 11595
rect 14934 11483 15143 11484
rect 14930 11468 15143 11483
rect 17255 11483 17308 11489
rect 14930 11456 17255 11468
rect 14930 11440 14993 11456
rect 15115 11440 17255 11456
rect 14930 11381 14962 11440
rect 14915 11374 14973 11381
rect 15021 11374 15027 11428
rect 15080 11374 15087 11428
rect 17255 11418 17308 11424
rect 14915 11340 14927 11374
rect 14961 11340 14973 11374
rect 14915 11330 14973 11340
rect 14533 11196 14540 11256
rect 14592 11196 14599 11256
rect 14903 11240 14915 11298
rect 14976 11240 14988 11298
<< via1 >>
rect 16975 13051 17027 13103
rect 17185 12671 17237 12728
rect 15008 12421 15060 12473
rect 17115 12415 17167 12474
rect 14533 12035 14595 12103
rect 16906 12039 16958 12093
rect 14908 11800 14973 11812
rect 14908 11764 14926 11800
rect 14926 11764 14961 11800
rect 14961 11764 14973 11800
rect 14908 11752 14973 11764
rect 15027 11755 15079 11765
rect 15027 11721 15036 11755
rect 15036 11721 15070 11755
rect 15070 11721 15079 11755
rect 15027 11711 15079 11721
rect 17044 11637 17096 11698
rect 14540 11579 14592 11595
rect 14540 11543 14547 11579
rect 14547 11543 14583 11579
rect 14583 11543 14592 11579
rect 14540 11533 14592 11543
rect 15027 11418 15080 11428
rect 15027 11384 15037 11418
rect 15037 11384 15071 11418
rect 15071 11384 15080 11418
rect 15027 11374 15080 11384
rect 17255 11424 17308 11483
rect 14540 11240 14592 11256
rect 14540 11206 14549 11240
rect 14549 11206 14583 11240
rect 14583 11206 14592 11240
rect 14540 11196 14592 11206
rect 14915 11286 14976 11298
rect 14915 11252 14927 11286
rect 14927 11252 14961 11286
rect 14961 11252 14976 11286
rect 14915 11240 14976 11252
<< metal2 >>
rect 15002 12421 15008 12473
rect 15060 12421 15066 12473
rect 14533 12103 14595 12110
rect 14533 12028 14595 12035
rect 14548 11595 14582 12028
rect 14900 11752 14908 11812
rect 14973 11752 14986 11812
rect 15020 11765 15063 12421
rect 14531 11533 14540 11595
rect 14592 11533 14598 11595
rect 14549 11256 14582 11533
rect 14926 11298 14964 11752
rect 15020 11711 15027 11765
rect 15079 11711 15086 11765
rect 15037 11428 15070 11711
rect 15021 11374 15027 11428
rect 15080 11374 15087 11428
rect 14533 11196 14540 11256
rect 14592 11196 14599 11256
rect 14903 11240 14915 11298
rect 14976 11240 14988 11298
rect 16846 9072 16876 15110
rect 16916 12099 16946 15115
rect 16986 13109 17016 15115
rect 16975 13103 17027 13109
rect 16975 13045 17027 13051
rect 16906 12093 16958 12099
rect 16906 12033 16958 12039
rect 16916 9077 16946 12033
rect 16986 9077 17016 13045
rect 17056 11704 17086 15114
rect 17126 12480 17156 15113
rect 17196 12734 17226 15109
rect 17185 12728 17237 12734
rect 17185 12665 17237 12671
rect 17115 12474 17167 12480
rect 17115 12409 17167 12415
rect 17044 11698 17096 11704
rect 17044 11631 17096 11637
rect 17056 9076 17086 11631
rect 17126 9075 17156 12409
rect 17196 9071 17226 12665
rect 17266 11489 17296 15114
rect 17255 11483 17308 11489
rect 17255 11418 17308 11424
rect 17266 9076 17296 11418
use mux  mux_1
timestamp 1647510647
transform 0 -1 14945 1 0 11300
box -118 -152 220 422
use mux  mux_0
timestamp 1647510647
transform 0 -1 14944 1 0 11637
box -118 -152 220 422
use filter_p_m_fin  filter_p_m_fin_1
timestamp 1647895372
transform 1 0 5620 0 -1 21476
box -5284 -10468 28186 6398
use filter_p_m_fin  filter_p_m_fin_0
timestamp 1647895372
transform 1 0 5620 0 1 2680
box -5284 -10468 28186 6398
use filter_clkgen  filter_clkgen_0 ~/cochlea_latest/fossi_cochlea/mag/clkgen
timestamp 1647896663
transform 1 0 15039 0 1 11191
box -1895 666 1540 2096
<< labels >>
rlabel metal2 17283 9078 17283 9078 1 thresh_m
rlabel metal2 17071 9078 17071 9078 3 thresh_p
rlabel metal2 16862 9078 16862 9078 1 VDD
rlabel metal2 16930 9078 16930 9078 1 phi1
rlabel metal2 17001 9078 17001 9078 1 phi2
rlabel metal2 17139 9078 17139 9078 1 phi1b
rlabel metal2 17211 9078 17211 9078 1 phi2b
rlabel metal1 16579 13078 16579 13078 3 phi2
rlabel metal1 16557 12699 16557 12699 3 phi2b
rlabel metal1 16557 12447 16557 12447 3 phi1b
rlabel metal1 16579 12066 16579 12066 3 phi1
<< end >>
