magic
tech sky130B
magscale 1 2
timestamp 1654741520
<< nwell >>
rect -167 428 643 596
<< nmos >>
rect -30 79 0 163
rect 120 79 150 163
rect 237 79 267 163
rect 387 79 417 163
<< pmos >>
rect -30 464 0 548
rect 120 464 150 548
rect 237 464 267 548
rect 387 464 417 548
<< ndiff >>
rect -131 137 -30 163
rect -131 103 -91 137
rect -57 103 -30 137
rect -131 79 -30 103
rect 0 137 120 163
rect 0 103 42 137
rect 78 103 120 137
rect 0 79 120 103
rect 150 137 237 163
rect 150 103 176 137
rect 211 103 237 137
rect 150 79 237 103
rect 267 137 387 163
rect 267 103 309 137
rect 345 103 387 137
rect 267 79 387 103
rect 417 137 518 163
rect 417 103 444 137
rect 478 103 518 137
rect 417 79 518 103
<< pdiff >>
rect -131 524 -30 548
rect -131 490 -91 524
rect -57 490 -30 524
rect -131 464 -30 490
rect 0 524 120 548
rect 0 490 42 524
rect 78 490 120 524
rect 0 464 120 490
rect 150 524 237 548
rect 150 490 176 524
rect 211 490 237 524
rect 150 464 237 490
rect 267 524 387 548
rect 267 490 309 524
rect 345 490 387 524
rect 267 464 387 490
rect 417 524 518 548
rect 417 490 444 524
rect 478 490 518 524
rect 417 464 518 490
<< ndiffc >>
rect -91 103 -57 137
rect 42 103 78 137
rect 176 103 211 137
rect 309 103 345 137
rect 444 103 478 137
<< pdiffc >>
rect -91 490 -57 524
rect 42 490 78 524
rect 176 490 211 524
rect 309 490 345 524
rect 444 490 478 524
<< psubdiff >>
rect 518 137 606 163
rect 518 103 548 137
rect 582 103 606 137
rect 518 79 606 103
<< nsubdiff >>
rect 518 523 607 548
rect 518 489 556 523
rect 590 489 607 523
rect 518 464 607 489
<< psubdiffcont >>
rect 548 103 582 137
<< nsubdiffcont >>
rect 556 489 590 523
<< poly >>
rect -30 548 0 574
rect 120 548 150 574
rect 237 548 267 574
rect 387 548 417 574
rect -30 433 0 464
rect -35 427 0 433
rect 120 433 150 464
rect 237 433 267 464
rect 120 427 155 433
rect 232 427 267 433
rect 387 433 417 464
rect 387 427 422 433
rect -45 417 9 427
rect -45 383 -35 417
rect -1 383 9 417
rect -45 373 9 383
rect 111 417 165 427
rect 111 383 121 417
rect 155 383 165 417
rect 111 373 165 383
rect 222 417 276 427
rect 222 383 232 417
rect 266 383 276 417
rect 222 373 276 383
rect 378 417 432 427
rect 378 383 388 417
rect 422 383 432 417
rect 378 373 432 383
rect -35 367 -1 373
rect 121 367 155 373
rect 232 367 266 373
rect 388 367 422 373
rect 123 325 153 367
rect 390 325 420 367
rect -33 295 420 325
rect -33 253 -3 295
rect 234 253 264 295
rect -35 247 -1 253
rect 121 247 155 253
rect 232 247 266 253
rect 388 247 422 253
rect -45 237 9 247
rect -45 203 -35 237
rect -1 203 9 237
rect -45 193 9 203
rect 111 237 165 247
rect 111 203 121 237
rect 155 203 165 237
rect 111 193 165 203
rect 222 237 276 247
rect 222 203 232 237
rect 266 203 276 237
rect 222 193 276 203
rect 378 237 432 247
rect 378 203 388 237
rect 422 203 432 237
rect 378 193 432 203
rect -35 187 0 193
rect -30 163 0 187
rect 120 187 155 193
rect 232 187 267 193
rect 120 163 150 187
rect 237 163 267 187
rect 387 187 422 193
rect 387 163 417 187
rect -30 53 0 79
rect 120 53 150 79
rect 237 53 267 79
rect 387 53 417 79
<< polycont >>
rect -35 383 -1 417
rect 121 383 155 417
rect 232 383 266 417
rect 388 383 422 417
rect -35 203 -1 237
rect 121 203 155 237
rect 232 203 266 237
rect 388 203 422 237
<< locali >>
rect -99 524 -48 548
rect -99 490 -91 524
rect -57 490 -48 524
rect -99 474 -48 490
rect 34 524 86 548
rect 34 490 42 524
rect 78 490 86 524
rect 34 474 86 490
rect 168 524 219 548
rect 168 490 176 524
rect 211 490 219 524
rect 168 474 219 490
rect 301 524 353 548
rect 301 490 309 524
rect 345 490 353 524
rect 301 474 353 490
rect 435 524 486 548
rect 435 490 444 524
rect 478 490 486 524
rect 435 474 486 490
rect 556 523 590 539
rect 556 473 590 489
rect -35 417 -1 433
rect -35 327 -1 383
rect 121 417 155 433
rect 121 367 155 383
rect 232 417 266 433
rect 232 327 266 383
rect 388 417 422 433
rect 422 383 627 417
rect 388 367 422 383
rect -35 293 422 327
rect -35 237 -1 253
rect -35 187 -1 203
rect 121 237 155 293
rect 121 187 155 203
rect 232 237 266 253
rect 232 187 266 203
rect 388 237 422 293
rect 422 203 618 237
rect 388 187 422 203
rect -99 137 -48 153
rect -99 103 -91 137
rect -57 103 -48 137
rect -99 79 -48 103
rect 34 137 86 153
rect 34 103 42 137
rect 78 103 86 137
rect 34 79 86 103
rect 167 137 220 153
rect 167 103 176 137
rect 211 103 220 137
rect 167 79 220 103
rect 301 137 353 153
rect 301 103 309 137
rect 345 103 353 137
rect 301 79 353 103
rect 434 137 487 153
rect 434 103 444 137
rect 478 103 487 137
rect 434 79 487 103
rect 548 137 582 153
rect 548 87 582 103
rect -92 45 -58 79
rect 444 45 478 79
rect -92 11 478 45
<< viali >>
rect -91 490 -57 524
rect 42 490 78 524
rect 176 490 211 524
rect 309 490 345 524
rect 444 490 478 524
rect 556 489 590 523
rect -91 103 -57 137
rect 42 103 78 137
rect 176 103 211 137
rect 309 103 345 137
rect 444 103 478 137
rect 548 103 582 137
<< metal1 >>
rect -224 613 685 681
rect -99 534 -47 540
rect -99 475 -47 482
rect 34 533 86 539
rect 34 475 86 481
rect 167 534 220 540
rect 167 475 220 481
rect 301 533 353 539
rect 301 475 353 481
rect 434 534 487 540
rect 556 530 590 613
rect 549 523 597 530
rect 549 489 556 523
rect 590 489 597 523
rect 549 483 597 489
rect 434 475 487 481
rect 556 477 590 483
rect 42 474 78 475
rect 309 474 345 475
rect 34 379 86 385
rect 34 321 86 327
rect 295 207 301 259
rect 353 207 359 259
rect -100 146 -48 152
rect -103 103 -100 131
rect -100 88 -48 94
rect 34 146 86 152
rect 34 88 86 94
rect 167 146 220 153
rect 167 88 220 94
rect 301 146 353 152
rect 301 88 353 94
rect 434 146 487 153
rect 540 137 590 150
rect 540 103 548 137
rect 582 103 590 137
rect 540 95 590 103
rect 434 88 487 94
rect 548 -11 582 95
rect -224 -79 685 -11
<< via1 >>
rect -99 524 -47 534
rect -99 490 -91 524
rect -91 490 -57 524
rect -57 490 -47 524
rect -99 482 -47 490
rect 34 524 86 533
rect 34 490 42 524
rect 42 490 78 524
rect 78 490 86 524
rect 34 481 86 490
rect 167 524 220 534
rect 167 490 176 524
rect 176 490 211 524
rect 211 490 220 524
rect 167 481 220 490
rect 301 524 353 533
rect 301 490 309 524
rect 309 490 345 524
rect 345 490 353 524
rect 301 481 353 490
rect 434 524 487 534
rect 434 490 444 524
rect 444 490 478 524
rect 478 490 487 524
rect 434 481 487 490
rect 34 327 86 379
rect 301 207 353 259
rect -100 137 -48 146
rect -100 103 -91 137
rect -91 103 -57 137
rect -57 103 -48 137
rect -100 94 -48 103
rect 34 137 86 146
rect 34 103 42 137
rect 42 103 78 137
rect 78 103 86 137
rect 34 94 86 103
rect 167 137 220 146
rect 167 103 176 137
rect 176 103 211 137
rect 211 103 220 137
rect 167 94 220 103
rect 301 137 353 146
rect 301 103 309 137
rect 309 103 345 137
rect 345 103 353 137
rect 301 94 353 103
rect 434 137 487 146
rect 434 103 444 137
rect 444 103 478 137
rect 478 103 487 137
rect 434 94 487 103
<< metal2 >>
rect -99 534 -47 540
rect -99 476 -47 482
rect 34 533 86 539
rect -91 152 -57 476
rect 34 475 86 481
rect 167 534 220 540
rect 167 475 220 481
rect 301 533 353 539
rect 301 475 353 481
rect 434 534 487 540
rect 434 475 487 481
rect 43 385 77 475
rect 34 379 86 385
rect 34 321 86 327
rect 43 152 77 321
rect 176 291 211 475
rect 167 227 219 291
rect 310 259 344 475
rect 176 153 211 227
rect 295 207 301 259
rect 353 207 359 259
rect -100 146 -48 152
rect -100 88 -48 94
rect 34 146 86 152
rect 34 88 86 94
rect 167 146 220 153
rect 310 152 344 207
rect 444 153 478 475
rect 167 88 220 94
rect 301 146 353 152
rect 301 88 353 94
rect 434 146 487 153
rect 434 88 487 94
<< labels >>
rlabel metal1 -224 649 -224 649 7 VDD
rlabel metal1 -224 -43 -224 -43 7 GND
flabel metal2 34 321 86 385 0 FreeSans 160 0 0 0 out1
flabel metal2 295 207 359 259 0 FreeSans 160 0 0 0 out2
<< end >>
