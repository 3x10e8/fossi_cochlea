magic
tech sky130A
magscale 1 2
timestamp 1654479364
<< nwell >>
rect 1715 1373 2125 1605
<< nmos >>
rect 1230 1130 1260 1250
rect 1316 1130 1346 1250
rect 1403 1130 1433 1250
rect 1489 1130 1519 1250
rect 1576 1130 1606 1250
rect 1662 1130 1692 1250
rect 1749 1130 1779 1250
rect 1835 1130 1865 1250
rect 1922 1130 1952 1250
rect 2008 1130 2038 1250
rect 2095 1130 2125 1250
rect 2181 1130 2211 1250
rect 2268 1130 2298 1250
rect 2354 1130 2384 1250
rect 2441 1130 2471 1250
rect 2527 1130 2557 1250
rect 1230 690 1260 810
rect 1316 690 1346 810
rect 1403 690 1433 810
rect 1489 690 1519 810
rect 1576 690 1606 810
rect 1662 690 1692 810
rect 1749 690 1779 810
rect 1835 690 1865 810
rect 1922 690 1952 810
rect 2008 690 2038 810
rect 2095 690 2125 810
rect 2181 690 2211 810
rect 2268 690 2298 810
rect 2354 690 2384 810
rect 2441 690 2471 810
rect 2527 690 2557 810
<< pmos >>
rect 1829 1445 1859 1529
rect 1930 1445 1960 1529
<< ndiff >>
rect 1173 1238 1230 1250
rect 1173 1204 1185 1238
rect 1219 1204 1230 1238
rect 1173 1130 1230 1204
rect 1260 1176 1316 1250
rect 1260 1142 1271 1176
rect 1305 1142 1316 1176
rect 1260 1130 1316 1142
rect 1346 1238 1403 1250
rect 1346 1204 1358 1238
rect 1392 1204 1403 1238
rect 1346 1130 1403 1204
rect 1433 1176 1489 1250
rect 1433 1142 1444 1176
rect 1478 1142 1489 1176
rect 1433 1130 1489 1142
rect 1519 1238 1576 1250
rect 1519 1204 1531 1238
rect 1565 1204 1576 1238
rect 1519 1130 1576 1204
rect 1606 1176 1662 1250
rect 1606 1142 1617 1176
rect 1651 1142 1662 1176
rect 1606 1130 1662 1142
rect 1692 1238 1749 1250
rect 1692 1204 1704 1238
rect 1738 1204 1749 1238
rect 1692 1130 1749 1204
rect 1779 1176 1835 1250
rect 1779 1142 1790 1176
rect 1824 1142 1835 1176
rect 1779 1130 1835 1142
rect 1865 1238 1922 1250
rect 1865 1204 1877 1238
rect 1911 1204 1922 1238
rect 1865 1130 1922 1204
rect 1952 1176 2008 1250
rect 1952 1142 1963 1176
rect 1997 1142 2008 1176
rect 1952 1130 2008 1142
rect 2038 1238 2095 1250
rect 2038 1204 2050 1238
rect 2084 1204 2095 1238
rect 2038 1130 2095 1204
rect 2125 1176 2181 1250
rect 2125 1142 2136 1176
rect 2170 1142 2181 1176
rect 2125 1130 2181 1142
rect 2211 1238 2268 1250
rect 2211 1204 2223 1238
rect 2257 1204 2268 1238
rect 2211 1130 2268 1204
rect 2298 1176 2354 1250
rect 2298 1142 2309 1176
rect 2343 1142 2354 1176
rect 2298 1130 2354 1142
rect 2384 1238 2441 1250
rect 2384 1204 2396 1238
rect 2430 1204 2441 1238
rect 2384 1130 2441 1204
rect 2471 1176 2527 1250
rect 2471 1142 2482 1176
rect 2516 1142 2527 1176
rect 2471 1130 2527 1142
rect 2557 1238 2614 1250
rect 2557 1204 2569 1238
rect 2603 1204 2614 1238
rect 2557 1130 2614 1204
rect 1170 798 1230 810
rect 1170 764 1185 798
rect 1219 764 1230 798
rect 1170 690 1230 764
rect 1260 736 1316 810
rect 1260 702 1271 736
rect 1305 702 1316 736
rect 1260 690 1316 702
rect 1346 798 1403 810
rect 1346 764 1358 798
rect 1392 764 1403 798
rect 1346 690 1403 764
rect 1433 736 1489 810
rect 1433 702 1444 736
rect 1478 702 1489 736
rect 1433 690 1489 702
rect 1519 798 1576 810
rect 1519 764 1531 798
rect 1565 764 1576 798
rect 1519 690 1576 764
rect 1606 736 1662 810
rect 1606 702 1617 736
rect 1651 702 1662 736
rect 1606 690 1662 702
rect 1692 798 1749 810
rect 1692 764 1704 798
rect 1738 764 1749 798
rect 1692 690 1749 764
rect 1779 736 1835 810
rect 1779 702 1790 736
rect 1824 702 1835 736
rect 1779 690 1835 702
rect 1865 798 1922 810
rect 1865 764 1877 798
rect 1911 764 1922 798
rect 1865 690 1922 764
rect 1952 736 2008 810
rect 1952 702 1963 736
rect 1997 702 2008 736
rect 1952 690 2008 702
rect 2038 798 2095 810
rect 2038 764 2050 798
rect 2084 764 2095 798
rect 2038 690 2095 764
rect 2125 736 2181 810
rect 2125 702 2136 736
rect 2170 702 2181 736
rect 2125 690 2181 702
rect 2211 798 2268 810
rect 2211 764 2223 798
rect 2257 764 2268 798
rect 2211 690 2268 764
rect 2298 736 2354 810
rect 2298 702 2309 736
rect 2343 702 2354 736
rect 2298 690 2354 702
rect 2384 798 2441 810
rect 2384 764 2396 798
rect 2430 764 2441 798
rect 2384 690 2441 764
rect 2471 736 2527 810
rect 2471 702 2482 736
rect 2516 702 2527 736
rect 2471 690 2527 702
rect 2557 798 2618 810
rect 2557 764 2569 798
rect 2603 764 2618 798
rect 2557 690 2618 764
<< pdiff >>
rect 1763 1505 1829 1529
rect 1763 1471 1783 1505
rect 1817 1471 1829 1505
rect 1763 1445 1829 1471
rect 1859 1505 1930 1529
rect 1859 1471 1877 1505
rect 1911 1471 1930 1505
rect 1859 1445 1930 1471
rect 1960 1505 2020 1529
rect 1960 1471 1975 1505
rect 2009 1471 2020 1505
rect 1960 1445 2020 1471
<< ndiffc >>
rect 1185 1204 1219 1238
rect 1271 1142 1305 1176
rect 1358 1204 1392 1238
rect 1444 1142 1478 1176
rect 1531 1204 1565 1238
rect 1617 1142 1651 1176
rect 1704 1204 1738 1238
rect 1790 1142 1824 1176
rect 1877 1204 1911 1238
rect 1963 1142 1997 1176
rect 2050 1204 2084 1238
rect 2136 1142 2170 1176
rect 2223 1204 2257 1238
rect 2309 1142 2343 1176
rect 2396 1204 2430 1238
rect 2482 1142 2516 1176
rect 2569 1204 2603 1238
rect 1185 764 1219 798
rect 1271 702 1305 736
rect 1358 764 1392 798
rect 1444 702 1478 736
rect 1531 764 1565 798
rect 1617 702 1651 736
rect 1704 764 1738 798
rect 1790 702 1824 736
rect 1877 764 1911 798
rect 1963 702 1997 736
rect 2050 764 2084 798
rect 2136 702 2170 736
rect 2223 764 2257 798
rect 2309 702 2343 736
rect 2396 764 2430 798
rect 2482 702 2516 736
rect 2569 764 2603 798
<< pdiffc >>
rect 1783 1471 1817 1505
rect 1877 1471 1911 1505
rect 1975 1471 2009 1505
<< psubdiff >>
rect 1112 777 1170 810
rect 1112 743 1113 777
rect 1147 743 1170 777
rect 1112 690 1170 743
rect 2618 783 2691 810
rect 2618 749 2647 783
rect 2681 749 2691 783
rect 2618 690 2691 749
<< nsubdiff >>
rect 2020 1505 2089 1529
rect 2020 1471 2043 1505
rect 2077 1471 2089 1505
rect 2020 1445 2089 1471
<< psubdiffcont >>
rect 1113 743 1147 777
rect 2647 749 2681 783
<< nsubdiffcont >>
rect 2043 1471 2077 1505
<< poly >>
rect 1817 1610 1871 1620
rect 1811 1576 1827 1610
rect 1861 1576 1877 1610
rect 1817 1566 1871 1576
rect 1829 1529 1859 1566
rect 1930 1529 1960 1555
rect 1829 1419 1859 1445
rect 1930 1408 1960 1445
rect 1918 1398 1972 1408
rect 1912 1364 1928 1398
rect 1962 1364 1978 1398
rect 1918 1354 1972 1364
rect 1230 1250 1260 1276
rect 1316 1250 1346 1276
rect 1403 1250 1433 1276
rect 1489 1250 1519 1276
rect 1576 1250 1606 1276
rect 1662 1250 1692 1276
rect 1749 1250 1779 1276
rect 1835 1250 1865 1276
rect 1922 1250 1952 1276
rect 2008 1250 2038 1276
rect 2095 1250 2125 1276
rect 2181 1250 2211 1276
rect 2268 1250 2298 1276
rect 2354 1250 2384 1276
rect 2441 1250 2471 1276
rect 2527 1250 2557 1276
rect 1230 1104 1260 1130
rect 1316 1104 1346 1130
rect 1403 1104 1433 1130
rect 1489 1104 1519 1130
rect 1576 1104 1606 1130
rect 1662 1104 1692 1130
rect 1749 1104 1779 1130
rect 1835 1104 1865 1130
rect 1230 1084 1865 1104
rect 1230 1074 1245 1084
rect 1235 1050 1245 1074
rect 1280 1074 1865 1084
rect 1922 1104 1952 1130
rect 2008 1104 2038 1130
rect 2095 1104 2125 1130
rect 2181 1104 2211 1130
rect 2268 1104 2298 1130
rect 2354 1104 2384 1130
rect 2441 1104 2471 1130
rect 2527 1104 2557 1130
rect 1922 1074 2557 1104
rect 1280 1050 1290 1074
rect 1235 1034 1290 1050
rect 1778 1040 1788 1074
rect 1823 1040 1833 1074
rect 1778 1024 1833 1040
rect 1922 982 1952 1074
rect 1785 952 1952 982
rect 1235 890 1290 906
rect 1235 866 1245 890
rect 1230 856 1245 866
rect 1280 866 1290 890
rect 1785 866 1815 952
rect 1977 900 2032 916
rect 1977 866 1987 900
rect 2022 866 2032 900
rect 1280 856 1865 866
rect 1230 836 1865 856
rect 1230 810 1260 836
rect 1316 810 1346 836
rect 1403 810 1433 836
rect 1489 810 1519 836
rect 1576 810 1606 836
rect 1662 810 1692 836
rect 1749 810 1779 836
rect 1835 810 1865 836
rect 1922 836 2557 866
rect 1922 810 1952 836
rect 2008 810 2038 836
rect 2095 810 2125 836
rect 2181 810 2211 836
rect 2268 810 2298 836
rect 2354 810 2384 836
rect 2441 810 2471 836
rect 2527 810 2557 836
rect 1230 664 1260 690
rect 1316 664 1346 690
rect 1403 664 1433 690
rect 1489 664 1519 690
rect 1576 664 1606 690
rect 1662 664 1692 690
rect 1749 664 1779 690
rect 1835 664 1865 690
rect 1922 664 1952 690
rect 2008 664 2038 690
rect 2095 664 2125 690
rect 2181 664 2211 690
rect 2268 664 2298 690
rect 2354 664 2384 690
rect 2441 664 2471 690
rect 2527 664 2557 690
<< polycont >>
rect 1827 1576 1861 1610
rect 1928 1364 1962 1398
rect 1245 1050 1280 1084
rect 1788 1040 1823 1074
rect 1245 856 1280 890
rect 1987 866 2022 900
<< locali >>
rect 1811 1576 1827 1610
rect 1861 1576 2170 1610
rect 1783 1505 1817 1521
rect 1783 1398 1817 1471
rect 1877 1505 1911 1521
rect 1877 1455 1911 1471
rect 1975 1505 2009 1576
rect 1975 1455 2009 1471
rect 2043 1505 2077 1521
rect 2043 1455 2077 1471
rect 1783 1364 1928 1398
rect 1962 1364 1978 1398
rect 1185 1238 1219 1254
rect 1185 1188 1219 1204
rect 1358 1238 1392 1254
rect 1271 1176 1305 1192
rect 1358 1188 1392 1204
rect 1531 1238 1565 1254
rect 1271 1126 1305 1142
rect 1444 1176 1478 1192
rect 1531 1188 1565 1204
rect 1704 1238 1738 1254
rect 1444 1126 1478 1142
rect 1617 1176 1651 1192
rect 1704 1188 1738 1204
rect 1617 1126 1651 1142
rect 1790 1176 1824 1364
rect 1877 1238 1911 1254
rect 1877 1188 1911 1204
rect 2050 1238 2084 1254
rect 1790 1126 1824 1142
rect 1963 1176 1997 1192
rect 2050 1188 2084 1204
rect 1963 1126 1997 1142
rect 2136 1176 2170 1576
rect 2223 1238 2257 1254
rect 2223 1188 2257 1204
rect 2396 1238 2430 1254
rect 2136 1126 2170 1142
rect 2309 1176 2343 1192
rect 2396 1188 2430 1204
rect 2569 1238 2603 1254
rect 2309 1126 2343 1142
rect 2482 1176 2516 1192
rect 2569 1188 2603 1204
rect 2482 1126 2516 1142
rect 1229 1050 1245 1084
rect 1280 1050 1296 1084
rect 1772 1040 1788 1074
rect 1823 1040 1839 1074
rect 1788 900 1823 1040
rect 1229 856 1245 890
rect 1280 856 1296 890
rect 1788 866 1987 900
rect 2022 866 2038 900
rect 1185 798 1219 814
rect 1113 777 1147 793
rect 1185 748 1219 764
rect 1358 798 1392 814
rect 1113 727 1147 743
rect 1271 736 1305 752
rect 1358 748 1392 764
rect 1531 798 1565 814
rect 1271 686 1305 702
rect 1444 736 1478 752
rect 1531 748 1565 764
rect 1704 798 1738 814
rect 1444 686 1478 702
rect 1617 736 1651 752
rect 1704 748 1738 764
rect 1877 798 1911 814
rect 1617 686 1651 702
rect 1790 736 1824 752
rect 1877 748 1911 764
rect 2050 798 2084 814
rect 1790 686 1824 702
rect 1963 736 1997 752
rect 2050 748 2084 764
rect 2223 798 2257 814
rect 1963 686 1997 702
rect 2136 736 2170 752
rect 2223 748 2257 764
rect 2396 798 2430 814
rect 2136 686 2170 702
rect 2309 736 2343 752
rect 2396 748 2430 764
rect 2569 798 2603 814
rect 2309 686 2343 702
rect 2482 736 2516 752
rect 2569 748 2603 764
rect 2647 783 2681 799
rect 2647 733 2681 749
rect 2482 686 2516 702
<< viali >>
rect 1877 1471 1911 1505
rect 2043 1471 2077 1505
rect 1185 1204 1219 1238
rect 1358 1204 1392 1238
rect 1531 1204 1565 1238
rect 1271 1142 1305 1176
rect 1704 1204 1738 1238
rect 1444 1142 1478 1176
rect 1617 1142 1651 1176
rect 1877 1204 1911 1238
rect 2050 1204 2084 1238
rect 1790 1142 1824 1176
rect 1963 1142 1997 1176
rect 2223 1204 2257 1238
rect 2396 1204 2430 1238
rect 2136 1142 2170 1176
rect 2569 1204 2603 1238
rect 2309 1142 2343 1176
rect 2482 1142 2516 1176
rect 1245 1050 1280 1084
rect 1245 856 1280 890
rect 1113 743 1147 777
rect 1185 764 1219 798
rect 1358 764 1392 798
rect 1531 764 1565 798
rect 1271 702 1305 736
rect 1704 764 1738 798
rect 1444 702 1478 736
rect 1877 764 1911 798
rect 1617 702 1651 736
rect 2050 764 2084 798
rect 1790 702 1824 736
rect 2223 764 2257 798
rect 1963 702 1997 736
rect 2396 764 2430 798
rect 2136 702 2170 736
rect 2569 764 2603 798
rect 2309 702 2343 736
rect 2647 749 2681 783
rect 2482 702 2516 736
<< metal1 >>
rect 1050 1690 2782 1760
rect 1910 1517 1998 1690
rect 1871 1505 1998 1517
rect 2037 1505 2083 1511
rect 1871 1471 1877 1505
rect 1911 1471 2043 1505
rect 2077 1471 2089 1505
rect 1871 1465 1917 1471
rect 2037 1465 2083 1471
rect 1877 1244 1911 1465
rect 1173 1238 2615 1244
rect 1173 1204 1185 1238
rect 1219 1212 1358 1238
rect 1219 1204 1231 1212
rect 1173 1198 1231 1204
rect 1346 1204 1358 1212
rect 1392 1212 1531 1238
rect 1392 1204 1404 1212
rect 1346 1198 1404 1204
rect 1519 1204 1531 1212
rect 1565 1212 1704 1238
rect 1565 1204 1577 1212
rect 1519 1198 1577 1204
rect 1692 1204 1704 1212
rect 1738 1212 1877 1238
rect 1738 1204 1750 1212
rect 1692 1198 1750 1204
rect 1865 1204 1877 1212
rect 1911 1212 2050 1238
rect 1911 1204 1923 1212
rect 1865 1198 1923 1204
rect 2038 1204 2050 1212
rect 2084 1212 2223 1238
rect 2084 1204 2096 1212
rect 2038 1198 2096 1204
rect 2211 1204 2223 1212
rect 2257 1212 2396 1238
rect 2257 1204 2269 1212
rect 2211 1198 2269 1204
rect 2384 1204 2396 1212
rect 2430 1212 2569 1238
rect 2430 1204 2442 1212
rect 2384 1198 2442 1204
rect 2557 1204 2569 1212
rect 2603 1204 2615 1238
rect 2557 1198 2615 1204
rect 1259 1176 1320 1184
rect 1259 1142 1271 1176
rect 1305 1167 1320 1176
rect 1432 1176 1493 1184
rect 1432 1167 1444 1176
rect 1305 1142 1444 1167
rect 1478 1167 1493 1176
rect 1603 1167 1609 1184
rect 1478 1142 1609 1167
rect 1661 1167 1667 1184
rect 1778 1176 1839 1184
rect 1778 1167 1790 1176
rect 1661 1142 1790 1167
rect 1824 1142 1839 1176
rect 1951 1176 2012 1184
rect 1951 1167 1963 1176
rect 1259 1136 1609 1142
rect 1603 1132 1609 1136
rect 1661 1136 1839 1142
rect 1950 1142 1963 1167
rect 1997 1167 2012 1176
rect 2121 1167 2127 1184
rect 1997 1142 2127 1167
rect 2179 1167 2185 1184
rect 2297 1176 2358 1184
rect 2297 1167 2309 1176
rect 2179 1142 2309 1167
rect 2343 1167 2358 1176
rect 2470 1176 2531 1184
rect 2470 1167 2482 1176
rect 2343 1142 2482 1167
rect 2516 1167 2531 1176
rect 2516 1142 2614 1167
rect 1950 1136 2127 1142
rect 1661 1132 1667 1136
rect 2121 1132 2127 1136
rect 2179 1136 2614 1142
rect 2179 1132 2185 1136
rect 1603 1131 1667 1132
rect 1239 1084 1292 1090
rect 1050 1050 1245 1084
rect 1280 1050 1292 1084
rect 1239 1044 1292 1050
rect 2120 1016 2126 1068
rect 2178 1059 2184 1068
rect 2178 1025 2782 1059
rect 2178 1016 2184 1025
rect 1239 890 1286 896
rect 1604 894 1610 946
rect 1662 937 1668 946
rect 1662 903 2782 937
rect 1662 894 1668 903
rect 1050 856 1245 890
rect 1280 856 1292 890
rect 1239 850 1286 856
rect 1107 798 2687 804
rect 1107 777 1185 798
rect 1107 743 1113 777
rect 1147 764 1185 777
rect 1219 772 1358 798
rect 1219 764 1231 772
rect 1147 758 1231 764
rect 1346 764 1358 772
rect 1392 772 1531 798
rect 1392 764 1404 772
rect 1346 758 1404 764
rect 1519 764 1531 772
rect 1565 772 1704 798
rect 1565 764 1577 772
rect 1519 758 1577 764
rect 1692 764 1704 772
rect 1738 772 1877 798
rect 1738 764 1750 772
rect 1692 758 1750 764
rect 1865 764 1877 772
rect 1911 772 2050 798
rect 1911 764 1923 772
rect 1865 758 1923 764
rect 2038 764 2050 772
rect 2084 772 2223 798
rect 2084 764 2096 772
rect 2038 758 2096 764
rect 2211 764 2223 772
rect 2257 772 2396 798
rect 2257 764 2269 772
rect 2211 758 2269 764
rect 2384 764 2396 772
rect 2430 772 2569 798
rect 2430 764 2442 772
rect 2384 758 2442 764
rect 2557 764 2569 772
rect 2603 783 2687 798
rect 2603 764 2647 783
rect 2557 758 2647 764
rect 1147 743 1157 758
rect 1107 731 1157 743
rect 1259 736 1320 744
rect 1259 702 1271 736
rect 1305 727 1320 736
rect 1432 736 1493 744
rect 1432 727 1444 736
rect 1305 702 1444 727
rect 1478 727 1493 736
rect 1603 743 1667 744
rect 1603 727 1609 743
rect 1478 702 1609 727
rect 1661 727 1667 743
rect 1778 736 1839 744
rect 1778 727 1790 736
rect 1661 702 1790 727
rect 1824 702 1839 736
rect 1259 696 1609 702
rect 1603 691 1609 696
rect 1661 696 1839 702
rect 1661 691 1667 696
rect 1877 572 1911 758
rect 2639 749 2647 758
rect 2681 749 2687 783
rect 1951 736 2012 744
rect 2124 742 2185 744
rect 1951 727 1963 736
rect 1950 702 1963 727
rect 1997 727 2012 736
rect 2123 727 2129 742
rect 1997 702 2129 727
rect 2181 727 2187 742
rect 2297 736 2358 744
rect 2297 727 2309 736
rect 2181 702 2309 727
rect 2343 727 2358 736
rect 2470 736 2531 744
rect 2639 737 2687 749
rect 2470 727 2482 736
rect 2343 702 2482 727
rect 2516 702 2531 736
rect 1950 696 2129 702
rect 2123 690 2129 696
rect 2181 696 2531 702
rect 2181 690 2187 696
rect 1050 502 2782 572
<< via1 >>
rect 1609 1176 1661 1184
rect 1609 1142 1617 1176
rect 1617 1142 1651 1176
rect 1651 1142 1661 1176
rect 1609 1132 1661 1142
rect 2127 1176 2179 1184
rect 2127 1142 2136 1176
rect 2136 1142 2170 1176
rect 2170 1142 2179 1176
rect 2127 1132 2179 1142
rect 2126 1016 2178 1068
rect 1610 894 1662 946
rect 1609 736 1661 743
rect 1609 702 1617 736
rect 1617 702 1651 736
rect 1651 702 1661 736
rect 1609 691 1661 702
rect 2129 736 2181 742
rect 2129 702 2136 736
rect 2136 702 2170 736
rect 2170 702 2181 736
rect 2129 690 2181 702
<< metal2 >>
rect 1603 1132 1609 1184
rect 1661 1132 1667 1184
rect 2121 1132 2127 1184
rect 2179 1132 2185 1184
rect 1617 946 1651 1132
rect 2136 1068 2170 1132
rect 2120 1016 2126 1068
rect 2178 1016 2184 1068
rect 1604 894 1610 946
rect 1662 894 1668 946
rect 1617 743 1651 894
rect 1603 691 1609 743
rect 1661 691 1667 743
rect 2136 742 2170 1016
rect 2123 690 2129 742
rect 2181 690 2187 742
<< labels >>
flabel space 1910 1690 2001 1761 0 FreeSans 480 0 0 0 VDDA
flabel space 1850 502 1941 573 0 FreeSans 480 0 0 0 GND
flabel via1 2126 1016 2178 1068 0 FreeSans 160 0 0 0 out
flabel via1 1610 894 1662 946 0 FreeSans 160 0 0 0 outb
flabel metal1 1245 1050 1280 1084 0 FreeSans 160 0 0 0 in
flabel metal1 1245 856 1280 890 0 FreeSans 160 0 0 0 inb
rlabel metal1 2782 533 2782 533 3 GND
rlabel metal1 2782 1724 2782 1724 3 VDDA
<< end >>
