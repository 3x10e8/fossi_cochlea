magic
tech sky130A
timestamp 1647843721
<< metal1 >>
rect 5783 -1259 5809 -1256
rect 5596 -1285 5783 -1273
rect 5809 -1285 5862 -1273
rect 5596 -1287 5862 -1285
rect 5783 -1288 5809 -1287
rect 5747 -1304 5773 -1302
rect 5597 -1305 5872 -1304
rect 5597 -1318 5747 -1305
rect 5773 -1318 5872 -1305
rect 5747 -1334 5773 -1331
rect 5600 -1347 5626 -1344
rect 5158 -1367 5600 -1350
rect 5626 -1367 5872 -1350
rect 5600 -1376 5626 -1373
rect 5713 -1581 5739 -1578
rect 5597 -1599 5713 -1585
rect 5713 -1610 5739 -1607
rect 5817 -1581 5843 -1578
rect 5843 -1599 5861 -1585
rect 5817 -1610 5843 -1607
rect 5637 -1718 5663 -1715
rect 5596 -1744 5637 -1734
rect 5663 -1744 5859 -1734
rect 5596 -1748 5859 -1744
rect 5683 -1765 5709 -1762
rect 5597 -1780 5683 -1766
rect 5709 -1780 5861 -1766
rect 5683 -1794 5709 -1791
<< via1 >>
rect 5783 -1285 5809 -1259
rect 5747 -1331 5773 -1305
rect 5600 -1373 5626 -1347
rect 5713 -1607 5739 -1581
rect 5817 -1607 5843 -1581
rect 5637 -1744 5663 -1718
rect 5683 -1791 5709 -1765
<< metal2 >>
rect 5613 -1344 5628 3199
rect 5600 -1347 5628 -1344
rect 5626 -1373 5628 -1347
rect 5600 -1376 5628 -1373
rect 5648 -1715 5663 3199
rect 5637 -1718 5663 -1715
rect 5637 -1747 5663 -1744
rect 5642 -1748 5663 -1747
rect 5648 -4841 5663 -1748
rect 5683 -1762 5698 3199
rect 5718 -1578 5733 3199
rect 5753 -1302 5768 3199
rect 5788 -1256 5803 3199
rect 5783 -1259 5809 -1256
rect 5783 -1288 5809 -1285
rect 5747 -1305 5773 -1302
rect 5747 -1334 5773 -1331
rect 5713 -1581 5739 -1578
rect 5713 -1610 5739 -1607
rect 5683 -1765 5709 -1762
rect 5683 -1794 5709 -1791
rect 5753 -4840 5768 -1334
rect 5823 -1578 5838 3199
rect 5817 -1581 5843 -1578
rect 5817 -1610 5843 -1607
use fitler_cell  fitler_cell_1
timestamp 1647843682
transform -1 0 11449 0 1 0
box -2644 -4825 5604 3103
use fitler_cell  fitler_cell_0
timestamp 1647843682
transform 1 0 2 0 1 0
box -2644 -4825 5604 3103
<< end >>
