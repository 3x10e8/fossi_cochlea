magic
tech sky130A
magscale 1 2
timestamp 1654644556
<< obsli1 >>
rect 1104 2159 58880 27761
<< obsm1 >>
rect 1104 1912 58880 28212
<< metal2 >>
rect 2686 29200 2742 30000
rect 8114 29200 8170 30000
rect 13542 29200 13598 30000
rect 18970 29200 19026 30000
rect 24490 29200 24546 30000
rect 29918 29200 29974 30000
rect 35346 29200 35402 30000
rect 40774 29200 40830 30000
rect 46294 29200 46350 30000
rect 51722 29200 51778 30000
rect 57150 29200 57206 30000
rect 5998 0 6054 800
rect 17958 0 18014 800
rect 29918 0 29974 800
rect 41970 0 42026 800
rect 53930 0 53986 800
<< obsm2 >>
rect 1398 29144 2630 29889
rect 2798 29144 8058 29889
rect 8226 29144 13486 29889
rect 13654 29144 18914 29889
rect 19082 29144 24434 29889
rect 24602 29144 29862 29889
rect 30030 29144 35290 29889
rect 35458 29144 40718 29889
rect 40886 29144 46238 29889
rect 46406 29144 51666 29889
rect 51834 29144 57094 29889
rect 57262 29144 58218 29889
rect 1398 856 58218 29144
rect 1398 711 5942 856
rect 6110 711 17902 856
rect 18070 711 29862 856
rect 30030 711 41914 856
rect 42082 711 53874 856
rect 54042 711 58218 856
<< metal3 >>
rect 0 29112 800 29232
rect 59200 29112 60000 29232
rect 0 27480 800 27600
rect 59200 27344 60000 27464
rect 0 25984 800 26104
rect 59200 25576 60000 25696
rect 0 24352 800 24472
rect 59200 23808 60000 23928
rect 0 22720 800 22840
rect 59200 22040 60000 22160
rect 0 21224 800 21344
rect 59200 20272 60000 20392
rect 0 19592 800 19712
rect 59200 18504 60000 18624
rect 0 17960 800 18080
rect 59200 16736 60000 16856
rect 0 16464 800 16584
rect 0 14832 800 14952
rect 59200 14968 60000 15088
rect 0 13336 800 13456
rect 59200 13200 60000 13320
rect 0 11704 800 11824
rect 59200 11432 60000 11552
rect 0 10072 800 10192
rect 59200 9664 60000 9784
rect 0 8576 800 8696
rect 59200 7896 60000 8016
rect 0 6944 800 7064
rect 59200 6128 60000 6248
rect 0 5312 800 5432
rect 59200 4360 60000 4480
rect 0 3816 800 3936
rect 59200 2592 60000 2712
rect 0 2184 800 2304
rect 0 688 800 808
rect 59200 824 60000 944
<< obsm3 >>
rect 800 29312 59200 29885
rect 880 29032 59120 29312
rect 800 27680 59200 29032
rect 880 27544 59200 27680
rect 880 27400 59120 27544
rect 800 27264 59120 27400
rect 800 26184 59200 27264
rect 880 25904 59200 26184
rect 800 25776 59200 25904
rect 800 25496 59120 25776
rect 800 24552 59200 25496
rect 880 24272 59200 24552
rect 800 24008 59200 24272
rect 800 23728 59120 24008
rect 800 22920 59200 23728
rect 880 22640 59200 22920
rect 800 22240 59200 22640
rect 800 21960 59120 22240
rect 800 21424 59200 21960
rect 880 21144 59200 21424
rect 800 20472 59200 21144
rect 800 20192 59120 20472
rect 800 19792 59200 20192
rect 880 19512 59200 19792
rect 800 18704 59200 19512
rect 800 18424 59120 18704
rect 800 18160 59200 18424
rect 880 17880 59200 18160
rect 800 16936 59200 17880
rect 800 16664 59120 16936
rect 880 16656 59120 16664
rect 880 16384 59200 16656
rect 800 15168 59200 16384
rect 800 15032 59120 15168
rect 880 14888 59120 15032
rect 880 14752 59200 14888
rect 800 13536 59200 14752
rect 880 13400 59200 13536
rect 880 13256 59120 13400
rect 800 13120 59120 13256
rect 800 11904 59200 13120
rect 880 11632 59200 11904
rect 880 11624 59120 11632
rect 800 11352 59120 11624
rect 800 10272 59200 11352
rect 880 9992 59200 10272
rect 800 9864 59200 9992
rect 800 9584 59120 9864
rect 800 8776 59200 9584
rect 880 8496 59200 8776
rect 800 8096 59200 8496
rect 800 7816 59120 8096
rect 800 7144 59200 7816
rect 880 6864 59200 7144
rect 800 6328 59200 6864
rect 800 6048 59120 6328
rect 800 5512 59200 6048
rect 880 5232 59200 5512
rect 800 4560 59200 5232
rect 800 4280 59120 4560
rect 800 4016 59200 4280
rect 880 3736 59200 4016
rect 800 2792 59200 3736
rect 800 2512 59120 2792
rect 800 2384 59200 2512
rect 880 2104 59200 2384
rect 800 1024 59200 2104
rect 800 888 59120 1024
rect 880 744 59120 888
rect 880 715 59200 744
<< metal4 >>
rect 10576 2128 10896 27792
rect 20208 2128 20528 27792
rect 29840 2128 30160 27792
rect 39472 2128 39792 27792
rect 49104 2128 49424 27792
<< obsm4 >>
rect 15331 27872 46677 29885
rect 15331 2048 20128 27872
rect 20608 2048 29760 27872
rect 30240 2048 39392 27872
rect 39872 2048 46677 27872
rect 15331 1531 46677 2048
<< labels >>
rlabel metal2 s 29918 29200 29974 30000 6 cclk_I
port 1 nsew signal output
rlabel metal2 s 35346 29200 35402 30000 6 cclk_Q
port 2 nsew signal output
rlabel metal3 s 59200 2592 60000 2712 6 clk_master
port 3 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 clk_master_out
port 4 nsew signal output
rlabel metal3 s 59200 4360 60000 4480 6 clkdiv2
port 5 nsew signal input
rlabel metal2 s 13542 29200 13598 30000 6 comp_high_I
port 6 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 comp_high_Q
port 7 nsew signal input
rlabel metal2 s 2686 29200 2742 30000 6 cos_out
port 8 nsew signal output
rlabel metal2 s 24490 29200 24546 30000 6 cos_outb
port 9 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 div2out
port 10 nsew signal output
rlabel metal2 s 8114 29200 8170 30000 6 fb1_I
port 11 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 fb1_Q
port 12 nsew signal output
rlabel metal2 s 18970 29200 19026 30000 6 fb2_I
port 13 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 fb2_Q
port 14 nsew signal output
rlabel metal3 s 59200 7896 60000 8016 6 gray_clk_in[0]
port 15 nsew signal input
rlabel metal3 s 59200 9664 60000 9784 6 gray_clk_in[1]
port 16 nsew signal input
rlabel metal3 s 59200 11432 60000 11552 6 gray_clk_in[2]
port 17 nsew signal input
rlabel metal3 s 59200 13200 60000 13320 6 gray_clk_in[3]
port 18 nsew signal input
rlabel metal3 s 59200 14968 60000 15088 6 gray_clk_in[4]
port 19 nsew signal input
rlabel metal3 s 59200 16736 60000 16856 6 gray_clk_in[5]
port 20 nsew signal input
rlabel metal3 s 59200 18504 60000 18624 6 gray_clk_in[6]
port 21 nsew signal input
rlabel metal3 s 59200 20272 60000 20392 6 gray_clk_in[7]
port 22 nsew signal input
rlabel metal3 s 59200 22040 60000 22160 6 gray_clk_in[8]
port 23 nsew signal input
rlabel metal3 s 59200 23808 60000 23928 6 gray_clk_in[9]
port 24 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 gray_clk_out[10]
port 25 nsew signal output
rlabel metal3 s 0 6944 800 7064 6 gray_clk_out[1]
port 26 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 gray_clk_out[2]
port 27 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 gray_clk_out[3]
port 28 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 gray_clk_out[4]
port 29 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 gray_clk_out[5]
port 30 nsew signal output
rlabel metal3 s 0 14832 800 14952 6 gray_clk_out[6]
port 31 nsew signal output
rlabel metal3 s 0 16464 800 16584 6 gray_clk_out[7]
port 32 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 gray_clk_out[8]
port 33 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 gray_clk_out[9]
port 34 nsew signal output
rlabel metal3 s 59200 25576 60000 25696 6 no_ones_below_in[0]
port 35 nsew signal input
rlabel metal3 s 59200 27344 60000 27464 6 no_ones_below_in[1]
port 36 nsew signal input
rlabel metal3 s 59200 29112 60000 29232 6 no_ones_below_in[2]
port 37 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 no_ones_below_out[0]
port 38 nsew signal output
rlabel metal3 s 0 24352 800 24472 6 no_ones_below_out[1]
port 39 nsew signal output
rlabel metal3 s 0 25984 800 26104 6 no_ones_below_out[2]
port 40 nsew signal output
rlabel metal2 s 40774 29200 40830 30000 6 phi1b_dig_I
port 41 nsew signal input
rlabel metal2 s 46294 29200 46350 30000 6 phi1b_dig_Q
port 42 nsew signal input
rlabel metal2 s 51722 29200 51778 30000 6 read_out_I[0]
port 43 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 read_out_I[1]
port 44 nsew signal output
rlabel metal2 s 57150 29200 57206 30000 6 read_out_Q[0]
port 45 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 read_out_Q[1]
port 46 nsew signal output
rlabel metal3 s 59200 824 60000 944 6 rstb
port 47 nsew signal input
rlabel metal3 s 0 688 800 808 6 rstb_out
port 48 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 sin_out
port 49 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 sin_outb
port 50 nsew signal output
rlabel metal3 s 59200 6128 60000 6248 6 ud_en
port 51 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 ud_en_out
port 52 nsew signal output
rlabel metal4 s 10576 2128 10896 27792 6 vccd1
port 53 nsew power input
rlabel metal4 s 29840 2128 30160 27792 6 vccd1
port 53 nsew power input
rlabel metal4 s 49104 2128 49424 27792 6 vccd1
port 53 nsew power input
rlabel metal4 s 20208 2128 20528 27792 6 vssd1
port 54 nsew ground input
rlabel metal4 s 39472 2128 39792 27792 6 vssd1
port 54 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 60000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3160784
string GDS_FILE /Volumes/export/isn/ishan/fossi_cochlea/openlane/wrapper_cell/runs/wrapper_cell/results/finishing/wrapper_cell.magic.gds
string GDS_START 407630
<< end >>

