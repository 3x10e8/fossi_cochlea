magic
tech sky130A
magscale 1 2
timestamp 1654305936
<< metal2 >>
rect -10241 27926 -10232 27982
rect -10176 27926 -10167 27982
rect -8477 27925 -8468 27981
rect -8412 27925 -8403 27981
rect 1579 27689 1588 27745
rect 1644 27689 1653 27745
rect 2946 27690 2955 27746
rect 3011 27690 3020 27746
rect 8562 27410 8614 27558
rect 8391 27354 8400 27410
rect 8456 27402 8614 27410
rect 9509 27402 9556 27562
rect 8456 27354 9556 27402
rect 8611 27353 9556 27354
<< via2 >>
rect -10232 27926 -10176 27982
rect -8468 27925 -8412 27981
rect 1588 27689 1644 27745
rect 2955 27690 3011 27746
rect 8400 27354 8456 27410
<< metal3 >>
rect -10241 27982 -9936 27987
rect -10241 27926 -10232 27982
rect -10176 27926 -9936 27982
rect -10241 27921 -9936 27926
rect -8710 27981 -8402 27986
rect -8710 27925 -8468 27981
rect -8412 27925 -8402 27981
rect -8710 27920 -8402 27925
rect 1579 27745 1799 27750
rect 1579 27689 1588 27745
rect 1644 27689 1799 27745
rect 1579 27684 1799 27689
rect 2816 27746 3036 27751
rect 2816 27690 2955 27746
rect 3011 27690 3036 27746
rect 2816 27685 3036 27690
rect 2780 27565 2828 27579
rect -9711 27215 -9529 27517
rect 2771 27156 2832 27565
rect 8391 27410 8465 27415
rect 8391 27409 8400 27410
rect 8293 27354 8400 27409
rect 8456 27354 8465 27410
rect 8293 27349 8465 27354
rect 8293 27213 8353 27349
rect 1351 26290 2784 26410
rect 1351 26205 2100 26290
rect 2190 26205 2784 26290
rect 1351 26090 2784 26205
rect 1362 22684 2795 22810
rect 1362 22599 2097 22684
rect 2187 22599 2795 22684
rect 1362 22490 2795 22599
rect 1369 19230 2802 19332
rect 1369 19145 2120 19230
rect 2210 19145 2802 19230
rect 1369 19012 2802 19145
rect 1360 15756 2793 15879
rect 1360 15671 2082 15756
rect 2172 15671 2793 15756
rect 1360 15559 2793 15671
rect 1367 12270 2800 12381
rect 1367 12185 2089 12270
rect 2179 12185 2800 12270
rect 1367 12061 2800 12185
rect 1373 8782 2806 8906
rect 1373 8697 2060 8782
rect 2150 8697 2806 8782
rect 1373 8586 2806 8697
rect 1365 5333 2798 5457
rect 1365 5248 2062 5333
rect 2152 5248 2798 5333
rect 1365 5137 2798 5248
rect 1358 1828 2791 1935
rect 1358 1743 2042 1828
rect 2132 1743 2791 1828
rect 1358 1615 2791 1743
<< via3 >>
rect 2100 26205 2190 26290
rect 2097 22599 2187 22684
rect 2120 19145 2210 19230
rect 2082 15671 2172 15756
rect 2089 12185 2179 12270
rect 2060 8697 2150 8782
rect 2062 5248 2152 5333
rect 2042 1743 2132 1828
<< metal4 >>
rect -10135 28126 -9830 28198
rect -8751 28126 -8490 28198
rect -8137 28126 -8023 28198
rect -8083 27118 -8023 28126
rect 1126 27890 1314 27962
rect 1681 27890 1785 27962
rect 2835 27890 2915 27962
rect 3290 27890 3373 27962
rect 1126 27227 1286 27890
rect 3295 27202 3373 27890
rect 8089 27748 8294 27820
rect 8658 27748 8735 27820
rect 9371 27748 9466 27820
rect 8089 27222 8249 27748
rect 9834 27220 9992 27820
<< via4 >>
rect 2024 26290 2277 26368
rect 2024 26205 2100 26290
rect 2100 26205 2190 26290
rect 2190 26205 2277 26290
rect 2024 26131 2277 26205
rect 2021 22684 2274 22762
rect 2021 22599 2097 22684
rect 2097 22599 2187 22684
rect 2187 22599 2274 22684
rect 2021 22525 2274 22599
rect 2044 19230 2297 19308
rect 2044 19145 2120 19230
rect 2120 19145 2210 19230
rect 2210 19145 2297 19230
rect 2044 19071 2297 19145
rect 2006 15756 2259 15834
rect 2006 15671 2082 15756
rect 2082 15671 2172 15756
rect 2172 15671 2259 15756
rect 2006 15597 2259 15671
rect 2013 12270 2266 12348
rect 2013 12185 2089 12270
rect 2089 12185 2179 12270
rect 2179 12185 2266 12270
rect 2013 12111 2266 12185
rect 1984 8782 2237 8860
rect 1984 8697 2060 8782
rect 2060 8697 2150 8782
rect 2150 8697 2237 8782
rect 1984 8623 2237 8697
rect 1986 5333 2239 5411
rect 1986 5248 2062 5333
rect 2062 5248 2152 5333
rect 2152 5248 2239 5333
rect 1986 5174 2239 5248
rect 1966 1828 2219 1906
rect 1966 1743 2042 1828
rect 2042 1743 2132 1828
rect 2132 1743 2219 1828
rect 1966 1669 2219 1743
<< metal5 >>
rect 1351 26368 2784 26410
rect 1351 26131 2024 26368
rect 2277 26131 2784 26368
rect 1351 26090 2784 26131
rect 1362 22762 2795 22810
rect 1362 22525 2021 22762
rect 2274 22525 2795 22762
rect 1362 22490 2795 22525
rect 1369 19308 2802 19332
rect 1369 19071 2044 19308
rect 2297 19071 2802 19308
rect 1369 19012 2802 19071
rect 1360 15834 2793 15879
rect 1360 15597 2006 15834
rect 2259 15597 2793 15834
rect 1360 15559 2793 15597
rect 1367 12348 2800 12381
rect 1367 12111 2013 12348
rect 2266 12111 2800 12348
rect 1367 12061 2800 12111
rect 1373 8860 2806 8906
rect 1373 8623 1984 8860
rect 2237 8623 2806 8860
rect 1373 8586 2806 8623
rect 1365 5411 2798 5457
rect 1365 5174 1986 5411
rect 2239 5174 2798 5411
rect 1365 5137 2798 5174
rect 1358 1906 2791 1935
rect 1358 1669 1966 1906
rect 2219 1669 2791 1906
rect 1358 1615 2791 1669
use cap_3pF_8x1  cap_3pF_8x1_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654300736
transform 0 -1 11832 1 0 3532
box -2794 0 23698 2104
use cap_6pF_8x2  cap_6pF_8x2_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654300736
transform 0 -1 8353 1 0 3532
box -2794 0 23698 5588
use cap_10fF  cap_10fF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654300736
transform 0 -1 9349 1 0 27529
box -28 -28 708 628
use cap_12pF  cap_12pF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654300736
transform 0 -1 -1404 1 0 3558
box -2820 -2794 23672 9762
use cap_20fF  cap_20fF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654300736
transform 0 -1 2809 1 0 27514
box -28 -28 828 1028
use cap_40fF  cap_40fF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654300736
transform 0 -1 -8732 1 0 27498
box -28 -28 1368 1228
use cmos_switch_fin  cmos_switch_0
timestamp 1654304341
transform 1 0 -10337 0 1 28009
box -175 -88 205 381
use cmos_switch_fin  cmos_switch_1
timestamp 1654304341
transform -1 0 -8307 0 1 28009
box -175 -88 205 381
use cmos_switch_fin  cmos_switch_2
timestamp 1654304341
transform 1 0 1483 0 1 27773
box -175 -88 205 381
use cmos_switch_fin  cmos_switch_3
timestamp 1654304341
transform -1 0 3116 0 1 27773
box -175 -88 205 381
use cmos_switch_fin  cmos_switch_4
timestamp 1654304341
transform 1 0 8455 0 1 27631
box -175 -88 205 381
use cmos_switch_fin  cmos_switch_5
timestamp 1654304341
transform -1 0 9665 0 1 27631
box -175 -88 205 381
<< end >>
