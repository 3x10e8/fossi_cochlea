magic
tech sky130A
magscale 1 2
timestamp 1649299711
<< locali >>
rect 106 -2734 348 -2700
<< viali >>
rect 72 -2734 106 -2700
<< metal1 >>
rect 10938 -2522 10990 -2516
rect 9582 -2574 10938 -2546
rect 10990 -2574 11724 -2546
rect 9596 -2636 10340 -2608
rect 10392 -2636 11744 -2608
rect 10340 -2666 10392 -2660
rect 11500 -2688 11552 -2682
rect 66 -2700 112 -2694
rect -9764 -2734 72 -2700
rect 106 -2734 118 -2700
rect 9560 -2734 11500 -2700
rect 66 -2740 112 -2734
rect 11552 -2734 11744 -2700
rect 11500 -2746 11552 -2740
rect 9736 -3156 9788 -3150
rect 9596 -3198 9736 -3170
rect 9736 -3214 9788 -3208
rect 11238 -3158 11290 -3152
rect 11290 -3198 11722 -3170
rect 11238 -3216 11290 -3210
rect 10038 -3444 10090 -3438
rect 9596 -3496 10038 -3468
rect 10090 -3496 11718 -3468
rect 9588 -3560 10640 -3532
rect 10692 -3560 11722 -3532
rect 10640 -3590 10692 -3584
rect 20278 -10354 27410 -10282
rect 12244 -10504 12296 -10498
rect 12244 -10562 12296 -10556
rect 20292 -10672 27424 -10600
<< via1 >>
rect 10938 -2574 10990 -2522
rect 10340 -2660 10392 -2608
rect 11500 -2740 11552 -2688
rect 9736 -3208 9788 -3156
rect 11238 -3210 11290 -3158
rect 10038 -3496 10090 -3444
rect 10640 -3584 10692 -3532
rect 12244 -10556 12296 -10504
rect 17782 -10840 17848 -10774
<< metal2 >>
rect 1386 15012 10414 15112
rect 1532 9546 10116 9646
rect 9714 -3156 9814 -3118
rect 9714 -3208 9736 -3156
rect 9788 -3208 9814 -3156
rect 9714 -17722 9814 -3208
rect 10014 -3444 10114 9546
rect 10014 -3496 10038 -3444
rect 10090 -3496 10114 -3444
rect 10014 -9628 10114 -3496
rect 10314 -2608 10414 15012
rect 10314 -2660 10340 -2608
rect 10392 -2660 10414 -2608
rect 10014 -9712 10118 -9628
rect 10314 -9650 10414 -2660
rect 10056 -10040 10118 -9712
rect 10298 -9712 10414 -9650
rect 10614 15024 19642 15124
rect 10614 -3532 10714 15024
rect 10614 -3584 10640 -3532
rect 10692 -3584 10714 -3532
rect 10614 -9712 10714 -3584
rect 10914 9638 11014 9640
rect 10914 9538 19498 9638
rect 10914 -2522 11014 9538
rect 10914 -2574 10938 -2522
rect 10990 -2574 11014 -2522
rect 10914 -9712 11014 -2574
rect 11494 -2688 11556 -2682
rect 11494 -2740 11500 -2688
rect 11552 -2740 11556 -2688
rect 11214 -3158 11314 -3122
rect 11214 -3210 11238 -3158
rect 11290 -3210 11314 -3158
rect 10298 -10062 10360 -9712
rect 11214 -17722 11314 -3210
rect 11494 -10182 11556 -2740
rect 12222 -10504 12322 -10484
rect 12222 -10556 12244 -10504
rect 12296 -10556 12322 -10504
rect 12222 -17726 12322 -10556
rect 17710 -10756 17958 -10692
rect 17710 -10846 17776 -10756
rect 17858 -10846 17958 -10756
rect 17710 -10860 17958 -10846
<< via2 >>
rect 17776 -10774 17858 -10756
rect 17776 -10840 17782 -10774
rect 17782 -10840 17848 -10774
rect 17848 -10840 17858 -10774
rect 17776 -10846 17858 -10840
<< metal3 >>
rect -5284 5705 -5096 12132
rect 17692 -10756 17976 -9528
rect 17692 -10846 17776 -10756
rect 17858 -10846 17976 -10756
rect 17692 -10868 17976 -10846
<< metal4 >>
rect -9666 6002 -6364 6210
rect 27668 6110 41764 6190
rect 10388 -9590 11786 -9508
rect 9182 -10504 9246 -9602
rect 10388 -10478 10456 -9590
rect 9182 -10570 10126 -10504
use comparator_final  comparator_final_0
timestamp 1647895372
transform 1 0 10662 0 1 -10434
box -574 -430 9642 401
use fitler_cell  fitler_cell_0
timestamp 1647840975
transform 1 0 -1596 0 1 0
box -5288 -9650 11208 6206
use fitler_cell  fitler_cell_1
timestamp 1647840975
transform -1 0 22898 0 1 0
box -5288 -9650 11208 6206
<< labels >>
rlabel metal1 -9764 -2718 -9764 -2718 7 vdd
port 23 w power bidirectional
rlabel metal1 27410 -10318 27410 -10318 1 polxevent
port 24 n
rlabel metal1 27424 -10638 27424 -10638 1 events
port 25 n
rlabel metal2 12274 -17726 12274 -17726 1 compout
port 26 n
rlabel metal2 11264 -17722 11264 -17722 5 vbotm
port 27 s
rlabel metal2 9770 -17722 9770 -17722 5 vbotp
port 28 s
rlabel metal2 1532 9594 1532 9594 7 phi1
port 29 w
rlabel metal2 1386 15056 1386 15056 7 phi1b
port 30 w
rlabel metal2 19642 15074 19642 15074 3 phi2
port 31 e
rlabel metal2 19498 9592 19498 9592 3 phi2b
port 32 e
rlabel metal4 -9666 6106 -9666 6106 7 inp
port 33 w
rlabel metal3 -5184 12132 -5184 12132 1 gnd
port 34 n
rlabel metal4 41764 6150 41764 6150 3 inm
port 35 e
<< end >>
