* SPICE3 file created from /home/soumil/Desktop/cmos_reram/level_up_shifter.ext - technology: sky130B

.subckt x/home/soumil/Desktop/cmos_reram/level_up_shifter in out outb vssd1 vccd1
+ vdda1
X0 vssd1 a_0_n1540# out vssd1 sky130_fd_pr__nfet_g5v0d10v5 ad=9e+11p pd=5.8e+06u as=4.5e+11p ps=2.9e+06u w=1e+06u l=500000u
X1 outb in vssd1 vssd1 sky130_fd_pr__nfet_g5v0d10v5 ad=4.5e+11p pd=2.9e+06u as=0p ps=0u w=1e+06u l=500000u
X2 vdda1 outb out vdda1 sky130_fd_pr__pfet_g5v0d10v5 ad=9e+11p pd=5.8e+06u as=4.5e+11p ps=2.9e+06u w=1e+06u l=500000u
X3 vdda1 a_0_n1540# outb vssd1 sky130_fd_pr__nfet_g5v0d10v5 ad=1.15e+12p pd=6.3e+06u as=0p ps=0u w=1e+06u l=500000u
X4 vccd1 in a_0_n1540# vccd1 sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=150000u
X5 out in vdda1 vssd1 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X6 a_0_n1540# in vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=150000u
X7 outb out vdda1 vdda1 sky130_fd_pr__pfet_g5v0d10v5 ad=4.5e+11p pd=2.9e+06u as=0p ps=0u w=1e+06u l=500000u
.ends

