magic
tech sky130A
timestamp 1647810894
<< nwell >>
rect -256 -3 226 82
<< pmos >>
rect -209 17 -194 59
rect -165 17 -150 59
rect 0 17 15 59
rect 44 17 59 59
rect 88 17 103 59
rect 132 17 147 59
<< nmoslvt >>
rect -215 -133 -200 -91
rect -162 -133 -147 -91
rect -52 -133 -37 -91
rect 0 -133 15 -91
rect 44 -133 59 -91
rect 88 -133 103 -91
rect 132 -133 147 -91
<< ndiff >>
rect -252 -102 -215 -91
rect -252 -119 -248 -102
rect -231 -119 -215 -102
rect -252 -133 -215 -119
rect -200 -102 -162 -91
rect -200 -119 -189 -102
rect -172 -119 -162 -102
rect -200 -133 -162 -119
rect -147 -102 -110 -91
rect -147 -119 -131 -102
rect -114 -119 -110 -102
rect -147 -133 -110 -119
rect -79 -102 -52 -91
rect -79 -119 -75 -102
rect -58 -119 -52 -102
rect -79 -133 -52 -119
rect -37 -108 0 -91
rect -37 -125 -30 -108
rect -13 -125 0 -108
rect -37 -133 0 -125
rect 15 -102 44 -91
rect 15 -119 21 -102
rect 38 -119 44 -102
rect 15 -133 44 -119
rect 59 -102 88 -91
rect 59 -119 65 -102
rect 82 -119 88 -102
rect 59 -133 88 -119
rect 103 -102 132 -91
rect 103 -119 109 -102
rect 126 -119 132 -102
rect 103 -133 132 -119
rect 147 -102 177 -91
rect 147 -119 153 -102
rect 170 -119 177 -102
rect 147 -133 177 -119
<< pdiff >>
rect -238 48 -209 59
rect -238 31 -232 48
rect -215 31 -209 48
rect -238 17 -209 31
rect -194 48 -165 59
rect -194 31 -188 48
rect -171 31 -165 48
rect -194 17 -165 31
rect -150 48 -123 59
rect -150 31 -144 48
rect -127 31 -123 48
rect -150 17 -123 31
rect -27 48 0 59
rect -27 31 -23 48
rect -6 31 0 48
rect -27 17 0 31
rect 15 48 44 59
rect 15 31 21 48
rect 38 31 44 48
rect 15 17 44 31
rect 59 48 88 59
rect 59 31 65 48
rect 82 31 88 48
rect 59 17 88 31
rect 103 48 132 59
rect 103 31 109 48
rect 126 31 132 48
rect 103 17 132 31
rect 147 48 177 59
rect 147 31 153 48
rect 170 31 177 48
rect 147 17 177 31
<< ndiffc >>
rect -248 -119 -231 -102
rect -189 -119 -172 -102
rect -131 -119 -114 -102
rect -75 -119 -58 -102
rect -30 -125 -13 -108
rect 21 -119 38 -102
rect 65 -119 82 -102
rect 109 -119 126 -102
rect 153 -119 170 -102
<< pdiffc >>
rect -232 31 -215 48
rect -188 31 -171 48
rect -144 31 -127 48
rect -23 31 -6 48
rect 21 31 38 48
rect 65 31 82 48
rect 109 31 126 48
rect 153 31 170 48
<< psubdiff >>
rect 177 -103 208 -91
rect 177 -120 191 -103
rect 177 -133 208 -120
<< nsubdiff >>
rect 177 46 208 59
rect 177 29 191 46
rect 177 17 208 29
<< psubdiffcont >>
rect 191 -120 208 -103
<< nsubdiffcont >>
rect 191 29 208 46
<< poly >>
rect 75 115 108 123
rect 75 98 83 115
rect 100 113 108 115
rect 100 98 147 113
rect 75 93 108 98
rect -209 59 -194 72
rect -165 59 -150 72
rect 0 59 15 72
rect 44 59 59 72
rect 88 59 103 72
rect 132 59 147 98
rect -77 42 -35 50
rect -77 25 -72 42
rect -55 25 -35 42
rect -77 17 -35 25
rect -209 7 -194 17
rect -165 7 -150 17
rect -209 -8 -102 7
rect -50 6 -35 17
rect 0 6 15 17
rect -123 -13 -86 -8
rect -50 -9 15 6
rect -123 -15 -85 -13
rect -118 -23 -85 -15
rect -102 -30 -85 -23
rect -102 -35 -50 -30
rect -223 -45 -191 -36
rect -223 -62 -216 -45
rect -199 -62 -191 -45
rect -223 -70 -191 -62
rect -170 -45 -139 -36
rect -170 -62 -163 -45
rect -146 -62 -139 -45
rect -170 -70 -139 -62
rect -102 -52 -76 -35
rect -59 -52 -50 -35
rect 44 -39 59 17
rect 88 1 103 17
rect 132 4 147 17
rect 84 -7 111 1
rect 84 -24 89 -7
rect 106 -24 111 -7
rect 84 -32 111 -24
rect -102 -57 -50 -52
rect 36 -42 59 -39
rect 36 -50 63 -42
rect -215 -91 -200 -70
rect -162 -91 -147 -70
rect -215 -146 -200 -133
rect -162 -146 -147 -133
rect -102 -141 -87 -57
rect 36 -67 41 -50
rect 58 -67 63 -50
rect 36 -75 63 -67
rect -52 -91 -37 -78
rect 0 -91 15 -78
rect 44 -91 59 -75
rect 88 -91 103 -32
rect 152 -47 179 -39
rect 152 -57 157 -47
rect 132 -64 157 -57
rect 174 -64 179 -47
rect 132 -72 179 -64
rect 132 -91 147 -72
rect -52 -141 -37 -133
rect -102 -156 -37 -141
rect 0 -167 15 -133
rect 44 -146 59 -133
rect 88 -146 103 -133
rect 132 -167 147 -133
rect 0 -182 147 -167
<< polycont >>
rect 83 98 100 115
rect -72 25 -55 42
rect -216 -62 -199 -45
rect -163 -62 -146 -45
rect -76 -52 -59 -35
rect 89 -24 106 -7
rect 41 -67 58 -50
rect 157 -64 174 -47
<< locali >>
rect -286 134 -268 151
rect -251 134 -232 151
rect -215 134 -196 151
rect -179 134 -160 151
rect -143 134 -124 151
rect -107 134 -88 151
rect -71 134 -52 151
rect -35 134 -16 151
rect 1 134 20 151
rect 37 134 56 151
rect 73 134 92 151
rect 109 134 128 151
rect 145 134 164 151
rect 181 134 200 151
rect 217 134 236 151
rect 253 134 268 151
rect -188 56 -171 134
rect -140 115 108 117
rect -140 100 83 115
rect -140 56 -123 100
rect 75 98 83 100
rect 100 98 108 115
rect 75 90 108 98
rect -252 48 -211 56
rect -252 31 -232 48
rect -215 31 -211 48
rect -252 23 -211 31
rect -192 48 -167 56
rect -192 31 -188 48
rect -171 31 -167 48
rect -192 23 -167 31
rect -148 55 -123 56
rect -148 48 -109 55
rect -148 31 -144 48
rect -127 31 -109 48
rect -148 23 -109 31
rect -252 -94 -235 23
rect -216 -45 -199 -36
rect -216 -70 -199 -62
rect -163 -45 -146 -36
rect -163 -70 -146 -62
rect -126 -94 -109 23
rect -75 42 -52 50
rect -75 25 -72 42
rect -55 25 -52 42
rect -75 17 -52 25
rect -27 48 -2 56
rect -27 31 -23 48
rect -6 31 -2 48
rect -27 23 -2 31
rect 17 48 42 56
rect 17 31 21 48
rect 38 31 42 48
rect 17 23 42 31
rect 61 48 88 56
rect 61 31 65 48
rect 82 31 88 48
rect 61 23 88 31
rect 105 48 130 56
rect 105 31 109 48
rect 126 31 130 48
rect 105 23 130 31
rect 149 48 174 56
rect 149 31 153 48
rect 170 31 174 48
rect 149 23 174 31
rect 191 46 208 134
rect -27 -7 -10 23
rect 89 -7 106 1
rect 153 -2 170 23
rect 191 21 208 29
rect -27 -24 89 -7
rect -84 -52 -76 -35
rect -59 -52 -51 -35
rect 7 -94 24 -24
rect 89 -32 106 -24
rect 123 -19 170 -2
rect 41 -50 58 -42
rect 123 -50 140 -19
rect 58 -67 140 -50
rect 41 -75 58 -67
rect 110 -74 140 -67
rect 157 -47 174 -39
rect 157 -72 174 -64
rect 110 -94 127 -74
rect -252 -102 -227 -94
rect -252 -119 -248 -102
rect -231 -119 -227 -102
rect -252 -127 -227 -119
rect -193 -102 -168 -94
rect -193 -119 -189 -102
rect -172 -119 -168 -102
rect -193 -127 -168 -119
rect -135 -102 -109 -94
rect -135 -119 -131 -102
rect -114 -111 -109 -102
rect -78 -102 -54 -94
rect -114 -119 -110 -111
rect -135 -127 -110 -119
rect -78 -119 -75 -102
rect -58 -119 -54 -102
rect -78 -127 -54 -119
rect -33 -108 -10 -100
rect -33 -125 -30 -108
rect -13 -125 -10 -108
rect 7 -102 42 -94
rect 7 -111 21 -102
rect -190 -145 -173 -127
rect -78 -145 -61 -127
rect -33 -133 -10 -125
rect 17 -119 21 -111
rect 38 -119 42 -102
rect 17 -127 42 -119
rect 61 -102 86 -94
rect 61 -119 65 -102
rect 82 -119 86 -102
rect 61 -127 86 -119
rect 105 -102 130 -94
rect 105 -119 109 -102
rect 126 -119 130 -102
rect 105 -127 130 -119
rect 149 -102 174 -94
rect 149 -119 153 -102
rect 170 -119 174 -102
rect 149 -127 174 -119
rect 191 -103 208 -94
rect -190 -162 -61 -145
rect -27 -182 -10 -133
rect 66 -182 83 -127
rect 154 -182 171 -127
rect 191 -182 208 -120
rect -286 -199 -196 -182
rect -179 -199 -160 -182
rect -143 -199 -124 -182
rect -107 -199 -88 -182
rect -71 -199 -52 -182
rect -35 -199 -16 -182
rect 1 -199 20 -182
rect 37 -199 56 -182
rect 73 -199 92 -182
rect 109 -199 128 -182
rect 145 -199 164 -182
rect 181 -199 200 -182
rect 217 -199 236 -182
rect 253 -199 268 -182
<< viali >>
rect -268 134 -251 151
rect -232 134 -215 151
rect -196 134 -179 151
rect -160 134 -143 151
rect -124 134 -107 151
rect -88 134 -71 151
rect -52 134 -35 151
rect -16 134 1 151
rect 20 134 37 151
rect 56 134 73 151
rect 92 134 109 151
rect 128 134 145 151
rect 164 134 181 151
rect 200 134 217 151
rect 236 134 253 151
rect -232 31 -215 48
rect -72 25 -55 42
rect 65 31 82 48
rect -196 -199 -179 -182
rect -160 -199 -143 -182
rect -124 -199 -107 -182
rect -88 -199 -71 -182
rect -52 -199 -35 -182
rect -16 -199 1 -182
rect 20 -199 37 -182
rect 56 -199 73 -182
rect 92 -199 109 -182
rect 128 -199 145 -182
rect 164 -199 181 -182
rect 200 -199 217 -182
rect 236 -199 253 -182
<< metal1 >>
rect -286 151 268 167
rect -286 134 -268 151
rect -251 134 -232 151
rect -215 134 -196 151
rect -179 134 -160 151
rect -143 134 -124 151
rect -107 134 -88 151
rect -71 134 -52 151
rect -35 134 -16 151
rect 1 134 20 151
rect 37 134 56 151
rect 73 134 92 151
rect 109 134 128 151
rect 145 134 164 151
rect 181 134 200 151
rect 217 134 236 151
rect 253 134 268 151
rect -286 118 268 134
rect -238 49 -211 52
rect 65 51 82 118
rect -238 48 -52 49
rect -238 31 -232 48
rect -215 42 -52 48
rect -215 31 -72 42
rect -238 30 -72 31
rect -238 27 -211 30
rect -75 25 -72 30
rect -55 25 -52 42
rect 62 48 85 51
rect 62 31 65 48
rect 82 31 85 48
rect 62 25 85 31
rect -75 18 -52 25
rect -286 -182 268 -166
rect -286 -199 -196 -182
rect -179 -199 -160 -182
rect -143 -199 -124 -182
rect -107 -199 -88 -182
rect -71 -199 -52 -182
rect -35 -199 -16 -182
rect 1 -199 20 -182
rect 37 -199 56 -182
rect 73 -199 92 -182
rect 109 -199 128 -182
rect 145 -199 164 -182
rect 181 -199 200 -182
rect 217 -199 236 -182
rect 253 -199 268 -182
rect -286 -215 268 -199
<< labels >>
rlabel locali 268 -189 268 -189 3 GND
rlabel locali 268 142 268 142 3 VDD
flabel polycont 89 -24 106 -7 0 FreeSans 56 0 0 0 high
flabel polycont 41 -67 58 -50 0 FreeSans 56 0 0 0 low
flabel polycont 157 -64 174 -47 0 FreeSans 56 0 0 0 phi1b
flabel polycont -76 -52 -59 -35 0 FreeSans 56 0 0 0 phi1
rlabel locali -51 -44 -51 -44 3 phi1
rlabel locali 118 56 118 56 1 pfete
rlabel locali 30 56 30 56 1 pfetw
rlabel locali 118 -94 118 -94 1 low
rlabel locali 30 -94 30 -94 1 high
rlabel locali 165 -39 165 -39 1 phi1b
rlabel locali -104 -145 -104 -145 1 tail
rlabel locali -155 -37 -155 -37 1 inm
flabel polycont -163 -62 -146 -45 0 FreeSans 56 0 0 0 inm
flabel polycont -216 -62 -199 -45 0 FreeSans 56 0 0 0 inp
rlabel locali -207 -36 -207 -36 1 inp
rlabel locali -235 -20 -235 -20 3 FP
rlabel locali -126 -23 -126 -23 7 FN
<< end >>
