magic
tech sky130B
magscale 1 2
timestamp 1661195607
<< error_s >>
rect 25556 33422 25620 33506
rect 25620 33358 25724 33422
rect 26207 33110 26213 33116
rect 26253 33110 26259 33116
rect 26201 33104 26265 33110
rect 26207 33064 26259 33104
rect 26201 33058 26265 33064
rect 26207 33052 26213 33058
rect 26253 33052 26259 33058
rect 25260 32821 25311 32871
rect 26208 32636 26214 32642
rect 26254 32636 26260 32642
rect 26202 32630 26266 32636
rect 26208 32590 26260 32630
rect 26202 32584 26266 32590
rect 26208 32578 26214 32584
rect 26254 32578 26260 32584
rect 25563 32328 25569 32334
rect 25609 32328 25615 32334
rect 25557 32322 25621 32328
rect 25563 32282 25615 32322
rect 25557 32276 25621 32282
rect 25563 32270 25569 32276
rect 25609 32270 25615 32276
rect 21130 29440 21136 29446
rect 21176 29440 21182 29446
rect 26894 29440 26900 29446
rect 26940 29440 26946 29446
rect 21124 29434 21188 29440
rect 26888 29434 26952 29440
rect 21130 29394 21182 29434
rect 26894 29394 26946 29434
rect 21124 29388 21188 29394
rect 26888 29388 26952 29394
rect 21130 29382 21136 29388
rect 21176 29382 21182 29388
rect 26894 29382 26900 29388
rect 26940 29382 26946 29388
rect 22202 28666 22240 28717
rect 25820 28683 25861 28717
rect 494 26616 500 26622
rect 540 26616 546 26622
rect 1188 26621 1194 26627
rect 1234 26621 1240 26627
rect 46836 26621 46842 26627
rect 46882 26621 46888 26627
rect 488 26610 552 26616
rect 1182 26615 1246 26621
rect 46830 26615 46894 26621
rect 47530 26616 47536 26622
rect 47576 26616 47582 26622
rect 494 26570 546 26610
rect 488 26564 552 26570
rect 751 26568 785 26602
rect 494 26558 500 26564
rect 540 26558 546 26564
rect 931 26552 965 26602
rect 1188 26575 1240 26615
rect 46836 26575 46888 26615
rect 47524 26610 47588 26616
rect 1182 26569 1246 26575
rect 46830 26569 46894 26575
rect 1188 26563 1194 26569
rect 1234 26563 1240 26569
rect 46836 26563 46842 26569
rect 46882 26563 46888 26569
rect 47111 26552 47145 26602
rect 47291 26568 47325 26602
rect 47530 26570 47582 26610
rect 47524 26564 47588 26570
rect 47530 26558 47536 26564
rect 47576 26558 47582 26564
<< nwell >>
rect 25556 33358 25620 33422
<< psubdiff >>
rect 25260 32821 25311 32871
<< locali >>
rect 25260 32821 25311 32871
rect 22218 28813 22252 29386
rect 25824 28777 25858 29363
<< viali >>
rect 22218 29386 22252 29420
<< metal1 >>
rect 18170 37076 22434 37136
rect 18170 36702 18230 37076
rect 19566 36760 19660 36766
rect 19370 36754 21090 36760
rect 19370 36702 19586 36754
rect 19642 36744 21090 36754
rect 19642 36702 21208 36744
rect 19370 36698 21208 36702
rect 22374 36698 22434 37076
rect 20892 36666 21208 36698
rect 20892 36664 20998 36666
rect 19338 36202 21126 36216
rect 19338 36182 21206 36202
rect 19338 36130 21112 36182
rect 21164 36130 21206 36182
rect 19338 36120 21206 36130
rect 21066 36106 21206 36120
rect 20892 35658 20998 35662
rect 18902 35642 21168 35658
rect 18902 35572 19574 35642
rect 19644 35572 21168 35642
rect 18902 35560 21168 35572
rect 18906 35456 19118 35560
rect 18914 33738 19088 35456
rect 24646 34222 24698 34228
rect 23265 34172 24646 34216
rect 24646 34164 24698 34170
rect 24403 33734 24455 33740
rect 23252 33685 24403 33729
rect 24403 33676 24455 33682
rect 23531 33365 24319 33444
rect 25556 33415 25620 33422
rect 25556 33363 25562 33415
rect 25614 33363 25620 33415
rect 25556 33358 25620 33363
rect 18114 33228 18616 33264
rect 19238 33236 19270 33244
rect 18114 33162 18126 33228
rect 18180 33162 18616 33228
rect 18114 33126 18616 33162
rect 19130 33154 19270 33236
rect 19238 32818 19270 33154
rect 24210 33113 24262 33119
rect 23256 33065 24210 33109
rect 24210 33055 24262 33061
rect 23547 32823 24335 32902
rect 25260 32821 25311 32871
rect 23757 32641 23810 32647
rect 23250 32597 23757 32641
rect 23810 32589 24300 32635
rect 23757 32583 24300 32589
rect 23789 32581 24300 32583
rect 23538 32271 24326 32350
rect 23593 32016 23646 32022
rect 23229 31959 23593 32016
rect 23645 31959 23646 32016
rect 23593 31953 23646 31959
rect 23225 31614 23277 31620
rect 23225 31447 23277 31453
rect 13786 30310 22323 30350
rect 25813 30311 25866 30350
rect 25881 30311 34418 30350
rect 25884 30310 34418 30311
rect 13796 30190 22333 30230
rect 22335 30190 22387 30230
rect 25686 30190 25738 30230
rect 25744 30190 34281 30230
rect 24402 30120 24456 30126
rect 24402 30068 24403 30120
rect 24455 30068 24456 30120
rect 24402 30062 24456 30068
rect 24645 29997 24697 30003
rect 24645 29939 24697 29945
rect 23758 29880 23810 29886
rect 23758 29822 23810 29828
rect 24209 29756 24261 29762
rect 24209 29698 24261 29704
rect 23593 28713 23645 28719
rect 22201 28666 23593 28711
rect 23645 28666 25876 28711
rect 23593 28654 23645 28661
rect 23224 28544 23276 28550
rect 22279 28496 23224 28541
rect 23276 28496 25793 28541
rect 23224 28486 23276 28492
rect 24645 28453 24697 28459
rect 23390 28447 23442 28453
rect 22206 28406 23390 28440
rect 23442 28406 24645 28440
rect 24697 28406 25871 28440
rect 24645 28395 24697 28401
rect 23390 28389 23442 28395
<< via1 >>
rect 19586 36702 19642 36754
rect 22490 36666 22548 36722
rect 21112 36130 21164 36182
rect 19574 35572 19644 35642
rect 22954 35580 23014 35638
rect 24646 34170 24698 34222
rect 24403 33682 24455 33734
rect 25562 33363 25614 33415
rect 18126 33162 18180 33228
rect 24210 33061 24262 33113
rect 26207 33058 26259 33110
rect 23757 32589 23810 32641
rect 26208 32584 26260 32636
rect 25563 32276 25615 32328
rect 23593 31959 23645 32016
rect 23225 31453 23277 31614
rect 24403 30068 24455 30120
rect 24645 29945 24697 29997
rect 23758 29828 23810 29880
rect 24209 29704 24261 29756
rect 23593 28661 23645 28713
rect 23224 28492 23276 28544
rect 23390 28395 23442 28447
rect 24645 28401 24697 28453
rect 24018 26706 24070 26758
<< metal2 >>
rect 19566 36754 19660 36766
rect 19566 36702 19586 36754
rect 19642 36702 19660 36754
rect 18114 33228 18190 35674
rect 19566 35642 19660 36702
rect 22476 36730 22562 36750
rect 22476 36660 22484 36730
rect 22552 36660 22562 36730
rect 22476 36650 22562 36660
rect 21090 36188 21186 36206
rect 21090 36124 21106 36188
rect 21168 36124 21186 36188
rect 21090 36106 21186 36124
rect 19566 35572 19574 35642
rect 19644 35572 19660 35642
rect 19566 35564 19660 35572
rect 22934 35644 23032 35658
rect 22934 35574 22948 35644
rect 23018 35574 23032 35644
rect 22934 35562 23032 35574
rect 24646 34222 24698 34228
rect 24646 34164 24698 34170
rect 24403 33734 24455 33740
rect 24403 33676 24455 33682
rect 18114 33162 18126 33228
rect 18180 33162 18190 33228
rect 18114 33140 18190 33162
rect 24210 33113 24262 33119
rect 24210 33055 24262 33061
rect 23757 32641 23810 32647
rect 23757 32583 23810 32589
rect 23593 32016 23646 32022
rect 23645 31959 23646 32016
rect 23593 31953 23646 31959
rect 23225 31614 23277 31620
rect 23225 31447 23277 31453
rect 21701 30758 21757 30767
rect 21701 30693 21757 30702
rect 21714 30481 21748 30693
rect 22096 30579 22130 30580
rect 22085 30570 22141 30579
rect 22085 30505 22141 30514
rect 21713 28443 21749 30481
rect 21713 28405 21922 28443
rect 22095 28442 22131 30505
rect 22202 28666 22240 28717
rect 23227 28551 23275 31447
rect 23594 28719 23644 31953
rect 23758 29880 23810 32583
rect 23758 29809 23810 29828
rect 24009 30958 24080 30970
rect 24009 30902 24017 30958
rect 24073 30902 24080 30958
rect 23593 28713 23645 28719
rect 23593 28654 23645 28661
rect 23224 28544 23276 28551
rect 23224 28486 23276 28492
rect 23390 28447 23442 28453
rect 23390 28389 23442 28395
rect 23400 26902 23434 28389
rect 24009 26758 24080 30902
rect 24211 29762 24260 33055
rect 24404 30126 24454 33676
rect 24402 30120 24456 30126
rect 24402 30068 24403 30120
rect 24455 30068 24456 30120
rect 24402 30062 24456 30068
rect 24404 30060 24454 30062
rect 24647 30003 24696 34164
rect 25560 33419 25618 33428
rect 25560 33352 25618 33361
rect 26195 33118 26275 33127
rect 26195 33055 26204 33118
rect 26266 33055 26275 33118
rect 26195 33046 26275 33055
rect 26206 32638 26262 32647
rect 26206 32573 26262 32582
rect 25557 32334 25619 32343
rect 25557 32263 25619 32272
rect 25935 30765 25991 30774
rect 25935 30700 25991 30709
rect 24645 29997 24697 30003
rect 24645 29939 24697 29945
rect 24647 29925 24696 29939
rect 24209 29756 24261 29762
rect 24209 29698 24261 29704
rect 25820 28683 25861 28717
rect 24645 28453 24697 28459
rect 25946 28432 25980 30700
rect 26315 30568 26371 30578
rect 26315 30503 26371 30512
rect 26328 28440 26362 30503
rect 26152 28403 26362 28440
rect 24645 28395 24697 28401
rect 24656 26902 24690 28395
rect 24009 26706 24018 26758
rect 24070 26706 24080 26758
rect 24009 26700 24080 26706
rect 46310 26270 47033 26314
rect 24015 26077 24071 26081
rect 46310 26064 46355 26270
rect 1063 26007 1751 26051
<< via2 >>
rect 22484 36722 22552 36730
rect 22484 36666 22490 36722
rect 22490 36666 22548 36722
rect 22548 36666 22552 36722
rect 22484 36660 22552 36666
rect 21106 36182 21168 36188
rect 21106 36130 21112 36182
rect 21112 36130 21164 36182
rect 21164 36130 21168 36182
rect 21106 36124 21168 36130
rect 22948 35638 23018 35644
rect 22948 35580 22954 35638
rect 22954 35580 23014 35638
rect 23014 35580 23018 35638
rect 22948 35574 23018 35580
rect 21701 30702 21757 30758
rect 22085 30514 22141 30570
rect 24017 30902 24073 30958
rect 25560 33415 25618 33419
rect 25560 33363 25562 33415
rect 25562 33363 25614 33415
rect 25614 33363 25618 33415
rect 25560 33361 25618 33363
rect 26204 33110 26266 33118
rect 26204 33058 26207 33110
rect 26207 33058 26259 33110
rect 26259 33058 26266 33110
rect 26204 33055 26266 33058
rect 26206 32636 26262 32638
rect 26206 32584 26208 32636
rect 26208 32584 26260 32636
rect 26260 32584 26262 32636
rect 26206 32582 26262 32584
rect 25557 32328 25619 32334
rect 25557 32276 25563 32328
rect 25563 32276 25615 32328
rect 25615 32276 25619 32328
rect 25557 32272 25619 32276
rect 25935 30709 25991 30765
rect 26315 30512 26371 30568
<< metal3 >>
rect 22478 36730 22560 36744
rect 22478 36660 22484 36730
rect 22552 36660 22560 36730
rect 21092 36188 21186 36210
rect 21092 36124 21106 36188
rect 21168 36124 21186 36188
rect 21092 33964 21186 36124
rect 22478 34504 22560 36660
rect 22934 35644 23032 35658
rect 22934 35574 22948 35644
rect 23018 35574 23032 35644
rect 22934 35562 23032 35574
rect 22944 33914 23018 35562
rect 25540 33422 25640 33439
rect 25540 33358 25556 33422
rect 25620 33358 25640 33422
rect 25540 33340 25640 33358
rect 26179 33127 26288 33144
rect 26179 33046 26195 33127
rect 26275 33046 26288 33127
rect 26179 33036 26288 33046
rect 26181 32644 26283 32660
rect 26181 32580 26201 32644
rect 26267 32580 26283 32644
rect 26181 32558 26283 32580
rect 25532 32344 25643 32357
rect 25530 32337 25643 32344
rect 25530 32268 25553 32337
rect 25623 32268 25643 32337
rect 25530 32238 25643 32268
rect 25530 30928 25641 32238
rect 21701 30758 21757 30767
rect 21701 30693 21757 30702
rect 25935 30765 25991 30774
rect 25935 30700 25991 30709
rect 22085 30570 22141 30579
rect 22085 30505 22141 30514
rect 26315 30568 26371 30578
rect 26315 30503 26371 30512
rect 23278 26637 23355 26642
rect 23278 26571 23284 26637
rect 23349 26571 23355 26637
rect 23278 26566 23355 26571
rect 24730 26636 24807 26642
rect 24730 26572 24737 26636
rect 24801 26572 24807 26636
rect 24730 26566 24807 26572
rect 24004 26083 24081 26092
rect 24004 26019 24010 26083
rect 24074 26019 24081 26083
rect 24004 26013 24081 26019
<< via3 >>
rect 25556 33419 25620 33422
rect 25556 33361 25560 33419
rect 25560 33361 25618 33419
rect 25618 33361 25620 33419
rect 25556 33358 25620 33361
rect 26195 33118 26275 33127
rect 26195 33055 26204 33118
rect 26204 33055 26266 33118
rect 26266 33055 26275 33118
rect 26195 33046 26275 33055
rect 26201 32638 26267 32644
rect 26201 32582 26206 32638
rect 26206 32582 26262 32638
rect 26262 32582 26267 32638
rect 26201 32580 26267 32582
rect 25553 32334 25623 32337
rect 25553 32272 25557 32334
rect 25557 32272 25619 32334
rect 25619 32272 25623 32334
rect 25553 32268 25623 32272
rect 18624 30895 18710 30971
rect 22940 29565 23014 29636
rect 22483 29373 22555 29445
rect 23284 26571 23349 26637
rect 24737 26572 24801 26636
rect 24010 26019 24074 26083
<< metal4 >>
rect 25550 33422 25625 33423
rect 25550 33358 25556 33422
rect 25620 33358 25625 33422
rect 25550 32337 25625 33358
rect 26179 33127 26288 33144
rect 26179 33121 26195 33127
rect 26043 33048 26195 33121
rect 25550 32268 25553 32337
rect 25623 32268 25625 32337
rect 25550 32266 25625 32268
rect 26044 31848 26111 33048
rect 26179 33046 26195 33048
rect 26275 33046 26288 33127
rect 26179 33036 26288 33046
rect 26181 32644 26510 32654
rect 26181 32580 26201 32644
rect 26267 32580 26510 32644
rect 26181 32553 26510 32580
rect 24241 31776 26111 31848
rect 18618 30971 18716 31605
rect 18618 30895 18624 30971
rect 18710 30895 18716 30971
rect 18618 30886 18716 30895
rect 22481 29445 22558 31276
rect 22933 29636 23019 31187
rect 22933 29565 22940 29636
rect 23014 29565 23019 29636
rect 22933 29532 23019 29565
rect 22481 29373 22483 29445
rect 22555 29373 22558 29445
rect 22481 29341 22558 29373
rect 24241 27210 24316 31776
rect 26444 31486 26508 32553
rect 23824 27124 24316 27210
rect 24737 31422 26508 31486
rect 23284 26642 23349 26769
rect 23278 26637 23355 26642
rect 23278 26571 23284 26637
rect 23349 26571 23355 26637
rect 23278 26566 23355 26571
rect 24010 26089 24076 27124
rect 24737 26642 24801 31422
rect 26444 31421 26508 31422
rect 24730 26636 24807 26642
rect 24730 26572 24737 26636
rect 24801 26572 24807 26636
rect 24730 26566 24807 26572
rect 24004 26083 24081 26089
rect 24004 26019 24010 26083
rect 24074 26019 24081 26083
rect 24004 26013 24081 26019
use comp_for_tapeout  comparator_0 comparator
timestamp 1654756920
transform 1 0 23898 0 1 26079
box -3794 -2465 4606 4342
use filter  filter_0 comparator
timestamp 1661195607
transform 1 0 1272 0 1 -2522
box -1298 2522 22766 33508
use filter  filter_1
timestamp 1661195607
transform -1 0 46804 0 1 -2522
box -1298 2522 22766 33508
use filter_clkgen  filter_clkgen_0 ~/Documents/fossi_cochlea/mag/final_designs/clkgen
timestamp 1654754240
transform 1 0 20194 0 1 33321
box -1661 -2136 3360 1229
use level_shifter_low  level_shifter_low_0 comparator
timestamp 1654753126
transform 1 0 24311 0 1 32844
box -71 -46 2139 722
use level_shifter_low  level_shifter_low_1
timestamp 1654753126
transform 1 0 24311 0 -1 32848
box -71 -46 2139 722
use level_up_shifter_d_a  level_up_shifter_d_a_0 ~/Documents/fossi_cochlea/mag/final_designs/level_up_shifter
timestamp 1654754240
transform 1 0 20716 0 1 35064
box 402 498 2794 1682
use level_up_shifter_d_a  level_up_shifter_d_a_1
timestamp 1654754240
transform -1 0 19792 0 1 35100
box 402 498 2794 1682
<< end >>
