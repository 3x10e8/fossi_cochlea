magic
tech sky130A
magscale 1 2
timestamp 1654749871
use filter_i_q  filter_i_q_0
timestamp 1654749871
transform 0 1 85685 -1 0 629236
box -30375 4022 18307 154222
use user_analog_project_wrapper_empty  user_analog_project_wrapper_empty_0 /Volumes/export/isn/abhinav/caravel_user_project_analog/mag
timestamp 1632839657
transform 1 0 0 0 1 0
box -800 -800 584800 704800
<< end >>
