magic
tech sky130A
magscale 1 2
timestamp 1647878126
<< nwell >>
rect -482 1810 -398 1978
rect -62 784 235 987
<< locali >>
rect -522 2030 -494 2064
rect -516 1364 -496 1398
<< viali >>
rect -1118 1681 -1084 1715
rect -1628 1623 -1594 1657
rect -580 1584 -545 1620
rect -322 1590 -288 1624
<< metal1 >>
rect -520 2064 -492 2096
rect -522 2030 -492 2064
rect -520 1998 -492 2030
rect -1782 1751 -1730 1757
rect -1136 1727 -1130 1728
rect -1730 1699 -1130 1727
rect -1782 1693 -1730 1699
rect -1136 1669 -1130 1699
rect -1071 1669 -1065 1728
rect -1640 1657 -1582 1669
rect -1640 1623 -1628 1657
rect -1594 1623 -1582 1657
rect -334 1638 -276 1642
rect -1640 1611 -1582 1623
rect -587 1636 -276 1638
rect -587 1620 -334 1636
rect -587 1584 -580 1620
rect -545 1584 -334 1620
rect -587 1578 -334 1584
rect -587 1572 -276 1578
rect -587 1570 -293 1572
rect -518 1398 -498 1430
rect 946 1412 1006 1418
rect -544 1364 -480 1398
rect -518 1332 -498 1364
rect 946 1344 1006 1350
rect 39 1128 248 1158
rect -921 1096 -887 1109
rect -921 1089 -874 1096
rect 39 1089 68 1128
rect -921 1059 68 1089
rect 108 1059 154 1080
<< via1 >>
rect -1782 1699 -1730 1751
rect -1130 1715 -1071 1728
rect -1130 1681 -1118 1715
rect -1118 1681 -1084 1715
rect -1084 1681 -1071 1715
rect -1130 1669 -1071 1681
rect -334 1624 -276 1636
rect -334 1590 -322 1624
rect -322 1590 -288 1624
rect -288 1590 -276 1624
rect -334 1578 -276 1590
rect 946 1350 1006 1412
rect -1816 1031 -1749 1084
<< metal2 >>
rect -1782 1751 -1730 1757
rect -1782 1693 -1730 1699
rect -1782 1090 -1752 1693
rect -1136 1669 -1130 1728
rect -1071 1669 -1065 1728
rect -334 1636 -276 1642
rect -334 1572 -276 1578
rect 946 1412 1006 1418
rect 946 1344 1006 1350
rect 236 1092 270 1142
rect -1816 1084 -1749 1090
rect -1816 1025 -1749 1031
rect 958 1028 992 1344
use cclkgen  cclkgen_0
timestamp 1647875723
transform 1 0 -1536 0 -1 1430
box -359 -1 1646 764
use sky130_fd_sc_lp__dlclkp_1  sky130_fd_sc_lp__dlclkp_1_0 ~/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1640761190
transform 1 0 -1857 0 1 1381
box -38 -49 1382 715
use phi2gen  phi2gen_0
timestamp 1647876791
transform 1 0 192 0 1 1332
box -702 -666 1348 764
<< end >>
