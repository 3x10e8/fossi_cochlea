magic
tech sky130A
timestamp 1654156678
use cap_10_10_x2  cap_10_10_x2_0
array 0 3 1098 0 3 1098
timestamp 1654156239
transform 1 0 54 0 1 53
box -57 -52 1041 1046
<< labels >>
flabel space -3 1 4389 4393 0 FreeSans 4000 0 0 0 6.4pF
<< end >>
