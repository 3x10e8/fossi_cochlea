magic
tech sky130B
magscale 1 2
timestamp 1663021196
<< obsli1 >>
rect 1104 2159 382812 21777
<< obsm1 >>
rect 1104 1640 382971 22160
<< metal2 >>
rect 5998 23200 6054 24000
rect 13910 23200 13966 24000
rect 21822 23200 21878 24000
rect 29734 23200 29790 24000
rect 37646 23200 37702 24000
rect 45558 23200 45614 24000
rect 53470 23200 53526 24000
rect 61382 23200 61438 24000
rect 69294 23200 69350 24000
rect 77206 23200 77262 24000
rect 85118 23200 85174 24000
rect 93030 23200 93086 24000
rect 100942 23200 100998 24000
rect 108854 23200 108910 24000
rect 116766 23200 116822 24000
rect 124678 23200 124734 24000
rect 132590 23200 132646 24000
rect 140502 23200 140558 24000
rect 148414 23200 148470 24000
rect 156326 23200 156382 24000
rect 164238 23200 164294 24000
rect 172150 23200 172206 24000
rect 180062 23200 180118 24000
rect 187974 23200 188030 24000
rect 195886 23200 195942 24000
rect 203798 23200 203854 24000
rect 211710 23200 211766 24000
rect 219622 23200 219678 24000
rect 227534 23200 227590 24000
rect 235446 23200 235502 24000
rect 243358 23200 243414 24000
rect 251270 23200 251326 24000
rect 259182 23200 259238 24000
rect 267094 23200 267150 24000
rect 275006 23200 275062 24000
rect 282918 23200 282974 24000
rect 290830 23200 290886 24000
rect 298742 23200 298798 24000
rect 306654 23200 306710 24000
rect 314566 23200 314622 24000
rect 322478 23200 322534 24000
rect 330390 23200 330446 24000
rect 338302 23200 338358 24000
rect 346214 23200 346270 24000
rect 354126 23200 354182 24000
rect 362038 23200 362094 24000
rect 369950 23200 370006 24000
rect 377862 23200 377918 24000
rect 5998 0 6054 800
rect 13910 0 13966 800
rect 21822 0 21878 800
rect 29734 0 29790 800
rect 37646 0 37702 800
rect 45558 0 45614 800
rect 53470 0 53526 800
rect 61382 0 61438 800
rect 69294 0 69350 800
rect 77206 0 77262 800
rect 85118 0 85174 800
rect 93030 0 93086 800
rect 100942 0 100998 800
rect 108854 0 108910 800
rect 116766 0 116822 800
rect 124678 0 124734 800
rect 132590 0 132646 800
rect 140502 0 140558 800
rect 148414 0 148470 800
rect 156326 0 156382 800
rect 164238 0 164294 800
rect 172150 0 172206 800
rect 180062 0 180118 800
rect 187974 0 188030 800
rect 195886 0 195942 800
rect 203798 0 203854 800
rect 211710 0 211766 800
rect 219622 0 219678 800
rect 227534 0 227590 800
rect 235446 0 235502 800
rect 243358 0 243414 800
rect 251270 0 251326 800
rect 259182 0 259238 800
rect 267094 0 267150 800
rect 275006 0 275062 800
rect 282918 0 282974 800
rect 290830 0 290886 800
rect 298742 0 298798 800
rect 306654 0 306710 800
rect 314566 0 314622 800
rect 322478 0 322534 800
rect 330390 0 330446 800
rect 338302 0 338358 800
rect 346214 0 346270 800
rect 354126 0 354182 800
rect 362038 0 362094 800
rect 369950 0 370006 800
rect 377862 0 377918 800
<< obsm2 >>
rect 1582 23144 5942 23338
rect 6110 23144 13854 23338
rect 14022 23144 21766 23338
rect 21934 23144 29678 23338
rect 29846 23144 37590 23338
rect 37758 23144 45502 23338
rect 45670 23144 53414 23338
rect 53582 23144 61326 23338
rect 61494 23144 69238 23338
rect 69406 23144 77150 23338
rect 77318 23144 85062 23338
rect 85230 23144 92974 23338
rect 93142 23144 100886 23338
rect 101054 23144 108798 23338
rect 108966 23144 116710 23338
rect 116878 23144 124622 23338
rect 124790 23144 132534 23338
rect 132702 23144 140446 23338
rect 140614 23144 148358 23338
rect 148526 23144 156270 23338
rect 156438 23144 164182 23338
rect 164350 23144 172094 23338
rect 172262 23144 180006 23338
rect 180174 23144 187918 23338
rect 188086 23144 195830 23338
rect 195998 23144 203742 23338
rect 203910 23144 211654 23338
rect 211822 23144 219566 23338
rect 219734 23144 227478 23338
rect 227646 23144 235390 23338
rect 235558 23144 243302 23338
rect 243470 23144 251214 23338
rect 251382 23144 259126 23338
rect 259294 23144 267038 23338
rect 267206 23144 274950 23338
rect 275118 23144 282862 23338
rect 283030 23144 290774 23338
rect 290942 23144 298686 23338
rect 298854 23144 306598 23338
rect 306766 23144 314510 23338
rect 314678 23144 322422 23338
rect 322590 23144 330334 23338
rect 330502 23144 338246 23338
rect 338414 23144 346158 23338
rect 346326 23144 354070 23338
rect 354238 23144 361982 23338
rect 362150 23144 369894 23338
rect 370062 23144 377806 23338
rect 377974 23144 382965 23338
rect 1582 856 382965 23144
rect 1582 734 5942 856
rect 6110 734 13854 856
rect 14022 734 21766 856
rect 21934 734 29678 856
rect 29846 734 37590 856
rect 37758 734 45502 856
rect 45670 734 53414 856
rect 53582 734 61326 856
rect 61494 734 69238 856
rect 69406 734 77150 856
rect 77318 734 85062 856
rect 85230 734 92974 856
rect 93142 734 100886 856
rect 101054 734 108798 856
rect 108966 734 116710 856
rect 116878 734 124622 856
rect 124790 734 132534 856
rect 132702 734 140446 856
rect 140614 734 148358 856
rect 148526 734 156270 856
rect 156438 734 164182 856
rect 164350 734 172094 856
rect 172262 734 180006 856
rect 180174 734 187918 856
rect 188086 734 195830 856
rect 195998 734 203742 856
rect 203910 734 211654 856
rect 211822 734 219566 856
rect 219734 734 227478 856
rect 227646 734 235390 856
rect 235558 734 243302 856
rect 243470 734 251214 856
rect 251382 734 259126 856
rect 259294 734 267038 856
rect 267206 734 274950 856
rect 275118 734 282862 856
rect 283030 734 290774 856
rect 290942 734 298686 856
rect 298854 734 306598 856
rect 306766 734 314510 856
rect 314678 734 322422 856
rect 322590 734 330334 856
rect 330502 734 338246 856
rect 338414 734 346158 856
rect 346326 734 354070 856
rect 354238 734 361982 856
rect 362150 734 369894 856
rect 370062 734 377806 856
rect 377974 734 382965 856
<< metal3 >>
rect 0 22040 800 22160
rect 0 18640 800 18760
rect 0 15240 800 15360
rect 0 11840 800 11960
rect 0 8440 800 8560
rect 0 5040 800 5160
rect 0 1640 800 1760
<< obsm3 >>
rect 880 21960 382969 22133
rect 800 18840 382969 21960
rect 880 18560 382969 18840
rect 800 15440 382969 18560
rect 880 15160 382969 15440
rect 800 12040 382969 15160
rect 880 11760 382969 12040
rect 800 8640 382969 11760
rect 880 8360 382969 8640
rect 800 5240 382969 8360
rect 880 4960 382969 5240
rect 800 1840 382969 4960
rect 880 1667 382969 1840
<< metal4 >>
rect 48657 2128 48977 21808
rect 96370 2128 96690 21808
rect 144084 2128 144404 21808
rect 191797 2128 192117 21808
rect 239511 2128 239831 21808
rect 287224 2128 287544 21808
rect 334938 2128 335258 21808
rect 382651 2128 382971 21808
<< obsm4 >>
rect 110275 2483 144004 21317
rect 144484 2483 191717 21317
rect 192197 2483 239431 21317
rect 239911 2483 287144 21317
rect 287624 2483 334858 21317
rect 335338 2483 367205 21317
<< labels >>
rlabel metal2 s 13910 23200 13966 24000 6 cclk_I[0]
port 1 nsew signal output
rlabel metal2 s 61382 23200 61438 24000 6 cclk_I[1]
port 2 nsew signal output
rlabel metal2 s 108854 23200 108910 24000 6 cclk_I[2]
port 3 nsew signal output
rlabel metal2 s 156326 23200 156382 24000 6 cclk_I[3]
port 4 nsew signal output
rlabel metal2 s 203798 23200 203854 24000 6 cclk_I[4]
port 5 nsew signal output
rlabel metal2 s 251270 23200 251326 24000 6 cclk_I[5]
port 6 nsew signal output
rlabel metal2 s 298742 23200 298798 24000 6 cclk_I[6]
port 7 nsew signal output
rlabel metal2 s 346214 23200 346270 24000 6 cclk_I[7]
port 8 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 cclk_Q[0]
port 9 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 cclk_Q[1]
port 10 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 cclk_Q[2]
port 11 nsew signal output
rlabel metal2 s 156326 0 156382 800 6 cclk_Q[3]
port 12 nsew signal output
rlabel metal2 s 203798 0 203854 800 6 cclk_Q[4]
port 13 nsew signal output
rlabel metal2 s 251270 0 251326 800 6 cclk_Q[5]
port 14 nsew signal output
rlabel metal2 s 298742 0 298798 800 6 cclk_Q[6]
port 15 nsew signal output
rlabel metal2 s 346214 0 346270 800 6 cclk_Q[7]
port 16 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 clk_master
port 17 nsew signal input
rlabel metal2 s 21822 23200 21878 24000 6 clkdiv2_I[0]
port 18 nsew signal output
rlabel metal2 s 69294 23200 69350 24000 6 clkdiv2_I[1]
port 19 nsew signal output
rlabel metal2 s 116766 23200 116822 24000 6 clkdiv2_I[2]
port 20 nsew signal output
rlabel metal2 s 164238 23200 164294 24000 6 clkdiv2_I[3]
port 21 nsew signal output
rlabel metal2 s 211710 23200 211766 24000 6 clkdiv2_I[4]
port 22 nsew signal output
rlabel metal2 s 259182 23200 259238 24000 6 clkdiv2_I[5]
port 23 nsew signal output
rlabel metal2 s 306654 23200 306710 24000 6 clkdiv2_I[6]
port 24 nsew signal output
rlabel metal2 s 354126 23200 354182 24000 6 clkdiv2_I[7]
port 25 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 clkdiv2_Q[0]
port 26 nsew signal output
rlabel metal2 s 69294 0 69350 800 6 clkdiv2_Q[1]
port 27 nsew signal output
rlabel metal2 s 116766 0 116822 800 6 clkdiv2_Q[2]
port 28 nsew signal output
rlabel metal2 s 164238 0 164294 800 6 clkdiv2_Q[3]
port 29 nsew signal output
rlabel metal2 s 211710 0 211766 800 6 clkdiv2_Q[4]
port 30 nsew signal output
rlabel metal2 s 259182 0 259238 800 6 clkdiv2_Q[5]
port 31 nsew signal output
rlabel metal2 s 306654 0 306710 800 6 clkdiv2_Q[6]
port 32 nsew signal output
rlabel metal2 s 354126 0 354182 800 6 clkdiv2_Q[7]
port 33 nsew signal output
rlabel metal2 s 29734 23200 29790 24000 6 comp_high_I[0]
port 34 nsew signal input
rlabel metal2 s 77206 23200 77262 24000 6 comp_high_I[1]
port 35 nsew signal input
rlabel metal2 s 124678 23200 124734 24000 6 comp_high_I[2]
port 36 nsew signal input
rlabel metal2 s 172150 23200 172206 24000 6 comp_high_I[3]
port 37 nsew signal input
rlabel metal2 s 219622 23200 219678 24000 6 comp_high_I[4]
port 38 nsew signal input
rlabel metal2 s 267094 23200 267150 24000 6 comp_high_I[5]
port 39 nsew signal input
rlabel metal2 s 314566 23200 314622 24000 6 comp_high_I[6]
port 40 nsew signal input
rlabel metal2 s 362038 23200 362094 24000 6 comp_high_I[7]
port 41 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 comp_high_Q[0]
port 42 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 comp_high_Q[1]
port 43 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 comp_high_Q[2]
port 44 nsew signal input
rlabel metal2 s 172150 0 172206 800 6 comp_high_Q[3]
port 45 nsew signal input
rlabel metal2 s 219622 0 219678 800 6 comp_high_Q[4]
port 46 nsew signal input
rlabel metal2 s 267094 0 267150 800 6 comp_high_Q[5]
port 47 nsew signal input
rlabel metal2 s 314566 0 314622 800 6 comp_high_Q[6]
port 48 nsew signal input
rlabel metal2 s 362038 0 362094 800 6 comp_high_Q[7]
port 49 nsew signal input
rlabel metal2 s 45558 23200 45614 24000 6 cos_out[0]
port 50 nsew signal output
rlabel metal2 s 93030 23200 93086 24000 6 cos_out[1]
port 51 nsew signal output
rlabel metal2 s 140502 23200 140558 24000 6 cos_out[2]
port 52 nsew signal output
rlabel metal2 s 187974 23200 188030 24000 6 cos_out[3]
port 53 nsew signal output
rlabel metal2 s 235446 23200 235502 24000 6 cos_out[4]
port 54 nsew signal output
rlabel metal2 s 282918 23200 282974 24000 6 cos_out[5]
port 55 nsew signal output
rlabel metal2 s 330390 23200 330446 24000 6 cos_out[6]
port 56 nsew signal output
rlabel metal2 s 377862 23200 377918 24000 6 cos_out[7]
port 57 nsew signal output
rlabel metal2 s 5998 23200 6054 24000 6 fb1_I[0]
port 58 nsew signal output
rlabel metal2 s 53470 23200 53526 24000 6 fb1_I[1]
port 59 nsew signal output
rlabel metal2 s 100942 23200 100998 24000 6 fb1_I[2]
port 60 nsew signal output
rlabel metal2 s 148414 23200 148470 24000 6 fb1_I[3]
port 61 nsew signal output
rlabel metal2 s 195886 23200 195942 24000 6 fb1_I[4]
port 62 nsew signal output
rlabel metal2 s 243358 23200 243414 24000 6 fb1_I[5]
port 63 nsew signal output
rlabel metal2 s 290830 23200 290886 24000 6 fb1_I[6]
port 64 nsew signal output
rlabel metal2 s 338302 23200 338358 24000 6 fb1_I[7]
port 65 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 fb1_Q[0]
port 66 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 fb1_Q[1]
port 67 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 fb1_Q[2]
port 68 nsew signal output
rlabel metal2 s 148414 0 148470 800 6 fb1_Q[3]
port 69 nsew signal output
rlabel metal2 s 195886 0 195942 800 6 fb1_Q[4]
port 70 nsew signal output
rlabel metal2 s 243358 0 243414 800 6 fb1_Q[5]
port 71 nsew signal output
rlabel metal2 s 290830 0 290886 800 6 fb1_Q[6]
port 72 nsew signal output
rlabel metal2 s 338302 0 338358 800 6 fb1_Q[7]
port 73 nsew signal output
rlabel metal2 s 37646 23200 37702 24000 6 phi1b_dig_I[0]
port 74 nsew signal input
rlabel metal2 s 85118 23200 85174 24000 6 phi1b_dig_I[1]
port 75 nsew signal input
rlabel metal2 s 132590 23200 132646 24000 6 phi1b_dig_I[2]
port 76 nsew signal input
rlabel metal2 s 180062 23200 180118 24000 6 phi1b_dig_I[3]
port 77 nsew signal input
rlabel metal2 s 227534 23200 227590 24000 6 phi1b_dig_I[4]
port 78 nsew signal input
rlabel metal2 s 275006 23200 275062 24000 6 phi1b_dig_I[5]
port 79 nsew signal input
rlabel metal2 s 322478 23200 322534 24000 6 phi1b_dig_I[6]
port 80 nsew signal input
rlabel metal2 s 369950 23200 370006 24000 6 phi1b_dig_I[7]
port 81 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 phi1b_dig_Q[0]
port 82 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 phi1b_dig_Q[1]
port 83 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 phi1b_dig_Q[2]
port 84 nsew signal input
rlabel metal2 s 180062 0 180118 800 6 phi1b_dig_Q[3]
port 85 nsew signal input
rlabel metal2 s 227534 0 227590 800 6 phi1b_dig_Q[4]
port 86 nsew signal input
rlabel metal2 s 275006 0 275062 800 6 phi1b_dig_Q[5]
port 87 nsew signal input
rlabel metal2 s 322478 0 322534 800 6 phi1b_dig_Q[6]
port 88 nsew signal input
rlabel metal2 s 369950 0 370006 800 6 phi1b_dig_Q[7]
port 89 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 read_out_I[0]
port 90 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 read_out_I[1]
port 91 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 read_out_Q[0]
port 92 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 read_out_Q[1]
port 93 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 rstb
port 94 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 sin_out[0]
port 95 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 sin_out[1]
port 96 nsew signal output
rlabel metal2 s 140502 0 140558 800 6 sin_out[2]
port 97 nsew signal output
rlabel metal2 s 187974 0 188030 800 6 sin_out[3]
port 98 nsew signal output
rlabel metal2 s 235446 0 235502 800 6 sin_out[4]
port 99 nsew signal output
rlabel metal2 s 282918 0 282974 800 6 sin_out[5]
port 100 nsew signal output
rlabel metal2 s 330390 0 330446 800 6 sin_out[6]
port 101 nsew signal output
rlabel metal2 s 377862 0 377918 800 6 sin_out[7]
port 102 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 ud_en
port 103 nsew signal input
rlabel metal4 s 48657 2128 48977 21808 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 144084 2128 144404 21808 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 239511 2128 239831 21808 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 334938 2128 335258 21808 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 96370 2128 96690 21808 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 191797 2128 192117 21808 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 287224 2128 287544 21808 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 382651 2128 382971 21808 6 vssd1
port 105 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 384000 24000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15155838
string GDS_FILE /local_disk/fossi_cochlea/openlane/digital_unison/runs/22_09_12_15_14/results/signoff/digital_unison.magic.gds
string GDS_START 644014
<< end >>

