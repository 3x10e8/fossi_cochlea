VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital_unison
  CLASS BLOCK ;
  FOREIGN digital_unison ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 250.000 ;
  PIN cclk_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END cclk_I[0]
  PIN cclk_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END cclk_I[1]
  PIN cclk_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 246.000 203.230 250.000 ;
    END
  END cclk_Q[0]
  PIN cclk_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 119.040 300.000 119.640 ;
    END
  END cclk_Q[1]
  PIN clk_master
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END clk_master
  PIN clkdiv2_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 246.000 177.470 250.000 ;
    END
  END clkdiv2_I[0]
  PIN clkdiv2_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END clkdiv2_I[1]
  PIN clkdiv2_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 246.000 64.770 250.000 ;
    END
  END clkdiv2_Q[0]
  PIN clkdiv2_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 176.840 300.000 177.440 ;
    END
  END clkdiv2_Q[1]
  PIN comp_high_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END comp_high_I[0]
  PIN comp_high_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 246.000 286.950 250.000 ;
    END
  END comp_high_I[1]
  PIN comp_high_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 207.440 300.000 208.040 ;
    END
  END comp_high_Q[0]
  PIN comp_high_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 246.000 93.750 250.000 ;
    END
  END comp_high_Q[1]
  PIN cos_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END cos_out[0]
  PIN cos_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 30.640 300.000 31.240 ;
    END
  END cos_out[1]
  PIN cos_outb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END cos_outb[0]
  PIN cos_outb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 146.240 300.000 146.840 ;
    END
  END cos_outb[1]
  PIN fb1_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END fb1_I[0]
  PIN fb1_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END fb1_I[1]
  PIN fb1_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 246.000 232.210 250.000 ;
    END
  END fb1_Q[0]
  PIN fb1_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END fb1_Q[1]
  PIN fb2_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END fb2_I[0]
  PIN fb2_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 246.000 39.010 250.000 ;
    END
  END fb2_I[1]
  PIN fb2_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END fb2_Q[0]
  PIN fb2_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 246.000 261.190 250.000 ;
    END
  END fb2_Q[1]
  PIN phi1b_dig_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 0.040 300.000 0.640 ;
    END
  END phi1b_dig_I[0]
  PIN phi1b_dig_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END phi1b_dig_I[1]
  PIN phi1b_dig_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END phi1b_dig_Q[0]
  PIN phi1b_dig_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END phi1b_dig_Q[1]
  PIN read_out_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 61.240 300.000 61.840 ;
    END
  END read_out_I[0]
  PIN read_out_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END read_out_I[1]
  PIN read_out_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END read_out_Q[0]
  PIN read_out_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 234.640 300.000 235.240 ;
    END
  END read_out_Q[1]
  PIN rstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 246.000 119.510 250.000 ;
    END
  END rstb
  PIN sin_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 246.000 148.490 250.000 ;
    END
  END sin_out[0]
  PIN sin_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END sin_out[1]
  PIN sin_outb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END sin_outb[0]
  PIN sin_outb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 246.000 10.030 250.000 ;
    END
  END sin_outb[1]
  PIN ud_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 88.440 300.000 89.040 ;
    END
  END ud_en
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 236.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 236.725 ;
      LAYER met1 ;
        RECT 0.070 2.760 299.390 244.080 ;
      LAYER met2 ;
        RECT 0.090 245.720 9.470 246.570 ;
        RECT 10.310 245.720 38.450 246.570 ;
        RECT 39.290 245.720 64.210 246.570 ;
        RECT 65.050 245.720 93.190 246.570 ;
        RECT 94.030 245.720 118.950 246.570 ;
        RECT 119.790 245.720 147.930 246.570 ;
        RECT 148.770 245.720 176.910 246.570 ;
        RECT 177.750 245.720 202.670 246.570 ;
        RECT 203.510 245.720 231.650 246.570 ;
        RECT 232.490 245.720 260.630 246.570 ;
        RECT 261.470 245.720 286.390 246.570 ;
        RECT 287.230 245.720 299.360 246.570 ;
        RECT 0.090 4.280 299.360 245.720 ;
        RECT 0.650 0.155 25.570 4.280 ;
        RECT 26.410 0.155 54.550 4.280 ;
        RECT 55.390 0.155 80.310 4.280 ;
        RECT 81.150 0.155 109.290 4.280 ;
        RECT 110.130 0.155 138.270 4.280 ;
        RECT 139.110 0.155 164.030 4.280 ;
        RECT 164.870 0.155 193.010 4.280 ;
        RECT 193.850 0.155 218.770 4.280 ;
        RECT 219.610 0.155 247.750 4.280 ;
        RECT 248.590 0.155 276.730 4.280 ;
        RECT 277.570 0.155 299.360 4.280 ;
      LAYER met3 ;
        RECT 0.065 235.640 298.935 248.700 ;
        RECT 0.065 234.240 295.600 235.640 ;
        RECT 0.065 232.240 298.935 234.240 ;
        RECT 4.400 230.840 298.935 232.240 ;
        RECT 0.065 208.440 298.935 230.840 ;
        RECT 0.065 207.040 295.600 208.440 ;
        RECT 0.065 205.040 298.935 207.040 ;
        RECT 4.400 203.640 298.935 205.040 ;
        RECT 0.065 177.840 298.935 203.640 ;
        RECT 0.065 176.440 295.600 177.840 ;
        RECT 0.065 174.440 298.935 176.440 ;
        RECT 4.400 173.040 298.935 174.440 ;
        RECT 0.065 147.240 298.935 173.040 ;
        RECT 4.400 145.840 295.600 147.240 ;
        RECT 0.065 120.040 298.935 145.840 ;
        RECT 0.065 118.640 295.600 120.040 ;
        RECT 0.065 116.640 298.935 118.640 ;
        RECT 4.400 115.240 298.935 116.640 ;
        RECT 0.065 89.440 298.935 115.240 ;
        RECT 0.065 88.040 295.600 89.440 ;
        RECT 0.065 86.040 298.935 88.040 ;
        RECT 4.400 84.640 298.935 86.040 ;
        RECT 0.065 62.240 298.935 84.640 ;
        RECT 0.065 60.840 295.600 62.240 ;
        RECT 0.065 58.840 298.935 60.840 ;
        RECT 4.400 57.440 298.935 58.840 ;
        RECT 0.065 31.640 298.935 57.440 ;
        RECT 0.065 30.240 295.600 31.640 ;
        RECT 0.065 28.240 298.935 30.240 ;
        RECT 4.400 26.840 298.935 28.240 ;
        RECT 0.065 1.040 298.935 26.840 ;
        RECT 0.065 0.175 295.600 1.040 ;
      LAYER met4 ;
        RECT 2.135 237.280 288.585 248.705 ;
        RECT 2.135 10.240 20.640 237.280 ;
        RECT 23.040 10.240 97.440 237.280 ;
        RECT 99.840 10.240 174.240 237.280 ;
        RECT 176.640 10.240 251.040 237.280 ;
        RECT 253.440 10.240 288.585 237.280 ;
        RECT 2.135 1.535 288.585 10.240 ;
  END
END digital_unison
END LIBRARY

