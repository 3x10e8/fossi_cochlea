magic
tech sky130A
magscale 1 2
timestamp 1654657422
<< metal3 >>
rect -710 2655 2678 2688
rect -710 -217 -677 2655
rect 281 2397 1997 2655
rect -419 2366 2387 2397
rect -419 1541 -388 2366
rect -68 1541 2036 2046
rect 2356 1541 2387 2366
rect -419 1221 2387 1541
rect -419 376 -388 1221
rect -68 376 2036 1221
rect 2356 376 2387 1221
rect -419 56 2387 376
rect -419 -217 -388 56
rect -68 -58 2036 56
rect -68 -60 276 -58
rect -710 -366 -388 -217
rect -44 -366 276 -60
rect 824 -366 1144 -58
rect 1692 -60 2036 -58
rect 1692 -366 2012 -60
rect 2356 -217 2387 56
rect 2645 -217 2678 2655
rect 2356 -366 2678 -217
<< via3 >>
rect -677 2397 281 2655
rect 1997 2397 2645 2655
rect -677 -217 -419 2397
rect 2387 -217 2645 2397
<< mimcap >>
rect -16 1786 1984 1994
rect -16 202 192 1786
rect 336 1066 912 1642
rect 1056 1066 1632 1642
rect 336 346 912 922
rect 1056 346 1632 922
rect 1776 202 1984 1786
rect -16 -6 1984 202
<< mimcapcontact >>
rect 192 1642 1776 1786
rect 192 1066 336 1642
rect 912 1066 1056 1642
rect 1632 1066 1776 1642
rect 192 922 1776 1066
rect 192 346 336 922
rect 912 346 1056 922
rect 1632 346 1776 922
rect 192 202 1776 346
<< metal4 >>
rect -685 2662 -412 2686
rect -708 2389 -684 2662
rect 281 2390 282 2662
rect 1996 2390 1997 2662
rect -44 1942 2012 2022
rect -45 1786 2012 1942
rect -45 1782 192 1786
rect -44 1074 192 1782
rect -45 914 192 1074
rect 336 1066 912 1642
rect 1056 1066 1632 1642
rect -44 206 192 914
rect 336 346 912 922
rect 1056 346 1632 922
rect -45 202 192 206
rect 1776 202 2012 1786
rect -45 46 2012 202
rect -44 -34 2012 46
rect -684 -366 -412 -217
rect 36 -366 196 -34
rect 904 -366 1064 -34
rect 1772 -366 1932 -34
rect 2380 -366 2652 -217
<< via4 >>
rect -684 2655 281 2662
rect -684 -217 -677 2655
rect -677 2397 281 2655
rect -677 -217 -419 2397
rect -419 2390 281 2397
rect 1997 2655 2652 2662
rect 1997 2397 2645 2655
rect 1997 2390 2387 2397
rect -419 -217 -412 2390
rect 2380 -217 2387 2390
rect 2387 -217 2645 2397
rect 2645 -217 2652 2655
<< mimcap2 >>
rect -16 1812 1984 1994
rect -16 1576 166 1812
rect 402 1576 516 1812
rect 752 1576 866 1812
rect 1102 1576 1216 1812
rect 1452 1576 1566 1812
rect 1802 1576 1984 1812
rect -16 1462 1984 1576
rect -16 1226 166 1462
rect 402 1226 866 1462
rect 1102 1226 1566 1462
rect 1802 1226 1984 1462
rect -16 1112 1984 1226
rect -16 876 166 1112
rect 402 876 516 1112
rect 752 876 866 1112
rect 1102 876 1216 1112
rect 1452 876 1566 1112
rect 1802 876 1984 1112
rect -16 762 1984 876
rect -16 526 166 762
rect 402 526 866 762
rect 1102 526 1566 762
rect 1802 526 1984 762
rect -16 412 1984 526
rect -16 176 166 412
rect 402 176 516 412
rect 752 176 866 412
rect 1102 176 1216 412
rect 1452 176 1566 412
rect 1802 176 1984 412
rect -16 -6 1984 176
<< mimcap2contact >>
rect 166 1576 402 1812
rect 516 1576 752 1812
rect 866 1576 1102 1812
rect 1216 1576 1452 1812
rect 1566 1576 1802 1812
rect 166 1226 402 1462
rect 866 1226 1102 1462
rect 1566 1226 1802 1462
rect 166 876 402 1112
rect 516 876 752 1112
rect 866 876 1102 1112
rect 1216 876 1452 1112
rect 1566 876 1802 1112
rect 166 526 402 762
rect 866 526 1102 762
rect 1566 526 1802 762
rect 166 176 402 412
rect 516 176 752 412
rect 866 176 1102 412
rect 1216 176 1452 412
rect 1566 176 1802 412
<< metal5 >>
rect -708 2662 2676 2686
rect -708 -217 -684 2662
rect 281 2390 1997 2662
rect -412 2366 2380 2390
rect -412 1541 -388 2366
rect -68 1812 2036 2046
rect -68 1576 166 1812
rect 402 1576 516 1812
rect 752 1576 866 1812
rect 1102 1576 1216 1812
rect 1452 1576 1566 1812
rect 1802 1576 2036 1812
rect -68 1541 2036 1576
rect 2356 1541 2380 2366
rect -412 1462 2380 1541
rect -412 1226 166 1462
rect 402 1226 866 1462
rect 1102 1226 1566 1462
rect 1802 1226 2380 1462
rect -412 1221 2380 1226
rect -412 376 -388 1221
rect -68 1112 2036 1221
rect -68 876 166 1112
rect 402 876 516 1112
rect 752 876 866 1112
rect 1102 876 1216 1112
rect 1452 876 1566 1112
rect 1802 876 2036 1112
rect -68 762 2036 876
rect -68 526 166 762
rect 402 526 866 762
rect 1102 526 1566 762
rect 1802 526 2036 762
rect -68 412 2036 526
rect -68 376 166 412
rect -412 176 166 376
rect 402 176 516 412
rect 752 176 866 412
rect 1102 176 1216 412
rect 1452 176 1566 412
rect 1802 376 2036 412
rect 2356 376 2380 1221
rect 1802 176 2380 376
rect -412 56 2380 176
rect -412 -217 -388 56
rect -68 -58 2036 56
rect -68 -60 276 -58
rect -708 -366 -388 -217
rect -44 -366 276 -60
rect 824 -366 1144 -58
rect 1692 -60 2036 -58
rect 1692 -366 2012 -60
rect 2356 -217 2380 56
rect 2652 -217 2676 2662
rect 2356 -366 2676 -217
<< end >>
