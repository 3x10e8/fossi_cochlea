magic
tech sky130A
timestamp 1654236220
use cap_10_10__side_x2  cap_10_10__side_x2_0
timestamp 1654233531
transform 1 0 -1363 0 1 2116
box -34 -374 1363 1368
use cap_10_10__side_x2  cap_10_10__side_x2_1
timestamp 1654233531
transform 1 0 -1363 0 1 374
box -34 -374 1363 1368
use cap_10_10__side_x2  cap_10_10__side_x2_2
timestamp 1654233531
transform 0 -1 1368 1 0 -1363
box -34 -374 1363 1368
use cap_10_10__side_x2  cap_10_10__side_x2_3
timestamp 1654233531
transform 0 -1 3110 1 0 -1363
box -34 -374 1363 1368
use cap_10_10__side_x2  cap_10_10__side_x2_4
timestamp 1654233531
transform -1 0 4847 0 -1 1368
box -34 -374 1363 1368
use cap_10_10__side_x2  cap_10_10__side_x2_5
timestamp 1654233531
transform -1 0 4847 0 -1 3110
box -34 -374 1363 1368
use cap_10_10__side_x2  cap_10_10__side_x2_6
timestamp 1654233531
transform 0 1 2116 -1 0 4847
box -34 -374 1363 1368
use cap_10_10__side_x2  cap_10_10__side_x2_7
timestamp 1654233531
transform 0 1 374 -1 0 4847
box -34 -374 1363 1368
use cap_10_10_edge_x2  cap_10_10_edge_x2_0
timestamp 1654233587
transform 0 1 -1368 -1 0 4847
box -34 -29 1363 1368
use cap_10_10_edge_x2  cap_10_10_edge_x2_1
timestamp 1654233587
transform -1 0 4847 0 -1 4852
box -34 -29 1363 1368
use cap_10_10_edge_x2  cap_10_10_edge_x2_2
timestamp 1654233587
transform 0 -1 4852 1 0 -1363
box -34 -29 1363 1368
use cap_10_10_edge_x2  cap_10_10_edge_x2_3
timestamp 1654233587
transform 1 0 -1363 0 1 -1368
box -34 -29 1363 1368
use cap_10_10_x2  cap_10_10_x2_0
array 0 1 1742 0 1 1742
timestamp 1654233242
transform 1 0 379 0 1 374
box -379 -374 1363 1368
<< end >>
