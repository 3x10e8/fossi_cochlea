magic
tech sky130B
magscale 1 2
timestamp 1663910114
<< metal1 >>
rect 406162 36972 406274 36978
rect 406162 36872 406168 36972
rect 406268 36872 407704 36972
rect 406162 36866 406274 36872
rect 406462 32994 406575 33000
rect 406462 32893 406468 32994
rect 406569 32893 407704 32994
rect 406462 32887 406575 32893
rect 407366 28900 407372 29000
rect 407472 28900 407704 29000
rect 407066 24900 407072 25000
rect 407172 24900 407704 25000
rect 406766 20900 406772 21000
rect 406872 20900 407704 21000
rect 406466 16900 406472 17000
rect 406572 16900 407704 17000
rect 406166 12900 406172 13000
rect 406272 12900 407700 13000
<< via1 >>
rect 406168 36872 406268 36972
rect 406468 32893 406569 32994
rect 407372 28900 407472 29000
rect 407072 24900 407172 25000
rect 406772 20900 406872 21000
rect 406472 16900 406572 17000
rect 406172 12900 406272 13000
<< metal2 >>
rect 5078 35378 5134 36978
rect 13542 35378 13598 36978
rect 22006 35378 22062 36978
rect 30470 35378 30526 36978
rect 38934 35378 38990 36978
rect 47398 35378 47454 36978
rect 55862 35378 55918 36978
rect 64326 35378 64382 36978
rect 72790 35378 72846 36978
rect 81254 35378 81310 36978
rect 89718 35378 89774 36978
rect 98182 35378 98238 36978
rect 106646 35378 106702 36978
rect 115110 35378 115166 36978
rect 123574 35378 123630 36978
rect 132038 35378 132094 36978
rect 140502 35378 140558 36978
rect 148966 35378 149022 36978
rect 157430 35378 157486 36978
rect 165894 35378 165950 36978
rect 174358 35378 174414 36978
rect 182822 35378 182878 36978
rect 191286 35378 191342 36978
rect 199750 35378 199806 36978
rect 208214 35378 208270 36978
rect 216678 35378 216734 36978
rect 225142 35378 225198 36978
rect 233606 35378 233662 36978
rect 242070 35378 242126 36978
rect 250534 35378 250590 36978
rect 258998 35378 259054 36978
rect 267462 35378 267518 36978
rect 275926 35378 275982 36978
rect 284390 35378 284446 36978
rect 292854 35378 292910 36978
rect 301318 35378 301374 36978
rect 309782 35378 309838 36978
rect 318246 35378 318302 36978
rect 326710 35378 326766 36978
rect 335174 35378 335230 36978
rect 343638 35378 343694 36978
rect 352102 35378 352158 36978
rect 360566 35378 360622 36978
rect 369030 35378 369086 36978
rect 377494 35378 377550 36978
rect 385958 35378 386014 36978
rect 394422 35378 394478 36978
rect 402886 35378 402942 36978
rect 406162 36972 406274 36978
rect 406162 36872 406168 36972
rect 406268 36872 406274 36972
rect 406162 36866 406274 36872
rect 406168 31573 406268 36866
rect 406462 32994 406575 33000
rect 406462 32893 406468 32994
rect 406569 32893 406575 32994
rect 406462 32887 406575 32893
rect 406168 31483 406173 31573
rect 406263 31483 406268 31573
rect 406168 31478 406268 31483
rect 406468 32010 406569 32887
rect 406173 31474 406263 31478
rect 406468 31373 406568 32010
rect 406468 31283 406473 31373
rect 406563 31283 406568 31373
rect 406468 31278 406568 31283
rect 406473 31274 406563 31278
rect 407377 30824 407467 30828
rect 407372 30819 407472 30824
rect 407372 30729 407377 30819
rect 407467 30729 407472 30819
rect 407077 30624 407167 30628
rect 407072 30619 407172 30624
rect 407072 30529 407077 30619
rect 407167 30529 407172 30619
rect 406777 30424 406867 30428
rect 406772 30419 406872 30424
rect 406772 30329 406777 30419
rect 406867 30329 406872 30419
rect 406477 29487 406567 29491
rect 406472 29482 406572 29487
rect 406472 29392 406477 29482
rect 406567 29392 406572 29482
rect 406168 29291 406276 29300
rect 406168 29201 406177 29291
rect 406267 29201 406276 29291
rect 406168 29196 406276 29201
rect 406172 13000 406272 29196
rect 406472 17000 406572 29392
rect 406772 21000 406872 30329
rect 407072 25000 407172 30529
rect 407372 29000 407472 30729
rect 407372 28894 407472 28900
rect 407072 24894 407172 24900
rect 406772 20894 406872 20900
rect 406472 16894 406572 16900
rect 406172 12894 406272 12900
<< via2 >>
rect 406173 31483 406263 31573
rect 406473 31283 406563 31373
rect 407377 30729 407467 30819
rect 407077 30529 407167 30619
rect 406777 30329 406867 30419
rect 406477 29392 406567 29482
rect 406177 29201 406267 29291
<< metal3 >>
rect 406168 31573 406268 31578
rect 406168 31483 406173 31573
rect 406263 31483 406268 31573
rect 406168 31478 406268 31483
rect 406170 31373 406568 31378
rect 406170 31283 406473 31373
rect 406563 31283 406568 31373
rect 406170 31278 406568 31283
rect 406172 30819 407472 30824
rect 406172 30729 407377 30819
rect 407467 30729 407472 30819
rect 406172 30724 407472 30729
rect 406172 30619 407172 30624
rect 406172 30529 407077 30619
rect 407167 30529 407172 30619
rect 406172 30524 407172 30529
rect 406168 30419 406872 30424
rect 406168 30329 406777 30419
rect 406867 30329 406872 30419
rect 406168 30324 406872 30329
rect 406154 29482 406572 29487
rect 406154 29392 406477 29482
rect 406567 29392 406572 29482
rect 406154 29387 406572 29392
rect 406172 29291 406272 29296
rect 406172 29201 406177 29291
rect 406267 29201 406272 29291
rect 406172 29196 406272 29201
use filter_p_m  filter_p_m_0
array 0 7 50784 0 0 13945
timestamp 1663891137
transform 1 0 26 0 1 -162
box -26 -328 50758 37140
<< labels >>
flabel metal2 5078 35378 5134 36978 1 FreeSans 1600 0 0 0 fb1[0]
port 1 n default input
flabel metal2 55862 35378 55918 36978 1 FreeSans 1600 0 0 0 fb1[1]
port 2 n default input
flabel metal2 106646 35378 106702 36978 1 FreeSans 1600 0 0 0 fb1[2]
port 3 n default input
flabel metal2 157430 35378 157486 36978 1 FreeSans 1600 0 0 0 fb1[3]
port 4 n default input
flabel metal2 208214 35378 208270 36978 1 FreeSans 1600 0 0 0 fb1[4]
port 5 n default input
flabel metal2 258998 35378 259054 36978 1 FreeSans 1600 0 0 0 fb1[5]
port 6 n default input
flabel metal2 309782 35378 309838 36978 1 FreeSans 1600 0 0 0 fb1[6]
port 7 n default input
flabel metal2 360566 35378 360622 36978 1 FreeSans 1600 0 0 0 fb1[7]
port 8 n default input
flabel metal2 13542 35378 13598 36978 1 FreeSans 1600 0 0 0 cclk[0]
port 9 n default input
flabel metal2 64326 35378 64382 36978 1 FreeSans 1600 0 0 0 cclk[1]
port 10 n default input
flabel metal2 115110 35378 115166 36978 1 FreeSans 1600 0 0 0 cclk[2]
port 11 n default input
flabel metal2 165894 35378 165950 36978 1 FreeSans 1600 0 0 0 cclk[3]
port 12 n default input
flabel metal2 216678 35378 216734 36978 1 FreeSans 1600 0 0 0 cclk[4]
port 13 n default input
flabel metal2 267462 35378 267518 36978 1 FreeSans 1600 0 0 0 cclk[5]
port 14 n default input
flabel metal2 318246 35378 318302 36978 1 FreeSans 1600 0 0 0 cclk[6]
port 15 n default input
flabel metal2 369030 35378 369086 36978 1 FreeSans 1600 0 0 0 cclk[7]
port 16 n default input
flabel metal2 22006 35378 22062 36978 1 FreeSans 1600 0 0 0 div2[0]
port 17 n default input
flabel metal2 72790 35378 72846 36978 1 FreeSans 1600 0 0 0 div2[1]
port 18 n default input
flabel metal2 123574 35378 123630 36978 1 FreeSans 1600 0 0 0 div2[2]
port 19 n default input
flabel metal2 174358 35378 174414 36978 1 FreeSans 1600 0 0 0 div2[3]
port 20 n default input
flabel metal2 225142 35378 225198 36978 1 FreeSans 1600 0 0 0 div2[4]
port 21 n default input
flabel metal2 275926 35378 275982 36978 1 FreeSans 1600 0 0 0 div2[5]
port 22 n default input
flabel metal2 326710 35378 326766 36978 1 FreeSans 1600 0 0 0 div2[6]
port 23 n default input
flabel metal2 377494 35378 377550 36978 1 FreeSans 1600 0 0 0 div2[7]
port 24 n default input
flabel metal2 30470 35378 30526 36978 1 FreeSans 1600 0 0 0 high_buf[0]
port 25 n default output
flabel metal2 81254 35378 81310 36978 1 FreeSans 1600 0 0 0 high_buf[1]
port 26 n default output
flabel metal2 132038 35378 132094 36978 1 FreeSans 1600 0 0 0 high_buf[2]
port 27 n default output
flabel metal2 182822 35378 182878 36978 1 FreeSans 1600 0 0 0 high_buf[3]
port 28 n default output
flabel metal2 233606 35378 233662 36978 1 FreeSans 1600 0 0 0 high_buf[4]
port 29 n default output
flabel metal2 284390 35378 284446 36978 1 FreeSans 1600 0 0 0 high_buf[5]
port 30 n default output
flabel metal2 335174 35378 335230 36978 1 FreeSans 1600 0 0 0 high_buf[6]
port 31 n default output
flabel metal2 385958 35378 386014 36978 1 FreeSans 1600 0 0 0 high_buf[7]
port 32 n default output
flabel metal2 38934 35378 38990 36978 1 FreeSans 1600 0 0 0 phi1b_dig[0]
port 33 n default output
flabel metal2 89718 35378 89774 36978 1 FreeSans 1600 0 0 0 phi1b_dig[1]
port 34 n default output
flabel metal2 140502 35378 140558 36978 1 FreeSans 1600 0 0 0 phi1b_dig[2]
port 35 n default output
flabel metal2 191286 35378 191342 36978 1 FreeSans 1600 0 0 0 phi1b_dig[3]
port 36 n default output
flabel metal2 242070 35378 242126 36978 1 FreeSans 1600 0 0 0 phi1b_dig[4]
port 37 n default output
flabel metal2 292854 35378 292910 36978 1 FreeSans 1600 0 0 0 phi1b_dig[5]
port 38 n default output
flabel metal2 343638 35378 343694 36978 1 FreeSans 1600 0 0 0 phi1b_dig[6]
port 39 n default output
flabel metal2 394422 35378 394478 36978 1 FreeSans 1600 0 0 0 phi1b_dig[7]
port 40 n default output
flabel metal2 47398 35378 47454 36978 1 FreeSans 1600 0 0 0 lo[0]
port 41 n default input
flabel metal2 98182 35378 98238 36978 1 FreeSans 1600 0 0 0 lo[1]
port 42 n default input
flabel metal2 148966 35378 149022 36978 1 FreeSans 1600 0 0 0 lo[2]
port 43 n default input
flabel metal2 199750 35378 199806 36978 1 FreeSans 1600 0 0 0 lo[3]
port 44 n default input
flabel metal2 250534 35378 250590 36978 1 FreeSans 1600 0 0 0 lo[4]
port 45 n default input
flabel metal2 301318 35378 301374 36978 1 FreeSans 1600 0 0 0 lo[5]
port 46 n default input
flabel metal2 352102 35378 352158 36978 1 FreeSans 1600 0 0 0 lo[6]
port 47 n default input
flabel metal2 402886 35378 402942 36978 1 FreeSans 1600 0 0 0 lo[7]
port 48 n default input
flabel metal1 406268 36872 407704 36972 1 FreeSans 1600 0 0 0 vnb
port 49 n default bidirectional
flabel metal1 406569 32893 407704 32994 1 FreeSans 1600 0 0 0 vpb
port 50 n default bidirectional
flabel metal1 407472 28900 407704 29000 1 FreeSans 1600 0 0 0 vccd1
port 51 n power bidirectional
flabel metal1 407172 24900 407704 25000 1 FreeSans 1600 0 0 0 th1
port 52 n default bidirectional
flabel metal1 406872 20900 407704 21000 1 FreeSans 1600 0 0 0 th2
port 53 n default bidirectional
flabel metal1 406572 16900 407704 17000 1 FreeSans 1600 0 0 0 vssd1
port 54 n ground bidirectional
flabel metal1 406272 12900 407700 13000 1 FreeSans 1600 0 0 0 vdda1
port 55 n power bidirectional
<< end >>
