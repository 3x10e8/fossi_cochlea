magic
tech sky130B
magscale 1 2
timestamp 1663630899
<< nwell >>
rect 1267 724 1597 1115
rect 1283 9 1613 29
rect 2073 28 3298 349
rect 1106 -173 1613 9
rect 1283 -362 1613 -173
rect -1589 -721 -1083 -534
rect 2236 -1050 3294 -795
<< poly >>
rect -1492 -385 -1355 -349
rect -1492 -989 -1355 -953
<< viali >>
rect 73 291 107 325
rect 72 -1663 106 -1629
<< metal1 >>
rect 635 1128 884 1224
rect 1378 1203 1434 1214
rect 1378 1151 1380 1203
rect 1432 1151 1434 1203
rect 1378 1140 1434 1151
rect 2299 1203 2355 1214
rect 2299 1151 2301 1203
rect 2353 1151 2355 1203
rect 2299 1140 2355 1151
rect 3217 1205 3273 1216
rect 3217 1153 3219 1205
rect 3271 1153 3273 1205
rect 3217 1142 3273 1153
rect -1661 450 -1078 468
rect -1661 398 -1546 450
rect -1494 398 -1078 450
rect -1661 371 -1078 398
rect 635 371 731 1128
rect 3032 784 3080 968
rect 906 705 962 716
rect 906 653 908 705
rect 960 653 962 705
rect 906 642 962 653
rect 1813 661 1869 672
rect 1813 609 1815 661
rect 1867 609 1869 661
rect 1813 598 1869 609
rect 2759 660 2815 671
rect 2759 608 2761 660
rect 2813 608 2815 660
rect 2759 597 2815 608
rect 59 334 124 337
rect 59 282 66 334
rect 118 282 124 334
rect 3032 296 3080 480
rect 59 278 124 282
rect 1378 116 1434 127
rect 1378 64 1380 116
rect 1432 64 1434 116
rect 1378 53 1434 64
rect 2300 114 2356 125
rect 2300 62 2302 114
rect 2354 62 2356 114
rect 2300 51 2356 62
rect 3216 114 3272 125
rect 3216 62 3218 114
rect 3270 62 3272 114
rect 3216 51 3272 62
rect -1090 -100 -1038 -94
rect -1638 -158 -1636 -126
rect -1592 -158 -1590 -126
rect -1090 -158 -1038 -152
rect 3031 -304 3082 -120
rect -1540 -396 -1476 -338
rect 912 -398 968 -387
rect 912 -408 914 -398
rect 860 -450 914 -408
rect 966 -450 968 -398
rect 860 -461 968 -450
rect 1840 -428 1896 -417
rect 860 -621 966 -461
rect 1840 -480 1842 -428
rect 1894 -480 1896 -428
rect 1840 -491 1896 -480
rect 2761 -428 2817 -417
rect 2761 -480 2763 -428
rect 2815 -480 2817 -428
rect 2761 -491 2817 -480
rect -1644 -706 -1590 -624
rect -1550 -639 -1498 -633
rect -1550 -697 -1498 -691
rect -692 -717 -446 -621
rect 723 -717 966 -621
rect 3031 -792 3082 -608
rect 1377 -974 1433 -963
rect 1377 -1026 1379 -974
rect 1431 -1026 1433 -974
rect 1377 -1037 1433 -1026
rect 2299 -972 2355 -961
rect 2299 -1024 2301 -972
rect 2353 -1024 2355 -972
rect 2299 -1035 2355 -1024
rect 3218 -972 3274 -961
rect 3218 -1024 3220 -972
rect 3272 -1024 3274 -972
rect 3218 -1035 3274 -1024
rect -1087 -1183 -1035 -1177
rect -1087 -1241 -1035 -1235
rect 3031 -1392 3082 -1208
rect 917 -1479 973 -1468
rect 917 -1531 919 -1479
rect 971 -1531 973 -1479
rect 917 -1542 973 -1531
rect 1837 -1517 1893 -1506
rect 1837 -1569 1839 -1517
rect 1891 -1569 1893 -1517
rect 1837 -1580 1893 -1569
rect 2759 -1517 2815 -1506
rect 2759 -1569 2761 -1517
rect 2813 -1569 2815 -1517
rect 2759 -1580 2815 -1569
rect 59 -1621 122 -1619
rect 57 -1673 63 -1621
rect 115 -1673 122 -1621
rect 59 -1674 122 -1673
rect 694 -2040 790 -1709
rect 1286 -1837 1962 -1799
rect 3031 -1880 3082 -1696
rect 694 -2136 887 -2040
rect 1378 -2061 1434 -2050
rect 1378 -2113 1380 -2061
rect 1432 -2113 1434 -2061
rect 1378 -2124 1434 -2113
rect 2302 -2061 2358 -2050
rect 2302 -2113 2304 -2061
rect 2356 -2113 2358 -2061
rect 2302 -2124 2358 -2113
rect 3216 -2061 3272 -2050
rect 3216 -2113 3218 -2061
rect 3270 -2113 3272 -2061
rect 3216 -2124 3272 -2113
<< via1 >>
rect 1380 1151 1432 1203
rect 2301 1151 2353 1203
rect 3219 1153 3271 1205
rect -1546 398 -1494 450
rect 908 653 960 705
rect 1815 609 1867 661
rect 2761 608 2813 660
rect 66 325 118 334
rect 66 291 73 325
rect 73 291 107 325
rect 107 291 118 325
rect 66 282 118 291
rect 1380 64 1432 116
rect 2302 62 2354 114
rect 3218 62 3270 114
rect -1090 -152 -1038 -100
rect 914 -450 966 -398
rect 1842 -480 1894 -428
rect 2763 -480 2815 -428
rect -1550 -691 -1498 -639
rect 1379 -1026 1431 -974
rect 2301 -1024 2353 -972
rect 3220 -1024 3272 -972
rect -1087 -1235 -1035 -1183
rect 919 -1531 971 -1479
rect 1839 -1569 1891 -1517
rect 2761 -1569 2813 -1517
rect 63 -1629 115 -1621
rect 63 -1663 72 -1629
rect 72 -1663 106 -1629
rect 106 -1663 115 -1629
rect 63 -1673 115 -1663
rect -1551 -1786 -1496 -1729
rect 1380 -2113 1432 -2061
rect 2304 -2113 2356 -2061
rect 3218 -2113 3270 -2061
<< metal2 >>
rect 1378 1205 1434 1214
rect 1378 1140 1434 1149
rect 2299 1205 2355 1214
rect 2299 1140 2355 1149
rect 3217 1207 3273 1216
rect 3217 1142 3273 1151
rect 906 707 962 716
rect 906 642 962 651
rect 1813 663 1869 672
rect 1813 598 1869 607
rect 998 491 1007 547
rect 1063 491 1072 547
rect -1548 452 -1492 461
rect -1548 387 -1492 396
rect 55 280 64 336
rect 120 280 129 336
rect -1092 -98 -1036 -89
rect -1092 -163 -1036 -154
rect 912 -396 968 -387
rect 912 -461 968 -452
rect -465 -594 -456 -538
rect -400 -594 -391 -538
rect 998 -597 1007 -541
rect 1063 -597 1072 -541
rect -1552 -637 -1496 -628
rect -1552 -702 -1496 -693
rect -692 -632 -544 -621
rect -692 -706 -686 -632
rect -554 -706 -544 -632
rect 1282 -700 1317 373
rect 1378 118 1434 127
rect 1378 53 1434 62
rect 1904 -322 1939 751
rect 2759 662 2815 671
rect 2759 597 2815 606
rect 2300 116 2356 125
rect 2300 51 2356 60
rect 3216 116 3272 125
rect 3216 51 3272 60
rect 1840 -426 1896 -417
rect 1840 -491 1896 -482
rect 2761 -426 2817 -417
rect 2761 -491 2817 -482
rect -692 -717 -544 -706
rect -1089 -1181 -1033 -1172
rect -1089 -1246 -1033 -1237
rect 917 -1477 973 -1468
rect 917 -1542 973 -1533
rect 52 -1675 61 -1619
rect 117 -1675 126 -1619
rect 998 -1685 1007 -1628
rect 1063 -1685 1072 -1628
rect -1554 -1726 -1494 -1717
rect -1554 -1799 -1494 -1790
rect 1284 -1799 1314 -700
rect 1377 -972 1433 -963
rect 1377 -1037 1433 -1028
rect 2299 -970 2355 -961
rect 2299 -1035 2355 -1026
rect 3218 -970 3274 -961
rect 3218 -1035 3274 -1026
rect 1837 -1515 1893 -1506
rect 1837 -1580 1893 -1571
rect 2759 -1515 2815 -1506
rect 2759 -1580 2815 -1571
rect 1378 -2059 1434 -2050
rect 1378 -2124 1434 -2115
rect 2302 -2059 2358 -2050
rect 2302 -2124 2358 -2115
rect 3216 -2059 3272 -2050
rect 3216 -2124 3272 -2115
<< via2 >>
rect 1378 1203 1434 1205
rect 1378 1151 1380 1203
rect 1380 1151 1432 1203
rect 1432 1151 1434 1203
rect 1378 1149 1434 1151
rect 2299 1203 2355 1205
rect 2299 1151 2301 1203
rect 2301 1151 2353 1203
rect 2353 1151 2355 1203
rect 2299 1149 2355 1151
rect 3217 1205 3273 1207
rect 3217 1153 3219 1205
rect 3219 1153 3271 1205
rect 3271 1153 3273 1205
rect 3217 1151 3273 1153
rect 906 705 962 707
rect 906 653 908 705
rect 908 653 960 705
rect 960 653 962 705
rect 906 651 962 653
rect 1813 661 1869 663
rect 1813 609 1815 661
rect 1815 609 1867 661
rect 1867 609 1869 661
rect 1813 607 1869 609
rect 1007 491 1063 547
rect -1548 450 -1492 452
rect -1548 398 -1546 450
rect -1546 398 -1494 450
rect -1494 398 -1492 450
rect -1548 396 -1492 398
rect 64 334 120 336
rect 64 282 66 334
rect 66 282 118 334
rect 118 282 120 334
rect 64 280 120 282
rect -1092 -100 -1036 -98
rect -1092 -152 -1090 -100
rect -1090 -152 -1038 -100
rect -1038 -152 -1036 -100
rect -1092 -154 -1036 -152
rect 912 -398 968 -396
rect 912 -450 914 -398
rect 914 -450 966 -398
rect 966 -450 968 -398
rect 912 -452 968 -450
rect -456 -594 -400 -538
rect 1007 -597 1063 -541
rect -1552 -639 -1496 -637
rect -1552 -691 -1550 -639
rect -1550 -691 -1498 -639
rect -1498 -691 -1496 -639
rect -1552 -693 -1496 -691
rect -686 -706 -554 -632
rect 1378 116 1434 118
rect 1378 64 1380 116
rect 1380 64 1432 116
rect 1432 64 1434 116
rect 1378 62 1434 64
rect 2759 660 2815 662
rect 2759 608 2761 660
rect 2761 608 2813 660
rect 2813 608 2815 660
rect 2759 606 2815 608
rect 2300 114 2356 116
rect 2300 62 2302 114
rect 2302 62 2354 114
rect 2354 62 2356 114
rect 2300 60 2356 62
rect 3216 114 3272 116
rect 3216 62 3218 114
rect 3218 62 3270 114
rect 3270 62 3272 114
rect 3216 60 3272 62
rect 1840 -428 1896 -426
rect 1840 -480 1842 -428
rect 1842 -480 1894 -428
rect 1894 -480 1896 -428
rect 1840 -482 1896 -480
rect 2761 -428 2817 -426
rect 2761 -480 2763 -428
rect 2763 -480 2815 -428
rect 2815 -480 2817 -428
rect 2761 -482 2817 -480
rect -1089 -1183 -1033 -1181
rect -1089 -1235 -1087 -1183
rect -1087 -1235 -1035 -1183
rect -1035 -1235 -1033 -1183
rect -1089 -1237 -1033 -1235
rect 917 -1479 973 -1477
rect 917 -1531 919 -1479
rect 919 -1531 971 -1479
rect 971 -1531 973 -1479
rect 917 -1533 973 -1531
rect 61 -1621 117 -1619
rect 61 -1673 63 -1621
rect 63 -1673 115 -1621
rect 115 -1673 117 -1621
rect 61 -1675 117 -1673
rect 1007 -1685 1063 -1628
rect -1554 -1729 -1494 -1726
rect -1554 -1786 -1551 -1729
rect -1551 -1786 -1496 -1729
rect -1496 -1786 -1494 -1729
rect -1554 -1790 -1494 -1786
rect 1377 -974 1433 -972
rect 1377 -1026 1379 -974
rect 1379 -1026 1431 -974
rect 1431 -1026 1433 -974
rect 1377 -1028 1433 -1026
rect 2299 -972 2355 -970
rect 2299 -1024 2301 -972
rect 2301 -1024 2353 -972
rect 2353 -1024 2355 -972
rect 2299 -1026 2355 -1024
rect 3218 -972 3274 -970
rect 3218 -1024 3220 -972
rect 3220 -1024 3272 -972
rect 3272 -1024 3274 -972
rect 3218 -1026 3274 -1024
rect 1837 -1517 1893 -1515
rect 1837 -1569 1839 -1517
rect 1839 -1569 1891 -1517
rect 1891 -1569 1893 -1517
rect 1837 -1571 1893 -1569
rect 2759 -1517 2815 -1515
rect 2759 -1569 2761 -1517
rect 2761 -1569 2813 -1517
rect 2813 -1569 2815 -1517
rect 2759 -1571 2815 -1569
rect 1378 -2061 1434 -2059
rect 1378 -2113 1380 -2061
rect 1380 -2113 1432 -2061
rect 1432 -2113 1434 -2061
rect 1378 -2115 1434 -2113
rect 2302 -2061 2358 -2059
rect 2302 -2113 2304 -2061
rect 2304 -2113 2356 -2061
rect 2356 -2113 2358 -2061
rect 2302 -2115 2358 -2113
rect 3216 -2061 3272 -2059
rect 3216 -2113 3218 -2061
rect 3218 -2113 3270 -2061
rect 3270 -2113 3272 -2061
rect 3216 -2115 3272 -2113
<< metal3 >>
rect 1358 1209 1456 1227
rect 1358 1145 1374 1209
rect 1438 1145 1456 1209
rect 1358 1129 1456 1145
rect 2279 1209 2377 1227
rect 2279 1145 2295 1209
rect 2359 1145 2377 1209
rect 2279 1129 2377 1145
rect 3197 1211 3295 1229
rect 3197 1147 3213 1211
rect 3277 1147 3295 1211
rect 3197 1131 3295 1147
rect 886 711 984 729
rect 886 647 902 711
rect 966 647 984 711
rect 886 631 984 647
rect 1793 667 1891 685
rect 1793 603 1809 667
rect 1873 603 1891 667
rect 1793 587 1891 603
rect 2739 666 2837 684
rect 2739 602 2755 666
rect 2819 602 2837 666
rect 2739 586 2837 602
rect 999 547 1070 568
rect 999 491 1007 547
rect 1063 491 1070 547
rect -1569 456 -1471 471
rect -1569 392 -1552 456
rect -1488 392 -1471 456
rect -1569 373 -1471 392
rect 55 340 151 341
rect 999 340 1070 491
rect 55 336 1070 340
rect 55 280 64 336
rect 120 280 1070 336
rect 55 275 1070 280
rect 1358 122 1456 140
rect 1358 58 1374 122
rect 1438 58 1456 122
rect 1358 42 1456 58
rect 2280 120 2378 138
rect 2280 56 2296 120
rect 2360 56 2378 120
rect 2280 40 2378 56
rect 3196 120 3294 138
rect 3196 56 3212 120
rect 3276 56 3294 120
rect 3196 40 3294 56
rect -1113 -94 -1015 -79
rect -1113 -158 -1096 -94
rect -1032 -158 -1015 -94
rect -1113 -177 -1015 -158
rect 892 -392 990 -374
rect 892 -456 908 -392
rect 972 -456 990 -392
rect 892 -472 990 -456
rect 1820 -422 1918 -404
rect 1820 -486 1836 -422
rect 1900 -486 1918 -422
rect 1820 -502 1918 -486
rect 2741 -422 2839 -404
rect 2741 -486 2757 -422
rect 2821 -486 2839 -422
rect 2741 -502 2839 -486
rect -471 -535 -391 -533
rect 998 -535 1072 -534
rect -471 -538 1072 -535
rect -471 -594 -456 -538
rect -400 -541 1072 -538
rect -400 -594 1007 -541
rect -471 -597 1007 -594
rect 1063 -597 1072 -541
rect -471 -599 1072 -597
rect 998 -602 1072 -599
rect -1573 -633 -1475 -618
rect -1573 -697 -1556 -633
rect -1492 -697 -1475 -633
rect -1573 -716 -1475 -697
rect -692 -632 -544 -621
rect -692 -706 -686 -632
rect -554 -706 -544 -632
rect -692 -717 -544 -706
rect 1357 -968 1455 -950
rect 1357 -1032 1373 -968
rect 1437 -1032 1455 -968
rect 1357 -1048 1455 -1032
rect 2279 -966 2377 -948
rect 2279 -1030 2295 -966
rect 2359 -1030 2377 -966
rect 2279 -1046 2377 -1030
rect 3198 -966 3296 -948
rect 3198 -1030 3214 -966
rect 3278 -1030 3296 -966
rect 3198 -1046 3296 -1030
rect -1110 -1177 -1012 -1162
rect -1110 -1241 -1093 -1177
rect -1029 -1241 -1012 -1177
rect -1110 -1260 -1012 -1241
rect 897 -1473 995 -1455
rect 897 -1537 913 -1473
rect 977 -1537 995 -1473
rect 897 -1553 995 -1537
rect 1817 -1511 1915 -1493
rect 1817 -1575 1833 -1511
rect 1897 -1575 1915 -1511
rect 1817 -1591 1915 -1575
rect 2739 -1511 2837 -1493
rect 2739 -1575 2755 -1511
rect 2819 -1575 2837 -1511
rect 2739 -1591 2837 -1575
rect 52 -1616 126 -1614
rect 52 -1619 1073 -1616
rect 52 -1675 61 -1619
rect 117 -1628 1073 -1619
rect 117 -1675 1007 -1628
rect 52 -1680 1007 -1675
rect 997 -1685 1007 -1680
rect 1063 -1685 1073 -1628
rect 997 -1694 1073 -1685
rect -1583 -1726 -1458 -1695
rect -1583 -1790 -1556 -1726
rect -1492 -1790 -1458 -1726
rect -1583 -1820 -1458 -1790
rect 1358 -2055 1456 -2037
rect 1358 -2119 1374 -2055
rect 1438 -2119 1456 -2055
rect 1358 -2135 1456 -2119
rect 2282 -2055 2380 -2037
rect 2282 -2119 2298 -2055
rect 2362 -2119 2380 -2055
rect 2282 -2135 2380 -2119
rect 3196 -2055 3294 -2037
rect 3196 -2119 3212 -2055
rect 3276 -2119 3294 -2055
rect 3196 -2135 3294 -2119
<< via3 >>
rect 1374 1205 1438 1209
rect 1374 1149 1378 1205
rect 1378 1149 1434 1205
rect 1434 1149 1438 1205
rect 1374 1145 1438 1149
rect 2295 1205 2359 1209
rect 2295 1149 2299 1205
rect 2299 1149 2355 1205
rect 2355 1149 2359 1205
rect 2295 1145 2359 1149
rect 3213 1207 3277 1211
rect 3213 1151 3217 1207
rect 3217 1151 3273 1207
rect 3273 1151 3277 1207
rect 3213 1147 3277 1151
rect 902 707 966 711
rect 902 651 906 707
rect 906 651 962 707
rect 962 651 966 707
rect 902 647 966 651
rect 1809 663 1873 667
rect 1809 607 1813 663
rect 1813 607 1869 663
rect 1869 607 1873 663
rect 1809 603 1873 607
rect 2755 662 2819 666
rect 2755 606 2759 662
rect 2759 606 2815 662
rect 2815 606 2819 662
rect 2755 602 2819 606
rect -1552 452 -1488 456
rect -1552 396 -1548 452
rect -1548 396 -1492 452
rect -1492 396 -1488 452
rect -1552 392 -1488 396
rect 1374 118 1438 122
rect 1374 62 1378 118
rect 1378 62 1434 118
rect 1434 62 1438 118
rect 1374 58 1438 62
rect 2296 116 2360 120
rect 2296 60 2300 116
rect 2300 60 2356 116
rect 2356 60 2360 116
rect 2296 56 2360 60
rect 3212 116 3276 120
rect 3212 60 3216 116
rect 3216 60 3272 116
rect 3272 60 3276 116
rect 3212 56 3276 60
rect -1096 -98 -1032 -94
rect -1096 -154 -1092 -98
rect -1092 -154 -1036 -98
rect -1036 -154 -1032 -98
rect -1096 -158 -1032 -154
rect 908 -396 972 -392
rect 908 -452 912 -396
rect 912 -452 968 -396
rect 968 -452 972 -396
rect 908 -456 972 -452
rect 1836 -426 1900 -422
rect 1836 -482 1840 -426
rect 1840 -482 1896 -426
rect 1896 -482 1900 -426
rect 1836 -486 1900 -482
rect 2757 -426 2821 -422
rect 2757 -482 2761 -426
rect 2761 -482 2817 -426
rect 2817 -482 2821 -426
rect 2757 -486 2821 -482
rect -1556 -637 -1492 -633
rect -1556 -693 -1552 -637
rect -1552 -693 -1496 -637
rect -1496 -693 -1492 -637
rect -1556 -697 -1492 -693
rect -686 -706 -554 -632
rect 1373 -972 1437 -968
rect 1373 -1028 1377 -972
rect 1377 -1028 1433 -972
rect 1433 -1028 1437 -972
rect 1373 -1032 1437 -1028
rect 2295 -970 2359 -966
rect 2295 -1026 2299 -970
rect 2299 -1026 2355 -970
rect 2355 -1026 2359 -970
rect 2295 -1030 2359 -1026
rect 3214 -970 3278 -966
rect 3214 -1026 3218 -970
rect 3218 -1026 3274 -970
rect 3274 -1026 3278 -970
rect 3214 -1030 3278 -1026
rect -1093 -1181 -1029 -1177
rect -1093 -1237 -1089 -1181
rect -1089 -1237 -1033 -1181
rect -1033 -1237 -1029 -1181
rect -1093 -1241 -1029 -1237
rect 913 -1477 977 -1473
rect 913 -1533 917 -1477
rect 917 -1533 973 -1477
rect 973 -1533 977 -1477
rect 913 -1537 977 -1533
rect 1833 -1515 1897 -1511
rect 1833 -1571 1837 -1515
rect 1837 -1571 1893 -1515
rect 1893 -1571 1897 -1515
rect 1833 -1575 1897 -1571
rect 2755 -1515 2819 -1511
rect 2755 -1571 2759 -1515
rect 2759 -1571 2815 -1515
rect 2815 -1571 2819 -1515
rect 2755 -1575 2819 -1571
rect -1556 -1790 -1554 -1726
rect -1554 -1790 -1494 -1726
rect -1494 -1790 -1492 -1726
rect 1374 -2059 1438 -2055
rect 1374 -2115 1378 -2059
rect 1378 -2115 1434 -2059
rect 1434 -2115 1438 -2059
rect 1374 -2119 1438 -2115
rect 2298 -2059 2362 -2055
rect 2298 -2115 2302 -2059
rect 2302 -2115 2358 -2059
rect 2358 -2115 2362 -2059
rect 2298 -2119 2362 -2115
rect 3212 -2059 3276 -2055
rect 3212 -2115 3216 -2059
rect 3216 -2115 3272 -2059
rect 3272 -2115 3276 -2059
rect 3212 -2119 3276 -2115
<< metal4 >>
rect 898 711 984 1224
rect 898 647 902 711
rect 966 647 984 711
rect -1573 456 -1479 472
rect -1573 392 -1552 456
rect -1488 392 -1479 456
rect -1573 -633 -1479 392
rect -1573 -697 -1556 -633
rect -1492 -697 -1479 -633
rect -1573 -1726 -1479 -697
rect -1116 -94 -1022 -68
rect -1116 -158 -1096 -94
rect -1032 -158 -1022 -94
rect -1116 -621 -1022 -158
rect 898 -392 984 647
rect 898 -456 908 -392
rect 972 -456 984 -392
rect -1116 -632 -544 -621
rect -1116 -706 -686 -632
rect -554 -706 -544 -632
rect -1116 -717 -544 -706
rect -1116 -1177 -1022 -717
rect -1116 -1241 -1093 -1177
rect -1029 -1241 -1022 -1177
rect -1116 -1267 -1022 -1241
rect -1573 -1790 -1556 -1726
rect -1492 -1790 -1479 -1726
rect -1573 -1811 -1479 -1790
rect 898 -1473 984 -456
rect 898 -1537 913 -1473
rect 977 -1537 984 -1473
rect 898 -2136 984 -1537
rect 1357 1209 1443 1224
rect 1357 1145 1374 1209
rect 1438 1145 1443 1209
rect 1357 122 1443 1145
rect 1818 668 1904 1224
rect 1808 667 1904 668
rect 1808 603 1809 667
rect 1873 603 1904 667
rect 1808 602 1904 603
rect 1357 58 1374 122
rect 1438 58 1443 122
rect 1357 -968 1443 58
rect 1357 -1032 1373 -968
rect 1437 -1032 1443 -968
rect 1357 -2055 1443 -1032
rect 1357 -2119 1374 -2055
rect 1438 -2119 1443 -2055
rect 1357 -2136 1443 -2119
rect 1818 -422 1904 602
rect 1818 -486 1836 -422
rect 1900 -486 1904 -422
rect 1818 -1511 1904 -486
rect 1818 -1575 1833 -1511
rect 1897 -1575 1904 -1511
rect 1818 -2136 1904 -1575
rect 2279 1209 2365 1224
rect 2279 1145 2295 1209
rect 2359 1145 2365 1209
rect 2279 120 2365 1145
rect 2279 56 2296 120
rect 2360 56 2365 120
rect 2279 -966 2365 56
rect 2279 -1030 2295 -966
rect 2359 -1030 2365 -966
rect 2279 -2055 2365 -1030
rect 2279 -2119 2298 -2055
rect 2362 -2119 2365 -2055
rect 2279 -2136 2365 -2119
rect 2739 666 2825 1224
rect 2739 602 2755 666
rect 2819 602 2825 666
rect 2739 -422 2825 602
rect 2739 -486 2757 -422
rect 2821 -486 2825 -422
rect 2739 -1511 2825 -486
rect 2739 -1575 2755 -1511
rect 2819 -1575 2825 -1511
rect 2739 -2136 2825 -1575
rect 3195 1211 3281 1224
rect 3195 1147 3213 1211
rect 3277 1147 3281 1211
rect 3195 120 3281 1147
rect 3195 56 3212 120
rect 3276 56 3281 120
rect 3195 -966 3281 56
rect 3195 -1030 3214 -966
rect 3278 -1030 3281 -966
rect 3195 -2055 3281 -1030
rect 3195 -2119 3212 -2055
rect 3276 -2119 3281 -2055
rect 3195 -2136 3281 -2119
use cclkgen  cclkgen_0
timestamp 1662953364
transform 1 0 876 0 1 -2136
box 0 0 2484 1184
use cclkgen  cclkgen_1
timestamp 1662953364
transform 1 0 876 0 1 -2136
box 0 0 2484 1184
use level_up_shifter_d_a  level_up_shifter_d_a_0
timestamp 1662953364
transform 1 0 -2063 0 1 -1215
box 402 498 2794 1683
use level_up_shifter_d_a  level_up_shifter_d_a_1
timestamp 1662953364
transform 1 0 -2063 0 1 -1215
box 402 498 2794 1683
use level_up_shifter_d_a  level_up_shifter_d_a_2
timestamp 1662953364
transform 1 0 -2063 0 -1 -123
box 402 498 2794 1683
use level_up_shifter_d_a  level_up_shifter_d_a_3
timestamp 1662953364
transform 1 0 -2063 0 -1 -123
box 402 498 2794 1683
use phigen  phigen_0
timestamp 1662953364
transform 1 0 876 0 1 40
box 0 0 2484 1184
use phigen  phigen_1
timestamp 1662953364
transform 1 0 876 0 1 40
box 0 0 2484 1184
use phigen  phigen_2
timestamp 1662953364
transform 1 0 876 0 1 -1048
box 0 0 2484 1184
use phigen  phigen_3
timestamp 1662953364
transform 1 0 876 0 1 -1048
box 0 0 2484 1184
<< labels >>
rlabel metal4 2739 750 2739 750 7 GND
rlabel metal4 1438 1118 1438 1118 3 VCCD
flabel metal1 3032 296 3080 480 1 FreeSans 800 0 0 0 phi2b
port 3 n default output
flabel metal1 3032 784 3080 968 1 FreeSans 800 0 0 0 phi2
port 4 n default output
flabel metal1 3031 -792 3082 -608 1 FreeSans 800 0 0 0 phi1b
port 5 n default output
flabel metal1 3031 -304 3082 -120 1 FreeSans 800 0 0 0 phi1
port 6 n default output
flabel metal1 3031 -1880 3082 -1696 1 FreeSans 800 0 0 0 cclkb_ana
port 7 n default output
flabel metal1 3031 -1392 3082 -1208 1 FreeSans 800 0 0 0 cclk_ana
port 8 n default output
flabel metal1 -1494 371 -1078 468 1 FreeSans 800 0 0 0 vccd
port 14 n default bidirectional
flabel poly -1492 -385 -1355 -349 1 FreeSans 800 0 0 0 div2
port 15 n default input
flabel poly -1492 -989 -1355 -953 1 FreeSans 800 0 0 0 cclk
port 16 n default input
flabel metal4 -1116 -717 -686 -621 1 FreeSans 800 0 0 0 vssd
port 17 n default bidirectional
flabel metal1 635 371 731 1224 1 FreeSans 800 0 0 0 vdda
port 18 n
flabel metal2 1282 -700 1317 373 1 FreeSans 800 0 0 0 vnb
port 19 n default bidirectional
flabel metal2 1904 -322 1939 751 1 FreeSans 800 0 0 0 vpb
port 20 n default bidirectional
<< end >>
