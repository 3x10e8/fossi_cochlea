magic
tech sky130B
magscale 1 2
timestamp 1663820320
use analog_core_I  analog_core_I_0 final_designs
timestamp 1663814281
transform 1 0 0 0 1 25779
box 0 -1779 406272 35689
use analog_core_Q  analog_core_Q_0 final_designs
timestamp 1663814281
transform 1 0 0 0 1 -37140
box 0 -328 406272 37140
use digital_unison  digital_unison_0
timestamp 1663814281
transform 1 0 0 0 1 0
box 0 0 406984 24000
<< end >>
