magic
tech sky130A
magscale 1 2
timestamp 1654693435
<< locali >>
rect -341 29074 -307 29090
<< viali >>
rect -521 29090 -487 29124
rect -341 29090 -307 29124
<< metal1 >>
rect -652 33072 22693 33112
rect -652 32952 22693 32992
rect -348 32881 -296 32887
rect -637 32832 -348 32872
rect -296 32832 12524 32872
rect -348 32823 -296 32829
rect -530 32756 -478 32762
rect -637 32712 -530 32752
rect -478 32712 12524 32752
rect -530 32698 -478 32704
rect 2575 32635 2627 32641
rect -637 32592 2575 32632
rect 6151 32632 6203 32638
rect 13884 32637 13936 32643
rect 2627 32592 6151 32632
rect 2575 32577 2627 32583
rect 6203 32592 13884 32632
rect 6151 32574 6203 32580
rect 20033 32640 20085 32646
rect 13936 32592 20033 32632
rect 13884 32579 13936 32585
rect 20085 32592 20877 32632
rect 20033 32582 20085 32588
rect 13806 32523 13858 32529
rect 2488 32515 2540 32521
rect -637 32472 2488 32512
rect 6073 32516 6125 32522
rect 2540 32472 6073 32512
rect 2488 32457 2540 32463
rect 6125 32472 13806 32512
rect 19967 32512 20019 32516
rect 13858 32510 20877 32512
rect 13858 32472 19967 32510
rect 13806 32465 13858 32471
rect 6073 32458 6125 32464
rect 20019 32472 20877 32510
rect 19967 32452 20019 32458
rect 546 32399 598 32405
rect -637 32352 546 32392
rect 4807 32399 4859 32405
rect 598 32352 4807 32392
rect 546 32341 598 32347
rect 12299 32394 12351 32400
rect 4859 32352 12299 32392
rect 4807 32341 4859 32347
rect 18508 32392 18560 32398
rect 12351 32352 18508 32392
rect 12299 32336 12351 32342
rect 18560 32352 20877 32392
rect 18508 32334 18560 32340
rect 632 32283 684 32289
rect -637 32232 632 32272
rect 12385 32282 12437 32288
rect 4891 32276 4943 32282
rect 684 32232 4891 32272
rect 632 32225 684 32231
rect 4943 32232 12385 32272
rect 18595 32281 18647 32287
rect 12437 32232 18595 32272
rect 12385 32224 12437 32230
rect 18647 32232 20877 32272
rect 4891 32218 4943 32224
rect 18595 32223 18647 32229
rect 20932 31897 20993 31954
rect 20716 30585 20758 30925
rect 20634 30560 20953 30585
rect 20634 30290 20647 30560
rect 20937 30290 20953 30560
rect 20634 30273 20953 30290
rect -536 29136 -472 29142
rect -536 29084 -530 29136
rect -478 29084 -472 29136
rect -536 29074 -472 29084
rect -356 29134 -292 29142
rect -356 29082 -350 29134
rect -298 29082 -292 29134
rect -356 29074 -292 29082
rect 669 28265 710 28322
rect -93 28225 710 28265
<< via1 >>
rect -348 32829 -296 32881
rect -530 32704 -478 32756
rect 2575 32583 2627 32635
rect 6151 32580 6203 32632
rect 13884 32585 13936 32637
rect 20033 32588 20085 32640
rect 2488 32463 2540 32515
rect 6073 32464 6125 32516
rect 13806 32471 13858 32523
rect 19967 32458 20019 32510
rect 546 32347 598 32399
rect 4807 32347 4859 32399
rect 12299 32342 12351 32394
rect 18508 32340 18560 32392
rect 632 32231 684 32283
rect 4891 32224 4943 32276
rect 12385 32230 12437 32282
rect 18595 32229 18647 32281
rect 20647 30290 20937 30560
rect -530 29124 -478 29136
rect -530 29090 -521 29124
rect -521 29090 -487 29124
rect -487 29090 -478 29124
rect -530 29084 -478 29090
rect -350 29124 -298 29134
rect -350 29090 -341 29124
rect -341 29090 -307 29124
rect -307 29090 -298 29124
rect -350 29082 -298 29090
<< metal2 >>
rect -348 32881 -296 32887
rect -348 32823 -296 32829
rect -530 32756 -478 32762
rect -530 32698 -478 32704
rect -518 29142 -488 32698
rect -530 29136 -478 29142
rect -339 29140 -309 32823
rect 2575 32635 2627 32641
rect 2575 32577 2627 32583
rect 6151 32632 6203 32638
rect 2488 32515 2540 32521
rect 2488 32457 2540 32463
rect 546 32399 598 32405
rect 546 32341 598 32347
rect -530 29078 -478 29084
rect -350 29134 -298 29140
rect -350 29076 -298 29082
rect 557 28791 587 32341
rect 632 32283 684 32289
rect 632 32225 684 32231
rect 636 28791 666 32225
rect 2508 28790 2538 32457
rect 2587 28790 2617 32577
rect 6151 32574 6203 32580
rect 13884 32637 13936 32643
rect 13884 32579 13936 32585
rect 20033 32640 20085 32646
rect 20033 32582 20085 32588
rect 6073 32516 6125 32522
rect 6073 32458 6125 32464
rect 4807 32399 4859 32405
rect 4807 32341 4859 32347
rect 4817 28790 4847 32341
rect 4891 32276 4943 32282
rect 4891 32218 4943 32224
rect 4896 28790 4926 32218
rect 6078 28790 6108 32458
rect 6157 28790 6187 32574
rect 13806 32523 13858 32529
rect 13806 32465 13858 32471
rect 12299 32394 12351 32400
rect 12299 32336 12351 32342
rect 12307 28791 12337 32336
rect 12385 32282 12437 32288
rect 12385 32224 12437 32230
rect 12386 28791 12416 32224
rect 13816 28790 13846 32465
rect 13895 28790 13925 32579
rect 19967 32510 20019 32516
rect 19967 32452 20019 32458
rect 18508 32392 18560 32398
rect 18508 32334 18560 32340
rect 18517 28791 18547 32334
rect 18595 32281 18647 32287
rect 18595 32223 18647 32229
rect 18596 28790 18626 32223
rect 19968 28790 19998 32452
rect 20047 28790 20077 32582
rect 20634 30560 20953 30585
rect 20634 30290 20647 30560
rect 20937 30290 20953 30560
rect 20634 30273 20953 30290
rect -649 28654 -640 28710
rect -584 28654 -575 28710
rect -261 28387 -252 28443
rect -196 28387 -187 28443
rect 653 28308 662 28364
rect 718 28308 727 28364
rect 2447 28304 2456 28365
rect 2516 28304 2525 28365
rect 4921 28363 4977 28372
rect 4921 28298 4977 28307
rect 6027 28363 6083 28372
rect 6027 28298 6083 28307
rect 12410 28363 12467 28372
rect 12410 28296 12467 28305
rect 13764 28364 13821 28373
rect 13764 28298 13821 28307
rect 18616 28365 18677 28374
rect 18616 28297 18677 28306
rect 19917 28363 19974 28372
rect 19917 28298 19974 28307
<< via2 >>
rect 20647 30290 20937 30560
rect -640 28654 -584 28710
rect -252 28387 -196 28443
rect 662 28308 718 28364
rect 2456 28304 2516 28365
rect 4921 28307 4977 28363
rect 6027 28307 6083 28363
rect 12410 28305 12467 28363
rect 13764 28307 13821 28364
rect 18616 28306 18677 28365
rect 19917 28307 19974 28363
<< metal3 >>
rect -679 31880 25174 31980
rect 20634 30560 20954 30585
rect 20634 30290 20647 30560
rect 20937 30290 20954 30560
rect -661 28714 -563 28733
rect -661 28650 -644 28714
rect -580 28650 -563 28714
rect -661 28635 -563 28650
rect -273 28447 -175 28467
rect -273 28383 -256 28447
rect -192 28383 -175 28447
rect -273 28369 -175 28383
rect 1425 28369 1819 28730
rect 5385 28382 5570 28642
rect 4908 28370 5570 28382
rect 2447 28369 2528 28370
rect 649 28365 2528 28369
rect 649 28364 2456 28365
rect 649 28308 662 28364
rect 718 28308 2456 28364
rect 649 28304 2456 28308
rect 2516 28304 2528 28365
rect 649 28300 2528 28304
rect -900 27972 -580 28197
rect -1160 27929 -580 27972
rect -1160 27695 -1135 27929
rect -901 27695 -580 27929
rect -1160 27652 -580 27695
rect -260 27972 60 28204
rect -260 27929 320 27972
rect -260 27695 61 27929
rect 295 27695 320 27929
rect -260 27652 320 27695
rect -900 27609 60 27652
rect -900 27375 -579 27609
rect -261 27375 60 27609
rect -900 27332 60 27375
rect -1160 27289 -580 27332
rect -1160 27055 -1135 27289
rect -901 27055 -580 27289
rect -1160 27012 -580 27055
rect -260 27289 320 27332
rect -260 27055 61 27289
rect 295 27055 320 27289
rect -260 27012 320 27055
rect -900 26969 60 27012
rect -900 26735 -579 26969
rect -261 26735 60 26969
rect 1425 26937 1819 28300
rect 2447 28299 2528 28300
rect 4908 28363 6092 28370
rect 4908 28307 4921 28363
rect 4977 28307 6027 28363
rect 6083 28307 6092 28363
rect 4908 28297 6092 28307
rect 12398 28363 12483 28373
rect 12398 28305 12410 28363
rect 12467 28305 12483 28363
rect 4908 28273 5570 28297
rect 5385 26929 5570 28273
rect 12398 28095 12483 28305
rect 13091 28100 13365 28644
rect 13744 28364 13833 28378
rect 19174 28376 19276 28646
rect 13744 28307 13764 28364
rect 13821 28307 13833 28364
rect 13744 28100 13833 28307
rect 18602 28375 19276 28376
rect 18602 28365 19991 28375
rect 18602 28306 18616 28365
rect 18677 28363 19991 28365
rect 18677 28307 19917 28363
rect 19974 28307 19991 28363
rect 18677 28306 19991 28307
rect 18602 28297 19991 28306
rect 13091 28095 13834 28100
rect 12398 28034 13834 28095
rect 12398 28026 13365 28034
rect -900 26692 60 26735
rect -1160 26649 -580 26692
rect -1160 26415 -1135 26649
rect -901 26415 -580 26649
rect -1160 26372 -580 26415
rect -260 26649 320 26692
rect -260 26415 61 26649
rect 295 26415 320 26649
rect 12261 26560 12670 26880
rect 13091 26873 13365 28026
rect 18602 26975 18711 28297
rect 20634 26985 20954 30290
rect -260 26372 320 26415
rect -900 26329 60 26372
rect -900 26095 -579 26329
rect -261 26095 60 26329
rect -900 26052 60 26095
rect -1160 26009 -580 26052
rect -1160 25775 -1135 26009
rect -901 25775 -580 26009
rect -1160 25732 -580 25775
rect -260 26009 832 26052
rect -260 25775 61 26009
rect 295 25775 832 26009
rect -260 25732 832 25775
rect -900 25689 60 25732
rect -900 25455 -579 25689
rect -261 25455 60 25689
rect -900 25412 60 25455
rect -1160 25369 -580 25412
rect -1160 25135 -1135 25369
rect -901 25135 -580 25369
rect -1160 25092 -580 25135
rect -260 25369 320 25412
rect -260 25135 61 25369
rect 295 25135 320 25369
rect -260 25092 320 25135
rect 12240 25129 12692 25449
rect -900 25049 60 25092
rect -900 24815 -579 25049
rect -261 24815 60 25049
rect -900 24772 60 24815
rect -1160 24729 -580 24772
rect -1160 24495 -1135 24729
rect -901 24495 -580 24729
rect -1160 24452 -580 24495
rect -260 24729 890 24772
rect -260 24495 61 24729
rect 295 24495 890 24729
rect -260 24452 890 24495
rect -900 24409 60 24452
rect -900 24175 -579 24409
rect -261 24175 60 24409
rect -900 24132 60 24175
rect -1160 24089 -580 24132
rect -1160 23855 -1135 24089
rect -901 23855 -580 24089
rect -1160 23812 -580 23855
rect -260 24089 320 24132
rect -260 23855 61 24089
rect 295 23855 320 24089
rect 12248 24007 12658 24327
rect -260 23812 320 23855
rect -900 23769 60 23812
rect -900 23535 -579 23769
rect -261 23535 60 23769
rect -900 23492 60 23535
rect -1160 23449 -580 23492
rect -1160 23215 -1135 23449
rect -901 23215 -580 23449
rect -1160 23172 -580 23215
rect -260 23449 888 23492
rect -260 23215 61 23449
rect 295 23215 888 23449
rect -260 23172 888 23215
rect -900 23129 60 23172
rect -900 22895 -579 23129
rect -261 22895 60 23129
rect 12258 23112 12667 23432
rect -900 22852 60 22895
rect -1160 22809 -580 22852
rect -1160 22575 -1135 22809
rect -901 22575 -580 22809
rect -1160 22532 -580 22575
rect -260 22809 320 22852
rect -260 22575 61 22809
rect 295 22575 320 22809
rect -260 22532 320 22575
rect -900 22489 60 22532
rect -900 22255 -579 22489
rect -261 22255 60 22489
rect -900 22212 60 22255
rect 12249 22229 12658 22549
rect -1160 22169 -580 22212
rect -1160 21935 -1135 22169
rect -901 21935 -580 22169
rect -1160 21892 -580 21935
rect -260 22169 872 22212
rect -260 21935 61 22169
rect 295 21935 872 22169
rect -260 21892 872 21935
rect -900 21849 60 21892
rect -900 21615 -579 21849
rect -261 21615 60 21849
rect -900 21572 60 21615
rect -1160 21529 -580 21572
rect -1160 21295 -1135 21529
rect -901 21295 -580 21529
rect -1160 21252 -580 21295
rect -260 21529 320 21572
rect -260 21295 61 21529
rect 295 21295 320 21529
rect -260 21252 320 21295
rect -900 21209 60 21252
rect -900 20975 -579 21209
rect -261 20975 60 21209
rect -900 20932 60 20975
rect -1160 20889 -580 20932
rect -1160 20655 -1135 20889
rect -901 20655 -580 20889
rect -1160 20612 -580 20655
rect -260 20889 890 20932
rect -260 20655 61 20889
rect 295 20655 890 20889
rect -260 20612 890 20655
rect -900 20569 60 20612
rect -900 20335 -579 20569
rect -261 20335 60 20569
rect 12268 20525 12677 20845
rect -900 20292 60 20335
rect -1160 20249 -580 20292
rect -1160 20015 -1135 20249
rect -901 20015 -580 20249
rect -1160 19972 -580 20015
rect -260 20249 320 20292
rect -260 20015 61 20249
rect 295 20015 320 20249
rect -260 19972 320 20015
rect -900 19929 60 19972
rect -900 19695 -579 19929
rect -261 19695 60 19929
rect -900 19652 60 19695
rect -1160 19609 -580 19652
rect -1160 19375 -1135 19609
rect -901 19375 -580 19609
rect -1160 19332 -580 19375
rect -260 19609 894 19652
rect 12263 19643 12672 19963
rect -260 19375 61 19609
rect 295 19375 894 19609
rect -260 19332 894 19375
rect -900 19289 60 19332
rect -900 19055 -579 19289
rect -261 19055 60 19289
rect -900 19012 60 19055
rect -1160 18969 -580 19012
rect -1160 18735 -1135 18969
rect -901 18735 -580 18969
rect -1160 18692 -580 18735
rect -260 18969 320 19012
rect -260 18735 61 18969
rect 295 18735 320 18969
rect 12274 18746 12683 19066
rect -260 18692 320 18735
rect -900 18649 60 18692
rect -900 18415 -579 18649
rect -261 18415 60 18649
rect -900 18372 60 18415
rect -1160 18329 -580 18372
rect -1160 18095 -1135 18329
rect -901 18095 -580 18329
rect -1160 18052 -580 18095
rect -260 18329 909 18372
rect -260 18095 61 18329
rect 295 18095 909 18329
rect -260 18052 909 18095
rect -900 18009 60 18052
rect -900 17775 -579 18009
rect -261 17775 60 18009
rect -900 17732 60 17775
rect -1160 17689 -580 17732
rect -1160 17455 -1135 17689
rect -901 17455 -580 17689
rect -1160 17412 -580 17455
rect -260 17689 320 17732
rect -260 17455 61 17689
rect 295 17455 320 17689
rect -260 17412 320 17455
rect -900 17369 60 17412
rect -900 17135 -579 17369
rect -261 17135 60 17369
rect -900 17092 60 17135
rect -1160 17049 -580 17092
rect -1160 16815 -1135 17049
rect -901 16815 -580 17049
rect -1160 16772 -580 16815
rect -260 17049 906 17092
rect 12263 17053 12672 17373
rect -260 16815 61 17049
rect 295 16815 906 17049
rect -260 16772 906 16815
rect -900 16729 60 16772
rect -900 16495 -579 16729
rect -261 16495 60 16729
rect -900 16452 60 16495
rect -1160 16409 -580 16452
rect -1160 16175 -1135 16409
rect -901 16175 -580 16409
rect -1160 16132 -580 16175
rect -260 16409 320 16452
rect -260 16175 61 16409
rect 295 16175 320 16409
rect -260 16132 320 16175
rect 12269 16155 12678 16475
rect -900 16089 60 16132
rect -900 15855 -579 16089
rect -261 15855 60 16089
rect -900 15812 60 15855
rect -1160 15769 -580 15812
rect -1160 15535 -1135 15769
rect -901 15535 -580 15769
rect -1160 15492 -580 15535
rect -260 15769 879 15812
rect -260 15535 61 15769
rect 295 15535 879 15769
rect -260 15492 879 15535
rect -900 15449 60 15492
rect -900 15215 -579 15449
rect -261 15215 60 15449
rect 12272 15262 12681 15582
rect -900 15172 60 15215
rect -1160 15129 -580 15172
rect -1160 14895 -1135 15129
rect -901 14895 -580 15129
rect -1160 14852 -580 14895
rect -260 15129 320 15172
rect -260 14895 61 15129
rect 295 14895 320 15129
rect -260 14852 320 14895
rect -900 14809 60 14852
rect -900 14575 -579 14809
rect -261 14575 60 14809
rect -900 14532 60 14575
rect -1160 14489 -580 14532
rect -1160 14255 -1135 14489
rect -901 14255 -580 14489
rect -1160 14212 -580 14255
rect -260 14489 879 14532
rect -260 14255 61 14489
rect 295 14255 879 14489
rect -260 14212 879 14255
rect -900 14169 60 14212
rect -900 13935 -579 14169
rect -261 13935 60 14169
rect -900 13892 60 13935
rect -1160 13849 -580 13892
rect -1160 13615 -1135 13849
rect -901 13615 -580 13849
rect -1160 13572 -580 13615
rect -260 13849 320 13892
rect -260 13615 61 13849
rect 295 13615 320 13849
rect -260 13572 320 13615
rect -900 13529 60 13572
rect 12277 13566 12686 13886
rect -900 13295 -579 13529
rect -261 13295 60 13529
rect -900 13252 60 13295
rect -1160 13209 -580 13252
rect -1160 12975 -1135 13209
rect -901 12975 -580 13209
rect -1160 12932 -580 12975
rect -260 13209 866 13252
rect -260 12975 61 13209
rect 295 12975 866 13209
rect -260 12932 866 12975
rect -900 12889 60 12932
rect -900 12655 -579 12889
rect -261 12655 60 12889
rect 12272 12673 12681 12993
rect -900 12612 60 12655
rect -1160 12569 -580 12612
rect -1160 12335 -1135 12569
rect -901 12335 -580 12569
rect -1160 12292 -580 12335
rect -260 12569 320 12612
rect -260 12335 61 12569
rect 295 12335 320 12569
rect -260 12292 320 12335
rect -900 12249 60 12292
rect -900 12015 -579 12249
rect -261 12015 60 12249
rect -900 11972 60 12015
rect -1160 11929 -580 11972
rect -1160 11695 -1135 11929
rect -901 11695 -580 11929
rect -1160 11652 -580 11695
rect -260 11929 863 11972
rect -260 11695 61 11929
rect 295 11695 863 11929
rect 12278 11778 12687 12098
rect -260 11652 863 11695
rect -900 11609 60 11652
rect -900 11375 -579 11609
rect -261 11375 60 11609
rect -900 11332 60 11375
rect -1160 11289 -580 11332
rect -1160 11055 -1135 11289
rect -901 11055 -580 11289
rect -1160 11012 -580 11055
rect -260 11289 320 11332
rect -260 11055 61 11289
rect 295 11055 320 11289
rect -260 11012 320 11055
rect -900 10969 60 11012
rect -900 10735 -579 10969
rect -261 10735 60 10969
rect -900 10692 60 10735
rect -1160 10649 -580 10692
rect -1160 10415 -1135 10649
rect -901 10415 -580 10649
rect -1160 10372 -580 10415
rect -260 10649 882 10692
rect -260 10415 61 10649
rect 295 10415 882 10649
rect -260 10372 882 10415
rect -900 10329 60 10372
rect -900 10095 -579 10329
rect -261 10095 60 10329
rect -900 10052 60 10095
rect 12276 10080 12685 10400
rect -1160 10009 -580 10052
rect -1160 9775 -1135 10009
rect -901 9775 -580 10009
rect -1160 9732 -580 9775
rect -260 10009 320 10052
rect -260 9775 61 10009
rect 295 9775 320 10009
rect -260 9732 320 9775
rect -900 9689 60 9732
rect -900 9455 -579 9689
rect -261 9455 60 9689
rect -900 9412 60 9455
rect -1160 9369 -580 9412
rect -1160 9135 -1135 9369
rect -901 9135 -580 9369
rect -1160 9092 -580 9135
rect -260 9369 798 9412
rect -260 9135 61 9369
rect 295 9135 798 9369
rect 12273 9187 12682 9507
rect -260 9092 798 9135
rect -900 9049 60 9092
rect -900 8815 -579 9049
rect -261 8815 60 9049
rect -900 8772 60 8815
rect -1160 8729 -580 8772
rect -1160 8495 -1135 8729
rect -901 8495 -580 8729
rect -1160 8452 -580 8495
rect -260 8729 320 8772
rect -260 8495 61 8729
rect 295 8495 320 8729
rect -260 8452 320 8495
rect -900 8409 60 8452
rect -900 8175 -579 8409
rect -261 8175 60 8409
rect 12269 8295 12671 8615
rect -900 8132 60 8175
rect -1160 8089 -580 8132
rect -1160 7855 -1135 8089
rect -901 7855 -580 8089
rect -1160 7812 -580 7855
rect -260 8089 865 8132
rect -260 7855 61 8089
rect 295 7855 865 8089
rect -260 7812 865 7855
rect -900 7769 60 7812
rect -900 7535 -579 7769
rect -261 7535 60 7769
rect -900 7492 60 7535
rect -1160 7449 -580 7492
rect -1160 7215 -1135 7449
rect -901 7215 -580 7449
rect -1160 7172 -580 7215
rect -260 7449 320 7492
rect -260 7215 61 7449
rect 295 7215 320 7449
rect -260 7172 320 7215
rect -900 7129 60 7172
rect -900 6895 -579 7129
rect -261 6895 60 7129
rect -900 6852 60 6895
rect -1160 6809 -580 6852
rect -1160 6575 -1135 6809
rect -901 6575 -580 6809
rect -1160 6532 -580 6575
rect -260 6809 901 6852
rect -260 6575 61 6809
rect 295 6575 901 6809
rect 12271 6599 12673 6919
rect -260 6532 901 6575
rect -900 6489 60 6532
rect -900 6255 -579 6489
rect -261 6255 60 6489
rect -900 6212 60 6255
rect -1160 6169 -580 6212
rect -1160 5935 -1135 6169
rect -901 5935 -580 6169
rect -1160 5892 -580 5935
rect -260 6169 320 6212
rect -260 5935 61 6169
rect 295 5935 320 6169
rect -260 5892 320 5935
rect -900 5849 60 5892
rect -900 5615 -579 5849
rect -261 5615 60 5849
rect 12275 5705 12677 6025
rect -900 5572 60 5615
rect -1160 5529 -580 5572
rect -1160 5295 -1135 5529
rect -901 5295 -580 5529
rect -1160 5252 -580 5295
rect -900 4692 -580 5252
rect -260 5529 838 5572
rect -260 5295 61 5529
rect 295 5295 838 5529
rect -260 5252 838 5295
rect -260 4692 60 5252
rect 12267 4811 12669 5131
rect -845 4621 -636 4627
rect -845 4432 -839 4621
rect -642 4432 -636 4621
rect -845 3035 -636 4432
rect -204 4621 5 4627
rect -204 4432 -198 4621
rect -1 4432 5 4621
rect -204 3676 5 4432
rect 642 3977 962 4002
rect 642 3743 685 3977
rect 919 3743 962 3977
rect 642 3742 962 3743
rect 1282 3977 1602 4591
rect 1282 3743 1325 3977
rect 1559 3743 1602 3977
rect 1282 3742 1602 3743
rect 1922 3977 2242 4002
rect 1922 3743 1965 3977
rect 2199 3743 2242 3977
rect 1922 3742 2242 3743
rect 2562 3977 2882 4589
rect 2562 3743 2605 3977
rect 2839 3743 2882 3977
rect 2562 3742 2882 3743
rect 3202 3977 3522 4002
rect 3202 3743 3245 3977
rect 3479 3743 3522 3977
rect 3202 3742 3522 3743
rect 3842 3977 4162 4592
rect 3842 3743 3885 3977
rect 4119 3743 4162 3977
rect 3842 3742 4162 3743
rect 4482 3977 4802 4002
rect 4482 3743 4525 3977
rect 4759 3743 4802 3977
rect 4482 3742 4802 3743
rect 5122 3977 5442 4590
rect 5122 3743 5165 3977
rect 5399 3743 5442 3977
rect 5122 3742 5442 3743
rect 5762 3977 6082 4002
rect 5762 3743 5805 3977
rect 6039 3743 6082 3977
rect 5762 3742 6082 3743
rect 6402 3977 6722 4591
rect 6402 3743 6445 3977
rect 6679 3743 6722 3977
rect 6402 3742 6722 3743
rect 7042 3977 7362 4002
rect 7042 3743 7085 3977
rect 7319 3743 7362 3977
rect 7042 3742 7362 3743
rect 7682 3977 8002 4590
rect 7682 3743 7725 3977
rect 7959 3743 8002 3977
rect 7682 3742 8002 3743
rect 8322 3977 8642 4002
rect 8322 3743 8365 3977
rect 8599 3743 8642 3977
rect 8322 3742 8642 3743
rect 8962 3977 9282 4591
rect 8962 3743 9005 3977
rect 9239 3743 9282 3977
rect 8962 3742 9282 3743
rect 9602 3977 9922 4002
rect 9602 3743 9645 3977
rect 9879 3743 9922 3977
rect 9602 3742 9922 3743
rect 10242 3977 10562 4592
rect 10242 3743 10285 3977
rect 10519 3743 10562 3977
rect 10242 3742 10562 3743
rect 10882 3977 11202 4002
rect 10882 3743 10925 3977
rect 11159 3743 11202 3977
rect 10882 3742 11202 3743
rect 11522 3977 11842 4592
rect 11522 3743 11565 3977
rect 11799 3743 11842 3977
rect 11522 3742 11842 3743
rect 12162 3977 12482 4002
rect 12162 3743 12205 3977
rect 12439 3743 12482 3977
rect 12162 3742 12482 3743
rect 12802 3977 13122 4591
rect 12802 3743 12845 3977
rect 13079 3743 13122 3977
rect 12802 3742 13122 3743
rect 13442 3977 13762 4002
rect 13442 3743 13485 3977
rect 13719 3743 13762 3977
rect 13442 3742 13762 3743
rect 14082 3977 14402 4002
rect 14082 3743 14125 3977
rect 14359 3743 14402 3977
rect 14082 3742 14402 3743
rect 14722 3977 15042 4002
rect 14722 3743 14765 3977
rect 14999 3743 15042 3977
rect 14722 3742 15042 3743
rect 15362 3977 15682 4590
rect 15362 3743 15405 3977
rect 15639 3743 15682 3977
rect 15362 3742 15682 3743
rect 16002 3977 16322 4002
rect 16002 3743 16045 3977
rect 16279 3743 16322 3977
rect 16002 3742 16322 3743
rect 16642 3977 16962 4592
rect 16642 3743 16685 3977
rect 16919 3743 16962 3977
rect 16642 3742 16962 3743
rect 17282 3977 17602 4002
rect 17282 3743 17325 3977
rect 17559 3743 17602 3977
rect 17282 3742 17602 3743
rect 17922 3977 18242 4589
rect 17922 3743 17965 3977
rect 18199 3743 18242 3977
rect 17922 3742 18242 3743
rect 18562 3977 18882 4002
rect 18562 3743 18605 3977
rect 18839 3743 18882 3977
rect 18562 3742 18882 3743
rect 19202 3977 19522 4002
rect 19202 3743 19245 3977
rect 19479 3743 19522 3977
rect 19202 3742 19522 3743
rect 19842 3977 20162 4002
rect 19842 3743 19885 3977
rect 20119 3743 20162 3977
rect 19842 3742 20162 3743
rect 20482 3977 20802 4002
rect 20482 3743 20525 3977
rect 20759 3743 20802 3977
rect 20482 3742 20802 3743
rect 21122 3977 21442 4002
rect 21122 3743 21165 3977
rect 21399 3743 21442 3977
rect 21122 3742 21442 3743
rect 21762 3977 22082 4002
rect 21762 3743 21805 3977
rect 22039 3743 22082 3977
rect 21762 3742 22082 3743
rect -204 3487 -198 3676
rect -1 3487 5 3676
rect -204 3483 5 3487
rect 70 3422 22766 3742
rect 322 3421 642 3422
rect 322 3103 365 3421
rect 599 3103 642 3421
rect 322 3102 642 3103
rect 962 3421 1282 3422
rect 962 3103 1005 3421
rect 1239 3103 1282 3421
rect 962 3102 1282 3103
rect 1602 3421 1922 3422
rect 1602 3103 1645 3421
rect 1879 3103 1922 3421
rect 1602 3102 1922 3103
rect 2242 3421 2562 3422
rect 2242 3103 2285 3421
rect 2519 3103 2562 3421
rect 2242 3102 2562 3103
rect 2882 3421 3202 3422
rect 2882 3103 2925 3421
rect 3159 3103 3202 3421
rect 2882 3102 3202 3103
rect 3522 3421 3842 3422
rect 3522 3103 3565 3421
rect 3799 3103 3842 3421
rect 3522 3102 3842 3103
rect 4162 3421 4482 3422
rect 4162 3103 4205 3421
rect 4439 3103 4482 3421
rect 4162 3102 4482 3103
rect 4802 3421 5122 3422
rect 4802 3103 4845 3421
rect 5079 3103 5122 3421
rect 4802 3102 5122 3103
rect 5442 3421 5762 3422
rect 5442 3103 5485 3421
rect 5719 3103 5762 3421
rect 5442 3102 5762 3103
rect 6082 3421 6402 3422
rect 6082 3103 6125 3421
rect 6359 3103 6402 3421
rect 6082 3102 6402 3103
rect 6722 3421 7042 3422
rect 6722 3103 6765 3421
rect 6999 3103 7042 3421
rect 6722 3102 7042 3103
rect 7362 3421 7682 3422
rect 7362 3103 7405 3421
rect 7639 3103 7682 3421
rect 7362 3102 7682 3103
rect 8002 3421 8322 3422
rect 8002 3103 8045 3421
rect 8279 3103 8322 3421
rect 8002 3102 8322 3103
rect 8642 3421 8962 3422
rect 8642 3103 8685 3421
rect 8919 3103 8962 3421
rect 8642 3102 8962 3103
rect 9282 3421 9602 3422
rect 9282 3103 9325 3421
rect 9559 3103 9602 3421
rect 9282 3102 9602 3103
rect 9922 3421 10242 3422
rect 9922 3103 9965 3421
rect 10199 3103 10242 3421
rect 9922 3102 10242 3103
rect 10562 3421 10882 3422
rect 10562 3103 10605 3421
rect 10839 3103 10882 3421
rect 10562 3102 10882 3103
rect 11202 3421 11522 3422
rect 11202 3103 11245 3421
rect 11479 3103 11522 3421
rect 11202 3102 11522 3103
rect 11842 3421 12162 3422
rect 11842 3103 11885 3421
rect 12119 3103 12162 3421
rect 11842 3102 12162 3103
rect 12482 3421 12802 3422
rect 12482 3103 12525 3421
rect 12759 3103 12802 3421
rect 12482 3102 12802 3103
rect 13122 3421 13442 3422
rect 13122 3103 13165 3421
rect 13399 3103 13442 3421
rect 13122 3102 13442 3103
rect 13762 3421 14082 3422
rect 13762 3103 13805 3421
rect 14039 3103 14082 3421
rect 13762 3102 14082 3103
rect 14402 3421 14722 3422
rect 14402 3103 14445 3421
rect 14679 3103 14722 3421
rect 14402 3102 14722 3103
rect 15042 3421 15362 3422
rect 15042 3103 15085 3421
rect 15319 3103 15362 3421
rect 15042 3102 15362 3103
rect 15682 3421 16002 3422
rect 15682 3103 15725 3421
rect 15959 3103 16002 3421
rect 15682 3102 16002 3103
rect 16322 3421 16642 3422
rect 16322 3103 16365 3421
rect 16599 3103 16642 3421
rect 16322 3102 16642 3103
rect 16962 3421 17282 3422
rect 16962 3103 17005 3421
rect 17239 3103 17282 3421
rect 16962 3102 17282 3103
rect 17602 3421 17922 3422
rect 17602 3103 17645 3421
rect 17879 3103 17922 3421
rect 17602 3102 17922 3103
rect 18242 3421 18562 3422
rect 18242 3103 18285 3421
rect 18519 3103 18562 3421
rect 18242 3102 18562 3103
rect 18882 3421 19202 3422
rect 18882 3103 18925 3421
rect 19159 3103 19202 3421
rect 18882 3102 19202 3103
rect 19522 3421 19842 3422
rect 19522 3103 19565 3421
rect 19799 3103 19842 3421
rect 19522 3102 19842 3103
rect 20162 3421 20482 3422
rect 20162 3103 20205 3421
rect 20439 3103 20482 3421
rect 20162 3102 20482 3103
rect 20802 3421 21122 3422
rect 20802 3103 20845 3421
rect 21079 3103 21122 3421
rect 20802 3102 21122 3103
rect 21442 3421 21762 3422
rect 21442 3103 21485 3421
rect 21719 3103 21762 3421
rect 21442 3102 21762 3103
rect 22082 3421 22402 3422
rect 22082 3103 22125 3421
rect 22359 3103 22402 3421
rect 22082 3102 22402 3103
rect -845 2846 -839 3035
rect -642 2846 -636 3035
rect -845 2842 -636 2846
rect -571 2782 22766 3102
rect 642 2781 962 2782
rect 642 2547 685 2781
rect 919 2547 962 2781
rect 642 2522 962 2547
rect 1282 2781 1602 2782
rect 1282 2547 1325 2781
rect 1559 2547 1602 2781
rect 1282 2522 1602 2547
rect 1922 2781 2242 2782
rect 1922 2547 1965 2781
rect 2199 2547 2242 2781
rect 1922 2522 2242 2547
rect 2562 2781 2882 2782
rect 2562 2547 2605 2781
rect 2839 2547 2882 2781
rect 2562 2522 2882 2547
rect 3202 2781 3522 2782
rect 3202 2547 3245 2781
rect 3479 2547 3522 2781
rect 3202 2522 3522 2547
rect 3842 2781 4162 2782
rect 3842 2547 3885 2781
rect 4119 2547 4162 2781
rect 3842 2522 4162 2547
rect 4482 2781 4802 2782
rect 4482 2547 4525 2781
rect 4759 2547 4802 2781
rect 4482 2522 4802 2547
rect 5122 2781 5442 2782
rect 5122 2547 5165 2781
rect 5399 2547 5442 2781
rect 5122 2522 5442 2547
rect 5762 2781 6082 2782
rect 5762 2547 5805 2781
rect 6039 2547 6082 2781
rect 5762 2522 6082 2547
rect 6402 2781 6722 2782
rect 6402 2547 6445 2781
rect 6679 2547 6722 2781
rect 6402 2522 6722 2547
rect 7042 2781 7362 2782
rect 7042 2547 7085 2781
rect 7319 2547 7362 2781
rect 7042 2522 7362 2547
rect 7682 2781 8002 2782
rect 7682 2547 7725 2781
rect 7959 2547 8002 2781
rect 7682 2522 8002 2547
rect 8322 2781 8642 2782
rect 8322 2547 8365 2781
rect 8599 2547 8642 2781
rect 8322 2522 8642 2547
rect 8962 2781 9282 2782
rect 8962 2547 9005 2781
rect 9239 2547 9282 2781
rect 8962 2522 9282 2547
rect 9602 2781 9922 2782
rect 9602 2547 9645 2781
rect 9879 2547 9922 2781
rect 9602 2522 9922 2547
rect 10242 2781 10562 2782
rect 10242 2547 10285 2781
rect 10519 2547 10562 2781
rect 10242 2522 10562 2547
rect 10882 2781 11202 2782
rect 10882 2547 10925 2781
rect 11159 2547 11202 2781
rect 10882 2522 11202 2547
rect 11522 2781 11842 2782
rect 11522 2547 11565 2781
rect 11799 2547 11842 2781
rect 11522 2522 11842 2547
rect 12162 2781 12482 2782
rect 12162 2547 12205 2781
rect 12439 2547 12482 2781
rect 12162 2522 12482 2547
rect 12802 2781 13122 2782
rect 12802 2547 12845 2781
rect 13079 2547 13122 2781
rect 12802 2522 13122 2547
rect 13442 2781 13762 2782
rect 13442 2547 13485 2781
rect 13719 2547 13762 2781
rect 13442 2522 13762 2547
rect 14082 2781 14402 2782
rect 14082 2547 14125 2781
rect 14359 2547 14402 2781
rect 14082 2522 14402 2547
rect 14722 2781 15042 2782
rect 14722 2547 14765 2781
rect 14999 2547 15042 2781
rect 14722 2522 15042 2547
rect 15362 2781 15682 2782
rect 15362 2547 15405 2781
rect 15639 2547 15682 2781
rect 15362 2522 15682 2547
rect 16002 2781 16322 2782
rect 16002 2547 16045 2781
rect 16279 2547 16322 2781
rect 16002 2522 16322 2547
rect 16642 2781 16962 2782
rect 16642 2547 16685 2781
rect 16919 2547 16962 2781
rect 16642 2522 16962 2547
rect 17282 2781 17602 2782
rect 17282 2547 17325 2781
rect 17559 2547 17602 2781
rect 17282 2522 17602 2547
rect 17922 2781 18242 2782
rect 17922 2547 17965 2781
rect 18199 2547 18242 2781
rect 17922 2522 18242 2547
rect 18562 2781 18882 2782
rect 18562 2547 18605 2781
rect 18839 2547 18882 2781
rect 18562 2522 18882 2547
rect 19202 2781 19522 2782
rect 19202 2547 19245 2781
rect 19479 2547 19522 2781
rect 19202 2522 19522 2547
rect 19842 2781 20162 2782
rect 19842 2547 19885 2781
rect 20119 2547 20162 2781
rect 19842 2522 20162 2547
rect 20482 2781 20802 2782
rect 20482 2547 20525 2781
rect 20759 2547 20802 2781
rect 20482 2522 20802 2547
rect 21122 2781 21442 2782
rect 21122 2547 21165 2781
rect 21399 2547 21442 2781
rect 21122 2522 21442 2547
rect 21762 2781 22082 2782
rect 21762 2547 21805 2781
rect 22039 2547 22082 2781
rect 21762 2522 22082 2547
<< via3 >>
rect 20647 30290 20937 30560
rect -644 28710 -580 28714
rect -644 28654 -640 28710
rect -640 28654 -584 28710
rect -584 28654 -580 28710
rect -644 28650 -580 28654
rect -256 28443 -192 28447
rect -256 28387 -252 28443
rect -252 28387 -196 28443
rect -196 28387 -192 28443
rect -256 28383 -192 28387
rect -1135 27695 -901 27929
rect 61 27695 295 27929
rect -579 27375 -261 27609
rect -1135 27055 -901 27289
rect 61 27055 295 27289
rect -579 26735 -261 26969
rect -1135 26415 -901 26649
rect 61 26415 295 26649
rect -579 26095 -261 26329
rect -1135 25775 -901 26009
rect 61 25775 295 26009
rect -579 25455 -261 25689
rect -1135 25135 -901 25369
rect 61 25135 295 25369
rect -579 24815 -261 25049
rect -1135 24495 -901 24729
rect 61 24495 295 24729
rect -579 24175 -261 24409
rect -1135 23855 -901 24089
rect 61 23855 295 24089
rect -579 23535 -261 23769
rect -1135 23215 -901 23449
rect 61 23215 295 23449
rect -579 22895 -261 23129
rect -1135 22575 -901 22809
rect 61 22575 295 22809
rect -579 22255 -261 22489
rect -1135 21935 -901 22169
rect 61 21935 295 22169
rect -579 21615 -261 21849
rect -1135 21295 -901 21529
rect 61 21295 295 21529
rect -579 20975 -261 21209
rect -1135 20655 -901 20889
rect 61 20655 295 20889
rect -579 20335 -261 20569
rect -1135 20015 -901 20249
rect 61 20015 295 20249
rect -579 19695 -261 19929
rect -1135 19375 -901 19609
rect 61 19375 295 19609
rect -579 19055 -261 19289
rect -1135 18735 -901 18969
rect 61 18735 295 18969
rect -579 18415 -261 18649
rect -1135 18095 -901 18329
rect 61 18095 295 18329
rect -579 17775 -261 18009
rect -1135 17455 -901 17689
rect 61 17455 295 17689
rect -579 17135 -261 17369
rect -1135 16815 -901 17049
rect 61 16815 295 17049
rect -579 16495 -261 16729
rect -1135 16175 -901 16409
rect 61 16175 295 16409
rect -579 15855 -261 16089
rect -1135 15535 -901 15769
rect 61 15535 295 15769
rect -579 15215 -261 15449
rect -1135 14895 -901 15129
rect 61 14895 295 15129
rect -579 14575 -261 14809
rect -1135 14255 -901 14489
rect 61 14255 295 14489
rect -579 13935 -261 14169
rect -1135 13615 -901 13849
rect 61 13615 295 13849
rect -579 13295 -261 13529
rect -1135 12975 -901 13209
rect 61 12975 295 13209
rect -579 12655 -261 12889
rect -1135 12335 -901 12569
rect 61 12335 295 12569
rect -579 12015 -261 12249
rect -1135 11695 -901 11929
rect 61 11695 295 11929
rect -579 11375 -261 11609
rect -1135 11055 -901 11289
rect 61 11055 295 11289
rect -579 10735 -261 10969
rect -1135 10415 -901 10649
rect 61 10415 295 10649
rect -579 10095 -261 10329
rect -1135 9775 -901 10009
rect 61 9775 295 10009
rect -579 9455 -261 9689
rect -1135 9135 -901 9369
rect 61 9135 295 9369
rect -579 8815 -261 9049
rect -1135 8495 -901 8729
rect 61 8495 295 8729
rect -579 8175 -261 8409
rect -1135 7855 -901 8089
rect 61 7855 295 8089
rect -579 7535 -261 7769
rect -1135 7215 -901 7449
rect 61 7215 295 7449
rect -579 6895 -261 7129
rect -1135 6575 -901 6809
rect 61 6575 295 6809
rect -579 6255 -261 6489
rect -1135 5935 -901 6169
rect 61 5935 295 6169
rect -579 5615 -261 5849
rect -1135 5295 -901 5529
rect 61 5295 295 5529
rect -839 4432 -642 4621
rect -198 4432 -1 4621
rect 685 3743 919 3977
rect 1325 3743 1559 3977
rect 1965 3743 2199 3977
rect 2605 3743 2839 3977
rect 3245 3743 3479 3977
rect 3885 3743 4119 3977
rect 4525 3743 4759 3977
rect 5165 3743 5399 3977
rect 5805 3743 6039 3977
rect 6445 3743 6679 3977
rect 7085 3743 7319 3977
rect 7725 3743 7959 3977
rect 8365 3743 8599 3977
rect 9005 3743 9239 3977
rect 9645 3743 9879 3977
rect 10285 3743 10519 3977
rect 10925 3743 11159 3977
rect 11565 3743 11799 3977
rect 12205 3743 12439 3977
rect 12845 3743 13079 3977
rect 13485 3743 13719 3977
rect 14125 3743 14359 3977
rect 14765 3743 14999 3977
rect 15405 3743 15639 3977
rect 16045 3743 16279 3977
rect 16685 3743 16919 3977
rect 17325 3743 17559 3977
rect 17965 3743 18199 3977
rect 18605 3743 18839 3977
rect 19245 3743 19479 3977
rect 19885 3743 20119 3977
rect 20525 3743 20759 3977
rect 21165 3743 21399 3977
rect 21805 3743 22039 3977
rect -198 3487 -1 3676
rect 365 3103 599 3421
rect 1005 3103 1239 3421
rect 1645 3103 1879 3421
rect 2285 3103 2519 3421
rect 2925 3103 3159 3421
rect 3565 3103 3799 3421
rect 4205 3103 4439 3421
rect 4845 3103 5079 3421
rect 5485 3103 5719 3421
rect 6125 3103 6359 3421
rect 6765 3103 6999 3421
rect 7405 3103 7639 3421
rect 8045 3103 8279 3421
rect 8685 3103 8919 3421
rect 9325 3103 9559 3421
rect 9965 3103 10199 3421
rect 10605 3103 10839 3421
rect 11245 3103 11479 3421
rect 11885 3103 12119 3421
rect 12525 3103 12759 3421
rect 13165 3103 13399 3421
rect 13805 3103 14039 3421
rect 14445 3103 14679 3421
rect 15085 3103 15319 3421
rect 15725 3103 15959 3421
rect 16365 3103 16599 3421
rect 17005 3103 17239 3421
rect 17645 3103 17879 3421
rect 18285 3103 18519 3421
rect 18925 3103 19159 3421
rect 19565 3103 19799 3421
rect 20205 3103 20439 3421
rect 20845 3103 21079 3421
rect 21485 3103 21719 3421
rect 22125 3103 22359 3421
rect -839 2846 -642 3035
rect 685 2547 919 2781
rect 1325 2547 1559 2781
rect 1965 2547 2199 2781
rect 2605 2547 2839 2781
rect 3245 2547 3479 2781
rect 3885 2547 4119 2781
rect 4525 2547 4759 2781
rect 5165 2547 5399 2781
rect 5805 2547 6039 2781
rect 6445 2547 6679 2781
rect 7085 2547 7319 2781
rect 7725 2547 7959 2781
rect 8365 2547 8599 2781
rect 9005 2547 9239 2781
rect 9645 2547 9879 2781
rect 10285 2547 10519 2781
rect 10925 2547 11159 2781
rect 11565 2547 11799 2781
rect 12205 2547 12439 2781
rect 12845 2547 13079 2781
rect 13485 2547 13719 2781
rect 14125 2547 14359 2781
rect 14765 2547 14999 2781
rect 15405 2547 15639 2781
rect 16045 2547 16279 2781
rect 16685 2547 16919 2781
rect 17325 2547 17559 2781
rect 17965 2547 18199 2781
rect 18605 2547 18839 2781
rect 19245 2547 19479 2781
rect 19885 2547 20119 2781
rect 20525 2547 20759 2781
rect 21165 2547 21399 2781
rect 21805 2547 22039 2781
<< metal4 >>
rect 20634 30560 20953 30585
rect 20634 30290 20647 30560
rect 20937 30290 20953 30560
rect 20634 30273 20953 30290
rect -840 28714 -577 28721
rect -840 28650 -644 28714
rect -580 28650 -577 28714
rect -840 28648 -577 28650
rect -840 4621 -641 28648
rect 787 28498 1165 28789
rect 2122 28587 2269 28740
rect 5134 28587 5245 28680
rect 2122 28515 2395 28587
rect 2788 28519 2947 28587
rect 2659 28518 2947 28519
rect -273 28447 0 28462
rect -273 28383 -256 28447
rect -192 28383 0 28447
rect 2658 28436 2947 28518
rect 5050 28515 5245 28587
rect 5798 28587 5906 28678
rect 12691 28587 12825 28710
rect 13535 28637 13657 28731
rect 5798 28515 5961 28587
rect 6347 28540 6576 28587
rect 5798 28513 5906 28515
rect 6259 28436 6576 28540
rect -273 28369 0 28383
rect -840 4432 -839 4621
rect -642 4432 -641 4621
rect -840 4431 -641 4432
rect -199 4621 0 28369
rect 2839 26338 2947 28436
rect 6456 26234 6576 28436
rect 10976 28515 12155 28587
rect 12539 28515 12825 28587
rect 13595 28587 13657 28637
rect 18909 28587 19055 28680
rect 13595 28515 13716 28587
rect 14087 28515 14820 28587
rect 10976 26339 11163 28515
rect 12691 28514 12825 28515
rect 12261 26560 12670 26880
rect 14686 26343 14820 28515
rect 17493 28515 18364 28587
rect 18747 28515 19055 28587
rect 17493 26336 17670 28515
rect 18909 28510 19055 28515
rect 19534 28587 19645 28663
rect 19534 28515 19885 28587
rect 20252 28521 20378 28587
rect 19534 28512 19645 28515
rect 20117 28436 20378 28521
rect 20253 26313 20378 28436
rect 12240 25129 12692 25449
rect 12248 24007 12658 24327
rect 12258 23112 12667 23432
rect 12249 22229 12658 22549
rect 12268 20525 12677 20845
rect 12263 19643 12672 19963
rect 12274 18746 12683 19066
rect 12263 17053 12672 17373
rect 12269 16155 12678 16475
rect 12272 15262 12681 15582
rect 12277 13566 12686 13886
rect 12272 12673 12681 12993
rect 12278 11778 12687 12098
rect 12276 10080 12685 10400
rect 12273 9187 12682 9507
rect 12269 8295 12671 8615
rect 12271 6599 12673 6919
rect 12275 5705 12677 6025
rect 12267 4811 12669 5131
rect -199 4432 -198 4621
rect -1 4432 0 4621
rect -199 4431 0 4432
rect -900 3676 22766 3682
rect -900 3487 -198 3676
rect -1 3487 22766 3676
rect -900 3483 22766 3487
rect -900 3035 22766 3041
rect -900 2846 -839 3035
rect -642 2846 22766 3035
rect -900 2842 22766 2846
<< via4 >>
rect 20659 30300 20895 30537
rect -1136 27929 -900 27930
rect -1136 27695 -1135 27929
rect -1135 27695 -901 27929
rect -901 27695 -900 27929
rect -1136 27694 -900 27695
rect -1136 27289 -900 27290
rect -1136 27055 -1135 27289
rect -1135 27055 -901 27289
rect -901 27055 -900 27289
rect -1136 27054 -900 27055
rect -1136 26649 -900 26650
rect -1136 26415 -1135 26649
rect -1135 26415 -901 26649
rect -901 26415 -900 26649
rect -1136 26414 -900 26415
rect -1136 26009 -900 26010
rect -1136 25775 -1135 26009
rect -1135 25775 -901 26009
rect -901 25775 -900 26009
rect -1136 25774 -900 25775
rect -1136 25369 -900 25370
rect -1136 25135 -1135 25369
rect -1135 25135 -901 25369
rect -901 25135 -900 25369
rect -1136 25134 -900 25135
rect -1136 24729 -900 24730
rect -1136 24495 -1135 24729
rect -1135 24495 -901 24729
rect -901 24495 -900 24729
rect -1136 24494 -900 24495
rect -1136 24089 -900 24090
rect -1136 23855 -1135 24089
rect -1135 23855 -901 24089
rect -901 23855 -900 24089
rect -1136 23854 -900 23855
rect -1136 23449 -900 23450
rect -1136 23215 -1135 23449
rect -1135 23215 -901 23449
rect -901 23215 -900 23449
rect -1136 23214 -900 23215
rect -1136 22809 -900 22810
rect -1136 22575 -1135 22809
rect -1135 22575 -901 22809
rect -901 22575 -900 22809
rect -1136 22574 -900 22575
rect -1136 22169 -900 22170
rect -1136 21935 -1135 22169
rect -1135 21935 -901 22169
rect -901 21935 -900 22169
rect -1136 21934 -900 21935
rect -1136 21529 -900 21530
rect -1136 21295 -1135 21529
rect -1135 21295 -901 21529
rect -901 21295 -900 21529
rect -1136 21294 -900 21295
rect -1136 20889 -900 20890
rect -1136 20655 -1135 20889
rect -1135 20655 -901 20889
rect -901 20655 -900 20889
rect -1136 20654 -900 20655
rect -1136 20249 -900 20250
rect -1136 20015 -1135 20249
rect -1135 20015 -901 20249
rect -901 20015 -900 20249
rect -1136 20014 -900 20015
rect -1136 19609 -900 19610
rect -1136 19375 -1135 19609
rect -1135 19375 -901 19609
rect -901 19375 -900 19609
rect -1136 19374 -900 19375
rect -1136 18969 -900 18970
rect -1136 18735 -1135 18969
rect -1135 18735 -901 18969
rect -901 18735 -900 18969
rect -1136 18734 -900 18735
rect -1136 18329 -900 18330
rect -1136 18095 -1135 18329
rect -1135 18095 -901 18329
rect -901 18095 -900 18329
rect -1136 18094 -900 18095
rect -1136 17689 -900 17690
rect -1136 17455 -1135 17689
rect -1135 17455 -901 17689
rect -901 17455 -900 17689
rect -1136 17454 -900 17455
rect -1136 17049 -900 17050
rect -1136 16815 -1135 17049
rect -1135 16815 -901 17049
rect -901 16815 -900 17049
rect -1136 16814 -900 16815
rect -1136 16409 -900 16410
rect -1136 16175 -1135 16409
rect -1135 16175 -901 16409
rect -901 16175 -900 16409
rect -1136 16174 -900 16175
rect -1136 15769 -900 15770
rect -1136 15535 -1135 15769
rect -1135 15535 -901 15769
rect -901 15535 -900 15769
rect -1136 15534 -900 15535
rect -1136 15129 -900 15130
rect -1136 14895 -1135 15129
rect -1135 14895 -901 15129
rect -901 14895 -900 15129
rect -1136 14894 -900 14895
rect -1136 14489 -900 14490
rect -1136 14255 -1135 14489
rect -1135 14255 -901 14489
rect -901 14255 -900 14489
rect -1136 14254 -900 14255
rect -1136 13849 -900 13850
rect -1136 13615 -1135 13849
rect -1135 13615 -901 13849
rect -901 13615 -900 13849
rect -1136 13614 -900 13615
rect -1136 13209 -900 13210
rect -1136 12975 -1135 13209
rect -1135 12975 -901 13209
rect -901 12975 -900 13209
rect -1136 12974 -900 12975
rect -1136 12569 -900 12570
rect -1136 12335 -1135 12569
rect -1135 12335 -901 12569
rect -901 12335 -900 12569
rect -1136 12334 -900 12335
rect -1136 11929 -900 11930
rect -1136 11695 -1135 11929
rect -1135 11695 -901 11929
rect -901 11695 -900 11929
rect -1136 11694 -900 11695
rect -1136 11289 -900 11290
rect -1136 11055 -1135 11289
rect -1135 11055 -901 11289
rect -901 11055 -900 11289
rect -1136 11054 -900 11055
rect -1136 10649 -900 10650
rect -1136 10415 -1135 10649
rect -1135 10415 -901 10649
rect -901 10415 -900 10649
rect -1136 10414 -900 10415
rect -1136 10009 -900 10010
rect -1136 9775 -1135 10009
rect -1135 9775 -901 10009
rect -901 9775 -900 10009
rect -1136 9774 -900 9775
rect -1136 9369 -900 9370
rect -1136 9135 -1135 9369
rect -1135 9135 -901 9369
rect -901 9135 -900 9369
rect -1136 9134 -900 9135
rect -1136 8729 -900 8730
rect -1136 8495 -1135 8729
rect -1135 8495 -901 8729
rect -901 8495 -900 8729
rect -1136 8494 -900 8495
rect -1136 8089 -900 8090
rect -1136 7855 -1135 8089
rect -1135 7855 -901 8089
rect -901 7855 -900 8089
rect -1136 7854 -900 7855
rect -1136 7449 -900 7450
rect -1136 7215 -1135 7449
rect -1135 7215 -901 7449
rect -901 7215 -900 7449
rect -1136 7214 -900 7215
rect -1136 6809 -900 6810
rect -1136 6575 -1135 6809
rect -1135 6575 -901 6809
rect -901 6575 -900 6809
rect -1136 6574 -900 6575
rect -1136 6169 -900 6170
rect -1136 5935 -1135 6169
rect -1135 5935 -901 6169
rect -901 5935 -900 6169
rect -1136 5934 -900 5935
rect -1136 5529 -900 5530
rect -1136 5295 -1135 5529
rect -1135 5295 -901 5529
rect -901 5295 -900 5529
rect -1136 5294 -900 5295
rect -580 27609 -260 27610
rect -580 27375 -579 27609
rect -579 27375 -261 27609
rect -261 27375 -260 27609
rect -580 27374 -260 27375
rect -580 26969 -260 26970
rect -580 26735 -579 26969
rect -579 26735 -261 26969
rect -261 26735 -260 26969
rect -580 26734 -260 26735
rect -580 26329 -260 26330
rect -580 26095 -579 26329
rect -579 26095 -261 26329
rect -261 26095 -260 26329
rect -580 26094 -260 26095
rect -580 25689 -260 25690
rect -580 25455 -579 25689
rect -579 25455 -261 25689
rect -261 25455 -260 25689
rect -580 25454 -260 25455
rect -580 25049 -260 25050
rect -580 24815 -579 25049
rect -579 24815 -261 25049
rect -261 24815 -260 25049
rect -580 24814 -260 24815
rect -580 24409 -260 24410
rect -580 24175 -579 24409
rect -579 24175 -261 24409
rect -261 24175 -260 24409
rect -580 24174 -260 24175
rect -580 23769 -260 23770
rect -580 23535 -579 23769
rect -579 23535 -261 23769
rect -261 23535 -260 23769
rect -580 23534 -260 23535
rect -580 23129 -260 23130
rect -580 22895 -579 23129
rect -579 22895 -261 23129
rect -261 22895 -260 23129
rect -580 22894 -260 22895
rect -580 22489 -260 22490
rect -580 22255 -579 22489
rect -579 22255 -261 22489
rect -261 22255 -260 22489
rect -580 22254 -260 22255
rect -580 21849 -260 21850
rect -580 21615 -579 21849
rect -579 21615 -261 21849
rect -261 21615 -260 21849
rect -580 21614 -260 21615
rect -580 21209 -260 21210
rect -580 20975 -579 21209
rect -579 20975 -261 21209
rect -261 20975 -260 21209
rect -580 20974 -260 20975
rect -580 20569 -260 20570
rect -580 20335 -579 20569
rect -579 20335 -261 20569
rect -261 20335 -260 20569
rect -580 20334 -260 20335
rect -580 19929 -260 19930
rect -580 19695 -579 19929
rect -579 19695 -261 19929
rect -261 19695 -260 19929
rect -580 19694 -260 19695
rect -580 19289 -260 19290
rect -580 19055 -579 19289
rect -579 19055 -261 19289
rect -261 19055 -260 19289
rect -580 19054 -260 19055
rect -580 18649 -260 18650
rect -580 18415 -579 18649
rect -579 18415 -261 18649
rect -261 18415 -260 18649
rect -580 18414 -260 18415
rect -580 18009 -260 18010
rect -580 17775 -579 18009
rect -579 17775 -261 18009
rect -261 17775 -260 18009
rect -580 17774 -260 17775
rect -580 17369 -260 17370
rect -580 17135 -579 17369
rect -579 17135 -261 17369
rect -261 17135 -260 17369
rect -580 17134 -260 17135
rect -580 16729 -260 16730
rect -580 16495 -579 16729
rect -579 16495 -261 16729
rect -261 16495 -260 16729
rect -580 16494 -260 16495
rect -580 16089 -260 16090
rect -580 15855 -579 16089
rect -579 15855 -261 16089
rect -261 15855 -260 16089
rect -580 15854 -260 15855
rect -580 15449 -260 15450
rect -580 15215 -579 15449
rect -579 15215 -261 15449
rect -261 15215 -260 15449
rect -580 15214 -260 15215
rect -580 14809 -260 14810
rect -580 14575 -579 14809
rect -579 14575 -261 14809
rect -261 14575 -260 14809
rect -580 14574 -260 14575
rect -580 14169 -260 14170
rect -580 13935 -579 14169
rect -579 13935 -261 14169
rect -261 13935 -260 14169
rect -580 13934 -260 13935
rect -580 13529 -260 13530
rect -580 13295 -579 13529
rect -579 13295 -261 13529
rect -261 13295 -260 13529
rect -580 13294 -260 13295
rect -580 12889 -260 12890
rect -580 12655 -579 12889
rect -579 12655 -261 12889
rect -261 12655 -260 12889
rect -580 12654 -260 12655
rect -580 12249 -260 12250
rect -580 12015 -579 12249
rect -579 12015 -261 12249
rect -261 12015 -260 12249
rect -580 12014 -260 12015
rect -580 11609 -260 11610
rect -580 11375 -579 11609
rect -579 11375 -261 11609
rect -261 11375 -260 11609
rect -580 11374 -260 11375
rect -580 10969 -260 10970
rect -580 10735 -579 10969
rect -579 10735 -261 10969
rect -261 10735 -260 10969
rect -580 10734 -260 10735
rect -580 10329 -260 10330
rect -580 10095 -579 10329
rect -579 10095 -261 10329
rect -261 10095 -260 10329
rect -580 10094 -260 10095
rect -580 9689 -260 9690
rect -580 9455 -579 9689
rect -579 9455 -261 9689
rect -261 9455 -260 9689
rect -580 9454 -260 9455
rect -580 9049 -260 9050
rect -580 8815 -579 9049
rect -579 8815 -261 9049
rect -261 8815 -260 9049
rect -580 8814 -260 8815
rect -580 8409 -260 8410
rect -580 8175 -579 8409
rect -579 8175 -261 8409
rect -261 8175 -260 8409
rect -580 8174 -260 8175
rect -580 7769 -260 7770
rect -580 7535 -579 7769
rect -579 7535 -261 7769
rect -261 7535 -260 7769
rect -580 7534 -260 7535
rect -580 7129 -260 7130
rect -580 6895 -579 7129
rect -579 6895 -261 7129
rect -261 6895 -260 7129
rect -580 6894 -260 6895
rect -580 6489 -260 6490
rect -580 6255 -579 6489
rect -579 6255 -261 6489
rect -261 6255 -260 6489
rect -580 6254 -260 6255
rect -580 5849 -260 5850
rect -580 5615 -579 5849
rect -579 5615 -261 5849
rect -261 5615 -260 5849
rect -580 5614 -260 5615
rect 60 27929 296 27930
rect 60 27695 61 27929
rect 61 27695 295 27929
rect 295 27695 296 27929
rect 60 27694 296 27695
rect 60 27289 296 27290
rect 60 27055 61 27289
rect 61 27055 295 27289
rect 295 27055 296 27289
rect 60 27054 296 27055
rect 60 26649 296 26650
rect 60 26415 61 26649
rect 61 26415 295 26649
rect 295 26415 296 26649
rect 60 26414 296 26415
rect 60 26009 296 26010
rect 60 25775 61 26009
rect 61 25775 295 26009
rect 295 25775 296 26009
rect 60 25774 296 25775
rect 60 25369 296 25370
rect 60 25135 61 25369
rect 61 25135 295 25369
rect 295 25135 296 25369
rect 60 25134 296 25135
rect 60 24729 296 24730
rect 60 24495 61 24729
rect 61 24495 295 24729
rect 295 24495 296 24729
rect 60 24494 296 24495
rect 60 24089 296 24090
rect 60 23855 61 24089
rect 61 23855 295 24089
rect 295 23855 296 24089
rect 60 23854 296 23855
rect 60 23449 296 23450
rect 60 23215 61 23449
rect 61 23215 295 23449
rect 295 23215 296 23449
rect 60 23214 296 23215
rect 60 22809 296 22810
rect 60 22575 61 22809
rect 61 22575 295 22809
rect 295 22575 296 22809
rect 60 22574 296 22575
rect 60 22169 296 22170
rect 60 21935 61 22169
rect 61 21935 295 22169
rect 295 21935 296 22169
rect 60 21934 296 21935
rect 60 21529 296 21530
rect 60 21295 61 21529
rect 61 21295 295 21529
rect 295 21295 296 21529
rect 60 21294 296 21295
rect 60 20889 296 20890
rect 60 20655 61 20889
rect 61 20655 295 20889
rect 295 20655 296 20889
rect 60 20654 296 20655
rect 60 20249 296 20250
rect 60 20015 61 20249
rect 61 20015 295 20249
rect 295 20015 296 20249
rect 60 20014 296 20015
rect 60 19609 296 19610
rect 60 19375 61 19609
rect 61 19375 295 19609
rect 295 19375 296 19609
rect 60 19374 296 19375
rect 60 18969 296 18970
rect 60 18735 61 18969
rect 61 18735 295 18969
rect 295 18735 296 18969
rect 60 18734 296 18735
rect 60 18329 296 18330
rect 60 18095 61 18329
rect 61 18095 295 18329
rect 295 18095 296 18329
rect 60 18094 296 18095
rect 60 17689 296 17690
rect 60 17455 61 17689
rect 61 17455 295 17689
rect 295 17455 296 17689
rect 60 17454 296 17455
rect 60 17049 296 17050
rect 60 16815 61 17049
rect 61 16815 295 17049
rect 295 16815 296 17049
rect 60 16814 296 16815
rect 60 16409 296 16410
rect 60 16175 61 16409
rect 61 16175 295 16409
rect 295 16175 296 16409
rect 60 16174 296 16175
rect 60 15769 296 15770
rect 60 15535 61 15769
rect 61 15535 295 15769
rect 295 15535 296 15769
rect 60 15534 296 15535
rect 60 15129 296 15130
rect 60 14895 61 15129
rect 61 14895 295 15129
rect 295 14895 296 15129
rect 60 14894 296 14895
rect 60 14489 296 14490
rect 60 14255 61 14489
rect 61 14255 295 14489
rect 295 14255 296 14489
rect 60 14254 296 14255
rect 60 13849 296 13850
rect 60 13615 61 13849
rect 61 13615 295 13849
rect 295 13615 296 13849
rect 60 13614 296 13615
rect 60 13209 296 13210
rect 60 12975 61 13209
rect 61 12975 295 13209
rect 295 12975 296 13209
rect 60 12974 296 12975
rect 60 12569 296 12570
rect 60 12335 61 12569
rect 61 12335 295 12569
rect 295 12335 296 12569
rect 60 12334 296 12335
rect 60 11929 296 11930
rect 60 11695 61 11929
rect 61 11695 295 11929
rect 295 11695 296 11929
rect 60 11694 296 11695
rect 60 11289 296 11290
rect 60 11055 61 11289
rect 61 11055 295 11289
rect 295 11055 296 11289
rect 60 11054 296 11055
rect 60 10649 296 10650
rect 60 10415 61 10649
rect 61 10415 295 10649
rect 295 10415 296 10649
rect 60 10414 296 10415
rect 60 10009 296 10010
rect 60 9775 61 10009
rect 61 9775 295 10009
rect 295 9775 296 10009
rect 60 9774 296 9775
rect 60 9369 296 9370
rect 60 9135 61 9369
rect 61 9135 295 9369
rect 295 9135 296 9369
rect 60 9134 296 9135
rect 60 8729 296 8730
rect 60 8495 61 8729
rect 61 8495 295 8729
rect 295 8495 296 8729
rect 60 8494 296 8495
rect 60 8089 296 8090
rect 60 7855 61 8089
rect 61 7855 295 8089
rect 295 7855 296 8089
rect 60 7854 296 7855
rect 60 7449 296 7450
rect 60 7215 61 7449
rect 61 7215 295 7449
rect 295 7215 296 7449
rect 60 7214 296 7215
rect 60 6809 296 6810
rect 60 6575 61 6809
rect 61 6575 295 6809
rect 295 6575 296 6809
rect 60 6574 296 6575
rect 60 6169 296 6170
rect 60 5935 61 6169
rect 61 5935 295 6169
rect 295 5935 296 6169
rect 60 5934 296 5935
rect 60 5529 296 5530
rect 60 5295 61 5529
rect 61 5295 295 5529
rect 295 5295 296 5529
rect 60 5294 296 5295
rect 684 3977 920 3978
rect 684 3743 685 3977
rect 685 3743 919 3977
rect 919 3743 920 3977
rect 684 3742 920 3743
rect 1324 3977 1560 3978
rect 1324 3743 1325 3977
rect 1325 3743 1559 3977
rect 1559 3743 1560 3977
rect 1324 3742 1560 3743
rect 1964 3977 2200 3978
rect 1964 3743 1965 3977
rect 1965 3743 2199 3977
rect 2199 3743 2200 3977
rect 1964 3742 2200 3743
rect 2604 3977 2840 3978
rect 2604 3743 2605 3977
rect 2605 3743 2839 3977
rect 2839 3743 2840 3977
rect 2604 3742 2840 3743
rect 3244 3977 3480 3978
rect 3244 3743 3245 3977
rect 3245 3743 3479 3977
rect 3479 3743 3480 3977
rect 3244 3742 3480 3743
rect 3884 3977 4120 3978
rect 3884 3743 3885 3977
rect 3885 3743 4119 3977
rect 4119 3743 4120 3977
rect 3884 3742 4120 3743
rect 4524 3977 4760 3978
rect 4524 3743 4525 3977
rect 4525 3743 4759 3977
rect 4759 3743 4760 3977
rect 4524 3742 4760 3743
rect 5164 3977 5400 3978
rect 5164 3743 5165 3977
rect 5165 3743 5399 3977
rect 5399 3743 5400 3977
rect 5164 3742 5400 3743
rect 5804 3977 6040 3978
rect 5804 3743 5805 3977
rect 5805 3743 6039 3977
rect 6039 3743 6040 3977
rect 5804 3742 6040 3743
rect 6444 3977 6680 3978
rect 6444 3743 6445 3977
rect 6445 3743 6679 3977
rect 6679 3743 6680 3977
rect 6444 3742 6680 3743
rect 7084 3977 7320 3978
rect 7084 3743 7085 3977
rect 7085 3743 7319 3977
rect 7319 3743 7320 3977
rect 7084 3742 7320 3743
rect 7724 3977 7960 3978
rect 7724 3743 7725 3977
rect 7725 3743 7959 3977
rect 7959 3743 7960 3977
rect 7724 3742 7960 3743
rect 8364 3977 8600 3978
rect 8364 3743 8365 3977
rect 8365 3743 8599 3977
rect 8599 3743 8600 3977
rect 8364 3742 8600 3743
rect 9004 3977 9240 3978
rect 9004 3743 9005 3977
rect 9005 3743 9239 3977
rect 9239 3743 9240 3977
rect 9004 3742 9240 3743
rect 9644 3977 9880 3978
rect 9644 3743 9645 3977
rect 9645 3743 9879 3977
rect 9879 3743 9880 3977
rect 9644 3742 9880 3743
rect 10284 3977 10520 3978
rect 10284 3743 10285 3977
rect 10285 3743 10519 3977
rect 10519 3743 10520 3977
rect 10284 3742 10520 3743
rect 10924 3977 11160 3978
rect 10924 3743 10925 3977
rect 10925 3743 11159 3977
rect 11159 3743 11160 3977
rect 10924 3742 11160 3743
rect 11564 3977 11800 3978
rect 11564 3743 11565 3977
rect 11565 3743 11799 3977
rect 11799 3743 11800 3977
rect 11564 3742 11800 3743
rect 12204 3977 12440 3978
rect 12204 3743 12205 3977
rect 12205 3743 12439 3977
rect 12439 3743 12440 3977
rect 12204 3742 12440 3743
rect 12844 3977 13080 3978
rect 12844 3743 12845 3977
rect 12845 3743 13079 3977
rect 13079 3743 13080 3977
rect 12844 3742 13080 3743
rect 13484 3977 13720 3978
rect 13484 3743 13485 3977
rect 13485 3743 13719 3977
rect 13719 3743 13720 3977
rect 13484 3742 13720 3743
rect 14124 3977 14360 3978
rect 14124 3743 14125 3977
rect 14125 3743 14359 3977
rect 14359 3743 14360 3977
rect 14124 3742 14360 3743
rect 14764 3977 15000 3978
rect 14764 3743 14765 3977
rect 14765 3743 14999 3977
rect 14999 3743 15000 3977
rect 14764 3742 15000 3743
rect 15404 3977 15640 3978
rect 15404 3743 15405 3977
rect 15405 3743 15639 3977
rect 15639 3743 15640 3977
rect 15404 3742 15640 3743
rect 16044 3977 16280 3978
rect 16044 3743 16045 3977
rect 16045 3743 16279 3977
rect 16279 3743 16280 3977
rect 16044 3742 16280 3743
rect 16684 3977 16920 3978
rect 16684 3743 16685 3977
rect 16685 3743 16919 3977
rect 16919 3743 16920 3977
rect 16684 3742 16920 3743
rect 17324 3977 17560 3978
rect 17324 3743 17325 3977
rect 17325 3743 17559 3977
rect 17559 3743 17560 3977
rect 17324 3742 17560 3743
rect 17964 3977 18200 3978
rect 17964 3743 17965 3977
rect 17965 3743 18199 3977
rect 18199 3743 18200 3977
rect 17964 3742 18200 3743
rect 18604 3977 18840 3978
rect 18604 3743 18605 3977
rect 18605 3743 18839 3977
rect 18839 3743 18840 3977
rect 18604 3742 18840 3743
rect 19244 3977 19480 3978
rect 19244 3743 19245 3977
rect 19245 3743 19479 3977
rect 19479 3743 19480 3977
rect 19244 3742 19480 3743
rect 19884 3977 20120 3978
rect 19884 3743 19885 3977
rect 19885 3743 20119 3977
rect 20119 3743 20120 3977
rect 19884 3742 20120 3743
rect 20524 3977 20760 3978
rect 20524 3743 20525 3977
rect 20525 3743 20759 3977
rect 20759 3743 20760 3977
rect 20524 3742 20760 3743
rect 21164 3977 21400 3978
rect 21164 3743 21165 3977
rect 21165 3743 21399 3977
rect 21399 3743 21400 3977
rect 21164 3742 21400 3743
rect 21804 3977 22040 3978
rect 21804 3743 21805 3977
rect 21805 3743 22039 3977
rect 22039 3743 22040 3977
rect 21804 3742 22040 3743
rect 364 3421 600 3422
rect 364 3103 365 3421
rect 365 3103 599 3421
rect 599 3103 600 3421
rect 364 3102 600 3103
rect 1004 3421 1240 3422
rect 1004 3103 1005 3421
rect 1005 3103 1239 3421
rect 1239 3103 1240 3421
rect 1004 3102 1240 3103
rect 1644 3421 1880 3422
rect 1644 3103 1645 3421
rect 1645 3103 1879 3421
rect 1879 3103 1880 3421
rect 1644 3102 1880 3103
rect 2284 3421 2520 3422
rect 2284 3103 2285 3421
rect 2285 3103 2519 3421
rect 2519 3103 2520 3421
rect 2284 3102 2520 3103
rect 2924 3421 3160 3422
rect 2924 3103 2925 3421
rect 2925 3103 3159 3421
rect 3159 3103 3160 3421
rect 2924 3102 3160 3103
rect 3564 3421 3800 3422
rect 3564 3103 3565 3421
rect 3565 3103 3799 3421
rect 3799 3103 3800 3421
rect 3564 3102 3800 3103
rect 4204 3421 4440 3422
rect 4204 3103 4205 3421
rect 4205 3103 4439 3421
rect 4439 3103 4440 3421
rect 4204 3102 4440 3103
rect 4844 3421 5080 3422
rect 4844 3103 4845 3421
rect 4845 3103 5079 3421
rect 5079 3103 5080 3421
rect 4844 3102 5080 3103
rect 5484 3421 5720 3422
rect 5484 3103 5485 3421
rect 5485 3103 5719 3421
rect 5719 3103 5720 3421
rect 5484 3102 5720 3103
rect 6124 3421 6360 3422
rect 6124 3103 6125 3421
rect 6125 3103 6359 3421
rect 6359 3103 6360 3421
rect 6124 3102 6360 3103
rect 6764 3421 7000 3422
rect 6764 3103 6765 3421
rect 6765 3103 6999 3421
rect 6999 3103 7000 3421
rect 6764 3102 7000 3103
rect 7404 3421 7640 3422
rect 7404 3103 7405 3421
rect 7405 3103 7639 3421
rect 7639 3103 7640 3421
rect 7404 3102 7640 3103
rect 8044 3421 8280 3422
rect 8044 3103 8045 3421
rect 8045 3103 8279 3421
rect 8279 3103 8280 3421
rect 8044 3102 8280 3103
rect 8684 3421 8920 3422
rect 8684 3103 8685 3421
rect 8685 3103 8919 3421
rect 8919 3103 8920 3421
rect 8684 3102 8920 3103
rect 9324 3421 9560 3422
rect 9324 3103 9325 3421
rect 9325 3103 9559 3421
rect 9559 3103 9560 3421
rect 9324 3102 9560 3103
rect 9964 3421 10200 3422
rect 9964 3103 9965 3421
rect 9965 3103 10199 3421
rect 10199 3103 10200 3421
rect 9964 3102 10200 3103
rect 10604 3421 10840 3422
rect 10604 3103 10605 3421
rect 10605 3103 10839 3421
rect 10839 3103 10840 3421
rect 10604 3102 10840 3103
rect 11244 3421 11480 3422
rect 11244 3103 11245 3421
rect 11245 3103 11479 3421
rect 11479 3103 11480 3421
rect 11244 3102 11480 3103
rect 11884 3421 12120 3422
rect 11884 3103 11885 3421
rect 11885 3103 12119 3421
rect 12119 3103 12120 3421
rect 11884 3102 12120 3103
rect 12524 3421 12760 3422
rect 12524 3103 12525 3421
rect 12525 3103 12759 3421
rect 12759 3103 12760 3421
rect 12524 3102 12760 3103
rect 13164 3421 13400 3422
rect 13164 3103 13165 3421
rect 13165 3103 13399 3421
rect 13399 3103 13400 3421
rect 13164 3102 13400 3103
rect 13804 3421 14040 3422
rect 13804 3103 13805 3421
rect 13805 3103 14039 3421
rect 14039 3103 14040 3421
rect 13804 3102 14040 3103
rect 14444 3421 14680 3422
rect 14444 3103 14445 3421
rect 14445 3103 14679 3421
rect 14679 3103 14680 3421
rect 14444 3102 14680 3103
rect 15084 3421 15320 3422
rect 15084 3103 15085 3421
rect 15085 3103 15319 3421
rect 15319 3103 15320 3421
rect 15084 3102 15320 3103
rect 15724 3421 15960 3422
rect 15724 3103 15725 3421
rect 15725 3103 15959 3421
rect 15959 3103 15960 3421
rect 15724 3102 15960 3103
rect 16364 3421 16600 3422
rect 16364 3103 16365 3421
rect 16365 3103 16599 3421
rect 16599 3103 16600 3421
rect 16364 3102 16600 3103
rect 17004 3421 17240 3422
rect 17004 3103 17005 3421
rect 17005 3103 17239 3421
rect 17239 3103 17240 3421
rect 17004 3102 17240 3103
rect 17644 3421 17880 3422
rect 17644 3103 17645 3421
rect 17645 3103 17879 3421
rect 17879 3103 17880 3421
rect 17644 3102 17880 3103
rect 18284 3421 18520 3422
rect 18284 3103 18285 3421
rect 18285 3103 18519 3421
rect 18519 3103 18520 3421
rect 18284 3102 18520 3103
rect 18924 3421 19160 3422
rect 18924 3103 18925 3421
rect 18925 3103 19159 3421
rect 19159 3103 19160 3421
rect 18924 3102 19160 3103
rect 19564 3421 19800 3422
rect 19564 3103 19565 3421
rect 19565 3103 19799 3421
rect 19799 3103 19800 3421
rect 19564 3102 19800 3103
rect 20204 3421 20440 3422
rect 20204 3103 20205 3421
rect 20205 3103 20439 3421
rect 20439 3103 20440 3421
rect 20204 3102 20440 3103
rect 20844 3421 21080 3422
rect 20844 3103 20845 3421
rect 20845 3103 21079 3421
rect 21079 3103 21080 3421
rect 20844 3102 21080 3103
rect 21484 3421 21720 3422
rect 21484 3103 21485 3421
rect 21485 3103 21719 3421
rect 21719 3103 21720 3421
rect 21484 3102 21720 3103
rect 22124 3421 22360 3422
rect 22124 3103 22125 3421
rect 22125 3103 22359 3421
rect 22359 3103 22360 3421
rect 22124 3102 22360 3103
rect 684 2781 920 2782
rect 684 2547 685 2781
rect 685 2547 919 2781
rect 919 2547 920 2781
rect 684 2546 920 2547
rect 1324 2781 1560 2782
rect 1324 2547 1325 2781
rect 1325 2547 1559 2781
rect 1559 2547 1560 2781
rect 1324 2546 1560 2547
rect 1964 2781 2200 2782
rect 1964 2547 1965 2781
rect 1965 2547 2199 2781
rect 2199 2547 2200 2781
rect 1964 2546 2200 2547
rect 2604 2781 2840 2782
rect 2604 2547 2605 2781
rect 2605 2547 2839 2781
rect 2839 2547 2840 2781
rect 2604 2546 2840 2547
rect 3244 2781 3480 2782
rect 3244 2547 3245 2781
rect 3245 2547 3479 2781
rect 3479 2547 3480 2781
rect 3244 2546 3480 2547
rect 3884 2781 4120 2782
rect 3884 2547 3885 2781
rect 3885 2547 4119 2781
rect 4119 2547 4120 2781
rect 3884 2546 4120 2547
rect 4524 2781 4760 2782
rect 4524 2547 4525 2781
rect 4525 2547 4759 2781
rect 4759 2547 4760 2781
rect 4524 2546 4760 2547
rect 5164 2781 5400 2782
rect 5164 2547 5165 2781
rect 5165 2547 5399 2781
rect 5399 2547 5400 2781
rect 5164 2546 5400 2547
rect 5804 2781 6040 2782
rect 5804 2547 5805 2781
rect 5805 2547 6039 2781
rect 6039 2547 6040 2781
rect 5804 2546 6040 2547
rect 6444 2781 6680 2782
rect 6444 2547 6445 2781
rect 6445 2547 6679 2781
rect 6679 2547 6680 2781
rect 6444 2546 6680 2547
rect 7084 2781 7320 2782
rect 7084 2547 7085 2781
rect 7085 2547 7319 2781
rect 7319 2547 7320 2781
rect 7084 2546 7320 2547
rect 7724 2781 7960 2782
rect 7724 2547 7725 2781
rect 7725 2547 7959 2781
rect 7959 2547 7960 2781
rect 7724 2546 7960 2547
rect 8364 2781 8600 2782
rect 8364 2547 8365 2781
rect 8365 2547 8599 2781
rect 8599 2547 8600 2781
rect 8364 2546 8600 2547
rect 9004 2781 9240 2782
rect 9004 2547 9005 2781
rect 9005 2547 9239 2781
rect 9239 2547 9240 2781
rect 9004 2546 9240 2547
rect 9644 2781 9880 2782
rect 9644 2547 9645 2781
rect 9645 2547 9879 2781
rect 9879 2547 9880 2781
rect 9644 2546 9880 2547
rect 10284 2781 10520 2782
rect 10284 2547 10285 2781
rect 10285 2547 10519 2781
rect 10519 2547 10520 2781
rect 10284 2546 10520 2547
rect 10924 2781 11160 2782
rect 10924 2547 10925 2781
rect 10925 2547 11159 2781
rect 11159 2547 11160 2781
rect 10924 2546 11160 2547
rect 11564 2781 11800 2782
rect 11564 2547 11565 2781
rect 11565 2547 11799 2781
rect 11799 2547 11800 2781
rect 11564 2546 11800 2547
rect 12204 2781 12440 2782
rect 12204 2547 12205 2781
rect 12205 2547 12439 2781
rect 12439 2547 12440 2781
rect 12204 2546 12440 2547
rect 12844 2781 13080 2782
rect 12844 2547 12845 2781
rect 12845 2547 13079 2781
rect 13079 2547 13080 2781
rect 12844 2546 13080 2547
rect 13484 2781 13720 2782
rect 13484 2547 13485 2781
rect 13485 2547 13719 2781
rect 13719 2547 13720 2781
rect 13484 2546 13720 2547
rect 14124 2781 14360 2782
rect 14124 2547 14125 2781
rect 14125 2547 14359 2781
rect 14359 2547 14360 2781
rect 14124 2546 14360 2547
rect 14764 2781 15000 2782
rect 14764 2547 14765 2781
rect 14765 2547 14999 2781
rect 14999 2547 15000 2781
rect 14764 2546 15000 2547
rect 15404 2781 15640 2782
rect 15404 2547 15405 2781
rect 15405 2547 15639 2781
rect 15639 2547 15640 2781
rect 15404 2546 15640 2547
rect 16044 2781 16280 2782
rect 16044 2547 16045 2781
rect 16045 2547 16279 2781
rect 16279 2547 16280 2781
rect 16044 2546 16280 2547
rect 16684 2781 16920 2782
rect 16684 2547 16685 2781
rect 16685 2547 16919 2781
rect 16919 2547 16920 2781
rect 16684 2546 16920 2547
rect 17324 2781 17560 2782
rect 17324 2547 17325 2781
rect 17325 2547 17559 2781
rect 17559 2547 17560 2781
rect 17324 2546 17560 2547
rect 17964 2781 18200 2782
rect 17964 2547 17965 2781
rect 17965 2547 18199 2781
rect 18199 2547 18200 2781
rect 17964 2546 18200 2547
rect 18604 2781 18840 2782
rect 18604 2547 18605 2781
rect 18605 2547 18839 2781
rect 18839 2547 18840 2781
rect 18604 2546 18840 2547
rect 19244 2781 19480 2782
rect 19244 2547 19245 2781
rect 19245 2547 19479 2781
rect 19479 2547 19480 2781
rect 19244 2546 19480 2547
rect 19884 2781 20120 2782
rect 19884 2547 19885 2781
rect 19885 2547 20119 2781
rect 20119 2547 20120 2781
rect 19884 2546 20120 2547
rect 20524 2781 20760 2782
rect 20524 2547 20525 2781
rect 20525 2547 20759 2781
rect 20759 2547 20760 2781
rect 20524 2546 20760 2547
rect 21164 2781 21400 2782
rect 21164 2547 21165 2781
rect 21165 2547 21399 2781
rect 21399 2547 21400 2781
rect 21164 2546 21400 2547
rect 21804 2781 22040 2782
rect 21804 2547 21805 2781
rect 21805 2547 22039 2781
rect 22039 2547 22040 2781
rect 21804 2546 22040 2547
<< metal5 >>
rect 20634 30537 20954 30585
rect 20634 30300 20659 30537
rect 20895 30300 20954 30537
rect -900 27972 -580 28197
rect -1160 27930 -580 27972
rect -1160 27694 -1136 27930
rect -900 27694 -580 27930
rect -1160 27652 -580 27694
rect -260 27972 60 28204
rect -260 27930 320 27972
rect -260 27694 60 27930
rect 296 27694 320 27930
rect -260 27652 320 27694
rect -900 27610 60 27652
rect -900 27374 -580 27610
rect -260 27374 60 27610
rect -900 27332 60 27374
rect -1160 27290 -580 27332
rect -1160 27054 -1136 27290
rect -900 27054 -580 27290
rect -1160 27012 -580 27054
rect -260 27290 320 27332
rect -260 27054 60 27290
rect 296 27054 320 27290
rect -260 27012 320 27054
rect -900 26970 60 27012
rect 20634 26985 20954 30300
rect -900 26734 -580 26970
rect -260 26734 60 26970
rect -900 26692 60 26734
rect -1160 26650 -580 26692
rect -1160 26414 -1136 26650
rect -900 26414 -580 26650
rect -1160 26372 -580 26414
rect -260 26650 320 26692
rect -260 26414 60 26650
rect 296 26414 320 26650
rect 12261 26560 12670 26880
rect -260 26372 320 26414
rect -900 26330 60 26372
rect -900 26094 -580 26330
rect -260 26094 60 26330
rect -900 26052 60 26094
rect -1160 26010 -580 26052
rect -1160 25774 -1136 26010
rect -900 25774 -580 26010
rect -1160 25732 -580 25774
rect -260 26010 832 26052
rect -260 25774 60 26010
rect 296 25774 832 26010
rect -260 25732 832 25774
rect -900 25690 60 25732
rect -900 25454 -580 25690
rect -260 25454 60 25690
rect -900 25412 60 25454
rect -1160 25370 -580 25412
rect -1160 25134 -1136 25370
rect -900 25134 -580 25370
rect -1160 25092 -580 25134
rect -260 25370 320 25412
rect -260 25134 60 25370
rect 296 25134 320 25370
rect -260 25092 320 25134
rect 12240 25129 12692 25449
rect -900 25050 60 25092
rect -900 24814 -580 25050
rect -260 24814 60 25050
rect -900 24772 60 24814
rect -1160 24730 -580 24772
rect -1160 24494 -1136 24730
rect -900 24494 -580 24730
rect -1160 24452 -580 24494
rect -260 24730 890 24772
rect -260 24494 60 24730
rect 296 24494 890 24730
rect -260 24452 890 24494
rect -900 24410 60 24452
rect -900 24174 -580 24410
rect -260 24174 60 24410
rect -900 24132 60 24174
rect -1160 24090 -580 24132
rect -1160 23854 -1136 24090
rect -900 23854 -580 24090
rect -1160 23812 -580 23854
rect -260 24090 320 24132
rect -260 23854 60 24090
rect 296 23854 320 24090
rect 12248 24007 12657 24327
rect -260 23812 320 23854
rect -900 23770 60 23812
rect -900 23534 -580 23770
rect -260 23534 60 23770
rect -900 23492 60 23534
rect -1160 23450 -580 23492
rect -1160 23214 -1136 23450
rect -900 23214 -580 23450
rect -1160 23172 -580 23214
rect -260 23450 888 23492
rect -260 23214 60 23450
rect 296 23214 888 23450
rect -260 23172 888 23214
rect -900 23130 60 23172
rect -900 22894 -580 23130
rect -260 22894 60 23130
rect 12258 23112 12667 23432
rect -900 22852 60 22894
rect -1160 22810 -580 22852
rect -1160 22574 -1136 22810
rect -900 22574 -580 22810
rect -1160 22532 -580 22574
rect -260 22810 320 22852
rect -260 22574 60 22810
rect 296 22574 320 22810
rect -260 22532 320 22574
rect -900 22490 60 22532
rect -900 22254 -580 22490
rect -260 22254 60 22490
rect -900 22212 60 22254
rect 12249 22229 12658 22549
rect -1160 22170 -580 22212
rect -1160 21934 -1136 22170
rect -900 21934 -580 22170
rect -1160 21892 -580 21934
rect -260 22170 872 22212
rect -260 21934 60 22170
rect 296 21934 872 22170
rect -260 21892 872 21934
rect -900 21850 60 21892
rect -900 21614 -580 21850
rect -260 21614 60 21850
rect -900 21572 60 21614
rect -1160 21530 -580 21572
rect -1160 21294 -1136 21530
rect -900 21294 -580 21530
rect -1160 21252 -580 21294
rect -260 21530 320 21572
rect -260 21294 60 21530
rect 296 21294 320 21530
rect -260 21252 320 21294
rect -900 21210 60 21252
rect -900 20974 -580 21210
rect -260 20974 60 21210
rect -900 20932 60 20974
rect -1160 20890 -580 20932
rect -1160 20654 -1136 20890
rect -900 20654 -580 20890
rect -1160 20612 -580 20654
rect -260 20890 890 20932
rect -260 20654 60 20890
rect 296 20654 890 20890
rect -260 20612 890 20654
rect -900 20570 60 20612
rect -900 20334 -580 20570
rect -260 20334 60 20570
rect 12268 20525 12677 20845
rect -900 20292 60 20334
rect -1160 20250 -580 20292
rect -1160 20014 -1136 20250
rect -900 20014 -580 20250
rect -1160 19972 -580 20014
rect -260 20250 320 20292
rect -260 20014 60 20250
rect 296 20014 320 20250
rect -260 19972 320 20014
rect -900 19930 60 19972
rect -900 19694 -580 19930
rect -260 19694 60 19930
rect -900 19652 60 19694
rect -1160 19610 -580 19652
rect -1160 19374 -1136 19610
rect -900 19374 -580 19610
rect -1160 19332 -580 19374
rect -260 19610 894 19652
rect 12263 19643 12672 19963
rect -260 19374 60 19610
rect 296 19374 894 19610
rect -260 19332 894 19374
rect -900 19290 60 19332
rect -900 19054 -580 19290
rect -260 19054 60 19290
rect -900 19012 60 19054
rect -1160 18970 -580 19012
rect -1160 18734 -1136 18970
rect -900 18734 -580 18970
rect -1160 18692 -580 18734
rect -260 18970 320 19012
rect -260 18734 60 18970
rect 296 18734 320 18970
rect 12274 18746 12683 19066
rect -260 18692 320 18734
rect -900 18650 60 18692
rect -900 18414 -580 18650
rect -260 18414 60 18650
rect -900 18372 60 18414
rect -1160 18330 -580 18372
rect -1160 18094 -1136 18330
rect -900 18094 -580 18330
rect -1160 18052 -580 18094
rect -260 18330 909 18372
rect -260 18094 60 18330
rect 296 18094 909 18330
rect -260 18052 909 18094
rect -900 18010 60 18052
rect -900 17774 -580 18010
rect -260 17774 60 18010
rect -900 17732 60 17774
rect -1160 17690 -580 17732
rect -1160 17454 -1136 17690
rect -900 17454 -580 17690
rect -1160 17412 -580 17454
rect -260 17690 320 17732
rect -260 17454 60 17690
rect 296 17454 320 17690
rect -260 17412 320 17454
rect -900 17370 60 17412
rect -900 17134 -580 17370
rect -260 17134 60 17370
rect -900 17092 60 17134
rect -1160 17050 -580 17092
rect -1160 16814 -1136 17050
rect -900 16814 -580 17050
rect -1160 16772 -580 16814
rect -260 17050 906 17092
rect 12263 17053 12672 17373
rect -260 16814 60 17050
rect 296 16814 906 17050
rect -260 16772 906 16814
rect -900 16730 60 16772
rect -900 16494 -580 16730
rect -260 16494 60 16730
rect -900 16452 60 16494
rect -1160 16410 -580 16452
rect -1160 16174 -1136 16410
rect -900 16174 -580 16410
rect -1160 16132 -580 16174
rect -260 16410 320 16452
rect -260 16174 60 16410
rect 296 16174 320 16410
rect -260 16132 320 16174
rect 12269 16155 12678 16475
rect -900 16090 60 16132
rect -900 15854 -580 16090
rect -260 15854 60 16090
rect -900 15812 60 15854
rect -1160 15770 -580 15812
rect -1160 15534 -1136 15770
rect -900 15534 -580 15770
rect -1160 15492 -580 15534
rect -260 15770 879 15812
rect -260 15534 60 15770
rect 296 15534 879 15770
rect -260 15492 879 15534
rect -900 15450 60 15492
rect -900 15214 -580 15450
rect -260 15214 60 15450
rect 12272 15262 12681 15582
rect -900 15172 60 15214
rect -1160 15130 -580 15172
rect -1160 14894 -1136 15130
rect -900 14894 -580 15130
rect -1160 14852 -580 14894
rect -260 15130 320 15172
rect -260 14894 60 15130
rect 296 14894 320 15130
rect -260 14852 320 14894
rect -900 14810 60 14852
rect -900 14574 -580 14810
rect -260 14574 60 14810
rect -900 14532 60 14574
rect -1160 14490 -580 14532
rect -1160 14254 -1136 14490
rect -900 14254 -580 14490
rect -1160 14212 -580 14254
rect -260 14490 879 14532
rect -260 14254 60 14490
rect 296 14254 879 14490
rect -260 14212 879 14254
rect -900 14170 60 14212
rect -900 13934 -580 14170
rect -260 13934 60 14170
rect -900 13892 60 13934
rect -1160 13850 -580 13892
rect -1160 13614 -1136 13850
rect -900 13614 -580 13850
rect -1160 13572 -580 13614
rect -260 13850 320 13892
rect -260 13614 60 13850
rect 296 13614 320 13850
rect -260 13572 320 13614
rect -900 13530 60 13572
rect 12277 13566 12686 13886
rect -900 13294 -580 13530
rect -260 13294 60 13530
rect -900 13252 60 13294
rect -1160 13210 -580 13252
rect -1160 12974 -1136 13210
rect -900 12974 -580 13210
rect -1160 12932 -580 12974
rect -260 13210 866 13252
rect -260 12974 60 13210
rect 296 12974 866 13210
rect -260 12932 866 12974
rect -900 12890 60 12932
rect -900 12654 -580 12890
rect -260 12654 60 12890
rect 12272 12673 12681 12993
rect -900 12612 60 12654
rect -1160 12570 -580 12612
rect -1160 12334 -1136 12570
rect -900 12334 -580 12570
rect -1160 12292 -580 12334
rect -260 12570 320 12612
rect -260 12334 60 12570
rect 296 12334 320 12570
rect -260 12292 320 12334
rect -900 12250 60 12292
rect -900 12014 -580 12250
rect -260 12014 60 12250
rect -900 11972 60 12014
rect -1160 11930 -580 11972
rect -1160 11694 -1136 11930
rect -900 11694 -580 11930
rect -1160 11652 -580 11694
rect -260 11930 863 11972
rect -260 11694 60 11930
rect 296 11694 863 11930
rect 12278 11778 12687 12098
rect -260 11652 863 11694
rect -900 11610 60 11652
rect -900 11374 -580 11610
rect -260 11374 60 11610
rect -900 11332 60 11374
rect -1160 11290 -580 11332
rect -1160 11054 -1136 11290
rect -900 11054 -580 11290
rect -1160 11012 -580 11054
rect -260 11290 320 11332
rect -260 11054 60 11290
rect 296 11054 320 11290
rect -260 11012 320 11054
rect -900 10970 60 11012
rect -900 10734 -580 10970
rect -260 10734 60 10970
rect -900 10692 60 10734
rect -1160 10650 -580 10692
rect -1160 10414 -1136 10650
rect -900 10414 -580 10650
rect -1160 10372 -580 10414
rect -260 10650 882 10692
rect -260 10414 60 10650
rect 296 10414 882 10650
rect -260 10372 882 10414
rect -900 10330 60 10372
rect -900 10094 -580 10330
rect -260 10094 60 10330
rect -900 10052 60 10094
rect 12276 10080 12685 10400
rect -1160 10010 -580 10052
rect -1160 9774 -1136 10010
rect -900 9774 -580 10010
rect -1160 9732 -580 9774
rect -260 10010 320 10052
rect -260 9774 60 10010
rect 296 9774 320 10010
rect -260 9732 320 9774
rect -900 9690 60 9732
rect -900 9454 -580 9690
rect -260 9454 60 9690
rect -900 9412 60 9454
rect -1160 9370 -580 9412
rect -1160 9134 -1136 9370
rect -900 9134 -580 9370
rect -1160 9092 -580 9134
rect -260 9370 798 9412
rect -260 9134 60 9370
rect 296 9134 798 9370
rect 12273 9187 12682 9507
rect -260 9092 798 9134
rect -900 9050 60 9092
rect -900 8814 -580 9050
rect -260 8814 60 9050
rect -900 8772 60 8814
rect -1160 8730 -580 8772
rect -1160 8494 -1136 8730
rect -900 8494 -580 8730
rect -1160 8452 -580 8494
rect -260 8730 320 8772
rect -260 8494 60 8730
rect 296 8494 320 8730
rect -260 8452 320 8494
rect -900 8410 60 8452
rect -900 8174 -580 8410
rect -260 8174 60 8410
rect 12269 8295 12671 8615
rect -900 8132 60 8174
rect -1160 8090 -580 8132
rect -1160 7854 -1136 8090
rect -900 7854 -580 8090
rect -1160 7812 -580 7854
rect -260 8090 865 8132
rect -260 7854 60 8090
rect 296 7854 865 8090
rect -260 7812 865 7854
rect -900 7770 60 7812
rect -900 7534 -580 7770
rect -260 7534 60 7770
rect -900 7492 60 7534
rect -1160 7450 -580 7492
rect -1160 7214 -1136 7450
rect -900 7214 -580 7450
rect -1160 7172 -580 7214
rect -260 7450 320 7492
rect -260 7214 60 7450
rect 296 7214 320 7450
rect -260 7172 320 7214
rect -900 7130 60 7172
rect -900 6894 -580 7130
rect -260 6894 60 7130
rect -900 6852 60 6894
rect -1160 6810 -580 6852
rect -1160 6574 -1136 6810
rect -900 6574 -580 6810
rect -1160 6532 -580 6574
rect -260 6810 901 6852
rect -260 6574 60 6810
rect 296 6574 901 6810
rect 12271 6599 12673 6919
rect -260 6532 901 6574
rect -900 6490 60 6532
rect -900 6254 -580 6490
rect -260 6254 60 6490
rect -900 6212 60 6254
rect -1160 6170 -580 6212
rect -1160 5934 -1136 6170
rect -900 5934 -580 6170
rect -1160 5892 -580 5934
rect -260 6170 320 6212
rect -260 5934 60 6170
rect 296 5934 320 6170
rect -260 5892 320 5934
rect -900 5850 60 5892
rect -900 5614 -580 5850
rect -260 5614 60 5850
rect 12275 5705 12677 6025
rect -900 5572 60 5614
rect -1160 5530 -580 5572
rect -1160 5294 -1136 5530
rect -900 5294 -580 5530
rect -1160 5252 -580 5294
rect -900 3742 -580 5252
rect -260 5530 838 5572
rect -260 5294 60 5530
rect 296 5294 838 5530
rect -260 5252 838 5294
rect -260 3742 60 5252
rect 12267 4811 12669 5131
rect 642 3978 962 4002
rect 642 3742 684 3978
rect 920 3742 962 3978
rect 1282 3978 1602 4591
rect 1282 3742 1324 3978
rect 1560 3742 1602 3978
rect 1922 3978 2242 4002
rect 1922 3742 1964 3978
rect 2200 3742 2242 3978
rect 2562 3978 2882 4589
rect 2562 3742 2604 3978
rect 2840 3742 2882 3978
rect 3202 3978 3522 4002
rect 3202 3742 3244 3978
rect 3480 3742 3522 3978
rect 3842 3978 4162 4592
rect 3842 3742 3884 3978
rect 4120 3742 4162 3978
rect 4482 3978 4802 4002
rect 4482 3742 4524 3978
rect 4760 3742 4802 3978
rect 5122 3978 5442 4590
rect 5122 3742 5164 3978
rect 5400 3742 5442 3978
rect 5762 3978 6082 4002
rect 5762 3742 5804 3978
rect 6040 3742 6082 3978
rect 6402 3978 6722 4591
rect 6402 3742 6444 3978
rect 6680 3742 6722 3978
rect 7042 3978 7362 4002
rect 7042 3742 7084 3978
rect 7320 3742 7362 3978
rect 7682 3978 8002 4590
rect 7682 3742 7724 3978
rect 7960 3742 8002 3978
rect 8322 3978 8642 4002
rect 8322 3742 8364 3978
rect 8600 3742 8642 3978
rect 8962 3978 9282 4591
rect 8962 3742 9004 3978
rect 9240 3742 9282 3978
rect 9602 3978 9922 4002
rect 9602 3742 9644 3978
rect 9880 3742 9922 3978
rect 10242 3978 10562 4592
rect 10242 3742 10284 3978
rect 10520 3742 10562 3978
rect 10882 3978 11202 4002
rect 10882 3742 10924 3978
rect 11160 3742 11202 3978
rect 11522 3978 11842 4592
rect 11522 3742 11564 3978
rect 11800 3742 11842 3978
rect 12162 3978 12482 4002
rect 12162 3742 12204 3978
rect 12440 3742 12482 3978
rect 12802 3978 13122 4591
rect 12802 3742 12844 3978
rect 13080 3742 13122 3978
rect 13442 3978 13762 4002
rect 13442 3742 13484 3978
rect 13720 3742 13762 3978
rect 14082 3978 14402 4002
rect 14082 3742 14124 3978
rect 14360 3742 14402 3978
rect 14722 3978 15042 4002
rect 14722 3742 14764 3978
rect 15000 3742 15042 3978
rect 15362 3978 15682 4590
rect 15362 3742 15404 3978
rect 15640 3742 15682 3978
rect 16002 3978 16322 4002
rect 16002 3742 16044 3978
rect 16280 3742 16322 3978
rect 16642 3978 16962 4592
rect 16642 3742 16684 3978
rect 16920 3742 16962 3978
rect 17282 3978 17602 4002
rect 17282 3742 17324 3978
rect 17560 3742 17602 3978
rect 17922 3978 18242 4589
rect 17922 3742 17964 3978
rect 18200 3742 18242 3978
rect 18562 3978 18882 4002
rect 18562 3742 18604 3978
rect 18840 3742 18882 3978
rect 19202 3978 19522 4002
rect 19202 3742 19244 3978
rect 19480 3742 19522 3978
rect 19842 3978 20162 4002
rect 19842 3742 19884 3978
rect 20120 3742 20162 3978
rect 20482 3978 20802 4002
rect 20482 3742 20524 3978
rect 20760 3742 20802 3978
rect 21122 3978 21442 4002
rect 21122 3742 21164 3978
rect 21400 3742 21442 3978
rect 21762 3978 22082 4002
rect 21762 3742 21804 3978
rect 22040 3742 22082 3978
rect -900 3422 22766 3742
rect -900 3102 -580 3422
rect 322 3102 364 3422
rect 600 3102 642 3422
rect 962 3102 1004 3422
rect 1240 3102 1282 3422
rect 1602 3102 1644 3422
rect 1880 3102 1922 3422
rect 2242 3102 2284 3422
rect 2520 3102 2562 3422
rect 2882 3102 2924 3422
rect 3160 3102 3202 3422
rect 3522 3102 3564 3422
rect 3800 3102 3842 3422
rect 4162 3102 4204 3422
rect 4440 3102 4482 3422
rect 4802 3102 4844 3422
rect 5080 3102 5122 3422
rect 5442 3102 5484 3422
rect 5720 3102 5762 3422
rect 6082 3102 6124 3422
rect 6360 3102 6402 3422
rect 6722 3102 6764 3422
rect 7000 3102 7042 3422
rect 7362 3102 7404 3422
rect 7640 3102 7682 3422
rect 8002 3102 8044 3422
rect 8280 3102 8322 3422
rect 8642 3102 8684 3422
rect 8920 3102 8962 3422
rect 9282 3102 9324 3422
rect 9560 3102 9602 3422
rect 9922 3102 9964 3422
rect 10200 3102 10242 3422
rect 10562 3102 10604 3422
rect 10840 3102 10882 3422
rect 11202 3102 11244 3422
rect 11480 3102 11522 3422
rect 11842 3102 11884 3422
rect 12120 3102 12162 3422
rect 12482 3102 12524 3422
rect 12760 3102 12802 3422
rect 13122 3102 13164 3422
rect 13400 3102 13442 3422
rect 13762 3102 13804 3422
rect 14040 3102 14082 3422
rect 14402 3102 14444 3422
rect 14680 3102 14722 3422
rect 15042 3102 15084 3422
rect 15320 3102 15362 3422
rect 15682 3102 15724 3422
rect 15960 3102 16002 3422
rect 16322 3102 16364 3422
rect 16600 3102 16642 3422
rect 16962 3102 17004 3422
rect 17240 3102 17282 3422
rect 17602 3102 17644 3422
rect 17880 3102 17922 3422
rect 18242 3102 18284 3422
rect 18520 3102 18562 3422
rect 18882 3102 18924 3422
rect 19160 3102 19202 3422
rect 19522 3102 19564 3422
rect 19800 3102 19842 3422
rect 20162 3102 20204 3422
rect 20440 3102 20482 3422
rect 20802 3102 20844 3422
rect 21080 3102 21122 3422
rect 21442 3102 21484 3422
rect 21720 3102 21762 3422
rect 22082 3102 22124 3422
rect 22360 3102 22402 3422
rect -900 2782 22766 3102
rect 642 2546 684 2782
rect 920 2546 962 2782
rect 642 2522 962 2546
rect 1282 2546 1324 2782
rect 1560 2546 1602 2782
rect 1282 2522 1602 2546
rect 1922 2546 1964 2782
rect 2200 2546 2242 2782
rect 1922 2522 2242 2546
rect 2562 2546 2604 2782
rect 2840 2546 2882 2782
rect 2562 2522 2882 2546
rect 3202 2546 3244 2782
rect 3480 2546 3522 2782
rect 3202 2522 3522 2546
rect 3842 2546 3884 2782
rect 4120 2546 4162 2782
rect 3842 2522 4162 2546
rect 4482 2546 4524 2782
rect 4760 2546 4802 2782
rect 4482 2522 4802 2546
rect 5122 2546 5164 2782
rect 5400 2546 5442 2782
rect 5122 2522 5442 2546
rect 5762 2546 5804 2782
rect 6040 2546 6082 2782
rect 5762 2522 6082 2546
rect 6402 2546 6444 2782
rect 6680 2546 6722 2782
rect 6402 2522 6722 2546
rect 7042 2546 7084 2782
rect 7320 2546 7362 2782
rect 7042 2522 7362 2546
rect 7682 2546 7724 2782
rect 7960 2546 8002 2782
rect 7682 2522 8002 2546
rect 8322 2546 8364 2782
rect 8600 2546 8642 2782
rect 8322 2522 8642 2546
rect 8962 2546 9004 2782
rect 9240 2546 9282 2782
rect 8962 2522 9282 2546
rect 9602 2546 9644 2782
rect 9880 2546 9922 2782
rect 9602 2522 9922 2546
rect 10242 2546 10284 2782
rect 10520 2546 10562 2782
rect 10242 2522 10562 2546
rect 10882 2546 10924 2782
rect 11160 2546 11202 2782
rect 10882 2522 11202 2546
rect 11522 2546 11564 2782
rect 11800 2546 11842 2782
rect 11522 2522 11842 2546
rect 12162 2546 12204 2782
rect 12440 2546 12482 2782
rect 12162 2522 12482 2546
rect 12802 2546 12844 2782
rect 13080 2546 13122 2782
rect 12802 2522 13122 2546
rect 13442 2546 13484 2782
rect 13720 2546 13762 2782
rect 13442 2522 13762 2546
rect 14082 2546 14124 2782
rect 14360 2546 14402 2782
rect 14082 2522 14402 2546
rect 14722 2546 14764 2782
rect 15000 2546 15042 2782
rect 14722 2522 15042 2546
rect 15362 2546 15404 2782
rect 15640 2546 15682 2782
rect 15362 2522 15682 2546
rect 16002 2546 16044 2782
rect 16280 2546 16322 2782
rect 16002 2522 16322 2546
rect 16642 2546 16684 2782
rect 16920 2546 16962 2782
rect 16642 2522 16962 2546
rect 17282 2546 17324 2782
rect 17560 2546 17602 2782
rect 17282 2522 17602 2546
rect 17922 2546 17964 2782
rect 18200 2546 18242 2782
rect 17922 2522 18242 2546
rect 18562 2546 18604 2782
rect 18840 2546 18882 2782
rect 18562 2522 18882 2546
rect 19202 2546 19244 2782
rect 19480 2546 19522 2782
rect 19202 2522 19522 2546
rect 19842 2546 19884 2782
rect 20120 2546 20162 2782
rect 19842 2522 20162 2546
rect 20482 2546 20524 2782
rect 20760 2546 20802 2782
rect 20482 2522 20802 2546
rect 21122 2546 21164 2782
rect 21400 2546 21442 2782
rect 21122 2522 21442 2546
rect 21762 2546 21804 2782
rect 22040 2546 22082 2782
rect 21762 2522 22082 2546
use analog_mux  analog_mux_0
timestamp 1654693421
transform 1 0 20673 0 1 30912
box -239 -36 446 2223
use cap_3pF  cap_3pF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654658877
transform 0 1 16965 -1 0 20343
box -6669 2096 15759 5484
use cap_6pF  cap_6pF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654661395
transform 0 1 15305 -1 0 24342
box -2674 -2673 19758 3439
use cap_10fF  cap_10fF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654685434
transform 1 0 18937 0 1 28644
box -28 -28 708 628
use cap_10fF  cap_10fF_1
timestamp 1654685434
transform 1 0 5164 0 1 28662
box -28 -28 708 628
use cap_12pF  cap_12pF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654661395
transform 0 1 3438 -1 0 24342
box -2674 -2674 19758 8878
use cap_20fF  cap_20fF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654307754
transform 1 0 12735 0 1 28665
box -28 -28 828 1028
use cap_40fF  cap_40fF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654602114
transform 1 0 901 0 1 28672
box -28 -28 1368 1228
use cmos_switch  cmos_switch_0 ~/Documents/fossi_cochlea/mag/final_designs/switch
timestamp 1654685434
transform 1 0 557 0 1 28398
box -175 -95 235 3570
use cmos_switch  cmos_switch_1
timestamp 1654685434
transform -1 0 2617 0 1 28398
box -175 -95 235 3570
use cmos_switch  cmos_switch_2
timestamp 1654685434
transform 1 0 12307 0 1 28398
box -175 -95 235 3570
use cmos_switch  cmos_switch_3
timestamp 1654685434
transform -1 0 13925 0 1 28398
box -175 -95 235 3570
use cmos_switch  cmos_switch_4
timestamp 1654685434
transform 1 0 18517 0 1 28398
box -175 -95 235 3570
use cmos_switch  cmos_switch_5
timestamp 1654685434
transform -1 0 20077 0 1 28398
box -175 -95 235 3570
use cmos_switch  cmos_switch_6
timestamp 1654685434
transform 1 0 4817 0 1 28398
box -175 -95 235 3570
use cmos_switch  cmos_switch_7
timestamp 1654685434
transform -1 0 6187 0 1 28398
box -175 -95 235 3570
use mux  mux_0 ~/Documents/fossi_cochlea/mag/final_designs/mux
timestamp 1654666893
transform 0 -1 -104 1 0 28489
box -224 -79 685 681
<< labels >>
rlabel metal1 -637 32252 -637 32252 7 phi1
rlabel metal1 -637 32375 -637 32375 7 phi1b
rlabel metal1 -637 32494 -637 32494 7 phi2
rlabel metal1 -637 32612 -637 32612 7 phi2b
rlabel metal1 -637 32733 -637 32733 7 ctrl
rlabel metal1 -637 32852 -637 32852 7 ctrlb
<< end >>
