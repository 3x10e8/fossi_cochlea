VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO /local_disk/fossi_cochlea/mag/final_designs/filter_p_m
  CLASS BLOCK ;
  FOREIGN /local_disk/fossi_cochlea/mag/final_designs/filter_p_m ;
  ORIGIN 0.130 1.640 ;
  SIZE 253.920 BY 187.340 ;
  PIN th1
    DIRECTION INOUT ;
    ANTENNADIFFAREA 0.554400 ;
    PORT
      LAYER li1 ;
        RECT 109.395 143.815 109.670 144.195 ;
        RECT 129.695 143.775 129.995 144.195 ;
        RECT 109.395 141.900 109.670 142.280 ;
        RECT 129.695 141.900 129.995 142.320 ;
      LAYER mcon ;
        RECT 109.440 143.905 109.610 144.075 ;
        RECT 129.735 143.885 129.905 144.055 ;
        RECT 109.440 142.020 109.610 142.190 ;
        RECT 129.735 142.040 129.905 142.210 ;
      LAYER met1 ;
        RECT 109.400 144.135 109.660 144.155 ;
        RECT 109.380 143.865 109.670 144.135 ;
        RECT 129.700 144.115 129.960 144.140 ;
        RECT 109.400 143.835 109.660 143.865 ;
        RECT 109.440 142.250 109.610 143.835 ;
        RECT 129.675 143.825 129.965 144.115 ;
        RECT 129.700 143.820 129.960 143.825 ;
        RECT 129.735 142.270 129.905 143.820 ;
        RECT 109.380 141.960 109.670 142.250 ;
        RECT 129.675 141.980 129.965 142.270 ;
      LAYER via ;
        RECT 109.400 143.865 109.660 144.125 ;
        RECT 129.700 143.850 129.960 144.110 ;
      LAYER met2 ;
        RECT 108.505 153.465 108.785 153.835 ;
        RECT 129.675 153.500 129.955 153.870 ;
        RECT 108.570 152.405 108.740 153.465 ;
        RECT 108.565 144.075 108.745 152.405 ;
        RECT 109.400 144.075 109.660 144.155 ;
        RECT 129.730 144.140 129.900 153.500 ;
        RECT 108.565 143.905 109.660 144.075 ;
        RECT 108.565 142.215 108.745 143.905 ;
        RECT 109.400 143.835 109.660 143.905 ;
        RECT 129.700 143.820 129.960 144.140 ;
        RECT 108.565 142.025 109.610 142.215 ;
        RECT 129.730 142.160 129.900 143.820 ;
      LAYER via2 ;
        RECT 108.505 153.510 108.785 153.790 ;
        RECT 129.675 153.545 129.955 153.825 ;
      LAYER met3 ;
        RECT -0.130 153.430 253.790 153.930 ;
    END
  END th1
  PIN th2
    DIRECTION INOUT ;
    ANTENNADIFFAREA 0.554400 ;
    PORT
      LAYER li1 ;
        RECT 110.385 143.775 110.685 144.195 ;
        RECT 130.710 143.815 130.985 144.195 ;
        RECT 110.385 141.900 110.685 142.320 ;
        RECT 130.710 141.900 130.985 142.280 ;
      LAYER mcon ;
        RECT 110.475 143.885 110.645 144.055 ;
        RECT 130.770 143.905 130.940 144.075 ;
        RECT 110.475 142.040 110.645 142.210 ;
        RECT 130.770 142.020 130.940 142.190 ;
      LAYER met1 ;
        RECT 110.420 144.115 110.680 144.140 ;
        RECT 130.720 144.135 130.980 144.155 ;
        RECT 110.415 143.825 110.705 144.115 ;
        RECT 130.710 143.865 131.000 144.135 ;
        RECT 130.720 143.835 130.980 143.865 ;
        RECT 110.420 143.820 110.680 143.825 ;
        RECT 110.475 142.270 110.645 143.820 ;
        RECT 110.415 141.980 110.705 142.270 ;
        RECT 130.770 142.250 130.940 143.835 ;
        RECT 130.710 141.960 131.000 142.250 ;
      LAYER via ;
        RECT 110.420 143.850 110.680 144.110 ;
        RECT 130.720 143.865 130.980 144.125 ;
      LAYER met2 ;
        RECT 110.480 152.895 110.650 152.900 ;
        RECT 110.425 152.525 110.705 152.895 ;
        RECT 110.475 144.140 110.655 152.525 ;
        RECT 131.575 152.515 131.855 152.890 ;
        RECT 110.420 143.820 110.680 144.140 ;
        RECT 130.720 144.075 130.980 144.155 ;
        RECT 131.640 144.075 131.810 152.515 ;
        RECT 130.720 143.905 131.810 144.075 ;
        RECT 130.720 143.835 130.980 143.905 ;
        RECT 110.475 142.210 110.655 143.820 ;
        RECT 131.640 142.200 131.810 143.905 ;
        RECT 130.760 142.015 131.810 142.200 ;
      LAYER via2 ;
        RECT 110.425 152.570 110.705 152.850 ;
        RECT 131.575 152.560 131.855 152.840 ;
      LAYER met3 ;
        RECT -0.130 152.430 253.790 152.930 ;
    END
  END th2
  PIN vnb
    DIRECTION INOUT ;
    ANTENNAGATEAREA 0.907200 ;
    PORT
      LAYER li1 ;
        RECT 107.380 171.785 107.550 171.835 ;
        RECT 107.350 171.555 107.580 171.785 ;
        RECT 107.380 171.505 107.550 171.555 ;
        RECT 107.380 166.345 107.550 166.395 ;
        RECT 107.350 166.115 107.580 166.345 ;
        RECT 107.380 166.065 107.550 166.115 ;
        RECT 107.380 160.905 107.550 160.955 ;
        RECT 110.600 160.905 110.770 160.955 ;
        RECT 107.350 160.675 107.580 160.905 ;
        RECT 110.570 160.675 110.800 160.905 ;
        RECT 107.380 160.625 107.550 160.675 ;
        RECT 110.600 160.625 110.770 160.675 ;
      LAYER mcon ;
        RECT 107.380 171.585 107.550 171.755 ;
        RECT 107.380 166.145 107.550 166.315 ;
        RECT 107.380 160.705 107.550 160.875 ;
        RECT 110.600 160.705 110.770 160.875 ;
      LAYER met1 ;
        RECT 107.325 171.505 107.585 171.835 ;
        RECT 107.325 166.065 107.585 166.395 ;
        RECT 107.325 160.890 107.585 160.955 ;
        RECT 110.545 160.890 110.805 160.955 ;
        RECT 107.325 160.700 110.805 160.890 ;
        RECT 107.325 160.625 107.585 160.700 ;
        RECT 110.545 160.625 110.805 160.700 ;
      LAYER via ;
        RECT 107.325 171.540 107.585 171.800 ;
        RECT 107.325 166.100 107.585 166.360 ;
        RECT 107.325 160.660 107.585 160.920 ;
        RECT 110.545 160.660 110.805 160.920 ;
      LAYER met2 ;
        RECT 107.325 171.505 107.585 171.835 ;
        RECT 107.380 166.395 107.555 171.505 ;
        RECT 107.325 166.065 107.585 166.395 ;
        RECT 107.390 160.955 107.540 166.065 ;
        RECT 107.325 160.625 107.585 160.955 ;
        RECT 110.545 160.625 110.805 160.955 ;
        RECT 107.390 158.635 107.540 160.625 ;
        RECT 107.315 158.245 107.615 158.635 ;
      LAYER via2 ;
        RECT 107.315 158.290 107.615 158.590 ;
      LAYER met3 ;
        RECT -0.130 158.200 253.790 158.700 ;
    END
  END vnb
  PIN vpb
    DIRECTION INOUT ;
    ANTENNAGATEAREA 1.360800 ;
    PORT
      LAYER li1 ;
        RECT 110.495 173.470 110.665 173.800 ;
        RECT 110.495 168.030 110.665 168.360 ;
      LAYER mcon ;
        RECT 110.495 173.550 110.665 173.720 ;
        RECT 110.495 168.110 110.665 168.280 ;
      LAYER met1 ;
        RECT 110.405 173.470 110.760 173.760 ;
        RECT 110.405 168.280 110.760 168.320 ;
        RECT 111.510 168.280 111.830 168.325 ;
        RECT 110.405 168.110 111.830 168.280 ;
        RECT 110.405 168.030 110.760 168.110 ;
        RECT 111.510 168.065 111.830 168.110 ;
      LAYER via ;
        RECT 110.450 173.500 110.710 173.760 ;
        RECT 110.450 168.060 110.710 168.320 ;
        RECT 111.540 168.065 111.800 168.325 ;
      LAYER met2 ;
        RECT 110.420 173.500 110.740 173.760 ;
        RECT 110.490 168.320 110.665 173.500 ;
        RECT 110.420 168.060 110.740 168.320 ;
        RECT 111.540 168.035 111.800 168.355 ;
        RECT 111.585 157.615 111.755 168.035 ;
        RECT 111.520 157.225 111.820 157.615 ;
      LAYER via2 ;
        RECT 111.520 157.270 111.820 157.570 ;
      LAYER met3 ;
        RECT -0.130 157.200 253.790 157.700 ;
    END
  END vpb
  PIN inm
    DIRECTION INOUT ;
    ANTENNADIFFAREA 1.696800 ;
    PORT
      LAYER li1 ;
        RECT 3.100 132.010 3.470 132.265 ;
        RECT 5.075 132.225 5.445 132.270 ;
        RECT 234.935 132.225 235.305 132.270 ;
        RECT 5.075 132.055 5.785 132.225 ;
        RECT 5.075 132.005 5.445 132.055 ;
        RECT 3.100 129.340 3.470 129.595 ;
        RECT 5.075 129.545 5.445 129.595 ;
        RECT 5.615 129.545 5.785 132.055 ;
        RECT 5.075 129.375 5.785 129.545 ;
        RECT 234.595 132.055 235.305 132.225 ;
        RECT 234.595 129.545 234.765 132.055 ;
        RECT 234.935 132.005 235.305 132.055 ;
        RECT 236.910 132.010 237.280 132.265 ;
        RECT 234.935 129.545 235.305 129.595 ;
        RECT 234.595 129.375 235.305 129.545 ;
        RECT 5.075 129.340 5.445 129.375 ;
        RECT 234.935 129.340 235.305 129.375 ;
        RECT 236.910 129.340 237.280 129.595 ;
      LAYER mcon ;
        RECT 3.220 132.055 3.390 132.225 ;
        RECT 5.155 132.055 5.325 132.225 ;
        RECT 3.220 129.380 3.390 129.550 ;
        RECT 5.155 129.380 5.325 129.550 ;
        RECT 235.055 132.055 235.225 132.225 ;
        RECT 236.990 132.055 237.160 132.225 ;
        RECT 235.055 129.380 235.225 129.550 ;
        RECT 236.990 129.380 237.160 129.550 ;
      LAYER met1 ;
        RECT 3.140 132.005 3.465 132.270 ;
        RECT 5.075 132.005 5.400 132.270 ;
        RECT 234.980 132.005 235.305 132.270 ;
        RECT 236.915 132.005 237.240 132.270 ;
        RECT 3.140 129.340 3.465 129.600 ;
        RECT 5.080 129.335 5.400 129.595 ;
        RECT 234.980 129.335 235.300 129.595 ;
        RECT 236.915 129.340 237.240 129.600 ;
        RECT 5.185 129.320 5.325 129.335 ;
        RECT 235.055 129.320 235.195 129.335 ;
      LAYER via ;
        RECT 3.170 132.005 3.435 132.270 ;
        RECT 5.110 132.005 5.370 132.270 ;
        RECT 235.010 132.005 235.270 132.270 ;
        RECT 236.945 132.005 237.210 132.270 ;
        RECT 3.170 129.340 3.430 129.600 ;
        RECT 5.110 129.335 5.370 129.595 ;
        RECT 235.010 129.335 235.270 129.595 ;
        RECT 236.950 129.340 237.210 129.600 ;
      LAYER met2 ;
        RECT 3.140 132.225 3.465 132.270 ;
        RECT 5.075 132.225 5.400 132.270 ;
        RECT 3.140 132.055 5.400 132.225 ;
        RECT 3.140 132.005 3.465 132.055 ;
        RECT 5.075 132.005 5.400 132.055 ;
        RECT 234.980 132.225 235.305 132.270 ;
        RECT 236.915 132.225 237.240 132.270 ;
        RECT 234.980 132.055 237.240 132.225 ;
        RECT 234.980 132.005 235.305 132.055 ;
        RECT 236.915 132.005 237.240 132.055 ;
        RECT 3.140 129.550 3.460 129.600 ;
        RECT 5.055 129.550 5.425 129.605 ;
        RECT 3.140 129.380 5.425 129.550 ;
        RECT 3.140 129.340 3.460 129.380 ;
        RECT 5.055 129.325 5.425 129.380 ;
        RECT 234.955 129.550 235.325 129.605 ;
        RECT 236.920 129.550 237.240 129.600 ;
        RECT 234.955 129.380 237.240 129.550 ;
        RECT 234.955 129.325 235.325 129.380 ;
        RECT 236.920 129.340 237.240 129.380 ;
      LAYER via2 ;
        RECT 5.100 129.325 5.380 129.605 ;
        RECT 235.000 129.325 235.280 129.605 ;
      LAYER met3 ;
        RECT 4.995 129.235 5.485 129.725 ;
        RECT 234.895 129.235 235.385 129.725 ;
        RECT 5.340 4.805 6.385 10.525 ;
        RECT 233.995 4.805 235.040 10.525 ;
      LAYER via3 ;
        RECT 5.080 129.305 5.400 129.625 ;
        RECT 234.980 129.305 235.300 129.625 ;
        RECT 5.370 9.550 6.355 10.495 ;
        RECT 5.370 4.825 6.355 5.770 ;
        RECT 234.025 9.550 235.010 10.495 ;
        RECT 234.025 4.825 235.010 5.770 ;
      LAYER met4 ;
        RECT 4.995 129.235 6.360 129.700 ;
        RECT 5.365 9.545 6.360 129.235 ;
        RECT 234.020 129.235 235.385 129.700 ;
        RECT 234.020 9.545 235.015 129.235 ;
        RECT -0.130 4.805 253.790 5.800 ;
    END
  END inm
  PIN inp
    DIRECTION INOUT ;
    ANTENNADIFFAREA 0.730800 ;
    PORT
      LAYER li1 ;
        RECT 3.100 130.675 3.470 130.930 ;
        RECT 5.075 130.670 5.445 130.935 ;
        RECT 234.935 130.670 235.305 130.935 ;
        RECT 236.910 130.675 237.280 130.930 ;
      LAYER mcon ;
        RECT 3.220 130.715 3.390 130.890 ;
        RECT 5.155 130.715 5.325 130.890 ;
        RECT 235.055 130.715 235.225 130.890 ;
        RECT 236.990 130.715 237.160 130.890 ;
      LAYER met1 ;
        RECT 3.140 130.670 3.465 130.935 ;
        RECT 5.075 130.670 5.400 130.935 ;
        RECT 234.980 130.670 235.305 130.935 ;
        RECT 236.915 130.670 237.240 130.935 ;
      LAYER via ;
        RECT 3.170 130.670 3.435 130.935 ;
        RECT 5.110 130.670 5.370 130.935 ;
        RECT 235.010 130.670 235.270 130.935 ;
        RECT 236.945 130.670 237.210 130.935 ;
      LAYER met2 ;
        RECT 3.115 130.890 3.485 130.940 ;
        RECT 4.385 130.890 4.705 130.930 ;
        RECT 5.075 130.890 5.400 130.935 ;
        RECT 3.115 130.715 5.400 130.890 ;
        RECT 3.115 130.660 3.485 130.715 ;
        RECT 4.385 130.670 4.705 130.715 ;
        RECT 5.075 130.670 5.400 130.715 ;
        RECT 234.980 130.890 235.305 130.935 ;
        RECT 235.675 130.890 235.995 130.930 ;
        RECT 236.895 130.890 237.265 130.940 ;
        RECT 234.980 130.715 237.265 130.890 ;
        RECT 234.980 130.670 235.305 130.715 ;
        RECT 235.675 130.670 235.995 130.715 ;
        RECT 236.895 130.660 237.265 130.715 ;
      LAYER via2 ;
        RECT 3.160 130.660 3.440 130.940 ;
        RECT 236.940 130.660 237.220 130.940 ;
      LAYER met3 ;
        RECT 3.055 130.565 3.545 131.055 ;
        RECT 236.835 130.565 237.325 131.055 ;
        RECT 2.135 1.600 3.180 10.525 ;
        RECT 237.200 1.600 238.245 10.525 ;
      LAYER via3 ;
        RECT 3.140 130.640 3.460 130.960 ;
        RECT 236.920 130.640 237.240 130.960 ;
        RECT 2.165 9.550 3.150 10.495 ;
        RECT 2.165 1.620 3.150 2.565 ;
        RECT 237.230 9.550 238.215 10.495 ;
        RECT 237.230 1.620 238.215 2.565 ;
      LAYER met4 ;
        RECT 2.160 130.630 3.475 130.995 ;
        RECT 236.905 130.630 238.220 130.995 ;
        RECT 2.160 9.545 3.155 130.630 ;
        RECT 237.225 9.545 238.220 130.630 ;
        RECT -0.130 2.595 5.370 2.605 ;
        RECT -0.130 1.600 253.790 2.595 ;
    END
  END inp
  PIN cclk
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.302400 ;
    ANTENNADIFFAREA 0.493500 ;
    PORT
      LAYER li1 ;
        RECT 93.260 164.945 93.590 165.115 ;
        RECT 94.270 163.415 94.540 163.440 ;
        RECT 94.270 163.060 94.820 163.415 ;
        RECT 94.425 162.205 94.595 163.060 ;
        RECT 94.250 162.195 94.595 162.205 ;
        RECT 94.205 162.035 94.595 162.195 ;
        RECT 94.205 161.590 94.575 162.035 ;
        RECT 94.205 161.550 94.570 161.590 ;
      LAYER mcon ;
        RECT 93.340 164.945 93.510 165.115 ;
        RECT 94.320 163.150 94.740 163.320 ;
      LAYER met1 ;
        RECT 93.275 165.160 93.590 165.165 ;
        RECT 67.560 165.115 67.880 165.160 ;
        RECT 67.560 165.110 68.730 165.115 ;
        RECT 93.265 165.110 93.590 165.160 ;
        RECT 67.560 164.945 93.590 165.110 ;
        RECT 67.560 164.900 67.880 164.945 ;
        RECT 68.730 164.940 93.590 164.945 ;
        RECT 93.265 164.900 93.590 164.940 ;
        RECT 93.275 164.895 93.590 164.900 ;
        RECT 94.260 163.105 94.800 163.365 ;
      LAYER via ;
        RECT 67.590 164.900 67.850 165.160 ;
        RECT 93.295 164.900 93.555 165.160 ;
        RECT 94.320 163.105 94.740 163.365 ;
      LAYER met2 ;
        RECT 67.580 164.895 67.860 185.700 ;
        RECT 93.265 164.900 93.585 165.160 ;
        RECT 67.590 164.870 67.850 164.895 ;
        RECT 93.340 163.320 93.510 164.900 ;
        RECT 94.290 163.320 94.770 163.365 ;
        RECT 93.340 163.150 94.770 163.320 ;
        RECT 94.290 163.105 94.770 163.150 ;
    END
  END cclk
  PIN fb1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.302400 ;
    ANTENNADIFFAREA 0.493500 ;
    PORT
      LAYER li1 ;
        RECT 45.310 171.610 45.675 171.650 ;
        RECT 45.310 171.165 45.680 171.610 ;
        RECT 45.310 171.005 45.700 171.165 ;
        RECT 45.355 170.995 45.700 171.005 ;
        RECT 45.530 170.140 45.700 170.995 ;
        RECT 45.375 169.785 45.925 170.140 ;
        RECT 45.375 169.760 45.645 169.785 ;
        RECT 44.365 168.085 44.695 168.255 ;
      LAYER mcon ;
        RECT 45.425 169.880 45.845 170.050 ;
        RECT 44.445 168.085 44.615 168.255 ;
      LAYER met1 ;
        RECT 25.230 175.655 25.550 175.700 ;
        RECT 44.370 175.655 44.690 175.700 ;
        RECT 25.230 175.485 44.690 175.655 ;
        RECT 25.230 175.440 25.550 175.485 ;
        RECT 44.370 175.440 44.690 175.485 ;
        RECT 45.365 169.835 45.905 170.095 ;
        RECT 44.380 168.300 44.695 168.305 ;
        RECT 44.370 168.040 44.695 168.300 ;
        RECT 44.380 168.035 44.695 168.040 ;
      LAYER via ;
        RECT 25.260 175.440 25.520 175.700 ;
        RECT 44.400 175.440 44.660 175.700 ;
        RECT 45.425 169.835 45.845 170.095 ;
        RECT 44.400 168.040 44.660 168.300 ;
      LAYER met2 ;
        RECT 25.260 175.410 25.540 185.700 ;
        RECT 44.400 175.410 44.660 175.730 ;
        RECT 44.445 170.050 44.615 175.410 ;
        RECT 45.395 170.050 45.875 170.095 ;
        RECT 44.445 169.880 45.875 170.050 ;
        RECT 44.445 168.300 44.615 169.880 ;
        RECT 45.395 169.835 45.875 169.880 ;
        RECT 44.370 168.040 44.690 168.300 ;
    END
  END fb1
  PIN div2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.302400 ;
    ANTENNADIFFAREA 0.493500 ;
    PORT
      LAYER li1 ;
        RECT 94.205 171.490 94.570 171.530 ;
        RECT 94.205 171.045 94.575 171.490 ;
        RECT 94.205 170.885 94.595 171.045 ;
        RECT 94.250 170.875 94.595 170.885 ;
        RECT 94.425 170.020 94.595 170.875 ;
        RECT 94.270 169.665 94.820 170.020 ;
        RECT 94.270 169.640 94.540 169.665 ;
        RECT 93.260 167.965 93.590 168.135 ;
      LAYER mcon ;
        RECT 94.320 169.760 94.740 169.930 ;
        RECT 93.340 167.965 93.510 168.135 ;
      LAYER met1 ;
        RECT 94.350 177.305 94.670 177.380 ;
        RECT 109.880 177.305 110.200 177.350 ;
        RECT 94.350 177.135 110.200 177.305 ;
        RECT 94.350 177.060 94.670 177.135 ;
        RECT 109.880 177.090 110.200 177.135 ;
        RECT 94.260 169.715 94.800 169.975 ;
        RECT 93.270 168.180 93.590 168.195 ;
        RECT 93.265 167.920 93.590 168.180 ;
        RECT 93.270 167.905 93.590 167.920 ;
      LAYER via ;
        RECT 94.380 177.090 94.640 177.350 ;
        RECT 109.910 177.090 110.170 177.350 ;
        RECT 94.320 169.715 94.740 169.975 ;
        RECT 93.295 167.920 93.555 168.180 ;
      LAYER met2 ;
        RECT 94.350 177.060 94.670 177.380 ;
        RECT 109.900 177.080 110.180 185.700 ;
        RECT 109.910 177.060 110.170 177.080 ;
        RECT 94.425 169.975 94.595 177.060 ;
        RECT 94.290 169.930 94.770 169.975 ;
        RECT 93.340 169.760 94.770 169.930 ;
        RECT 93.340 168.180 93.510 169.760 ;
        RECT 94.290 169.715 94.770 169.760 ;
        RECT 93.265 167.920 93.585 168.180 ;
    END
  END div2
  PIN high_buf
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.310800 ;
    PORT
      LAYER li1 ;
        RECT 111.390 132.915 111.720 133.295 ;
        RECT 111.400 131.065 111.730 131.445 ;
      LAYER mcon ;
        RECT 111.470 132.965 111.640 133.255 ;
        RECT 111.480 131.115 111.650 131.405 ;
      LAYER met1 ;
        RECT 119.390 138.075 119.710 138.120 ;
        RECT 111.420 137.905 119.710 138.075 ;
        RECT 111.420 133.295 111.590 137.905 ;
        RECT 119.390 137.860 119.710 137.905 ;
        RECT 111.410 132.915 111.700 133.295 ;
        RECT 111.420 131.445 111.590 132.915 ;
        RECT 111.420 131.065 111.710 131.445 ;
      LAYER via ;
        RECT 119.420 137.860 119.680 138.120 ;
      LAYER met2 ;
        RECT 152.220 177.450 152.500 185.700 ;
        RECT 152.145 177.020 152.555 177.450 ;
        RECT 152.170 177.000 152.530 177.020 ;
        RECT 119.420 138.115 119.680 138.150 ;
        RECT 119.325 137.835 119.695 138.115 ;
        RECT 119.420 137.830 119.680 137.835 ;
      LAYER via2 ;
        RECT 152.170 177.045 152.530 177.405 ;
        RECT 119.370 137.835 119.650 138.115 ;
      LAYER met3 ;
        RECT 119.330 177.425 152.555 177.430 ;
        RECT 119.305 177.025 152.555 177.425 ;
        RECT 119.330 177.020 152.555 177.025 ;
        RECT 119.270 137.720 119.770 138.210 ;
      LAYER via3 ;
        RECT 119.335 177.025 119.735 177.425 ;
        RECT 119.355 137.800 119.720 138.165 ;
      LAYER met4 ;
        RECT 119.330 163.695 119.740 177.430 ;
        RECT 119.350 137.795 119.725 163.695 ;
    END
  END high_buf
  PIN phi1b_dig
    DIRECTION OUTPUT ;
    ANTENNAGATEAREA 1.680000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 127.935 166.795 128.265 167.255 ;
        RECT 128.775 166.795 129.105 167.255 ;
        RECT 129.615 166.795 129.945 167.255 ;
        RECT 130.455 166.795 130.785 167.255 ;
        RECT 127.340 166.605 131.310 166.795 ;
        RECT 127.340 166.015 127.685 166.605 ;
        RECT 130.990 166.015 131.310 166.605 ;
        RECT 127.340 165.845 131.310 166.015 ;
        RECT 127.935 165.045 128.265 165.845 ;
        RECT 128.775 165.045 129.105 165.845 ;
        RECT 129.615 165.045 129.945 165.845 ;
        RECT 130.455 165.045 130.785 165.845 ;
        RECT 116.510 132.680 116.680 133.315 ;
        RECT 123.760 132.680 123.930 133.315 ;
      LAYER mcon ;
        RECT 131.085 166.235 131.255 166.405 ;
        RECT 116.510 132.760 116.680 133.235 ;
        RECT 123.760 132.760 123.930 133.235 ;
      LAYER met1 ;
        RECT 131.900 166.485 132.280 166.515 ;
        RECT 130.920 166.165 132.280 166.485 ;
        RECT 131.900 166.135 132.280 166.165 ;
        RECT 116.510 133.265 116.680 133.295 ;
        RECT 123.760 133.265 123.930 133.295 ;
        RECT 116.480 133.175 116.710 133.265 ;
        RECT 123.730 133.175 123.960 133.265 ;
        RECT 116.465 133.085 116.725 133.175 ;
        RECT 123.715 133.085 123.975 133.175 ;
        RECT 116.400 132.945 116.735 133.085 ;
        RECT 123.705 132.945 124.040 133.085 ;
        RECT 116.465 132.855 116.725 132.945 ;
        RECT 123.715 132.855 123.975 132.945 ;
        RECT 116.480 132.730 116.710 132.855 ;
        RECT 123.730 132.730 123.960 132.855 ;
        RECT 116.510 132.700 116.680 132.730 ;
        RECT 123.760 132.700 123.930 132.730 ;
      LAYER via ;
        RECT 131.930 166.165 132.250 166.485 ;
        RECT 116.465 132.885 116.725 133.145 ;
        RECT 123.715 132.885 123.975 133.145 ;
      LAYER met2 ;
        RECT 131.900 166.135 132.280 166.515 ;
        RECT 131.930 160.210 132.250 166.135 ;
        RECT 169.690 160.595 170.010 177.340 ;
        RECT 194.540 177.330 194.820 185.700 ;
        RECT 194.530 176.940 194.830 177.330 ;
        RECT 169.670 160.240 170.030 160.595 ;
        RECT 116.455 132.835 116.735 133.205 ;
        RECT 123.705 132.830 123.985 133.200 ;
      LAYER via2 ;
        RECT 169.690 176.975 170.010 177.295 ;
        RECT 194.530 176.985 194.830 177.285 ;
        RECT 131.930 160.255 132.250 160.575 ;
        RECT 169.710 160.285 169.990 160.565 ;
        RECT 116.455 132.880 116.735 133.160 ;
        RECT 123.705 132.875 123.985 133.155 ;
      LAYER met3 ;
        RECT 169.665 177.295 170.035 177.320 ;
        RECT 194.505 177.295 194.855 177.310 ;
        RECT 169.665 176.975 194.855 177.295 ;
        RECT 169.665 176.950 170.035 176.975 ;
        RECT 194.505 176.960 194.855 176.975 ;
        RECT 131.905 160.585 132.275 160.600 ;
        RECT 169.685 160.585 170.015 160.590 ;
        RECT 123.655 160.265 170.015 160.585 ;
        RECT 131.905 160.230 132.275 160.265 ;
        RECT 169.685 160.260 170.015 160.265 ;
        RECT 116.390 133.165 116.775 133.210 ;
        RECT 123.650 133.165 124.035 133.210 ;
        RECT 116.390 132.865 124.035 133.165 ;
        RECT 116.390 132.830 116.775 132.865 ;
        RECT 123.650 132.830 124.035 132.865 ;
      LAYER via3 ;
        RECT 123.685 160.265 124.005 160.585 ;
        RECT 116.420 132.855 116.745 133.185 ;
        RECT 123.685 132.860 124.005 133.180 ;
      LAYER met4 ;
        RECT 123.680 160.260 124.010 160.590 ;
        RECT 116.420 133.210 116.745 133.845 ;
        RECT 123.685 133.210 124.005 160.260 ;
        RECT 116.390 132.830 116.775 133.210 ;
        RECT 123.650 132.830 124.035 133.210 ;
    END
  END phi1b_dig
  PIN lo
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.302400 ;
    ANTENNADIFFAREA 0.493500 ;
    PORT
      LAYER li1 ;
        RECT 195.845 171.610 196.210 171.650 ;
        RECT 195.840 171.165 196.210 171.610 ;
        RECT 195.820 171.005 196.210 171.165 ;
        RECT 195.820 170.995 196.165 171.005 ;
        RECT 195.820 170.140 195.990 170.995 ;
        RECT 195.595 169.785 196.145 170.140 ;
        RECT 195.875 169.760 196.145 169.785 ;
        RECT 196.825 168.085 197.155 168.255 ;
      LAYER mcon ;
        RECT 195.675 169.880 196.095 170.050 ;
        RECT 196.905 168.085 197.075 168.255 ;
      LAYER met1 ;
        RECT 195.615 169.835 196.155 170.095 ;
        RECT 196.825 168.300 197.140 168.305 ;
        RECT 196.825 168.040 197.150 168.300 ;
        RECT 196.825 168.035 197.140 168.040 ;
      LAYER via ;
        RECT 195.675 169.835 196.095 170.095 ;
        RECT 196.860 168.040 197.120 168.300 ;
      LAYER met2 ;
        RECT 196.840 174.580 197.140 174.970 ;
        RECT 236.860 174.960 237.140 185.700 ;
        RECT 236.840 174.625 237.140 174.960 ;
        RECT 236.850 174.590 237.130 174.625 ;
        RECT 195.645 170.050 196.125 170.095 ;
        RECT 196.905 170.050 197.075 174.580 ;
        RECT 195.645 169.880 197.075 170.050 ;
        RECT 195.645 169.835 196.125 169.880 ;
        RECT 196.905 168.300 197.075 169.880 ;
        RECT 196.830 168.040 197.150 168.300 ;
      LAYER via2 ;
        RECT 196.840 174.625 197.140 174.925 ;
        RECT 236.850 174.635 237.130 174.915 ;
      LAYER met3 ;
        RECT 196.815 174.925 197.165 174.950 ;
        RECT 236.825 174.925 237.155 174.940 ;
        RECT 196.815 174.625 237.155 174.925 ;
        RECT 196.815 174.600 197.165 174.625 ;
        RECT 236.825 174.610 237.155 174.625 ;
    END
  END lo
  PIN vdda
    DIRECTION INOUT ;
    ANTENNAGATEAREA 0.226800 ;
    ANTENNADIFFAREA 27.605099 ;
    PORT
      LAYER nwell ;
        RECT 107.305 175.455 108.955 175.460 ;
        RECT 111.335 175.455 117.440 175.530 ;
        RECT 107.305 175.145 117.440 175.455 ;
        RECT 105.710 174.465 117.440 175.145 ;
        RECT 105.710 174.460 112.260 174.465 ;
        RECT 105.710 173.770 111.380 174.460 ;
        RECT 105.710 173.505 108.955 173.770 ;
        RECT 105.710 173.495 107.470 173.505 ;
        RECT 50.335 170.445 52.385 171.605 ;
        RECT 99.230 170.325 101.280 171.485 ;
        RECT 107.385 170.015 109.035 170.030 ;
        RECT 111.335 170.025 117.460 171.630 ;
        RECT 111.335 170.015 117.440 170.025 ;
        RECT 107.385 169.930 117.440 170.015 ;
        RECT 106.500 169.705 117.440 169.930 ;
        RECT 105.710 169.025 117.440 169.705 ;
        RECT 105.710 169.020 112.260 169.025 ;
        RECT 105.710 168.330 111.380 169.020 ;
        RECT 121.275 168.815 125.795 170.900 ;
        RECT 189.135 170.445 191.185 171.605 ;
        RECT 105.710 168.075 109.035 168.330 ;
        RECT 105.710 168.055 107.470 168.075 ;
        RECT 111.905 165.120 117.440 166.185 ;
        RECT 99.230 161.595 101.280 162.755 ;
        RECT 105.710 162.615 107.470 164.265 ;
        RECT 108.930 162.615 110.690 164.265 ;
        RECT 112.150 163.585 117.440 165.120 ;
        RECT 121.275 164.120 125.795 166.205 ;
        RECT 111.905 159.680 117.440 160.745 ;
        RECT 109.100 143.590 111.510 144.435 ;
        RECT 128.870 143.590 131.280 144.435 ;
        RECT 2.860 129.000 3.700 133.050 ;
        RECT 8.675 130.190 10.070 131.030 ;
        RECT 18.520 130.190 19.915 131.030 ;
        RECT 29.975 130.190 31.370 131.030 ;
        RECT 36.370 130.190 37.765 131.030 ;
        RECT 67.425 130.190 68.820 131.030 ;
        RECT 75.060 130.190 76.455 131.030 ;
        RECT 98.475 130.190 99.870 131.030 ;
        RECT 105.820 130.190 107.215 131.030 ;
        RECT 133.165 130.190 134.560 131.030 ;
        RECT 140.510 130.190 141.905 131.030 ;
        RECT 163.925 130.190 165.320 131.030 ;
        RECT 171.560 130.190 172.955 131.030 ;
        RECT 202.615 130.190 204.010 131.030 ;
        RECT 209.010 130.190 210.405 131.030 ;
        RECT 220.465 130.190 221.860 131.030 ;
        RECT 230.310 130.190 231.705 131.030 ;
        RECT 236.680 129.000 237.520 133.050 ;
      LAYER li1 ;
        RECT 105.350 175.680 117.770 175.850 ;
        RECT 105.990 174.890 106.540 175.680 ;
        RECT 109.500 175.225 109.770 175.680 ;
        RECT 112.430 175.315 112.980 175.680 ;
        RECT 112.430 175.275 113.120 175.315 ;
        RECT 113.990 175.310 114.170 175.680 ;
        RECT 115.190 175.315 115.740 175.680 ;
        RECT 105.970 173.700 106.680 174.890 ;
        RECT 109.030 173.960 109.820 175.225 ;
        RECT 112.410 174.670 113.120 175.275 ;
        RECT 113.915 175.270 114.280 175.310 ;
        RECT 115.190 175.275 115.880 175.315 ;
        RECT 116.750 175.310 116.930 175.680 ;
        RECT 112.795 174.660 113.085 174.670 ;
        RECT 113.915 174.665 114.285 175.270 ;
        RECT 115.170 174.670 115.880 175.275 ;
        RECT 116.675 175.270 117.040 175.310 ;
        RECT 113.960 174.655 114.250 174.665 ;
        RECT 115.555 174.660 115.845 174.670 ;
        RECT 116.675 174.665 117.045 175.270 ;
        RECT 116.720 174.655 117.010 174.665 ;
        RECT 109.140 173.945 109.310 173.960 ;
        RECT 109.595 173.940 109.765 173.960 ;
        RECT 106.355 173.690 106.645 173.700 ;
        RECT 49.290 172.015 55.730 172.185 ;
        RECT 98.185 171.895 104.625 172.065 ;
        RECT 113.950 171.785 114.120 172.115 ;
        RECT 185.790 172.015 192.230 172.185 ;
        RECT 51.145 170.855 51.315 171.185 ;
        RECT 51.975 170.855 52.145 171.185 ;
        RECT 100.040 170.735 100.210 171.065 ;
        RECT 100.870 170.735 101.040 171.065 ;
        RECT 112.080 170.825 112.455 171.445 ;
        RECT 115.555 171.420 115.845 171.430 ;
        RECT 116.720 171.425 117.010 171.435 ;
        RECT 112.175 170.410 112.345 170.825 ;
        RECT 115.170 170.815 115.880 171.420 ;
        RECT 115.190 170.775 115.880 170.815 ;
        RECT 116.675 170.820 117.045 171.425 ;
        RECT 189.375 170.855 189.545 171.185 ;
        RECT 190.205 170.855 190.375 171.185 ;
        RECT 116.675 170.780 117.040 170.820 ;
        RECT 115.190 170.410 115.740 170.775 ;
        RECT 116.750 170.410 116.930 170.780 ;
        RECT 105.350 170.240 117.770 170.410 ;
        RECT 123.445 170.315 123.830 170.665 ;
        RECT 47.685 169.520 47.855 169.850 ;
        RECT 48.550 169.520 48.720 169.850 ;
        RECT 49.415 169.520 49.585 169.850 ;
        RECT 50.280 169.520 50.450 169.850 ;
        RECT 51.145 169.520 51.315 169.850 ;
        RECT 52.010 169.520 52.180 169.850 ;
        RECT 52.875 169.520 53.045 169.850 ;
        RECT 53.740 169.520 53.910 169.850 ;
        RECT 54.605 169.520 54.775 169.850 ;
        RECT 96.580 169.400 96.750 169.730 ;
        RECT 97.445 169.400 97.615 169.730 ;
        RECT 98.310 169.400 98.480 169.730 ;
        RECT 99.175 169.400 99.345 169.730 ;
        RECT 100.040 169.400 100.210 169.730 ;
        RECT 100.905 169.400 101.075 169.730 ;
        RECT 101.770 169.400 101.940 169.730 ;
        RECT 102.635 169.400 102.805 169.730 ;
        RECT 103.500 169.400 103.670 169.730 ;
        RECT 105.990 169.450 106.540 170.240 ;
        RECT 109.500 169.785 109.770 170.240 ;
        RECT 112.430 169.875 112.980 170.240 ;
        RECT 112.430 169.835 113.120 169.875 ;
        RECT 113.990 169.870 114.170 170.240 ;
        RECT 115.190 169.875 115.740 170.240 ;
        RECT 105.970 168.260 106.680 169.450 ;
        RECT 109.030 168.520 109.820 169.785 ;
        RECT 112.410 169.230 113.120 169.835 ;
        RECT 113.915 169.830 114.280 169.870 ;
        RECT 115.190 169.835 115.880 169.875 ;
        RECT 116.750 169.870 116.930 170.240 ;
        RECT 121.465 170.145 125.605 170.315 ;
        RECT 112.795 169.220 113.085 169.230 ;
        RECT 113.915 169.225 114.285 169.830 ;
        RECT 115.170 169.230 115.880 169.835 ;
        RECT 116.675 169.830 117.040 169.870 ;
        RECT 113.960 169.215 114.250 169.225 ;
        RECT 115.555 169.220 115.845 169.230 ;
        RECT 116.675 169.225 117.045 169.830 ;
        RECT 121.720 169.345 121.975 170.145 ;
        RECT 122.645 169.345 122.815 170.145 ;
        RECT 123.485 169.345 123.655 170.145 ;
        RECT 124.325 169.345 124.495 170.145 ;
        RECT 125.165 169.345 125.465 170.145 ;
        RECT 186.745 169.520 186.915 169.850 ;
        RECT 187.610 169.520 187.780 169.850 ;
        RECT 188.475 169.520 188.645 169.850 ;
        RECT 189.340 169.520 189.510 169.850 ;
        RECT 190.205 169.520 190.375 169.850 ;
        RECT 191.070 169.520 191.240 169.850 ;
        RECT 191.935 169.520 192.105 169.850 ;
        RECT 192.800 169.520 192.970 169.850 ;
        RECT 193.665 169.520 193.835 169.850 ;
        RECT 116.720 169.215 117.010 169.225 ;
        RECT 109.140 168.505 109.310 168.520 ;
        RECT 109.595 168.500 109.765 168.520 ;
        RECT 106.355 168.250 106.645 168.260 ;
        RECT 113.950 166.345 114.120 166.675 ;
        RECT 112.080 165.385 112.455 166.005 ;
        RECT 115.555 165.980 115.845 165.990 ;
        RECT 116.720 165.985 117.010 165.995 ;
        RECT 112.175 164.970 112.345 165.385 ;
        RECT 115.170 165.375 115.880 165.980 ;
        RECT 115.190 165.335 115.880 165.375 ;
        RECT 116.675 165.380 117.045 165.985 ;
        RECT 116.675 165.340 117.040 165.380 ;
        RECT 115.190 164.970 115.740 165.335 ;
        RECT 116.750 164.970 116.930 165.340 ;
        RECT 105.350 164.800 117.770 164.970 ;
        RECT 121.720 164.875 121.975 165.675 ;
        RECT 122.645 164.875 122.815 165.675 ;
        RECT 123.485 164.875 123.655 165.675 ;
        RECT 124.325 164.875 124.495 165.675 ;
        RECT 125.165 164.875 125.465 165.675 ;
        RECT 105.990 164.010 106.540 164.800 ;
        RECT 109.210 164.010 109.760 164.800 ;
        RECT 112.430 164.435 112.980 164.800 ;
        RECT 112.430 164.395 113.120 164.435 ;
        RECT 113.990 164.430 114.170 164.800 ;
        RECT 115.190 164.435 115.740 164.800 ;
        RECT 96.580 163.350 96.750 163.680 ;
        RECT 97.445 163.350 97.615 163.680 ;
        RECT 98.310 163.350 98.480 163.680 ;
        RECT 99.175 163.350 99.345 163.680 ;
        RECT 100.040 163.350 100.210 163.680 ;
        RECT 100.905 163.350 101.075 163.680 ;
        RECT 101.770 163.350 101.940 163.680 ;
        RECT 102.635 163.350 102.805 163.680 ;
        RECT 103.500 163.350 103.670 163.680 ;
        RECT 105.970 162.820 106.680 164.010 ;
        RECT 109.190 162.820 109.900 164.010 ;
        RECT 112.410 163.790 113.120 164.395 ;
        RECT 113.915 164.390 114.280 164.430 ;
        RECT 115.190 164.395 115.880 164.435 ;
        RECT 116.750 164.430 116.930 164.800 ;
        RECT 121.465 164.705 125.605 164.875 ;
        RECT 112.795 163.780 113.085 163.790 ;
        RECT 113.915 163.785 114.285 164.390 ;
        RECT 115.170 163.790 115.880 164.395 ;
        RECT 116.675 164.390 117.040 164.430 ;
        RECT 113.960 163.775 114.250 163.785 ;
        RECT 115.555 163.780 115.845 163.790 ;
        RECT 116.675 163.785 117.045 164.390 ;
        RECT 123.445 164.355 123.830 164.705 ;
        RECT 116.720 163.775 117.010 163.785 ;
        RECT 106.355 162.810 106.645 162.820 ;
        RECT 109.575 162.810 109.865 162.820 ;
        RECT 100.040 162.015 100.210 162.345 ;
        RECT 100.870 162.015 101.040 162.345 ;
        RECT 98.185 161.015 104.625 161.185 ;
        RECT 113.950 160.905 114.120 161.235 ;
        RECT 112.080 159.945 112.455 160.565 ;
        RECT 115.555 160.540 115.845 160.550 ;
        RECT 116.720 160.545 117.010 160.555 ;
        RECT 112.175 159.530 112.345 159.945 ;
        RECT 115.170 159.935 115.880 160.540 ;
        RECT 115.190 159.895 115.880 159.935 ;
        RECT 116.675 159.940 117.045 160.545 ;
        RECT 116.675 159.900 117.040 159.940 ;
        RECT 115.190 159.530 115.740 159.895 ;
        RECT 116.750 159.530 116.930 159.900 ;
        RECT 105.350 159.360 117.770 159.530 ;
        RECT 111.090 143.820 111.260 147.235 ;
        RECT 129.120 143.820 129.290 147.235 ;
        RECT 3.145 132.615 3.475 132.785 ;
        RECT 236.905 132.615 237.235 132.785 ;
        RECT 9.715 131.100 10.195 131.270 ;
        RECT 18.395 131.100 18.875 131.270 ;
        RECT 9.715 130.415 9.885 131.100 ;
        RECT 18.705 130.415 18.875 131.100 ;
        RECT 31.015 131.100 31.495 131.270 ;
        RECT 36.245 131.100 36.725 131.270 ;
        RECT 31.015 130.415 31.185 131.100 ;
        RECT 36.555 130.415 36.725 131.100 ;
        RECT 68.465 131.100 68.945 131.270 ;
        RECT 74.935 131.100 75.415 131.270 ;
        RECT 68.465 130.415 68.635 131.100 ;
        RECT 75.245 130.415 75.415 131.100 ;
        RECT 99.515 131.100 99.995 131.270 ;
        RECT 105.695 131.100 106.175 131.270 ;
        RECT 99.515 130.415 99.685 131.100 ;
        RECT 106.005 130.415 106.175 131.100 ;
        RECT 134.205 131.100 134.685 131.270 ;
        RECT 140.385 131.100 140.865 131.270 ;
        RECT 134.205 130.415 134.375 131.100 ;
        RECT 140.695 130.415 140.865 131.100 ;
        RECT 164.965 131.100 165.445 131.270 ;
        RECT 171.435 131.100 171.915 131.270 ;
        RECT 164.965 130.415 165.135 131.100 ;
        RECT 171.745 130.415 171.915 131.100 ;
        RECT 203.655 131.100 204.135 131.270 ;
        RECT 208.885 131.100 209.365 131.270 ;
        RECT 203.655 130.415 203.825 131.100 ;
        RECT 209.195 130.415 209.365 131.100 ;
        RECT 221.505 131.100 221.985 131.270 ;
        RECT 230.185 131.100 230.665 131.270 ;
        RECT 221.505 130.415 221.675 131.100 ;
        RECT 230.495 130.415 230.665 131.100 ;
      LAYER mcon ;
        RECT 105.495 175.680 105.665 175.850 ;
        RECT 105.955 175.680 106.125 175.850 ;
        RECT 106.415 175.680 106.585 175.850 ;
        RECT 106.875 175.680 107.045 175.850 ;
        RECT 107.335 175.680 107.505 175.850 ;
        RECT 107.795 175.680 107.965 175.850 ;
        RECT 108.255 175.680 108.425 175.850 ;
        RECT 108.715 175.680 108.885 175.850 ;
        RECT 109.175 175.680 109.345 175.850 ;
        RECT 109.635 175.680 109.805 175.850 ;
        RECT 110.095 175.680 110.265 175.850 ;
        RECT 110.555 175.680 110.725 175.850 ;
        RECT 111.015 175.680 111.185 175.850 ;
        RECT 111.475 175.680 111.645 175.850 ;
        RECT 111.935 175.680 112.105 175.850 ;
        RECT 112.395 175.680 112.565 175.850 ;
        RECT 112.855 175.680 113.025 175.850 ;
        RECT 113.315 175.680 113.485 175.850 ;
        RECT 113.775 175.680 113.945 175.850 ;
        RECT 114.235 175.680 114.405 175.850 ;
        RECT 114.695 175.680 114.865 175.850 ;
        RECT 115.155 175.680 115.325 175.850 ;
        RECT 115.615 175.680 115.785 175.850 ;
        RECT 116.075 175.680 116.245 175.850 ;
        RECT 116.535 175.680 116.705 175.850 ;
        RECT 116.995 175.680 117.165 175.850 ;
        RECT 117.455 175.680 117.625 175.850 ;
        RECT 49.435 172.015 49.605 172.185 ;
        RECT 49.895 172.015 50.065 172.185 ;
        RECT 50.355 172.015 50.525 172.185 ;
        RECT 50.815 172.015 50.985 172.185 ;
        RECT 51.275 172.015 51.445 172.185 ;
        RECT 51.735 172.015 51.905 172.185 ;
        RECT 52.195 172.015 52.365 172.185 ;
        RECT 52.655 172.015 52.825 172.185 ;
        RECT 53.115 172.015 53.285 172.185 ;
        RECT 53.575 172.015 53.745 172.185 ;
        RECT 54.035 172.015 54.205 172.185 ;
        RECT 54.495 172.015 54.665 172.185 ;
        RECT 54.955 172.015 55.125 172.185 ;
        RECT 55.415 172.015 55.585 172.185 ;
        RECT 98.330 171.895 98.500 172.065 ;
        RECT 98.790 171.895 98.960 172.065 ;
        RECT 99.250 171.895 99.420 172.065 ;
        RECT 99.710 171.895 99.880 172.065 ;
        RECT 100.170 171.895 100.340 172.065 ;
        RECT 100.630 171.895 100.800 172.065 ;
        RECT 101.090 171.895 101.260 172.065 ;
        RECT 101.550 171.895 101.720 172.065 ;
        RECT 102.010 171.895 102.180 172.065 ;
        RECT 102.470 171.895 102.640 172.065 ;
        RECT 102.930 171.895 103.100 172.065 ;
        RECT 103.390 171.895 103.560 172.065 ;
        RECT 103.850 171.895 104.020 172.065 ;
        RECT 104.310 171.895 104.480 172.065 ;
        RECT 113.950 171.865 114.120 172.035 ;
        RECT 185.935 172.015 186.105 172.185 ;
        RECT 186.395 172.015 186.565 172.185 ;
        RECT 186.855 172.015 187.025 172.185 ;
        RECT 187.315 172.015 187.485 172.185 ;
        RECT 187.775 172.015 187.945 172.185 ;
        RECT 188.235 172.015 188.405 172.185 ;
        RECT 188.695 172.015 188.865 172.185 ;
        RECT 189.155 172.015 189.325 172.185 ;
        RECT 189.615 172.015 189.785 172.185 ;
        RECT 190.075 172.015 190.245 172.185 ;
        RECT 190.535 172.015 190.705 172.185 ;
        RECT 190.995 172.015 191.165 172.185 ;
        RECT 191.455 172.015 191.625 172.185 ;
        RECT 191.915 172.015 192.085 172.185 ;
        RECT 51.145 170.935 51.315 171.105 ;
        RECT 51.975 170.935 52.145 171.105 ;
        RECT 100.040 170.815 100.210 170.985 ;
        RECT 100.870 170.815 101.040 170.985 ;
        RECT 189.375 170.935 189.545 171.105 ;
        RECT 190.205 170.935 190.375 171.105 ;
        RECT 105.495 170.240 105.665 170.410 ;
        RECT 105.955 170.240 106.125 170.410 ;
        RECT 106.415 170.240 106.585 170.410 ;
        RECT 106.875 170.240 107.045 170.410 ;
        RECT 107.335 170.240 107.505 170.410 ;
        RECT 107.795 170.240 107.965 170.410 ;
        RECT 108.255 170.240 108.425 170.410 ;
        RECT 108.715 170.240 108.885 170.410 ;
        RECT 109.175 170.240 109.345 170.410 ;
        RECT 109.635 170.240 109.805 170.410 ;
        RECT 110.095 170.240 110.265 170.410 ;
        RECT 110.555 170.240 110.725 170.410 ;
        RECT 111.015 170.240 111.185 170.410 ;
        RECT 111.475 170.240 111.645 170.410 ;
        RECT 111.935 170.240 112.105 170.410 ;
        RECT 112.395 170.240 112.565 170.410 ;
        RECT 112.855 170.240 113.025 170.410 ;
        RECT 113.315 170.240 113.485 170.410 ;
        RECT 113.775 170.240 113.945 170.410 ;
        RECT 114.235 170.240 114.405 170.410 ;
        RECT 114.695 170.240 114.865 170.410 ;
        RECT 115.155 170.240 115.325 170.410 ;
        RECT 115.615 170.240 115.785 170.410 ;
        RECT 116.075 170.240 116.245 170.410 ;
        RECT 116.535 170.240 116.705 170.410 ;
        RECT 116.995 170.240 117.165 170.410 ;
        RECT 117.455 170.240 117.625 170.410 ;
        RECT 47.685 169.600 47.855 169.770 ;
        RECT 48.550 169.600 48.720 169.770 ;
        RECT 49.415 169.600 49.585 169.770 ;
        RECT 50.280 169.600 50.450 169.770 ;
        RECT 51.145 169.600 51.315 169.770 ;
        RECT 52.010 169.600 52.180 169.770 ;
        RECT 52.875 169.600 53.045 169.770 ;
        RECT 53.740 169.600 53.910 169.770 ;
        RECT 54.605 169.600 54.775 169.770 ;
        RECT 96.580 169.480 96.750 169.650 ;
        RECT 97.445 169.480 97.615 169.650 ;
        RECT 98.310 169.480 98.480 169.650 ;
        RECT 99.175 169.480 99.345 169.650 ;
        RECT 100.040 169.480 100.210 169.650 ;
        RECT 100.905 169.480 101.075 169.650 ;
        RECT 101.770 169.480 101.940 169.650 ;
        RECT 102.635 169.480 102.805 169.650 ;
        RECT 103.500 169.480 103.670 169.650 ;
        RECT 121.610 170.145 121.780 170.315 ;
        RECT 122.070 170.145 122.240 170.315 ;
        RECT 122.530 170.145 122.700 170.315 ;
        RECT 122.990 170.145 123.160 170.315 ;
        RECT 123.450 170.145 123.620 170.315 ;
        RECT 123.910 170.145 124.080 170.315 ;
        RECT 124.370 170.145 124.540 170.315 ;
        RECT 124.830 170.145 125.000 170.315 ;
        RECT 125.290 170.145 125.460 170.315 ;
        RECT 186.745 169.600 186.915 169.770 ;
        RECT 187.610 169.600 187.780 169.770 ;
        RECT 188.475 169.600 188.645 169.770 ;
        RECT 189.340 169.600 189.510 169.770 ;
        RECT 190.205 169.600 190.375 169.770 ;
        RECT 191.070 169.600 191.240 169.770 ;
        RECT 191.935 169.600 192.105 169.770 ;
        RECT 192.800 169.600 192.970 169.770 ;
        RECT 193.665 169.600 193.835 169.770 ;
        RECT 113.950 166.425 114.120 166.595 ;
        RECT 105.495 164.800 105.665 164.970 ;
        RECT 105.955 164.800 106.125 164.970 ;
        RECT 106.415 164.800 106.585 164.970 ;
        RECT 106.875 164.800 107.045 164.970 ;
        RECT 107.335 164.800 107.505 164.970 ;
        RECT 107.795 164.800 107.965 164.970 ;
        RECT 108.255 164.800 108.425 164.970 ;
        RECT 108.715 164.800 108.885 164.970 ;
        RECT 109.175 164.800 109.345 164.970 ;
        RECT 109.635 164.800 109.805 164.970 ;
        RECT 110.095 164.800 110.265 164.970 ;
        RECT 110.555 164.800 110.725 164.970 ;
        RECT 111.015 164.800 111.185 164.970 ;
        RECT 111.475 164.800 111.645 164.970 ;
        RECT 111.935 164.800 112.105 164.970 ;
        RECT 112.395 164.800 112.565 164.970 ;
        RECT 112.855 164.800 113.025 164.970 ;
        RECT 113.315 164.800 113.485 164.970 ;
        RECT 113.775 164.800 113.945 164.970 ;
        RECT 114.235 164.800 114.405 164.970 ;
        RECT 114.695 164.800 114.865 164.970 ;
        RECT 115.155 164.800 115.325 164.970 ;
        RECT 115.615 164.800 115.785 164.970 ;
        RECT 116.075 164.800 116.245 164.970 ;
        RECT 116.535 164.800 116.705 164.970 ;
        RECT 116.995 164.800 117.165 164.970 ;
        RECT 117.455 164.800 117.625 164.970 ;
        RECT 96.580 163.430 96.750 163.600 ;
        RECT 97.445 163.430 97.615 163.600 ;
        RECT 98.310 163.430 98.480 163.600 ;
        RECT 99.175 163.430 99.345 163.600 ;
        RECT 100.040 163.430 100.210 163.600 ;
        RECT 100.905 163.430 101.075 163.600 ;
        RECT 101.770 163.430 101.940 163.600 ;
        RECT 102.635 163.430 102.805 163.600 ;
        RECT 103.500 163.430 103.670 163.600 ;
        RECT 121.610 164.705 121.780 164.875 ;
        RECT 122.070 164.705 122.240 164.875 ;
        RECT 122.530 164.705 122.700 164.875 ;
        RECT 122.990 164.705 123.160 164.875 ;
        RECT 123.450 164.705 123.620 164.875 ;
        RECT 123.910 164.705 124.080 164.875 ;
        RECT 124.370 164.705 124.540 164.875 ;
        RECT 124.830 164.705 125.000 164.875 ;
        RECT 125.290 164.705 125.460 164.875 ;
        RECT 100.040 162.095 100.210 162.265 ;
        RECT 100.870 162.095 101.040 162.265 ;
        RECT 98.330 161.015 98.500 161.185 ;
        RECT 98.790 161.015 98.960 161.185 ;
        RECT 99.250 161.015 99.420 161.185 ;
        RECT 99.710 161.015 99.880 161.185 ;
        RECT 100.170 161.015 100.340 161.185 ;
        RECT 100.630 161.015 100.800 161.185 ;
        RECT 101.090 161.015 101.260 161.185 ;
        RECT 101.550 161.015 101.720 161.185 ;
        RECT 102.010 161.015 102.180 161.185 ;
        RECT 102.470 161.015 102.640 161.185 ;
        RECT 102.930 161.015 103.100 161.185 ;
        RECT 103.390 161.015 103.560 161.185 ;
        RECT 103.850 161.015 104.020 161.185 ;
        RECT 104.310 161.015 104.480 161.185 ;
        RECT 113.950 160.985 114.120 161.155 ;
        RECT 105.495 159.360 105.665 159.530 ;
        RECT 105.955 159.360 106.125 159.530 ;
        RECT 106.415 159.360 106.585 159.530 ;
        RECT 106.875 159.360 107.045 159.530 ;
        RECT 107.335 159.360 107.505 159.530 ;
        RECT 107.795 159.360 107.965 159.530 ;
        RECT 108.255 159.360 108.425 159.530 ;
        RECT 108.715 159.360 108.885 159.530 ;
        RECT 109.175 159.360 109.345 159.530 ;
        RECT 109.635 159.360 109.805 159.530 ;
        RECT 110.095 159.360 110.265 159.530 ;
        RECT 110.555 159.360 110.725 159.530 ;
        RECT 111.015 159.360 111.185 159.530 ;
        RECT 111.475 159.360 111.645 159.530 ;
        RECT 111.935 159.360 112.105 159.530 ;
        RECT 112.395 159.360 112.565 159.530 ;
        RECT 112.855 159.360 113.025 159.530 ;
        RECT 113.315 159.360 113.485 159.530 ;
        RECT 113.775 159.360 113.945 159.530 ;
        RECT 114.235 159.360 114.405 159.530 ;
        RECT 114.695 159.360 114.865 159.530 ;
        RECT 115.155 159.360 115.325 159.530 ;
        RECT 115.615 159.360 115.785 159.530 ;
        RECT 116.075 159.360 116.245 159.530 ;
        RECT 116.535 159.360 116.705 159.530 ;
        RECT 116.995 159.360 117.165 159.530 ;
        RECT 117.455 159.360 117.625 159.530 ;
        RECT 111.090 146.930 111.260 147.100 ;
        RECT 129.120 146.930 129.290 147.100 ;
        RECT 3.225 132.615 3.395 132.785 ;
        RECT 236.985 132.615 237.155 132.785 ;
        RECT 10.025 131.100 10.195 131.270 ;
        RECT 31.325 131.100 31.495 131.270 ;
        RECT 68.775 131.100 68.945 131.270 ;
        RECT 99.825 131.100 99.995 131.270 ;
        RECT 134.515 131.100 134.685 131.270 ;
        RECT 165.275 131.100 165.445 131.270 ;
        RECT 203.965 131.100 204.135 131.270 ;
        RECT 221.815 131.100 221.985 131.270 ;
      LAYER met1 ;
        RECT 104.145 175.525 117.770 176.005 ;
        RECT 49.290 171.860 57.570 172.340 ;
        RECT 104.145 172.220 104.625 175.525 ;
        RECT 51.310 171.165 51.750 171.860 ;
        RECT 98.185 171.740 104.625 172.220 ;
        RECT 113.900 172.005 114.170 172.120 ;
        RECT 113.900 171.780 114.730 172.005 ;
        RECT 183.950 171.860 192.230 172.340 ;
        RECT 51.115 171.105 51.750 171.165 ;
        RECT 51.945 171.105 52.175 171.135 ;
        RECT 51.115 170.935 52.205 171.105 ;
        RECT 100.205 171.045 100.645 171.740 ;
        RECT 100.010 170.985 100.645 171.045 ;
        RECT 100.840 170.985 101.070 171.015 ;
        RECT 51.115 170.905 51.345 170.935 ;
        RECT 51.945 170.905 52.175 170.935 ;
        RECT 51.145 169.800 51.315 170.905 ;
        RECT 100.010 170.815 101.100 170.985 ;
        RECT 100.010 170.785 100.240 170.815 ;
        RECT 100.840 170.785 101.070 170.815 ;
        RECT 47.625 169.640 54.835 169.800 ;
        RECT 100.040 169.680 100.210 170.785 ;
        RECT 114.505 170.565 114.730 171.780 ;
        RECT 189.770 171.165 190.210 171.860 ;
        RECT 189.345 171.105 189.575 171.135 ;
        RECT 189.770 171.105 190.405 171.165 ;
        RECT 189.315 170.935 190.405 171.105 ;
        RECT 189.345 170.905 189.575 170.935 ;
        RECT 190.175 170.905 190.405 170.935 ;
        RECT 105.350 170.500 117.770 170.565 ;
        RECT 105.350 170.470 121.595 170.500 ;
        RECT 105.350 170.105 125.605 170.470 ;
        RECT 105.350 170.085 117.770 170.105 ;
        RECT 121.465 169.990 125.605 170.105 ;
        RECT 190.205 169.800 190.375 170.905 ;
        RECT 47.625 169.570 47.915 169.640 ;
        RECT 48.490 169.570 48.780 169.640 ;
        RECT 49.355 169.570 49.645 169.640 ;
        RECT 50.220 169.570 50.510 169.640 ;
        RECT 51.085 169.570 51.375 169.640 ;
        RECT 51.950 169.570 52.240 169.640 ;
        RECT 52.815 169.570 53.105 169.640 ;
        RECT 53.680 169.570 53.970 169.640 ;
        RECT 54.545 169.570 54.835 169.640 ;
        RECT 96.520 169.520 103.730 169.680 ;
        RECT 186.685 169.640 193.895 169.800 ;
        RECT 186.685 169.570 186.975 169.640 ;
        RECT 187.550 169.570 187.840 169.640 ;
        RECT 188.415 169.570 188.705 169.640 ;
        RECT 189.280 169.570 189.570 169.640 ;
        RECT 190.145 169.570 190.435 169.640 ;
        RECT 191.010 169.570 191.300 169.640 ;
        RECT 191.875 169.570 192.165 169.640 ;
        RECT 192.740 169.570 193.030 169.640 ;
        RECT 193.605 169.570 193.895 169.640 ;
        RECT 96.520 169.450 96.810 169.520 ;
        RECT 97.385 169.450 97.675 169.520 ;
        RECT 98.250 169.450 98.540 169.520 ;
        RECT 99.115 169.450 99.405 169.520 ;
        RECT 99.980 169.450 100.270 169.520 ;
        RECT 100.845 169.450 101.135 169.520 ;
        RECT 101.710 169.450 102.000 169.520 ;
        RECT 102.575 169.450 102.865 169.520 ;
        RECT 103.440 169.450 103.730 169.520 ;
        RECT 113.900 166.565 114.170 166.680 ;
        RECT 113.900 166.340 114.730 166.565 ;
        RECT 114.505 165.125 114.730 166.340 ;
        RECT 105.350 165.030 117.770 165.125 ;
        RECT 105.350 164.645 125.605 165.030 ;
        RECT 117.690 164.635 125.605 164.645 ;
        RECT 121.465 164.550 125.605 164.635 ;
        RECT 96.520 163.560 96.810 163.630 ;
        RECT 97.385 163.560 97.675 163.630 ;
        RECT 98.250 163.560 98.540 163.630 ;
        RECT 99.115 163.560 99.405 163.630 ;
        RECT 99.980 163.560 100.270 163.630 ;
        RECT 100.845 163.560 101.135 163.630 ;
        RECT 101.710 163.560 102.000 163.630 ;
        RECT 102.575 163.560 102.865 163.630 ;
        RECT 103.440 163.560 103.730 163.630 ;
        RECT 96.520 163.400 103.730 163.560 ;
        RECT 100.040 162.295 100.210 163.400 ;
        RECT 100.010 162.265 100.240 162.295 ;
        RECT 100.840 162.265 101.070 162.295 ;
        RECT 100.010 162.095 101.100 162.265 ;
        RECT 100.010 162.035 100.645 162.095 ;
        RECT 100.840 162.065 101.070 162.095 ;
        RECT 100.205 161.340 100.645 162.035 ;
        RECT 98.185 160.860 104.920 161.340 ;
        RECT 113.900 161.125 114.170 161.240 ;
        RECT 113.900 160.900 114.730 161.125 ;
        RECT 104.440 159.685 104.920 160.860 ;
        RECT 114.505 159.685 114.730 160.900 ;
        RECT 104.440 159.205 117.770 159.685 ;
        RECT 9.980 146.910 10.240 147.230 ;
        RECT 18.340 146.885 18.620 147.255 ;
        RECT 31.280 146.910 31.540 147.230 ;
        RECT 36.200 146.910 36.460 147.230 ;
        RECT 68.730 146.910 68.990 147.230 ;
        RECT 74.890 146.910 75.150 147.230 ;
        RECT 99.780 146.910 100.040 147.230 ;
        RECT 105.650 146.910 105.910 147.230 ;
        RECT 109.615 147.100 109.985 147.165 ;
        RECT 111.020 147.100 111.325 147.160 ;
        RECT 109.615 146.925 111.325 147.100 ;
        RECT 109.615 146.885 109.985 146.925 ;
        RECT 111.020 146.875 111.325 146.925 ;
        RECT 129.055 147.100 129.360 147.160 ;
        RECT 130.395 147.100 130.765 147.165 ;
        RECT 129.055 146.925 130.765 147.100 ;
        RECT 129.055 146.875 129.360 146.925 ;
        RECT 130.395 146.885 130.765 146.925 ;
        RECT 134.470 146.910 134.730 147.230 ;
        RECT 140.340 146.910 140.600 147.230 ;
        RECT 165.230 146.910 165.490 147.230 ;
        RECT 171.390 146.910 171.650 147.230 ;
        RECT 203.920 146.910 204.180 147.230 ;
        RECT 208.840 146.910 209.100 147.230 ;
        RECT 221.760 146.885 222.040 147.255 ;
        RECT 230.140 146.910 230.400 147.230 ;
        RECT 2.435 132.785 2.775 133.260 ;
        RECT 3.190 132.785 3.425 132.820 ;
        RECT 236.955 132.785 237.190 132.820 ;
        RECT 237.605 132.785 237.945 133.260 ;
        RECT 2.435 132.615 3.455 132.785 ;
        RECT 236.925 132.615 237.945 132.785 ;
        RECT 2.435 128.715 2.775 132.615 ;
        RECT 3.190 132.580 3.425 132.615 ;
        RECT 236.955 132.580 237.190 132.615 ;
        RECT 9.980 131.030 10.240 131.350 ;
        RECT 18.350 131.030 18.610 131.350 ;
        RECT 31.280 131.030 31.540 131.350 ;
        RECT 36.200 131.030 36.460 131.350 ;
        RECT 68.730 131.030 68.990 131.350 ;
        RECT 74.890 131.030 75.150 131.350 ;
        RECT 99.780 131.030 100.040 131.350 ;
        RECT 105.650 131.030 105.910 131.350 ;
        RECT 134.470 131.030 134.730 131.350 ;
        RECT 140.340 131.030 140.600 131.350 ;
        RECT 165.230 131.030 165.490 131.350 ;
        RECT 171.390 131.030 171.650 131.350 ;
        RECT 203.920 131.030 204.180 131.350 ;
        RECT 208.840 131.030 209.100 131.350 ;
        RECT 221.770 131.030 222.030 131.350 ;
        RECT 230.140 131.030 230.400 131.350 ;
        RECT 237.605 128.715 237.945 132.615 ;
      LAYER via ;
        RECT 107.870 175.640 108.130 175.900 ;
        RECT 112.475 175.640 112.735 175.900 ;
        RECT 117.065 175.650 117.325 175.910 ;
        RECT 56.380 171.880 57.540 172.320 ;
        RECT 183.980 171.880 185.140 172.320 ;
        RECT 107.870 170.205 108.130 170.465 ;
        RECT 112.480 170.195 112.740 170.455 ;
        RECT 117.060 170.195 117.320 170.455 ;
        RECT 107.865 164.755 108.125 165.015 ;
        RECT 112.475 164.765 112.735 165.025 ;
        RECT 117.070 164.765 117.330 165.025 ;
        RECT 107.870 159.320 108.130 159.580 ;
        RECT 112.490 159.320 112.750 159.580 ;
        RECT 117.060 159.320 117.320 159.580 ;
        RECT 9.980 146.940 10.240 147.200 ;
        RECT 18.350 146.940 18.610 147.200 ;
        RECT 31.280 146.940 31.540 147.200 ;
        RECT 36.200 146.940 36.460 147.200 ;
        RECT 68.730 146.940 68.990 147.200 ;
        RECT 74.890 146.940 75.150 147.200 ;
        RECT 99.780 146.940 100.040 147.200 ;
        RECT 105.650 146.940 105.910 147.200 ;
        RECT 109.660 146.885 109.940 147.165 ;
        RECT 130.440 146.885 130.720 147.165 ;
        RECT 134.470 146.940 134.730 147.200 ;
        RECT 140.340 146.940 140.600 147.200 ;
        RECT 165.230 146.940 165.490 147.200 ;
        RECT 171.390 146.940 171.650 147.200 ;
        RECT 203.920 146.940 204.180 147.200 ;
        RECT 208.840 146.940 209.100 147.200 ;
        RECT 221.770 146.940 222.030 147.200 ;
        RECT 230.140 146.940 230.400 147.200 ;
        RECT 2.470 132.820 2.730 133.080 ;
        RECT 237.650 132.820 237.910 133.080 ;
        RECT 9.980 131.060 10.240 131.320 ;
        RECT 18.350 131.060 18.610 131.320 ;
        RECT 31.280 131.060 31.540 131.320 ;
        RECT 36.200 131.060 36.460 131.320 ;
        RECT 68.730 131.060 68.990 131.320 ;
        RECT 74.890 131.060 75.150 131.320 ;
        RECT 99.780 131.060 100.040 131.320 ;
        RECT 105.650 131.060 105.910 131.320 ;
        RECT 134.470 131.060 134.730 131.320 ;
        RECT 140.340 131.060 140.600 131.320 ;
        RECT 165.230 131.060 165.490 131.320 ;
        RECT 171.390 131.060 171.650 131.320 ;
        RECT 203.920 131.060 204.180 131.320 ;
        RECT 208.840 131.060 209.100 131.320 ;
        RECT 221.770 131.060 222.030 131.320 ;
        RECT 230.140 131.060 230.400 131.320 ;
      LAYER met2 ;
        RECT 107.860 175.585 108.140 175.955 ;
        RECT 112.465 175.585 112.745 175.955 ;
        RECT 117.055 175.595 117.335 175.965 ;
        RECT 56.380 147.360 57.540 172.350 ;
        RECT 107.860 170.150 108.140 170.520 ;
        RECT 112.470 170.140 112.750 170.510 ;
        RECT 117.050 170.140 117.330 170.510 ;
        RECT 107.855 164.700 108.135 165.070 ;
        RECT 112.465 164.710 112.745 165.080 ;
        RECT 117.060 164.710 117.340 165.080 ;
        RECT 107.860 159.265 108.140 159.635 ;
        RECT 112.480 159.265 112.760 159.635 ;
        RECT 117.050 159.265 117.330 159.635 ;
        RECT 183.980 147.360 185.140 172.350 ;
        RECT 2.460 146.860 2.740 147.230 ;
        RECT 9.970 146.885 10.250 147.255 ;
        RECT 18.340 146.885 18.620 147.255 ;
        RECT 31.270 146.885 31.550 147.255 ;
        RECT 36.190 146.885 36.470 147.255 ;
        RECT 2.470 132.790 2.730 146.860 ;
        RECT 10.025 131.350 10.195 146.885 ;
        RECT 18.395 131.350 18.565 146.885 ;
        RECT 31.325 131.350 31.495 146.885 ;
        RECT 36.245 131.350 36.415 146.885 ;
        RECT 56.330 146.740 57.590 147.360 ;
        RECT 68.720 146.880 69.000 147.250 ;
        RECT 74.880 146.885 75.160 147.260 ;
        RECT 99.770 146.885 100.050 147.260 ;
        RECT 68.775 131.350 68.945 146.880 ;
        RECT 74.935 131.350 75.105 146.885 ;
        RECT 99.825 131.350 99.995 146.885 ;
        RECT 105.635 146.880 105.925 147.265 ;
        RECT 109.615 146.885 109.985 147.165 ;
        RECT 130.395 146.885 130.765 147.165 ;
        RECT 134.455 146.880 134.745 147.265 ;
        RECT 140.330 146.885 140.610 147.260 ;
        RECT 165.220 146.885 165.500 147.260 ;
        RECT 105.695 131.350 105.865 146.880 ;
        RECT 134.515 131.350 134.685 146.880 ;
        RECT 140.385 131.350 140.555 146.885 ;
        RECT 165.275 131.350 165.445 146.885 ;
        RECT 171.380 146.880 171.660 147.250 ;
        RECT 171.435 131.350 171.605 146.880 ;
        RECT 183.930 146.740 185.190 147.360 ;
        RECT 203.910 146.885 204.190 147.255 ;
        RECT 208.830 146.885 209.110 147.255 ;
        RECT 221.760 146.885 222.040 147.255 ;
        RECT 230.130 146.885 230.410 147.255 ;
        RECT 203.965 131.350 204.135 146.885 ;
        RECT 208.885 131.350 209.055 146.885 ;
        RECT 221.815 131.350 221.985 146.885 ;
        RECT 230.185 131.350 230.355 146.885 ;
        RECT 237.640 146.860 237.920 147.230 ;
        RECT 237.650 132.790 237.910 146.860 ;
        RECT 9.980 131.030 10.240 131.350 ;
        RECT 18.350 131.030 18.610 131.350 ;
        RECT 31.280 131.030 31.540 131.350 ;
        RECT 36.200 131.030 36.460 131.350 ;
        RECT 68.730 131.030 68.990 131.350 ;
        RECT 74.890 131.030 75.150 131.350 ;
        RECT 99.780 131.030 100.040 131.350 ;
        RECT 105.650 131.030 105.910 131.350 ;
        RECT 134.470 131.030 134.730 131.350 ;
        RECT 140.340 131.030 140.600 131.350 ;
        RECT 165.230 131.030 165.490 131.350 ;
        RECT 171.390 131.030 171.650 131.350 ;
        RECT 203.920 131.030 204.180 131.350 ;
        RECT 208.840 131.030 209.100 131.350 ;
        RECT 221.770 131.030 222.030 131.350 ;
        RECT 230.140 131.030 230.400 131.350 ;
      LAYER via2 ;
        RECT 107.860 175.630 108.140 175.910 ;
        RECT 112.465 175.630 112.745 175.910 ;
        RECT 117.055 175.640 117.335 175.920 ;
        RECT 107.860 170.195 108.140 170.475 ;
        RECT 112.470 170.185 112.750 170.465 ;
        RECT 117.050 170.185 117.330 170.465 ;
        RECT 107.855 164.745 108.135 165.025 ;
        RECT 112.465 164.755 112.745 165.035 ;
        RECT 117.060 164.755 117.340 165.035 ;
        RECT 107.860 159.310 108.140 159.590 ;
        RECT 112.480 159.310 112.760 159.590 ;
        RECT 117.050 159.310 117.330 159.590 ;
        RECT 2.460 146.905 2.740 147.185 ;
        RECT 9.970 146.930 10.250 147.210 ;
        RECT 18.340 146.930 18.620 147.210 ;
        RECT 31.270 146.930 31.550 147.210 ;
        RECT 36.190 146.930 36.470 147.210 ;
        RECT 56.380 146.790 57.540 147.280 ;
        RECT 68.720 146.925 69.000 147.205 ;
        RECT 74.880 146.930 75.160 147.210 ;
        RECT 99.770 146.930 100.050 147.210 ;
        RECT 105.635 146.925 105.925 147.220 ;
        RECT 109.660 146.885 109.940 147.165 ;
        RECT 130.440 146.885 130.720 147.165 ;
        RECT 134.455 146.925 134.745 147.220 ;
        RECT 140.330 146.930 140.610 147.210 ;
        RECT 165.220 146.930 165.500 147.210 ;
        RECT 171.380 146.925 171.660 147.205 ;
        RECT 183.980 146.790 185.140 147.280 ;
        RECT 203.910 146.930 204.190 147.210 ;
        RECT 208.830 146.930 209.110 147.210 ;
        RECT 221.760 146.930 222.040 147.210 ;
        RECT 230.130 146.930 230.410 147.210 ;
        RECT 237.640 146.905 237.920 147.185 ;
      LAYER met3 ;
        RECT 107.760 175.530 108.250 176.020 ;
        RECT 112.365 175.530 112.855 176.020 ;
        RECT 116.955 175.540 117.445 176.030 ;
        RECT 107.760 170.095 108.250 170.585 ;
        RECT 112.370 170.085 112.860 170.575 ;
        RECT 116.950 170.085 117.440 170.575 ;
        RECT 107.755 164.645 108.245 165.135 ;
        RECT 112.365 164.655 112.855 165.145 ;
        RECT 116.960 164.655 117.450 165.145 ;
        RECT 107.760 159.210 108.250 159.700 ;
        RECT 112.380 159.210 112.870 159.700 ;
        RECT 116.950 159.210 117.440 159.700 ;
        RECT 56.330 147.290 57.590 147.360 ;
        RECT 183.930 147.290 185.190 147.360 ;
        RECT -0.130 146.790 253.790 147.290 ;
        RECT 56.330 146.740 57.590 146.790 ;
        RECT 183.930 146.740 185.190 146.790 ;
      LAYER via3 ;
        RECT 107.840 175.610 108.160 175.930 ;
        RECT 112.445 175.610 112.765 175.930 ;
        RECT 117.035 175.620 117.355 175.940 ;
        RECT 107.840 170.175 108.160 170.495 ;
        RECT 112.450 170.165 112.770 170.485 ;
        RECT 117.030 170.165 117.350 170.485 ;
        RECT 107.835 164.725 108.155 165.045 ;
        RECT 112.445 164.735 112.765 165.055 ;
        RECT 117.040 164.735 117.360 165.055 ;
        RECT 107.840 159.290 108.160 159.610 ;
        RECT 112.460 159.290 112.780 159.610 ;
        RECT 117.030 159.290 117.350 159.610 ;
        RECT 112.415 146.865 112.775 147.225 ;
      LAYER met4 ;
        RECT 107.755 159.205 108.185 176.005 ;
        RECT 112.365 159.205 112.795 176.005 ;
        RECT 116.945 159.205 117.375 176.005 ;
        RECT 112.405 146.705 112.790 159.205 ;
    END
  END vdda
  PIN vssd
    DIRECTION INOUT ;
    ANTENNAGATEAREA 1.587600 ;
    ANTENNADIFFAREA 24.673849 ;
    PORT
      LAYER li1 ;
        RECT 112.405 173.865 112.635 173.880 ;
        RECT 112.855 173.865 113.085 173.890 ;
        RECT 112.405 173.860 113.085 173.865 ;
        RECT 115.165 173.865 115.395 173.880 ;
        RECT 115.615 173.865 115.845 173.890 ;
        RECT 115.165 173.860 115.845 173.865 ;
        RECT 112.405 173.450 113.130 173.860 ;
        RECT 115.165 173.450 115.890 173.860 ;
        RECT 112.405 173.430 113.085 173.450 ;
        RECT 115.165 173.430 115.845 173.450 ;
        RECT 112.405 173.425 112.905 173.430 ;
        RECT 115.165 173.425 115.665 173.430 ;
        RECT 112.435 173.130 112.905 173.425 ;
        RECT 115.195 173.130 115.665 173.425 ;
        RECT 105.350 172.960 117.770 173.130 ;
        RECT 106.490 171.420 106.665 172.960 ;
        RECT 105.965 171.395 106.195 171.410 ;
        RECT 106.415 171.395 106.665 171.420 ;
        RECT 109.400 171.525 109.570 172.960 ;
        RECT 112.775 172.645 112.945 172.960 ;
        RECT 115.195 172.665 115.665 172.960 ;
        RECT 115.165 172.660 115.665 172.665 ;
        RECT 112.675 172.230 113.025 172.645 ;
        RECT 115.165 172.640 115.845 172.660 ;
        RECT 115.165 172.230 115.890 172.640 ;
        RECT 115.165 172.225 115.845 172.230 ;
        RECT 115.165 172.210 115.395 172.225 ;
        RECT 115.615 172.200 115.845 172.225 ;
        RECT 113.145 171.625 113.315 171.955 ;
        RECT 109.400 171.405 109.815 171.525 ;
        RECT 105.965 171.390 106.665 171.395 ;
        RECT 105.965 170.980 106.690 171.390 ;
        RECT 109.035 171.205 109.815 171.405 ;
        RECT 109.535 171.105 109.815 171.205 ;
        RECT 105.965 170.960 106.645 170.980 ;
        RECT 105.965 170.955 106.495 170.960 ;
        RECT 45.125 170.470 45.295 170.800 ;
        RECT 94.020 170.350 94.190 170.680 ;
        RECT 196.225 170.470 196.395 170.800 ;
        RECT 44.655 169.780 45.005 170.195 ;
        RECT 44.755 169.465 44.925 169.780 ;
        RECT 93.550 169.660 93.900 170.075 ;
        RECT 196.515 169.780 196.865 170.195 ;
        RECT 43.770 169.295 46.990 169.465 ;
        RECT 93.650 169.345 93.820 169.660 ;
        RECT 196.595 169.465 196.765 169.780 ;
        RECT 44.415 169.000 44.885 169.295 ;
        RECT 92.665 169.175 95.885 169.345 ;
        RECT 194.530 169.295 197.750 169.465 ;
        RECT 44.385 168.995 44.885 169.000 ;
        RECT 44.385 168.975 45.065 168.995 ;
        RECT 44.385 168.565 45.110 168.975 ;
        RECT 93.310 168.880 93.780 169.175 ;
        RECT 196.635 169.000 197.105 169.295 ;
        RECT 196.635 168.995 197.135 169.000 ;
        RECT 196.455 168.975 197.135 168.995 ;
        RECT 93.280 168.875 93.780 168.880 ;
        RECT 93.280 168.855 93.960 168.875 ;
        RECT 44.385 168.560 45.065 168.565 ;
        RECT 44.385 168.545 44.615 168.560 ;
        RECT 44.835 168.535 45.065 168.560 ;
        RECT 93.280 168.445 94.005 168.855 ;
        RECT 196.410 168.565 197.135 168.975 ;
        RECT 196.455 168.560 197.135 168.565 ;
        RECT 196.455 168.535 196.685 168.560 ;
        RECT 196.905 168.545 197.135 168.560 ;
        RECT 93.280 168.440 93.960 168.445 ;
        RECT 93.280 168.425 93.510 168.440 ;
        RECT 93.730 168.415 93.960 168.440 ;
        RECT 112.405 168.425 112.635 168.440 ;
        RECT 112.855 168.425 113.085 168.450 ;
        RECT 112.405 168.420 113.085 168.425 ;
        RECT 115.165 168.425 115.395 168.440 ;
        RECT 115.615 168.425 115.845 168.450 ;
        RECT 115.165 168.420 115.845 168.425 ;
        RECT 112.405 168.010 113.130 168.420 ;
        RECT 115.165 168.010 115.890 168.420 ;
        RECT 112.405 167.990 113.085 168.010 ;
        RECT 115.165 167.990 115.845 168.010 ;
        RECT 112.405 167.985 112.905 167.990 ;
        RECT 115.165 167.985 115.665 167.990 ;
        RECT 112.435 167.690 112.905 167.985 ;
        RECT 115.195 167.690 115.665 167.985 ;
        RECT 47.325 167.215 47.495 167.545 ;
        RECT 47.685 167.320 47.855 167.650 ;
        RECT 48.550 167.320 48.720 167.650 ;
        RECT 49.415 167.320 49.585 167.650 ;
        RECT 50.280 167.320 50.450 167.650 ;
        RECT 51.145 167.320 51.315 167.650 ;
        RECT 52.010 167.320 52.180 167.650 ;
        RECT 52.875 167.320 53.045 167.650 ;
        RECT 53.740 167.320 53.910 167.650 ;
        RECT 54.605 167.320 54.775 167.650 ;
        RECT 54.995 166.745 55.165 167.575 ;
        RECT 96.220 167.095 96.390 167.425 ;
        RECT 96.580 167.200 96.750 167.530 ;
        RECT 97.445 167.200 97.615 167.530 ;
        RECT 98.310 167.200 98.480 167.530 ;
        RECT 99.175 167.200 99.345 167.530 ;
        RECT 100.040 167.200 100.210 167.530 ;
        RECT 100.905 167.200 101.075 167.530 ;
        RECT 101.770 167.200 101.940 167.530 ;
        RECT 102.635 167.200 102.805 167.530 ;
        RECT 103.500 167.200 103.670 167.530 ;
        RECT 105.350 167.520 117.770 167.690 ;
        RECT 121.720 167.595 121.975 168.055 ;
        RECT 122.645 167.595 122.815 168.055 ;
        RECT 123.485 167.595 123.655 168.055 ;
        RECT 124.325 167.595 124.495 168.055 ;
        RECT 125.165 167.595 125.470 168.055 ;
        RECT 49.740 166.575 55.730 166.745 ;
        RECT 103.890 166.625 104.060 167.455 ;
        RECT 98.635 166.455 104.625 166.625 ;
        RECT 96.220 165.655 96.390 165.985 ;
        RECT 96.580 165.550 96.750 165.880 ;
        RECT 97.445 165.550 97.615 165.880 ;
        RECT 98.310 165.550 98.480 165.880 ;
        RECT 99.175 165.550 99.345 165.880 ;
        RECT 100.040 165.550 100.210 165.880 ;
        RECT 100.905 165.550 101.075 165.880 ;
        RECT 101.770 165.550 101.940 165.880 ;
        RECT 102.635 165.550 102.805 165.880 ;
        RECT 103.500 165.550 103.670 165.880 ;
        RECT 103.890 165.625 104.060 166.455 ;
        RECT 106.490 165.980 106.665 167.520 ;
        RECT 105.965 165.955 106.195 165.970 ;
        RECT 106.415 165.955 106.665 165.980 ;
        RECT 109.400 166.085 109.570 167.520 ;
        RECT 112.775 167.205 112.945 167.520 ;
        RECT 115.195 167.225 115.665 167.520 ;
        RECT 121.465 167.425 125.605 167.595 ;
        RECT 115.165 167.220 115.665 167.225 ;
        RECT 112.675 166.790 113.025 167.205 ;
        RECT 115.165 167.200 115.845 167.220 ;
        RECT 115.165 166.790 115.890 167.200 ;
        RECT 121.720 166.965 121.975 167.425 ;
        RECT 122.645 166.965 122.815 167.425 ;
        RECT 123.485 166.965 123.655 167.425 ;
        RECT 124.325 166.965 124.495 167.425 ;
        RECT 125.165 166.965 125.470 167.425 ;
        RECT 126.300 167.050 126.555 167.970 ;
        RECT 127.510 167.595 127.765 168.055 ;
        RECT 128.435 167.595 128.605 168.055 ;
        RECT 129.275 167.595 129.445 168.055 ;
        RECT 130.115 167.595 130.285 168.055 ;
        RECT 130.955 167.595 131.260 168.055 ;
        RECT 127.255 167.425 131.395 167.595 ;
        RECT 127.510 166.965 127.765 167.425 ;
        RECT 128.435 166.965 128.605 167.425 ;
        RECT 129.275 166.965 129.445 167.425 ;
        RECT 130.115 166.965 130.285 167.425 ;
        RECT 130.955 166.965 131.260 167.425 ;
        RECT 115.165 166.785 115.845 166.790 ;
        RECT 115.165 166.770 115.395 166.785 ;
        RECT 115.615 166.760 115.845 166.785 ;
        RECT 186.355 166.745 186.525 167.575 ;
        RECT 186.745 167.320 186.915 167.650 ;
        RECT 187.610 167.320 187.780 167.650 ;
        RECT 188.475 167.320 188.645 167.650 ;
        RECT 189.340 167.320 189.510 167.650 ;
        RECT 190.205 167.320 190.375 167.650 ;
        RECT 191.070 167.320 191.240 167.650 ;
        RECT 191.935 167.320 192.105 167.650 ;
        RECT 192.800 167.320 192.970 167.650 ;
        RECT 193.665 167.320 193.835 167.650 ;
        RECT 194.025 167.215 194.195 167.545 ;
        RECT 185.790 166.575 191.780 166.745 ;
        RECT 113.145 166.185 113.315 166.515 ;
        RECT 109.400 165.965 109.815 166.085 ;
        RECT 105.965 165.950 106.665 165.955 ;
        RECT 105.965 165.540 106.690 165.950 ;
        RECT 109.035 165.765 109.815 165.965 ;
        RECT 109.535 165.665 109.815 165.765 ;
        RECT 105.965 165.520 106.645 165.540 ;
        RECT 105.965 165.515 106.495 165.520 ;
        RECT 93.280 164.640 93.510 164.655 ;
        RECT 93.730 164.640 93.960 164.665 ;
        RECT 93.280 164.635 93.960 164.640 ;
        RECT 93.280 164.225 94.005 164.635 ;
        RECT 93.280 164.205 93.960 164.225 ;
        RECT 93.280 164.200 93.780 164.205 ;
        RECT 93.310 163.905 93.780 164.200 ;
        RECT 92.665 163.735 95.885 163.905 ;
        RECT 93.650 163.420 93.820 163.735 ;
        RECT 93.550 163.005 93.900 163.420 ;
        RECT 112.405 162.985 112.635 163.000 ;
        RECT 112.855 162.985 113.085 163.010 ;
        RECT 112.405 162.980 113.085 162.985 ;
        RECT 115.165 162.985 115.395 163.000 ;
        RECT 115.615 162.985 115.845 163.010 ;
        RECT 115.165 162.980 115.845 162.985 ;
        RECT 94.020 162.400 94.190 162.730 ;
        RECT 112.405 162.570 113.130 162.980 ;
        RECT 115.165 162.570 115.890 162.980 ;
        RECT 112.405 162.550 113.085 162.570 ;
        RECT 115.165 162.550 115.845 162.570 ;
        RECT 112.405 162.545 112.905 162.550 ;
        RECT 115.165 162.545 115.665 162.550 ;
        RECT 112.435 162.250 112.905 162.545 ;
        RECT 115.195 162.250 115.665 162.545 ;
        RECT 105.350 162.080 117.770 162.250 ;
        RECT 106.490 160.540 106.665 162.080 ;
        RECT 109.710 160.540 109.885 162.080 ;
        RECT 112.775 161.765 112.945 162.080 ;
        RECT 115.195 161.785 115.665 162.080 ;
        RECT 115.165 161.780 115.665 161.785 ;
        RECT 112.675 161.350 113.025 161.765 ;
        RECT 115.165 161.760 115.845 161.780 ;
        RECT 115.165 161.350 115.890 161.760 ;
        RECT 115.165 161.345 115.845 161.350 ;
        RECT 115.165 161.330 115.395 161.345 ;
        RECT 115.615 161.320 115.845 161.345 ;
        RECT 113.145 160.745 113.315 161.075 ;
        RECT 105.965 160.515 106.195 160.530 ;
        RECT 106.415 160.515 106.665 160.540 ;
        RECT 105.965 160.510 106.665 160.515 ;
        RECT 109.185 160.515 109.415 160.530 ;
        RECT 109.635 160.515 109.885 160.540 ;
        RECT 109.185 160.510 109.885 160.515 ;
        RECT 105.965 160.100 106.690 160.510 ;
        RECT 109.185 160.100 109.910 160.510 ;
        RECT 105.965 160.080 106.645 160.100 ;
        RECT 109.185 160.080 109.865 160.100 ;
        RECT 105.965 160.075 106.495 160.080 ;
        RECT 109.185 160.075 109.715 160.080 ;
        RECT 116.920 134.695 117.250 134.865 ;
        RECT 123.200 134.695 123.530 134.865 ;
        RECT 117.000 134.510 117.170 134.695 ;
        RECT 123.280 134.510 123.450 134.695 ;
        RECT 116.830 134.245 117.330 134.510 ;
        RECT 123.110 134.245 123.610 134.510 ;
        RECT 5.075 132.575 5.405 132.745 ;
        RECT 234.975 132.575 235.305 132.745 ;
        RECT 111.920 131.065 112.270 131.445 ;
        RECT 113.080 131.065 113.430 131.445 ;
        RECT 114.240 131.065 114.590 131.445 ;
        RECT 115.400 131.340 115.750 131.445 ;
        RECT 124.690 131.345 125.040 131.445 ;
        RECT 115.400 131.165 116.215 131.340 ;
        RECT 124.225 131.170 125.040 131.345 ;
        RECT 115.400 131.065 115.750 131.165 ;
        RECT 124.690 131.065 125.040 131.170 ;
        RECT 125.850 131.065 126.200 131.445 ;
        RECT 127.010 131.065 127.360 131.445 ;
        RECT 128.170 131.065 128.520 131.445 ;
        RECT 9.725 128.985 9.895 129.810 ;
        RECT 18.695 128.985 18.865 129.810 ;
        RECT 31.025 128.985 31.195 129.810 ;
        RECT 36.545 128.985 36.715 129.810 ;
        RECT 68.475 128.985 68.645 129.810 ;
        RECT 75.235 128.985 75.405 129.810 ;
        RECT 99.525 128.985 99.695 129.810 ;
        RECT 105.995 128.985 106.165 129.810 ;
        RECT 115.970 129.695 117.330 129.960 ;
        RECT 123.110 129.695 124.470 129.960 ;
        RECT 134.215 128.985 134.385 129.810 ;
        RECT 140.685 128.985 140.855 129.810 ;
        RECT 164.975 128.985 165.145 129.810 ;
        RECT 171.735 128.985 171.905 129.810 ;
        RECT 203.665 128.985 203.835 129.810 ;
        RECT 209.185 128.985 209.355 129.810 ;
        RECT 221.515 128.985 221.685 129.810 ;
        RECT 230.485 128.985 230.655 129.810 ;
        RECT 119.970 125.495 120.470 125.760 ;
        RECT 120.140 125.310 120.310 125.495 ;
        RECT 120.060 125.140 120.390 125.310 ;
      LAYER mcon ;
        RECT 105.495 172.960 105.665 173.130 ;
        RECT 105.955 172.960 106.125 173.130 ;
        RECT 106.415 172.960 106.585 173.130 ;
        RECT 106.875 172.960 107.045 173.130 ;
        RECT 107.335 172.960 107.505 173.130 ;
        RECT 107.795 172.960 107.965 173.130 ;
        RECT 108.255 172.960 108.425 173.130 ;
        RECT 108.715 172.960 108.885 173.130 ;
        RECT 109.175 172.960 109.345 173.130 ;
        RECT 110.095 172.960 110.265 173.130 ;
        RECT 110.555 172.960 110.725 173.130 ;
        RECT 111.015 172.960 111.185 173.130 ;
        RECT 111.475 172.960 111.645 173.130 ;
        RECT 111.935 172.960 112.105 173.130 ;
        RECT 112.395 172.960 112.565 173.130 ;
        RECT 112.855 172.960 113.025 173.130 ;
        RECT 113.315 172.960 113.485 173.130 ;
        RECT 113.775 172.960 113.945 173.130 ;
        RECT 114.235 172.960 114.405 173.130 ;
        RECT 114.695 172.960 114.865 173.130 ;
        RECT 115.155 172.960 115.325 173.130 ;
        RECT 115.615 172.960 115.785 173.130 ;
        RECT 116.075 172.960 116.245 173.130 ;
        RECT 116.535 172.960 116.705 173.130 ;
        RECT 116.995 172.960 117.165 173.130 ;
        RECT 117.455 172.960 117.625 173.130 ;
        RECT 113.145 171.705 113.315 171.875 ;
        RECT 45.125 170.550 45.295 170.720 ;
        RECT 94.020 170.430 94.190 170.600 ;
        RECT 196.225 170.550 196.395 170.720 ;
        RECT 43.915 169.295 44.085 169.465 ;
        RECT 44.375 169.295 44.545 169.465 ;
        RECT 44.835 169.295 45.005 169.465 ;
        RECT 45.295 169.295 45.465 169.465 ;
        RECT 45.755 169.295 45.925 169.465 ;
        RECT 46.215 169.295 46.385 169.465 ;
        RECT 46.675 169.295 46.845 169.465 ;
        RECT 92.810 169.175 92.980 169.345 ;
        RECT 93.270 169.175 93.440 169.345 ;
        RECT 93.730 169.175 93.900 169.345 ;
        RECT 94.190 169.175 94.360 169.345 ;
        RECT 94.650 169.175 94.820 169.345 ;
        RECT 95.110 169.175 95.280 169.345 ;
        RECT 95.570 169.175 95.740 169.345 ;
        RECT 194.675 169.295 194.845 169.465 ;
        RECT 195.135 169.295 195.305 169.465 ;
        RECT 195.595 169.295 195.765 169.465 ;
        RECT 196.055 169.295 196.225 169.465 ;
        RECT 196.515 169.295 196.685 169.465 ;
        RECT 196.975 169.295 197.145 169.465 ;
        RECT 197.435 169.295 197.605 169.465 ;
        RECT 47.325 167.295 47.495 167.465 ;
        RECT 47.685 167.400 47.855 167.570 ;
        RECT 48.550 167.400 48.720 167.570 ;
        RECT 49.415 167.400 49.585 167.570 ;
        RECT 50.280 167.400 50.450 167.570 ;
        RECT 51.145 167.400 51.315 167.570 ;
        RECT 52.010 167.400 52.180 167.570 ;
        RECT 52.875 167.400 53.045 167.570 ;
        RECT 53.740 167.400 53.910 167.570 ;
        RECT 54.605 167.400 54.775 167.570 ;
        RECT 54.995 167.325 55.165 167.495 ;
        RECT 96.220 167.175 96.390 167.345 ;
        RECT 96.580 167.280 96.750 167.450 ;
        RECT 97.445 167.280 97.615 167.450 ;
        RECT 98.310 167.280 98.480 167.450 ;
        RECT 99.175 167.280 99.345 167.450 ;
        RECT 100.040 167.280 100.210 167.450 ;
        RECT 100.905 167.280 101.075 167.450 ;
        RECT 101.770 167.280 101.940 167.450 ;
        RECT 102.635 167.280 102.805 167.450 ;
        RECT 105.495 167.520 105.665 167.690 ;
        RECT 105.955 167.520 106.125 167.690 ;
        RECT 106.415 167.520 106.585 167.690 ;
        RECT 106.875 167.520 107.045 167.690 ;
        RECT 107.335 167.520 107.505 167.690 ;
        RECT 107.795 167.520 107.965 167.690 ;
        RECT 108.255 167.520 108.425 167.690 ;
        RECT 108.715 167.520 108.885 167.690 ;
        RECT 109.175 167.520 109.345 167.690 ;
        RECT 110.095 167.520 110.265 167.690 ;
        RECT 110.555 167.520 110.725 167.690 ;
        RECT 111.015 167.520 111.185 167.690 ;
        RECT 111.475 167.520 111.645 167.690 ;
        RECT 111.935 167.520 112.105 167.690 ;
        RECT 112.395 167.520 112.565 167.690 ;
        RECT 112.855 167.520 113.025 167.690 ;
        RECT 113.315 167.520 113.485 167.690 ;
        RECT 113.775 167.520 113.945 167.690 ;
        RECT 114.235 167.520 114.405 167.690 ;
        RECT 114.695 167.520 114.865 167.690 ;
        RECT 115.155 167.520 115.325 167.690 ;
        RECT 115.615 167.520 115.785 167.690 ;
        RECT 116.075 167.520 116.245 167.690 ;
        RECT 116.535 167.520 116.705 167.690 ;
        RECT 116.995 167.520 117.165 167.690 ;
        RECT 117.455 167.520 117.625 167.690 ;
        RECT 126.300 167.640 126.555 167.890 ;
        RECT 103.500 167.280 103.670 167.450 ;
        RECT 103.890 167.205 104.060 167.375 ;
        RECT 49.895 166.575 50.075 166.745 ;
        RECT 50.355 166.575 50.525 166.745 ;
        RECT 50.815 166.575 50.985 166.745 ;
        RECT 51.275 166.575 51.445 166.745 ;
        RECT 51.735 166.575 51.905 166.745 ;
        RECT 52.195 166.575 52.365 166.745 ;
        RECT 52.655 166.575 52.825 166.745 ;
        RECT 53.115 166.575 53.285 166.745 ;
        RECT 53.575 166.575 53.745 166.745 ;
        RECT 54.035 166.575 54.205 166.745 ;
        RECT 54.495 166.575 54.665 166.745 ;
        RECT 54.955 166.575 55.125 166.745 ;
        RECT 55.415 166.575 55.585 166.745 ;
        RECT 98.790 166.455 98.970 166.625 ;
        RECT 99.250 166.455 99.420 166.625 ;
        RECT 99.710 166.455 99.880 166.625 ;
        RECT 100.170 166.455 100.340 166.625 ;
        RECT 100.630 166.455 100.800 166.625 ;
        RECT 101.090 166.455 101.260 166.625 ;
        RECT 101.550 166.455 101.720 166.625 ;
        RECT 102.010 166.455 102.180 166.625 ;
        RECT 102.470 166.455 102.640 166.625 ;
        RECT 102.930 166.455 103.100 166.625 ;
        RECT 103.390 166.455 103.560 166.625 ;
        RECT 103.850 166.455 104.020 166.625 ;
        RECT 104.310 166.455 104.480 166.625 ;
        RECT 96.220 165.735 96.390 165.905 ;
        RECT 96.580 165.630 96.750 165.800 ;
        RECT 97.445 165.630 97.615 165.800 ;
        RECT 98.310 165.630 98.480 165.800 ;
        RECT 99.175 165.630 99.345 165.800 ;
        RECT 100.040 165.630 100.210 165.800 ;
        RECT 100.905 165.630 101.075 165.800 ;
        RECT 101.770 165.630 101.940 165.800 ;
        RECT 102.635 165.630 102.805 165.800 ;
        RECT 103.500 165.630 103.670 165.800 ;
        RECT 103.890 165.705 104.060 165.875 ;
        RECT 121.610 167.425 121.780 167.595 ;
        RECT 122.070 167.425 122.240 167.595 ;
        RECT 122.530 167.425 122.700 167.595 ;
        RECT 122.990 167.425 123.160 167.595 ;
        RECT 123.450 167.425 123.620 167.595 ;
        RECT 123.910 167.425 124.080 167.595 ;
        RECT 124.370 167.425 124.540 167.595 ;
        RECT 124.830 167.425 125.000 167.595 ;
        RECT 125.290 167.425 125.460 167.595 ;
        RECT 127.400 167.425 127.570 167.595 ;
        RECT 127.860 167.425 128.030 167.595 ;
        RECT 128.320 167.425 128.490 167.595 ;
        RECT 128.780 167.425 128.950 167.595 ;
        RECT 129.240 167.425 129.410 167.595 ;
        RECT 129.700 167.425 129.870 167.595 ;
        RECT 130.160 167.425 130.330 167.595 ;
        RECT 130.620 167.425 130.790 167.595 ;
        RECT 131.080 167.425 131.250 167.595 ;
        RECT 126.300 167.130 126.555 167.380 ;
        RECT 186.355 167.325 186.525 167.495 ;
        RECT 186.745 167.400 186.915 167.570 ;
        RECT 187.610 167.400 187.780 167.570 ;
        RECT 188.475 167.400 188.645 167.570 ;
        RECT 189.340 167.400 189.510 167.570 ;
        RECT 190.205 167.400 190.375 167.570 ;
        RECT 191.070 167.400 191.240 167.570 ;
        RECT 191.935 167.400 192.105 167.570 ;
        RECT 192.800 167.400 192.970 167.570 ;
        RECT 193.665 167.400 193.835 167.570 ;
        RECT 194.025 167.295 194.195 167.465 ;
        RECT 185.935 166.575 186.105 166.745 ;
        RECT 186.395 166.575 186.565 166.745 ;
        RECT 186.855 166.575 187.025 166.745 ;
        RECT 187.315 166.575 187.485 166.745 ;
        RECT 187.775 166.575 187.945 166.745 ;
        RECT 188.235 166.575 188.405 166.745 ;
        RECT 188.695 166.575 188.865 166.745 ;
        RECT 189.155 166.575 189.325 166.745 ;
        RECT 189.615 166.575 189.785 166.745 ;
        RECT 190.075 166.575 190.245 166.745 ;
        RECT 190.535 166.575 190.705 166.745 ;
        RECT 190.995 166.575 191.165 166.745 ;
        RECT 191.445 166.575 191.625 166.745 ;
        RECT 113.145 166.265 113.315 166.435 ;
        RECT 92.810 163.735 92.980 163.905 ;
        RECT 93.270 163.735 93.440 163.905 ;
        RECT 93.730 163.735 93.900 163.905 ;
        RECT 94.190 163.735 94.360 163.905 ;
        RECT 94.650 163.735 94.820 163.905 ;
        RECT 95.110 163.735 95.280 163.905 ;
        RECT 95.570 163.735 95.740 163.905 ;
        RECT 94.020 162.480 94.190 162.650 ;
        RECT 105.495 162.080 105.665 162.250 ;
        RECT 105.955 162.080 106.125 162.250 ;
        RECT 106.415 162.080 106.585 162.250 ;
        RECT 106.875 162.080 107.045 162.250 ;
        RECT 107.335 162.080 107.505 162.250 ;
        RECT 107.795 162.080 107.965 162.250 ;
        RECT 108.255 162.080 108.425 162.250 ;
        RECT 108.715 162.080 108.885 162.250 ;
        RECT 109.175 162.080 109.345 162.250 ;
        RECT 109.635 162.080 109.805 162.250 ;
        RECT 110.095 162.080 110.265 162.250 ;
        RECT 110.555 162.080 110.725 162.250 ;
        RECT 111.015 162.080 111.185 162.250 ;
        RECT 111.475 162.080 111.645 162.250 ;
        RECT 111.935 162.080 112.105 162.250 ;
        RECT 112.395 162.080 112.565 162.250 ;
        RECT 112.855 162.080 113.025 162.250 ;
        RECT 113.315 162.080 113.485 162.250 ;
        RECT 113.775 162.080 113.945 162.250 ;
        RECT 114.235 162.080 114.405 162.250 ;
        RECT 114.695 162.080 114.865 162.250 ;
        RECT 115.155 162.080 115.325 162.250 ;
        RECT 115.615 162.080 115.785 162.250 ;
        RECT 116.075 162.080 116.245 162.250 ;
        RECT 116.535 162.080 116.705 162.250 ;
        RECT 116.995 162.080 117.165 162.250 ;
        RECT 117.455 162.080 117.625 162.250 ;
        RECT 113.145 160.825 113.315 160.995 ;
        RECT 116.910 134.300 117.250 134.470 ;
        RECT 123.190 134.300 123.530 134.470 ;
        RECT 5.155 132.575 5.325 132.745 ;
        RECT 235.055 132.575 235.225 132.745 ;
        RECT 112.000 131.115 112.170 131.405 ;
        RECT 113.160 131.115 113.330 131.405 ;
        RECT 114.320 131.115 114.490 131.405 ;
        RECT 115.480 131.115 115.650 131.405 ;
        RECT 124.790 131.115 124.960 131.405 ;
        RECT 125.950 131.115 126.120 131.405 ;
        RECT 127.110 131.115 127.280 131.405 ;
        RECT 128.270 131.115 128.440 131.405 ;
        RECT 115.970 129.745 116.140 129.915 ;
        RECT 116.910 129.735 117.250 129.905 ;
        RECT 123.190 129.735 123.530 129.905 ;
        RECT 124.300 129.740 124.470 129.910 ;
        RECT 120.050 125.535 120.390 125.705 ;
      LAYER met1 ;
        RECT 105.500 173.285 105.780 173.465 ;
        RECT 105.350 172.805 117.770 173.285 ;
        RECT 113.045 171.935 113.240 172.805 ;
        RECT 113.045 171.645 113.365 171.935 ;
        RECT 45.055 170.735 45.345 170.780 ;
        RECT 43.895 170.535 45.345 170.735 ;
        RECT 196.175 170.735 196.465 170.780 ;
        RECT 93.950 170.615 94.240 170.660 ;
        RECT 43.895 169.650 44.115 170.535 ;
        RECT 45.055 170.490 45.345 170.535 ;
        RECT 43.210 169.620 44.115 169.650 ;
        RECT 92.790 170.415 94.240 170.615 ;
        RECT 196.175 170.535 197.625 170.735 ;
        RECT 196.175 170.490 196.465 170.535 ;
        RECT 43.210 169.140 46.990 169.620 ;
        RECT 92.790 169.500 93.010 170.415 ;
        RECT 93.950 170.370 94.240 170.415 ;
        RECT 197.405 169.650 197.625 170.535 ;
        RECT 197.405 169.620 198.310 169.650 ;
        RECT 92.665 169.460 95.885 169.500 ;
        RECT 96.190 169.460 96.350 169.500 ;
        RECT 43.210 169.110 44.060 169.140 ;
        RECT 92.665 169.050 96.350 169.460 ;
        RECT 194.530 169.140 198.310 169.620 ;
        RECT 197.460 169.110 198.310 169.140 ;
        RECT 92.665 169.020 95.885 169.050 ;
        RECT 47.295 167.450 55.195 167.600 ;
        RECT 47.295 167.445 52.240 167.450 ;
        RECT 47.295 167.440 49.645 167.445 ;
        RECT 47.295 167.370 47.915 167.440 ;
        RECT 48.490 167.370 48.780 167.440 ;
        RECT 49.355 167.370 49.645 167.440 ;
        RECT 50.220 167.440 52.240 167.445 ;
        RECT 50.220 167.370 50.510 167.440 ;
        RECT 51.085 167.370 51.375 167.440 ;
        RECT 51.950 167.370 52.240 167.440 ;
        RECT 52.815 167.440 55.195 167.450 ;
        RECT 52.815 167.400 53.105 167.440 ;
        RECT 52.835 167.370 53.105 167.400 ;
        RECT 53.680 167.370 53.970 167.440 ;
        RECT 54.545 167.370 55.195 167.440 ;
        RECT 47.295 167.235 47.545 167.370 ;
        RECT 51.145 166.900 51.315 167.370 ;
        RECT 54.955 167.265 55.195 167.370 ;
        RECT 96.190 167.480 96.350 169.050 ;
        RECT 105.530 167.845 105.810 167.950 ;
        RECT 105.270 167.790 117.770 167.845 ;
        RECT 105.270 167.750 121.675 167.790 ;
        RECT 126.245 167.750 126.600 167.985 ;
        RECT 96.190 167.330 104.090 167.480 ;
        RECT 96.190 167.325 101.135 167.330 ;
        RECT 96.190 167.320 98.540 167.325 ;
        RECT 96.190 167.250 96.810 167.320 ;
        RECT 97.385 167.250 97.675 167.320 ;
        RECT 98.250 167.250 98.540 167.320 ;
        RECT 99.115 167.320 101.135 167.325 ;
        RECT 99.115 167.250 99.405 167.320 ;
        RECT 99.980 167.250 100.270 167.320 ;
        RECT 100.845 167.250 101.135 167.320 ;
        RECT 101.710 167.320 104.090 167.330 ;
        RECT 101.710 167.280 102.000 167.320 ;
        RECT 101.730 167.250 102.000 167.280 ;
        RECT 102.575 167.250 102.865 167.320 ;
        RECT 103.440 167.250 104.090 167.320 ;
        RECT 96.190 167.115 96.440 167.250 ;
        RECT 49.615 166.420 55.730 166.900 ;
        RECT 100.040 166.780 100.210 167.250 ;
        RECT 103.850 167.145 104.090 167.250 ;
        RECT 105.270 167.395 131.395 167.750 ;
        RECT 105.270 167.365 117.770 167.395 ;
        RECT 105.270 166.780 105.800 167.365 ;
        RECT 97.510 166.300 105.800 166.780 ;
        RECT 113.045 166.495 113.240 167.365 ;
        RECT 121.465 167.270 131.395 167.395 ;
        RECT 186.325 167.450 194.225 167.600 ;
        RECT 186.325 167.440 188.705 167.450 ;
        RECT 186.325 167.370 186.975 167.440 ;
        RECT 187.550 167.370 187.840 167.440 ;
        RECT 188.415 167.400 188.705 167.440 ;
        RECT 189.280 167.445 194.225 167.450 ;
        RECT 189.280 167.440 191.300 167.445 ;
        RECT 188.415 167.370 188.685 167.400 ;
        RECT 189.280 167.370 189.570 167.440 ;
        RECT 190.145 167.370 190.435 167.440 ;
        RECT 191.010 167.370 191.300 167.440 ;
        RECT 191.875 167.440 194.225 167.445 ;
        RECT 191.875 167.370 192.165 167.440 ;
        RECT 192.740 167.370 193.030 167.440 ;
        RECT 193.605 167.370 194.225 167.440 ;
        RECT 126.245 167.035 126.600 167.270 ;
        RECT 186.325 167.265 186.565 167.370 ;
        RECT 190.205 166.900 190.375 167.370 ;
        RECT 193.975 167.235 194.225 167.370 ;
        RECT 96.190 165.830 96.440 165.965 ;
        RECT 100.040 165.830 100.210 166.300 ;
        RECT 113.045 166.205 113.365 166.495 ;
        RECT 185.790 166.420 191.905 166.900 ;
        RECT 103.850 165.830 104.090 165.935 ;
        RECT 96.190 165.760 96.810 165.830 ;
        RECT 97.385 165.760 97.675 165.830 ;
        RECT 98.250 165.760 98.540 165.830 ;
        RECT 96.190 165.755 98.540 165.760 ;
        RECT 99.115 165.760 99.405 165.830 ;
        RECT 99.980 165.760 100.270 165.830 ;
        RECT 100.845 165.760 101.135 165.830 ;
        RECT 101.730 165.800 102.000 165.830 ;
        RECT 99.115 165.755 101.135 165.760 ;
        RECT 96.190 165.750 101.135 165.755 ;
        RECT 101.710 165.760 102.000 165.800 ;
        RECT 102.575 165.760 102.865 165.830 ;
        RECT 103.440 165.760 104.090 165.830 ;
        RECT 101.710 165.750 104.090 165.760 ;
        RECT 96.190 165.600 104.090 165.750 ;
        RECT 92.665 163.580 95.885 164.060 ;
        RECT 92.790 162.665 93.010 163.580 ;
        RECT 93.950 162.665 94.240 162.710 ;
        RECT 92.790 162.465 94.240 162.665 ;
        RECT 93.950 162.420 94.240 162.465 ;
        RECT 105.555 162.405 105.835 162.545 ;
        RECT 105.350 161.925 117.770 162.405 ;
        RECT 113.045 161.055 113.240 161.925 ;
        RECT 113.045 160.765 113.365 161.055 ;
        RECT 116.950 142.200 117.210 142.265 ;
        RECT 123.225 142.200 123.485 142.295 ;
        RECT 111.030 142.030 129.355 142.200 ;
        RECT 116.950 141.945 117.210 142.030 ;
        RECT 123.225 141.975 123.485 142.030 ;
        RECT 116.880 134.470 117.280 134.515 ;
        RECT 123.160 134.470 123.560 134.515 ;
        RECT 116.850 134.300 117.310 134.470 ;
        RECT 123.130 134.300 123.590 134.470 ;
        RECT 116.880 134.255 117.280 134.300 ;
        RECT 123.160 134.255 123.560 134.300 ;
        RECT 5.090 132.745 5.365 132.785 ;
        RECT 5.895 132.745 6.235 133.260 ;
        RECT 5.090 132.575 6.235 132.745 ;
        RECT 5.090 132.535 5.365 132.575 ;
        RECT 5.895 128.715 6.235 132.575 ;
        RECT 234.145 132.745 234.485 133.260 ;
        RECT 235.015 132.745 235.290 132.785 ;
        RECT 234.145 132.575 235.290 132.745 ;
        RECT 111.940 131.025 112.230 131.445 ;
        RECT 113.100 131.025 113.390 131.445 ;
        RECT 114.260 131.025 114.550 131.445 ;
        RECT 115.420 131.025 115.710 131.445 ;
        RECT 124.730 131.025 125.020 131.445 ;
        RECT 125.890 131.025 126.180 131.445 ;
        RECT 127.050 131.025 127.340 131.445 ;
        RECT 128.210 131.025 128.500 131.445 ;
        RECT 111.930 130.915 112.250 131.025 ;
        RECT 113.090 130.915 113.410 131.025 ;
        RECT 114.250 130.915 114.570 131.025 ;
        RECT 115.410 130.915 115.730 131.025 ;
        RECT 111.885 130.880 115.730 130.915 ;
        RECT 124.710 130.895 125.030 131.025 ;
        RECT 125.870 130.895 126.190 131.025 ;
        RECT 127.030 130.895 127.350 131.025 ;
        RECT 128.190 130.895 128.510 131.025 ;
        RECT 124.710 130.880 128.750 130.895 ;
        RECT 111.885 130.725 116.140 130.880 ;
        RECT 115.970 129.960 116.140 130.725 ;
        RECT 124.300 130.725 128.750 130.880 ;
        RECT 124.300 129.960 124.470 130.725 ;
        RECT 115.910 129.695 116.200 129.960 ;
        RECT 9.645 128.925 9.965 129.215 ;
        RECT 18.625 128.925 18.945 129.215 ;
        RECT 30.945 128.925 31.265 129.215 ;
        RECT 36.475 128.925 36.795 129.215 ;
        RECT 68.395 128.925 68.715 129.215 ;
        RECT 75.165 128.925 75.485 129.215 ;
        RECT 99.445 128.925 99.765 129.215 ;
        RECT 105.925 128.925 106.245 129.215 ;
        RECT 9.705 128.715 9.910 128.925 ;
        RECT 5.895 128.515 9.910 128.715 ;
        RECT 115.970 125.720 116.140 129.695 ;
        RECT 116.850 129.690 117.310 129.950 ;
        RECT 123.130 129.690 123.590 129.950 ;
        RECT 124.240 129.695 124.530 129.960 ;
        RECT 120.020 125.720 120.420 125.735 ;
        RECT 124.300 125.720 124.470 129.695 ;
        RECT 134.135 128.925 134.455 129.215 ;
        RECT 140.615 128.925 140.935 129.215 ;
        RECT 164.895 128.925 165.215 129.215 ;
        RECT 171.665 128.925 171.985 129.215 ;
        RECT 203.585 128.925 203.905 129.215 ;
        RECT 209.115 128.925 209.435 129.215 ;
        RECT 221.435 128.925 221.755 129.215 ;
        RECT 230.415 128.925 230.735 129.215 ;
        RECT 230.470 128.715 230.675 128.925 ;
        RECT 234.145 128.715 234.485 132.575 ;
        RECT 235.015 132.535 235.290 132.575 ;
        RECT 230.470 128.515 234.485 128.715 ;
        RECT 115.970 125.530 124.470 125.720 ;
        RECT 120.020 125.505 120.420 125.530 ;
      LAYER via ;
        RECT 105.510 173.150 105.770 173.410 ;
        RECT 110.045 172.930 110.305 173.190 ;
        RECT 114.775 172.925 115.035 173.185 ;
        RECT 95.520 169.125 95.780 169.385 ;
        RECT 197.460 169.140 198.310 169.620 ;
        RECT 105.540 167.635 105.800 167.895 ;
        RECT 110.180 167.485 110.440 167.745 ;
        RECT 114.785 167.485 115.045 167.745 ;
        RECT 53.380 166.460 54.540 166.850 ;
        RECT 186.980 166.460 188.140 166.850 ;
        RECT 95.535 163.710 95.795 163.970 ;
        RECT 105.565 162.230 105.825 162.490 ;
        RECT 110.165 162.040 110.425 162.300 ;
        RECT 114.775 162.040 115.035 162.300 ;
        RECT 116.950 141.975 117.210 142.235 ;
        RECT 123.225 142.005 123.485 142.265 ;
        RECT 116.910 134.255 117.250 134.515 ;
        RECT 123.190 134.255 123.530 134.515 ;
        RECT 5.940 132.845 6.200 133.105 ;
        RECT 234.180 132.845 234.440 133.105 ;
        RECT 9.675 128.935 9.935 129.195 ;
        RECT 18.655 128.935 18.915 129.195 ;
        RECT 30.975 128.935 31.235 129.195 ;
        RECT 36.505 128.935 36.765 129.195 ;
        RECT 68.425 128.935 68.685 129.195 ;
        RECT 75.195 128.935 75.455 129.195 ;
        RECT 99.475 128.935 99.735 129.195 ;
        RECT 105.955 128.935 106.215 129.195 ;
        RECT 116.910 129.690 117.250 129.950 ;
        RECT 123.190 129.690 123.530 129.950 ;
        RECT 134.165 128.935 134.425 129.195 ;
        RECT 140.645 128.935 140.905 129.195 ;
        RECT 164.925 128.935 165.185 129.195 ;
        RECT 171.695 128.935 171.955 129.195 ;
        RECT 203.615 128.935 203.875 129.195 ;
        RECT 209.145 128.935 209.405 129.195 ;
        RECT 221.465 128.935 221.725 129.195 ;
        RECT 230.445 128.935 230.705 129.195 ;
      LAYER met2 ;
        RECT 105.500 173.095 105.780 173.465 ;
        RECT 110.035 172.875 110.315 173.245 ;
        RECT 114.765 172.870 115.045 173.240 ;
        RECT 43.210 148.290 44.060 169.650 ;
        RECT 95.510 169.070 95.790 169.440 ;
        RECT 105.530 167.580 105.810 167.950 ;
        RECT 110.170 167.430 110.450 167.800 ;
        RECT 114.775 167.430 115.055 167.800 ;
        RECT 5.930 147.845 6.210 148.215 ;
        RECT 5.940 132.815 6.200 147.845 ;
        RECT 43.000 147.700 44.260 148.290 ;
        RECT 53.380 148.280 54.540 166.900 ;
        RECT 97.510 166.300 98.250 166.780 ;
        RECT 95.525 163.655 95.805 164.025 ;
        RECT 105.555 162.175 105.835 162.545 ;
        RECT 110.155 161.985 110.435 162.355 ;
        RECT 114.765 161.985 115.045 162.355 ;
        RECT 186.980 148.280 188.140 166.900 ;
        RECT 197.460 148.290 198.310 169.650 ;
        RECT 53.330 147.700 54.590 148.280 ;
        RECT 116.950 148.205 117.210 148.220 ;
        RECT 123.170 148.205 123.430 148.220 ;
        RECT 116.940 147.835 117.220 148.205 ;
        RECT 123.160 147.835 123.440 148.205 ;
        RECT 116.950 141.945 117.210 147.835 ;
        RECT 123.170 142.295 123.430 147.835 ;
        RECT 186.930 147.700 188.190 148.280 ;
        RECT 197.260 147.700 198.520 148.290 ;
        RECT 234.170 147.845 234.450 148.215 ;
        RECT 123.170 141.975 123.485 142.295 ;
        RECT 117.000 134.515 117.170 141.945 ;
        RECT 123.280 134.515 123.450 141.975 ;
        RECT 116.880 134.255 117.280 134.515 ;
        RECT 123.160 134.255 123.560 134.515 ;
        RECT 117.000 129.980 117.160 134.255 ;
        RECT 123.280 129.980 123.440 134.255 ;
        RECT 234.180 132.815 234.440 147.845 ;
        RECT 116.910 129.660 117.250 129.980 ;
        RECT 123.190 129.660 123.530 129.980 ;
        RECT 9.675 129.210 9.935 129.225 ;
        RECT 18.655 129.215 18.915 129.225 ;
        RECT 9.625 128.930 9.995 129.210 ;
        RECT 9.675 128.905 9.935 128.930 ;
        RECT 18.595 128.910 18.985 129.215 ;
        RECT 18.655 128.905 18.915 128.910 ;
        RECT 30.965 128.880 31.245 129.250 ;
        RECT 36.495 128.880 36.775 129.250 ;
        RECT 68.410 128.870 68.695 129.250 ;
        RECT 75.180 128.880 75.465 129.255 ;
        RECT 99.440 128.875 99.745 129.260 ;
        RECT 105.945 128.880 106.230 129.250 ;
        RECT 134.150 128.880 134.435 129.250 ;
        RECT 140.635 128.875 140.940 129.260 ;
        RECT 164.915 128.880 165.200 129.255 ;
        RECT 171.685 128.870 171.970 129.250 ;
        RECT 203.605 128.880 203.885 129.250 ;
        RECT 209.135 128.880 209.415 129.250 ;
        RECT 221.465 129.215 221.725 129.225 ;
        RECT 221.395 128.910 221.785 129.215 ;
        RECT 230.445 129.210 230.705 129.225 ;
        RECT 230.385 128.930 230.755 129.210 ;
        RECT 221.465 128.905 221.725 128.910 ;
        RECT 230.445 128.905 230.705 128.930 ;
      LAYER via2 ;
        RECT 105.500 173.140 105.780 173.420 ;
        RECT 110.035 172.920 110.315 173.200 ;
        RECT 114.765 172.915 115.045 173.195 ;
        RECT 95.510 169.115 95.790 169.395 ;
        RECT 105.530 167.625 105.810 167.905 ;
        RECT 110.170 167.475 110.450 167.755 ;
        RECT 114.775 167.475 115.055 167.755 ;
        RECT 97.540 166.355 98.200 166.725 ;
        RECT 95.525 163.700 95.805 163.980 ;
        RECT 105.555 162.220 105.835 162.500 ;
        RECT 110.155 162.030 110.435 162.310 ;
        RECT 114.765 162.030 115.045 162.310 ;
        RECT 5.930 147.890 6.210 148.170 ;
        RECT 43.050 147.750 44.210 148.240 ;
        RECT 53.380 147.750 54.540 148.240 ;
        RECT 116.940 147.880 117.220 148.160 ;
        RECT 123.160 147.880 123.440 148.160 ;
        RECT 186.980 147.750 188.140 148.240 ;
        RECT 197.310 147.750 198.470 148.240 ;
        RECT 234.170 147.890 234.450 148.170 ;
        RECT 9.670 128.930 9.950 129.210 ;
        RECT 18.640 128.910 18.940 129.215 ;
        RECT 30.965 128.925 31.245 129.205 ;
        RECT 36.495 128.925 36.775 129.205 ;
        RECT 68.410 128.915 68.695 129.205 ;
        RECT 75.180 128.925 75.465 129.210 ;
        RECT 99.440 128.920 99.745 129.215 ;
        RECT 105.945 128.925 106.230 129.205 ;
        RECT 134.150 128.925 134.435 129.205 ;
        RECT 140.635 128.920 140.940 129.215 ;
        RECT 164.915 128.925 165.200 129.210 ;
        RECT 171.685 128.915 171.970 129.205 ;
        RECT 203.605 128.925 203.885 129.205 ;
        RECT 209.135 128.925 209.415 129.205 ;
        RECT 221.440 128.910 221.740 129.215 ;
        RECT 230.430 128.930 230.710 129.210 ;
      LAYER met3 ;
        RECT 105.400 173.040 105.890 173.530 ;
        RECT 109.935 172.820 110.425 173.310 ;
        RECT 114.665 172.815 115.155 173.305 ;
        RECT 95.405 169.000 95.895 169.490 ;
        RECT 105.430 167.525 105.920 168.015 ;
        RECT 110.070 167.375 110.560 167.865 ;
        RECT 114.675 167.375 115.165 167.865 ;
        RECT 97.510 166.300 98.250 166.780 ;
        RECT 95.420 163.585 95.910 164.075 ;
        RECT 105.455 162.120 105.945 162.610 ;
        RECT 110.055 161.930 110.545 162.420 ;
        RECT 114.665 161.930 115.155 162.420 ;
        RECT 43.000 148.245 44.260 148.290 ;
        RECT 53.330 148.245 54.590 148.280 ;
        RECT 186.930 148.245 188.190 148.280 ;
        RECT 197.260 148.245 198.520 148.290 ;
        RECT -0.130 147.745 253.790 148.245 ;
        RECT 43.000 147.700 44.260 147.745 ;
        RECT 53.330 147.700 54.590 147.745 ;
        RECT 186.930 147.700 188.190 147.745 ;
        RECT 197.260 147.700 198.520 147.745 ;
        RECT 10.725 130.610 17.705 136.890 ;
        RECT 13.485 129.235 15.455 130.610 ;
        RECT 32.040 130.560 35.720 133.840 ;
        RECT 69.895 130.575 74.175 135.855 ;
        RECT 33.285 129.300 34.210 130.560 ;
        RECT 30.900 129.240 34.210 129.300 ;
        RECT 18.595 129.235 19.000 129.240 ;
        RECT 9.605 128.890 19.000 129.235 ;
        RECT 1.860 127.250 3.460 128.375 ;
        RECT 0.560 125.650 3.460 127.250 ;
        RECT 5.060 127.250 6.660 128.410 ;
        RECT 5.060 125.650 7.960 127.250 ;
        RECT 1.860 124.050 6.660 125.650 ;
        RECT 0.560 122.450 3.460 124.050 ;
        RECT 5.060 122.450 7.960 124.050 ;
        RECT 13.485 122.470 15.455 128.890 ;
        RECT 18.595 128.885 19.000 128.890 ;
        RECT 30.900 128.875 36.820 129.240 ;
        RECT 30.900 128.755 34.210 128.875 ;
        RECT 33.285 122.470 34.210 128.755 ;
        RECT 68.350 127.865 68.775 129.255 ;
        RECT 71.815 127.890 73.185 130.575 ;
        RECT 100.905 130.470 104.585 133.750 ;
        RECT 135.795 130.470 139.475 133.750 ;
        RECT 166.205 130.575 170.485 135.855 ;
        RECT 75.080 127.890 75.525 129.280 ;
        RECT 102.230 129.270 102.740 130.470 ;
        RECT 99.370 129.265 102.740 129.270 ;
        RECT 137.640 129.270 138.150 130.470 ;
        RECT 137.640 129.265 141.010 129.270 ;
        RECT 99.370 128.875 106.315 129.265 ;
        RECT 134.065 128.875 141.010 129.265 ;
        RECT 71.815 127.865 75.530 127.890 ;
        RECT 68.350 127.560 75.530 127.865 ;
        RECT 68.350 127.520 73.185 127.560 ;
        RECT 71.815 122.470 73.185 127.520 ;
        RECT 99.370 122.470 99.915 128.875 ;
        RECT 140.465 122.470 141.010 128.875 ;
        RECT 164.855 127.890 165.300 129.280 ;
        RECT 167.195 127.890 168.565 130.575 ;
        RECT 204.660 130.560 208.340 133.840 ;
        RECT 222.675 130.610 229.655 136.890 ;
        RECT 206.170 129.300 207.095 130.560 ;
        RECT 164.850 127.865 168.565 127.890 ;
        RECT 171.605 127.865 172.030 129.255 ;
        RECT 206.170 129.240 209.480 129.300 ;
        RECT 203.560 128.875 209.480 129.240 ;
        RECT 221.380 129.235 221.785 129.240 ;
        RECT 224.925 129.235 226.895 130.610 ;
        RECT 221.380 128.890 230.775 129.235 ;
        RECT 221.380 128.885 221.785 128.890 ;
        RECT 164.850 127.560 172.030 127.865 ;
        RECT 167.195 127.520 172.030 127.560 ;
        RECT 206.170 128.755 209.480 128.875 ;
        RECT 167.195 122.470 168.565 127.520 ;
        RECT 206.170 122.470 207.095 128.755 ;
        RECT 224.925 122.470 226.895 128.890 ;
        RECT 233.720 127.250 235.320 128.410 ;
        RECT 232.420 125.650 235.320 127.250 ;
        RECT 236.920 127.250 238.520 128.375 ;
        RECT 236.920 125.650 239.820 127.250 ;
        RECT 233.720 124.050 238.520 125.650 ;
        RECT 1.860 120.850 6.660 122.450 ;
        RECT 10.180 121.790 67.940 122.470 ;
        RECT 69.520 121.790 100.080 122.470 ;
        RECT 10.180 120.860 100.080 121.790 ;
        RECT 0.560 119.250 3.460 120.850 ;
        RECT 5.060 119.250 7.960 120.850 ;
        RECT 10.180 119.250 11.790 120.860 ;
        RECT 13.800 119.250 15.400 120.860 ;
        RECT 18.065 119.250 19.670 120.860 ;
        RECT 22.330 119.250 23.930 120.860 ;
        RECT 1.860 117.650 6.660 119.250 ;
        RECT 10.180 119.130 23.930 119.250 ;
        RECT 26.990 119.250 28.590 120.860 ;
        RECT 31.460 119.250 33.060 120.860 ;
        RECT 35.930 119.250 37.530 120.860 ;
        RECT 26.990 119.130 37.530 119.250 ;
        RECT 40.590 119.250 42.190 120.860 ;
        RECT 45.060 119.250 46.660 120.860 ;
        RECT 49.530 119.250 51.130 120.860 ;
        RECT 40.590 119.130 51.130 119.250 ;
        RECT 54.190 119.250 55.790 120.860 ;
        RECT 58.655 119.250 60.255 120.860 ;
        RECT 63.120 119.250 64.720 120.860 ;
        RECT 54.190 119.130 64.720 119.250 ;
        RECT 10.180 118.850 64.720 119.130 ;
        RECT 66.330 120.190 71.130 120.860 ;
        RECT 66.330 118.850 67.940 120.190 ;
        RECT 10.180 117.650 67.940 118.850 ;
        RECT 0.560 116.050 3.460 117.650 ;
        RECT 5.060 116.050 11.790 117.650 ;
        RECT 1.860 114.450 6.660 116.050 ;
        RECT 10.180 114.785 11.790 116.050 ;
        RECT 13.400 117.530 67.940 117.650 ;
        RECT 13.400 114.790 23.920 117.530 ;
        RECT 27.000 114.790 37.520 117.530 ;
        RECT 40.600 114.790 51.120 117.530 ;
        RECT 54.200 117.250 67.940 117.530 ;
        RECT 54.200 114.790 64.720 117.250 ;
        RECT 13.400 114.785 64.720 114.790 ;
        RECT 10.180 114.585 64.720 114.785 ;
        RECT 66.330 114.635 67.940 117.250 ;
        RECT 69.520 119.250 71.130 120.190 ;
        RECT 73.140 119.250 74.740 120.860 ;
        RECT 77.405 119.250 79.010 120.860 ;
        RECT 81.670 119.250 83.270 120.860 ;
        RECT 69.520 119.130 83.270 119.250 ;
        RECT 86.330 119.250 87.930 120.860 ;
        RECT 90.795 119.250 92.395 120.860 ;
        RECT 95.260 119.250 96.860 120.860 ;
        RECT 86.330 119.130 96.860 119.250 ;
        RECT 69.520 118.850 96.860 119.130 ;
        RECT 98.470 118.850 100.080 120.860 ;
        RECT 69.520 117.650 100.080 118.850 ;
        RECT 69.520 114.785 71.130 117.650 ;
        RECT 72.740 117.530 100.080 117.650 ;
        RECT 72.740 114.790 83.260 117.530 ;
        RECT 86.340 117.250 100.080 117.530 ;
        RECT 86.340 114.790 96.860 117.250 ;
        RECT 72.740 114.785 96.860 114.790 ;
        RECT 69.520 114.635 96.860 114.785 ;
        RECT 66.330 114.585 96.860 114.635 ;
        RECT 98.470 114.585 100.080 117.250 ;
        RECT 0.560 112.850 3.460 114.450 ;
        RECT 5.060 112.850 7.960 114.450 ;
        RECT 10.180 113.190 100.080 114.585 ;
        RECT 10.180 113.185 23.920 113.190 ;
        RECT 1.860 111.250 6.660 112.850 ;
        RECT 10.180 111.250 11.790 113.185 ;
        RECT 0.560 109.650 3.460 111.250 ;
        RECT 5.060 110.320 11.790 111.250 ;
        RECT 13.400 110.450 23.920 113.185 ;
        RECT 27.000 110.450 37.520 113.190 ;
        RECT 40.600 110.450 51.120 113.190 ;
        RECT 54.200 113.185 83.260 113.190 ;
        RECT 54.200 113.035 71.130 113.185 ;
        RECT 54.200 112.980 67.940 113.035 ;
        RECT 54.200 110.450 64.720 112.980 ;
        RECT 13.400 110.320 64.720 110.450 ;
        RECT 66.330 110.320 67.940 112.980 ;
        RECT 5.060 109.650 67.940 110.320 ;
        RECT 1.860 108.050 6.660 109.650 ;
        RECT 10.180 109.025 67.940 109.650 ;
        RECT 69.520 110.320 71.130 113.035 ;
        RECT 72.740 110.450 83.260 113.185 ;
        RECT 86.340 112.980 100.080 113.190 ;
        RECT 86.340 110.450 96.860 112.980 ;
        RECT 72.740 110.320 96.860 110.450 ;
        RECT 98.470 110.320 100.080 112.980 ;
        RECT 69.520 109.025 100.080 110.320 ;
        RECT 10.180 108.850 100.080 109.025 ;
        RECT 10.180 108.730 23.930 108.850 ;
        RECT 10.180 108.720 15.120 108.730 ;
        RECT 0.560 106.450 3.460 108.050 ;
        RECT 5.060 106.450 7.960 108.050 ;
        RECT 1.860 104.850 6.660 106.450 ;
        RECT 10.180 105.660 11.790 108.720 ;
        RECT 13.520 105.660 15.120 108.720 ;
        RECT 10.180 105.650 15.120 105.660 ;
        RECT 17.860 105.650 19.460 108.730 ;
        RECT 22.200 108.720 23.930 108.730 ;
        RECT 26.990 108.730 37.530 108.850 ;
        RECT 26.990 108.720 28.720 108.730 ;
        RECT 22.200 105.660 23.800 108.720 ;
        RECT 27.120 105.660 28.720 108.720 ;
        RECT 22.200 105.650 23.930 105.660 ;
        RECT 10.180 105.530 23.930 105.650 ;
        RECT 26.990 105.650 28.720 105.660 ;
        RECT 31.460 105.650 33.060 108.730 ;
        RECT 35.800 108.720 37.530 108.730 ;
        RECT 40.590 108.730 51.130 108.850 ;
        RECT 40.590 108.720 42.320 108.730 ;
        RECT 35.800 105.660 37.400 108.720 ;
        RECT 40.720 105.660 42.320 108.720 ;
        RECT 35.800 105.650 37.530 105.660 ;
        RECT 26.990 105.530 37.530 105.650 ;
        RECT 40.590 105.650 42.320 105.660 ;
        RECT 45.060 105.650 46.660 108.730 ;
        RECT 49.400 108.720 51.130 108.730 ;
        RECT 54.190 108.730 83.270 108.850 ;
        RECT 54.190 108.720 55.920 108.730 ;
        RECT 49.400 105.660 51.000 108.720 ;
        RECT 54.320 105.660 55.920 108.720 ;
        RECT 49.400 105.650 51.130 105.660 ;
        RECT 40.590 105.530 51.130 105.650 ;
        RECT 54.190 105.650 55.920 105.660 ;
        RECT 58.660 105.650 60.260 108.730 ;
        RECT 63.000 108.720 74.460 108.730 ;
        RECT 63.000 105.660 64.600 108.720 ;
        RECT 66.330 107.425 71.130 108.720 ;
        RECT 66.330 105.660 67.940 107.425 ;
        RECT 63.000 105.650 67.940 105.660 ;
        RECT 54.190 105.530 67.940 105.650 ;
        RECT 10.180 104.850 67.940 105.530 ;
        RECT 0.560 103.250 3.460 104.850 ;
        RECT 5.060 104.550 67.940 104.850 ;
        RECT 69.520 105.660 71.130 107.425 ;
        RECT 72.860 105.660 74.460 108.720 ;
        RECT 69.520 105.650 74.460 105.660 ;
        RECT 77.200 105.650 78.800 108.730 ;
        RECT 81.540 108.720 83.270 108.730 ;
        RECT 86.330 108.730 100.080 108.850 ;
        RECT 86.330 108.720 88.060 108.730 ;
        RECT 81.540 105.660 83.140 108.720 ;
        RECT 86.460 105.660 88.060 108.720 ;
        RECT 81.540 105.650 83.270 105.660 ;
        RECT 69.520 105.530 83.270 105.650 ;
        RECT 86.330 105.650 88.060 105.660 ;
        RECT 90.800 105.650 92.400 108.730 ;
        RECT 95.140 108.720 100.080 108.730 ;
        RECT 95.140 105.660 96.740 108.720 ;
        RECT 98.470 105.660 100.080 108.720 ;
        RECT 95.140 105.650 100.080 105.660 ;
        RECT 86.330 105.530 100.080 105.650 ;
        RECT 69.520 104.550 100.080 105.530 ;
        RECT 5.060 104.060 100.080 104.550 ;
        RECT 5.060 103.250 11.790 104.060 ;
        RECT 1.860 101.650 6.660 103.250 ;
        RECT 0.560 100.050 3.460 101.650 ;
        RECT 5.060 100.050 7.960 101.650 ;
        RECT 10.180 101.190 11.790 103.250 ;
        RECT 13.400 103.930 64.720 104.060 ;
        RECT 13.400 101.190 23.920 103.930 ;
        RECT 27.000 101.190 37.520 103.930 ;
        RECT 40.600 101.190 51.120 103.930 ;
        RECT 54.200 101.190 64.720 103.930 ;
        RECT 66.330 102.950 71.130 104.060 ;
        RECT 66.330 101.190 67.940 102.950 ;
        RECT 10.180 100.135 67.940 101.190 ;
        RECT 69.520 101.190 71.130 102.950 ;
        RECT 72.740 103.930 96.860 104.060 ;
        RECT 72.740 101.190 83.260 103.930 ;
        RECT 86.340 101.190 96.860 103.930 ;
        RECT 98.470 101.190 100.080 104.060 ;
        RECT 69.520 100.135 100.080 101.190 ;
        RECT 1.860 98.450 6.660 100.050 ;
        RECT 10.180 99.590 100.080 100.135 ;
        RECT 10.180 98.450 11.790 99.590 ;
        RECT 0.560 96.850 3.460 98.450 ;
        RECT 5.060 96.850 11.790 98.450 ;
        RECT 1.860 95.250 6.660 96.850 ;
        RECT 10.180 96.720 11.790 96.850 ;
        RECT 13.400 96.850 23.920 99.590 ;
        RECT 27.000 96.850 37.520 99.590 ;
        RECT 40.600 96.850 51.120 99.590 ;
        RECT 54.200 96.850 64.720 99.590 ;
        RECT 13.400 96.720 64.720 96.850 ;
        RECT 66.330 98.535 71.130 99.590 ;
        RECT 66.330 96.720 67.940 98.535 ;
        RECT 10.180 95.250 67.940 96.720 ;
        RECT 0.560 93.650 3.460 95.250 ;
        RECT 5.060 93.650 7.960 95.250 ;
        RECT 10.180 95.130 23.930 95.250 ;
        RECT 10.180 95.120 15.120 95.130 ;
        RECT 1.860 92.050 6.660 93.650 ;
        RECT 10.180 92.060 11.790 95.120 ;
        RECT 13.520 92.060 15.120 95.120 ;
        RECT 10.180 92.050 15.120 92.060 ;
        RECT 17.860 92.050 19.460 95.130 ;
        RECT 22.200 95.120 23.930 95.130 ;
        RECT 26.990 95.130 37.530 95.250 ;
        RECT 26.990 95.120 28.720 95.130 ;
        RECT 22.200 92.060 23.800 95.120 ;
        RECT 27.120 92.060 28.720 95.120 ;
        RECT 22.200 92.050 23.930 92.060 ;
        RECT 0.560 90.450 3.460 92.050 ;
        RECT 5.060 91.930 23.930 92.050 ;
        RECT 26.990 92.050 28.720 92.060 ;
        RECT 31.460 92.050 33.060 95.130 ;
        RECT 35.800 95.120 37.530 95.130 ;
        RECT 40.590 95.130 51.130 95.250 ;
        RECT 40.590 95.120 42.320 95.130 ;
        RECT 35.800 92.060 37.400 95.120 ;
        RECT 40.720 92.060 42.320 95.120 ;
        RECT 35.800 92.050 37.530 92.060 ;
        RECT 26.990 91.930 37.530 92.050 ;
        RECT 40.590 92.050 42.320 92.060 ;
        RECT 45.060 92.050 46.660 95.130 ;
        RECT 49.400 95.120 51.130 95.130 ;
        RECT 54.190 95.130 67.940 95.250 ;
        RECT 54.190 95.120 55.920 95.130 ;
        RECT 49.400 92.060 51.000 95.120 ;
        RECT 54.320 92.060 55.920 95.120 ;
        RECT 49.400 92.050 51.130 92.060 ;
        RECT 40.590 91.930 51.130 92.050 ;
        RECT 54.190 92.050 55.920 92.060 ;
        RECT 58.660 92.050 60.260 95.130 ;
        RECT 63.000 95.120 67.940 95.130 ;
        RECT 63.000 92.060 64.600 95.120 ;
        RECT 66.330 92.060 67.940 95.120 ;
        RECT 63.000 92.050 67.940 92.060 ;
        RECT 54.190 91.930 67.940 92.050 ;
        RECT 5.060 91.615 67.940 91.930 ;
        RECT 69.520 96.720 71.130 98.535 ;
        RECT 72.740 96.850 83.260 99.590 ;
        RECT 86.340 96.850 96.860 99.590 ;
        RECT 72.740 96.720 96.860 96.850 ;
        RECT 98.470 96.720 100.080 99.590 ;
        RECT 69.520 95.250 100.080 96.720 ;
        RECT 69.520 95.130 83.270 95.250 ;
        RECT 69.520 95.120 74.460 95.130 ;
        RECT 69.520 92.060 71.130 95.120 ;
        RECT 72.860 92.060 74.460 95.120 ;
        RECT 69.520 92.050 74.460 92.060 ;
        RECT 77.200 92.050 78.800 95.130 ;
        RECT 81.540 95.120 83.270 95.130 ;
        RECT 86.330 95.130 100.080 95.250 ;
        RECT 86.330 95.120 88.060 95.130 ;
        RECT 81.540 92.060 83.140 95.120 ;
        RECT 86.460 92.060 88.060 95.120 ;
        RECT 81.540 92.050 83.270 92.060 ;
        RECT 69.520 91.930 83.270 92.050 ;
        RECT 86.330 92.050 88.060 92.060 ;
        RECT 90.800 92.050 92.400 95.130 ;
        RECT 95.140 95.120 100.080 95.130 ;
        RECT 95.140 92.060 96.740 95.120 ;
        RECT 98.470 92.060 100.080 95.120 ;
        RECT 95.140 92.050 100.080 92.060 ;
        RECT 86.330 91.930 100.080 92.050 ;
        RECT 69.520 91.615 100.080 91.930 ;
        RECT 5.060 90.460 100.080 91.615 ;
        RECT 5.060 90.450 11.790 90.460 ;
        RECT 1.860 88.850 6.660 90.450 ;
        RECT 0.560 87.250 3.460 88.850 ;
        RECT 5.060 87.250 7.960 88.850 ;
        RECT 10.180 87.590 11.790 90.450 ;
        RECT 13.400 90.330 64.720 90.460 ;
        RECT 13.400 87.590 23.920 90.330 ;
        RECT 27.000 87.590 37.520 90.330 ;
        RECT 40.600 87.590 51.120 90.330 ;
        RECT 54.200 87.590 64.720 90.330 ;
        RECT 66.330 90.015 71.130 90.460 ;
        RECT 66.330 87.590 67.940 90.015 ;
        RECT 1.860 85.650 6.660 87.250 ;
        RECT 10.180 87.205 67.940 87.590 ;
        RECT 69.520 87.590 71.130 90.015 ;
        RECT 72.740 90.330 96.860 90.460 ;
        RECT 72.740 87.590 83.260 90.330 ;
        RECT 86.340 87.590 96.860 90.330 ;
        RECT 98.470 87.590 100.080 90.460 ;
        RECT 69.520 87.205 100.080 87.590 ;
        RECT 10.180 85.990 100.080 87.205 ;
        RECT 10.180 85.650 11.790 85.990 ;
        RECT 0.560 84.050 3.460 85.650 ;
        RECT 5.060 84.050 11.790 85.650 ;
        RECT 1.860 82.450 6.660 84.050 ;
        RECT 10.180 83.120 11.790 84.050 ;
        RECT 13.400 83.250 23.920 85.990 ;
        RECT 27.000 83.250 37.520 85.990 ;
        RECT 40.600 83.250 51.120 85.990 ;
        RECT 54.200 83.250 64.720 85.990 ;
        RECT 13.400 83.120 64.720 83.250 ;
        RECT 66.330 85.605 71.130 85.990 ;
        RECT 66.330 83.120 67.940 85.605 ;
        RECT 10.180 82.720 67.940 83.120 ;
        RECT 69.520 83.120 71.130 85.605 ;
        RECT 72.740 83.250 83.260 85.990 ;
        RECT 86.340 83.250 96.860 85.990 ;
        RECT 72.740 83.120 96.860 83.250 ;
        RECT 98.470 83.120 100.080 85.990 ;
        RECT 69.520 82.720 100.080 83.120 ;
        RECT 0.560 80.850 3.460 82.450 ;
        RECT 5.060 80.850 7.960 82.450 ;
        RECT 10.180 81.650 100.080 82.720 ;
        RECT 10.180 81.530 23.930 81.650 ;
        RECT 10.180 81.520 15.120 81.530 ;
        RECT 1.860 79.250 6.660 80.850 ;
        RECT 10.180 79.250 11.790 81.520 ;
        RECT 0.560 77.650 3.460 79.250 ;
        RECT 5.060 78.460 11.790 79.250 ;
        RECT 13.520 78.460 15.120 81.520 ;
        RECT 5.060 78.450 15.120 78.460 ;
        RECT 17.860 78.450 19.460 81.530 ;
        RECT 22.200 81.520 23.930 81.530 ;
        RECT 26.990 81.530 37.530 81.650 ;
        RECT 26.990 81.520 28.720 81.530 ;
        RECT 22.200 78.460 23.800 81.520 ;
        RECT 27.120 78.460 28.720 81.520 ;
        RECT 22.200 78.450 23.930 78.460 ;
        RECT 5.060 78.330 23.930 78.450 ;
        RECT 26.990 78.450 28.720 78.460 ;
        RECT 31.460 78.450 33.060 81.530 ;
        RECT 35.800 81.520 37.530 81.530 ;
        RECT 40.590 81.530 51.130 81.650 ;
        RECT 40.590 81.520 42.320 81.530 ;
        RECT 35.800 78.460 37.400 81.520 ;
        RECT 40.720 78.460 42.320 81.520 ;
        RECT 35.800 78.450 37.530 78.460 ;
        RECT 26.990 78.330 37.530 78.450 ;
        RECT 40.590 78.450 42.320 78.460 ;
        RECT 45.060 78.450 46.660 81.530 ;
        RECT 49.400 81.520 51.130 81.530 ;
        RECT 54.190 81.530 83.270 81.650 ;
        RECT 54.190 81.520 55.920 81.530 ;
        RECT 49.400 78.460 51.000 81.520 ;
        RECT 54.320 78.460 55.920 81.520 ;
        RECT 49.400 78.450 51.130 78.460 ;
        RECT 40.590 78.330 51.130 78.450 ;
        RECT 54.190 78.450 55.920 78.460 ;
        RECT 58.660 78.450 60.260 81.530 ;
        RECT 63.000 81.520 74.460 81.530 ;
        RECT 63.000 78.460 64.600 81.520 ;
        RECT 66.330 81.120 71.130 81.520 ;
        RECT 66.330 78.460 67.940 81.120 ;
        RECT 63.000 78.450 67.940 78.460 ;
        RECT 54.190 78.330 67.940 78.450 ;
        RECT 5.060 77.650 67.940 78.330 ;
        RECT 1.860 76.050 6.660 77.650 ;
        RECT 10.180 76.860 67.940 77.650 ;
        RECT 0.560 74.450 3.460 76.050 ;
        RECT 5.060 74.450 7.960 76.050 ;
        RECT 1.860 72.850 6.660 74.450 ;
        RECT 10.180 73.990 11.790 76.860 ;
        RECT 13.400 76.730 64.720 76.860 ;
        RECT 13.400 73.990 23.920 76.730 ;
        RECT 27.000 73.990 37.520 76.730 ;
        RECT 40.600 73.990 51.120 76.730 ;
        RECT 54.200 73.990 64.720 76.730 ;
        RECT 66.330 74.255 67.940 76.860 ;
        RECT 69.520 78.460 71.130 81.120 ;
        RECT 72.860 78.460 74.460 81.520 ;
        RECT 69.520 78.450 74.460 78.460 ;
        RECT 77.200 78.450 78.800 81.530 ;
        RECT 81.540 81.520 83.270 81.530 ;
        RECT 86.330 81.530 100.080 81.650 ;
        RECT 86.330 81.520 88.060 81.530 ;
        RECT 81.540 78.460 83.140 81.520 ;
        RECT 86.460 78.460 88.060 81.520 ;
        RECT 81.540 78.450 83.270 78.460 ;
        RECT 69.520 78.330 83.270 78.450 ;
        RECT 86.330 78.450 88.060 78.460 ;
        RECT 90.800 78.450 92.400 81.530 ;
        RECT 95.140 81.520 100.080 81.530 ;
        RECT 95.140 78.460 96.740 81.520 ;
        RECT 98.470 78.460 100.080 81.520 ;
        RECT 95.140 78.450 100.080 78.460 ;
        RECT 86.330 78.330 100.080 78.450 ;
        RECT 69.520 76.860 100.080 78.330 ;
        RECT 69.520 74.255 71.130 76.860 ;
        RECT 66.330 73.990 71.130 74.255 ;
        RECT 72.740 76.730 96.860 76.860 ;
        RECT 72.740 73.990 83.260 76.730 ;
        RECT 86.340 73.990 96.860 76.730 ;
        RECT 98.470 73.990 100.080 76.860 ;
        RECT 10.180 72.850 100.080 73.990 ;
        RECT 0.560 71.250 3.460 72.850 ;
        RECT 5.060 72.655 100.080 72.850 ;
        RECT 5.060 72.390 67.940 72.655 ;
        RECT 5.060 71.250 11.790 72.390 ;
        RECT 1.860 69.650 6.660 71.250 ;
        RECT 0.560 68.050 3.460 69.650 ;
        RECT 5.060 68.050 7.960 69.650 ;
        RECT 10.180 69.520 11.790 71.250 ;
        RECT 13.400 69.650 23.920 72.390 ;
        RECT 27.000 69.650 37.520 72.390 ;
        RECT 40.600 69.650 51.120 72.390 ;
        RECT 54.200 69.650 64.720 72.390 ;
        RECT 13.400 69.520 64.720 69.650 ;
        RECT 66.330 69.765 67.940 72.390 ;
        RECT 69.520 72.390 100.080 72.655 ;
        RECT 69.520 69.765 71.130 72.390 ;
        RECT 66.330 69.520 71.130 69.765 ;
        RECT 72.740 69.650 83.260 72.390 ;
        RECT 86.340 69.650 96.860 72.390 ;
        RECT 72.740 69.520 96.860 69.650 ;
        RECT 98.470 69.520 100.080 72.390 ;
        RECT 10.180 68.165 100.080 69.520 ;
        RECT 10.180 68.050 67.940 68.165 ;
        RECT 1.860 66.450 6.660 68.050 ;
        RECT 10.180 67.930 23.930 68.050 ;
        RECT 10.180 67.920 15.120 67.930 ;
        RECT 10.180 66.450 11.790 67.920 ;
        RECT 0.560 64.850 3.460 66.450 ;
        RECT 5.060 64.860 11.790 66.450 ;
        RECT 13.520 64.860 15.120 67.920 ;
        RECT 5.060 64.850 15.120 64.860 ;
        RECT 17.860 64.850 19.460 67.930 ;
        RECT 22.200 67.920 23.930 67.930 ;
        RECT 26.990 67.930 37.530 68.050 ;
        RECT 26.990 67.920 28.720 67.930 ;
        RECT 22.200 64.860 23.800 67.920 ;
        RECT 27.120 64.860 28.720 67.920 ;
        RECT 22.200 64.850 23.930 64.860 ;
        RECT 1.860 63.250 6.660 64.850 ;
        RECT 10.180 64.730 23.930 64.850 ;
        RECT 26.990 64.850 28.720 64.860 ;
        RECT 31.460 64.850 33.060 67.930 ;
        RECT 35.800 67.920 37.530 67.930 ;
        RECT 40.590 67.930 51.130 68.050 ;
        RECT 40.590 67.920 42.320 67.930 ;
        RECT 35.800 64.860 37.400 67.920 ;
        RECT 40.720 64.860 42.320 67.920 ;
        RECT 35.800 64.850 37.530 64.860 ;
        RECT 26.990 64.730 37.530 64.850 ;
        RECT 40.590 64.850 42.320 64.860 ;
        RECT 45.060 64.850 46.660 67.930 ;
        RECT 49.400 67.920 51.130 67.930 ;
        RECT 54.190 67.930 67.940 68.050 ;
        RECT 54.190 67.920 55.920 67.930 ;
        RECT 49.400 64.860 51.000 67.920 ;
        RECT 54.320 64.860 55.920 67.920 ;
        RECT 49.400 64.850 51.130 64.860 ;
        RECT 40.590 64.730 51.130 64.850 ;
        RECT 54.190 64.850 55.920 64.860 ;
        RECT 58.660 64.850 60.260 67.930 ;
        RECT 63.000 67.920 67.940 67.930 ;
        RECT 63.000 64.860 64.600 67.920 ;
        RECT 66.330 65.300 67.940 67.920 ;
        RECT 69.520 68.050 100.080 68.165 ;
        RECT 69.520 67.930 83.270 68.050 ;
        RECT 69.520 67.920 74.460 67.930 ;
        RECT 69.520 65.300 71.130 67.920 ;
        RECT 66.330 64.860 71.130 65.300 ;
        RECT 72.860 64.860 74.460 67.920 ;
        RECT 63.000 64.850 74.460 64.860 ;
        RECT 77.200 64.850 78.800 67.930 ;
        RECT 81.540 67.920 83.270 67.930 ;
        RECT 86.330 67.930 100.080 68.050 ;
        RECT 86.330 67.920 88.060 67.930 ;
        RECT 81.540 64.860 83.140 67.920 ;
        RECT 86.460 64.860 88.060 67.920 ;
        RECT 81.540 64.850 83.270 64.860 ;
        RECT 54.190 64.730 83.270 64.850 ;
        RECT 86.330 64.850 88.060 64.860 ;
        RECT 90.800 64.850 92.400 67.930 ;
        RECT 95.140 67.920 100.080 67.930 ;
        RECT 95.140 64.860 96.740 67.920 ;
        RECT 98.470 64.860 100.080 67.920 ;
        RECT 95.140 64.850 100.080 64.860 ;
        RECT 86.330 64.730 100.080 64.850 ;
        RECT 10.180 63.700 100.080 64.730 ;
        RECT 10.180 63.260 67.940 63.700 ;
        RECT 0.560 61.650 3.460 63.250 ;
        RECT 5.060 61.650 7.960 63.250 ;
        RECT 1.860 60.050 6.660 61.650 ;
        RECT 10.180 60.390 11.790 63.260 ;
        RECT 13.400 63.130 64.720 63.260 ;
        RECT 13.400 60.390 23.920 63.130 ;
        RECT 27.000 60.390 37.520 63.130 ;
        RECT 40.600 60.390 51.120 63.130 ;
        RECT 54.200 60.390 64.720 63.130 ;
        RECT 66.330 60.390 67.940 63.260 ;
        RECT 10.180 60.050 67.940 60.390 ;
        RECT 0.560 58.450 3.460 60.050 ;
        RECT 5.060 58.790 67.940 60.050 ;
        RECT 5.060 58.450 11.790 58.790 ;
        RECT 1.860 56.850 6.660 58.450 ;
        RECT 0.560 55.250 3.460 56.850 ;
        RECT 5.060 55.250 7.960 56.850 ;
        RECT 10.180 55.920 11.790 58.450 ;
        RECT 13.400 56.050 23.920 58.790 ;
        RECT 27.000 56.050 37.520 58.790 ;
        RECT 40.600 56.050 51.120 58.790 ;
        RECT 54.200 56.050 64.720 58.790 ;
        RECT 13.400 55.920 64.720 56.050 ;
        RECT 66.330 56.820 67.940 58.790 ;
        RECT 69.520 63.260 100.080 63.700 ;
        RECT 69.520 60.390 71.130 63.260 ;
        RECT 72.740 63.130 96.860 63.260 ;
        RECT 72.740 60.390 83.260 63.130 ;
        RECT 86.340 60.390 96.860 63.130 ;
        RECT 98.470 60.390 100.080 63.260 ;
        RECT 69.520 58.790 100.080 60.390 ;
        RECT 69.520 56.820 71.130 58.790 ;
        RECT 66.330 55.920 71.130 56.820 ;
        RECT 72.740 56.050 83.260 58.790 ;
        RECT 86.340 56.050 96.860 58.790 ;
        RECT 72.740 55.920 96.860 56.050 ;
        RECT 98.470 55.920 100.080 58.790 ;
        RECT 1.860 53.650 6.660 55.250 ;
        RECT 10.180 55.220 100.080 55.920 ;
        RECT 10.180 54.450 67.940 55.220 ;
        RECT 10.180 54.330 23.930 54.450 ;
        RECT 10.180 54.320 15.120 54.330 ;
        RECT 10.180 53.650 11.790 54.320 ;
        RECT 0.560 52.050 3.460 53.650 ;
        RECT 5.060 52.050 11.790 53.650 ;
        RECT 1.860 50.450 6.660 52.050 ;
        RECT 10.180 51.260 11.790 52.050 ;
        RECT 13.520 51.260 15.120 54.320 ;
        RECT 10.180 51.250 15.120 51.260 ;
        RECT 17.860 51.250 19.460 54.330 ;
        RECT 22.200 54.320 23.930 54.330 ;
        RECT 26.990 54.330 37.530 54.450 ;
        RECT 26.990 54.320 28.720 54.330 ;
        RECT 22.200 51.260 23.800 54.320 ;
        RECT 27.120 51.260 28.720 54.320 ;
        RECT 22.200 51.250 23.930 51.260 ;
        RECT 10.180 51.130 23.930 51.250 ;
        RECT 26.990 51.250 28.720 51.260 ;
        RECT 31.460 51.250 33.060 54.330 ;
        RECT 35.800 54.320 37.530 54.330 ;
        RECT 40.590 54.330 51.130 54.450 ;
        RECT 40.590 54.320 42.320 54.330 ;
        RECT 35.800 51.260 37.400 54.320 ;
        RECT 40.720 51.260 42.320 54.320 ;
        RECT 35.800 51.250 37.530 51.260 ;
        RECT 26.990 51.130 37.530 51.250 ;
        RECT 40.590 51.250 42.320 51.260 ;
        RECT 45.060 51.250 46.660 54.330 ;
        RECT 49.400 54.320 51.130 54.330 ;
        RECT 54.190 54.330 67.940 54.450 ;
        RECT 54.190 54.320 55.920 54.330 ;
        RECT 49.400 51.260 51.000 54.320 ;
        RECT 54.320 51.260 55.920 54.320 ;
        RECT 49.400 51.250 51.130 51.260 ;
        RECT 40.590 51.130 51.130 51.250 ;
        RECT 54.190 51.250 55.920 51.260 ;
        RECT 58.660 51.250 60.260 54.330 ;
        RECT 63.000 54.320 67.940 54.330 ;
        RECT 63.000 51.260 64.600 54.320 ;
        RECT 66.330 52.355 67.940 54.320 ;
        RECT 69.520 54.450 100.080 55.220 ;
        RECT 69.520 54.330 83.270 54.450 ;
        RECT 69.520 54.320 74.460 54.330 ;
        RECT 69.520 52.355 71.130 54.320 ;
        RECT 66.330 51.260 71.130 52.355 ;
        RECT 72.860 51.260 74.460 54.320 ;
        RECT 63.000 51.250 74.460 51.260 ;
        RECT 77.200 51.250 78.800 54.330 ;
        RECT 81.540 54.320 83.270 54.330 ;
        RECT 86.330 54.330 100.080 54.450 ;
        RECT 86.330 54.320 88.060 54.330 ;
        RECT 81.540 51.260 83.140 54.320 ;
        RECT 86.460 51.260 88.060 54.320 ;
        RECT 81.540 51.250 83.270 51.260 ;
        RECT 54.190 51.130 83.270 51.250 ;
        RECT 86.330 51.250 88.060 51.260 ;
        RECT 90.800 51.250 92.400 54.330 ;
        RECT 95.140 54.320 100.080 54.330 ;
        RECT 95.140 51.260 96.740 54.320 ;
        RECT 98.470 51.260 100.080 54.320 ;
        RECT 95.140 51.250 100.080 51.260 ;
        RECT 86.330 51.130 100.080 51.250 ;
        RECT 10.180 50.755 100.080 51.130 ;
        RECT 0.560 48.850 3.460 50.450 ;
        RECT 5.060 48.850 7.960 50.450 ;
        RECT 10.180 49.660 67.940 50.755 ;
        RECT 1.860 47.250 6.660 48.850 ;
        RECT 10.180 47.250 11.790 49.660 ;
        RECT 0.560 45.650 3.460 47.250 ;
        RECT 5.060 46.790 11.790 47.250 ;
        RECT 13.400 49.530 64.720 49.660 ;
        RECT 13.400 46.790 23.920 49.530 ;
        RECT 27.000 46.790 37.520 49.530 ;
        RECT 40.600 46.790 51.120 49.530 ;
        RECT 54.200 46.790 64.720 49.530 ;
        RECT 66.330 47.880 67.940 49.660 ;
        RECT 69.520 49.660 100.080 50.755 ;
        RECT 69.520 47.880 71.130 49.660 ;
        RECT 66.330 46.790 71.130 47.880 ;
        RECT 72.740 49.530 96.860 49.660 ;
        RECT 72.740 46.790 83.260 49.530 ;
        RECT 86.340 46.790 96.860 49.530 ;
        RECT 98.470 46.790 100.080 49.660 ;
        RECT 5.060 46.280 100.080 46.790 ;
        RECT 5.060 45.650 67.940 46.280 ;
        RECT 1.860 44.050 6.660 45.650 ;
        RECT 10.180 45.190 67.940 45.650 ;
        RECT 0.560 42.450 3.460 44.050 ;
        RECT 5.060 42.450 7.960 44.050 ;
        RECT 1.860 40.850 6.660 42.450 ;
        RECT 10.180 42.320 11.790 45.190 ;
        RECT 13.400 42.450 23.920 45.190 ;
        RECT 27.000 42.450 37.520 45.190 ;
        RECT 40.600 42.450 51.120 45.190 ;
        RECT 54.200 42.450 64.720 45.190 ;
        RECT 13.400 42.320 64.720 42.450 ;
        RECT 66.330 42.320 67.940 45.190 ;
        RECT 10.180 40.850 67.940 42.320 ;
        RECT 0.560 39.250 3.460 40.850 ;
        RECT 5.060 40.730 23.930 40.850 ;
        RECT 5.060 40.720 15.120 40.730 ;
        RECT 5.060 39.250 11.790 40.720 ;
        RECT 1.860 37.650 6.660 39.250 ;
        RECT 10.180 37.660 11.790 39.250 ;
        RECT 13.520 37.660 15.120 40.720 ;
        RECT 10.180 37.650 15.120 37.660 ;
        RECT 17.860 37.650 19.460 40.730 ;
        RECT 22.200 40.720 23.930 40.730 ;
        RECT 26.990 40.730 37.530 40.850 ;
        RECT 26.990 40.720 28.720 40.730 ;
        RECT 22.200 37.660 23.800 40.720 ;
        RECT 27.120 37.660 28.720 40.720 ;
        RECT 22.200 37.650 23.930 37.660 ;
        RECT 0.560 36.050 3.460 37.650 ;
        RECT 5.060 36.050 7.960 37.650 ;
        RECT 10.180 37.530 23.930 37.650 ;
        RECT 26.990 37.650 28.720 37.660 ;
        RECT 31.460 37.650 33.060 40.730 ;
        RECT 35.800 40.720 37.530 40.730 ;
        RECT 40.590 40.730 51.130 40.850 ;
        RECT 40.590 40.720 42.320 40.730 ;
        RECT 35.800 37.660 37.400 40.720 ;
        RECT 40.720 37.660 42.320 40.720 ;
        RECT 35.800 37.650 37.530 37.660 ;
        RECT 26.990 37.530 37.530 37.650 ;
        RECT 40.590 37.650 42.320 37.660 ;
        RECT 45.060 37.650 46.660 40.730 ;
        RECT 49.400 40.720 51.130 40.730 ;
        RECT 54.190 40.730 67.940 40.850 ;
        RECT 54.190 40.720 55.920 40.730 ;
        RECT 49.400 37.660 51.000 40.720 ;
        RECT 54.320 37.660 55.920 40.720 ;
        RECT 49.400 37.650 51.130 37.660 ;
        RECT 40.590 37.530 51.130 37.650 ;
        RECT 54.190 37.650 55.920 37.660 ;
        RECT 58.660 37.650 60.260 40.730 ;
        RECT 63.000 40.720 67.940 40.730 ;
        RECT 63.000 37.660 64.600 40.720 ;
        RECT 66.330 39.390 67.940 40.720 ;
        RECT 69.520 45.190 100.080 46.280 ;
        RECT 69.520 42.320 71.130 45.190 ;
        RECT 72.740 42.450 83.260 45.190 ;
        RECT 86.340 42.450 96.860 45.190 ;
        RECT 72.740 42.320 96.860 42.450 ;
        RECT 98.470 42.320 100.080 45.190 ;
        RECT 69.520 40.850 100.080 42.320 ;
        RECT 69.520 40.730 83.270 40.850 ;
        RECT 69.520 40.720 74.460 40.730 ;
        RECT 69.520 39.390 71.130 40.720 ;
        RECT 66.330 37.790 71.130 39.390 ;
        RECT 66.330 37.660 67.940 37.790 ;
        RECT 63.000 37.650 67.940 37.660 ;
        RECT 54.190 37.530 67.940 37.650 ;
        RECT 10.180 36.060 67.940 37.530 ;
        RECT 1.860 34.450 6.660 36.050 ;
        RECT 10.180 34.450 11.790 36.060 ;
        RECT 0.560 32.850 3.460 34.450 ;
        RECT 5.060 33.190 11.790 34.450 ;
        RECT 13.400 35.930 64.720 36.060 ;
        RECT 13.400 33.190 23.920 35.930 ;
        RECT 27.000 33.190 37.520 35.930 ;
        RECT 40.600 33.190 51.120 35.930 ;
        RECT 54.200 33.190 64.720 35.930 ;
        RECT 66.330 34.925 67.940 36.060 ;
        RECT 69.520 37.660 71.130 37.790 ;
        RECT 72.860 37.660 74.460 40.720 ;
        RECT 69.520 37.650 74.460 37.660 ;
        RECT 77.200 37.650 78.800 40.730 ;
        RECT 81.540 40.720 83.270 40.730 ;
        RECT 86.330 40.730 100.080 40.850 ;
        RECT 86.330 40.720 88.060 40.730 ;
        RECT 81.540 37.660 83.140 40.720 ;
        RECT 86.460 37.660 88.060 40.720 ;
        RECT 81.540 37.650 83.270 37.660 ;
        RECT 69.520 37.530 83.270 37.650 ;
        RECT 86.330 37.650 88.060 37.660 ;
        RECT 90.800 37.650 92.400 40.730 ;
        RECT 95.140 40.720 100.080 40.730 ;
        RECT 95.140 37.660 96.740 40.720 ;
        RECT 98.470 37.660 100.080 40.720 ;
        RECT 95.140 37.650 100.080 37.660 ;
        RECT 86.330 37.530 100.080 37.650 ;
        RECT 69.520 36.060 100.080 37.530 ;
        RECT 69.520 34.925 71.130 36.060 ;
        RECT 66.330 33.325 71.130 34.925 ;
        RECT 66.330 33.190 67.940 33.325 ;
        RECT 5.060 32.850 67.940 33.190 ;
        RECT 1.860 31.250 6.660 32.850 ;
        RECT 10.180 31.590 67.940 32.850 ;
        RECT 0.560 29.650 3.460 31.250 ;
        RECT 5.060 29.650 7.960 31.250 ;
        RECT 1.860 28.050 6.660 29.650 ;
        RECT 10.180 28.720 11.790 31.590 ;
        RECT 13.400 28.850 23.920 31.590 ;
        RECT 27.000 28.850 37.520 31.590 ;
        RECT 40.600 28.850 51.120 31.590 ;
        RECT 54.200 28.850 64.720 31.590 ;
        RECT 13.400 28.720 64.720 28.850 ;
        RECT 66.330 30.465 67.940 31.590 ;
        RECT 69.520 33.190 71.130 33.325 ;
        RECT 72.740 35.930 96.860 36.060 ;
        RECT 72.740 33.190 83.260 35.930 ;
        RECT 86.340 33.190 96.860 35.930 ;
        RECT 98.470 33.190 100.080 36.060 ;
        RECT 69.520 31.590 100.080 33.190 ;
        RECT 69.520 30.465 71.130 31.590 ;
        RECT 66.330 28.865 71.130 30.465 ;
        RECT 66.330 28.720 67.940 28.865 ;
        RECT 10.180 28.050 67.940 28.720 ;
        RECT 0.560 26.450 3.460 28.050 ;
        RECT 5.060 27.250 67.940 28.050 ;
        RECT 5.060 27.130 23.930 27.250 ;
        RECT 5.060 27.120 15.120 27.130 ;
        RECT 5.060 26.450 11.790 27.120 ;
        RECT 1.860 24.850 6.660 26.450 ;
        RECT 0.560 23.250 3.460 24.850 ;
        RECT 5.060 23.250 7.960 24.850 ;
        RECT 10.180 24.060 11.790 26.450 ;
        RECT 13.520 24.060 15.120 27.120 ;
        RECT 10.180 24.050 15.120 24.060 ;
        RECT 17.860 24.050 19.460 27.130 ;
        RECT 22.200 27.120 23.930 27.130 ;
        RECT 26.990 27.130 37.530 27.250 ;
        RECT 26.990 27.120 28.720 27.130 ;
        RECT 22.200 24.060 23.800 27.120 ;
        RECT 27.120 24.060 28.720 27.120 ;
        RECT 22.200 24.050 23.930 24.060 ;
        RECT 10.180 23.930 23.930 24.050 ;
        RECT 26.990 24.050 28.720 24.060 ;
        RECT 31.460 24.050 33.060 27.130 ;
        RECT 35.800 27.120 37.530 27.130 ;
        RECT 40.590 27.130 51.130 27.250 ;
        RECT 40.590 27.120 42.320 27.130 ;
        RECT 35.800 24.060 37.400 27.120 ;
        RECT 40.720 24.060 42.320 27.120 ;
        RECT 35.800 24.050 37.530 24.060 ;
        RECT 26.990 23.930 37.530 24.050 ;
        RECT 40.590 24.050 42.320 24.060 ;
        RECT 45.060 24.050 46.660 27.130 ;
        RECT 49.400 27.120 51.130 27.130 ;
        RECT 54.190 27.130 67.940 27.250 ;
        RECT 54.190 27.120 55.920 27.130 ;
        RECT 49.400 24.060 51.000 27.120 ;
        RECT 54.320 24.060 55.920 27.120 ;
        RECT 49.400 24.050 51.130 24.060 ;
        RECT 40.590 23.930 51.130 24.050 ;
        RECT 54.190 24.050 55.920 24.060 ;
        RECT 58.660 24.050 60.260 27.130 ;
        RECT 63.000 27.120 67.940 27.130 ;
        RECT 63.000 24.060 64.600 27.120 ;
        RECT 66.330 24.060 67.940 27.120 ;
        RECT 63.000 24.050 67.940 24.060 ;
        RECT 54.190 23.930 67.940 24.050 ;
        RECT 1.860 21.650 6.660 23.250 ;
        RECT 10.180 22.460 67.940 23.930 ;
        RECT 10.180 21.650 11.790 22.460 ;
        RECT 0.560 20.050 3.460 21.650 ;
        RECT 5.060 20.050 11.790 21.650 ;
        RECT 1.860 18.450 6.660 20.050 ;
        RECT 10.180 19.800 11.790 20.050 ;
        RECT 13.400 22.330 64.720 22.460 ;
        RECT 13.400 19.800 23.920 22.330 ;
        RECT 10.180 19.590 23.920 19.800 ;
        RECT 27.000 19.590 37.520 22.330 ;
        RECT 40.600 19.590 51.120 22.330 ;
        RECT 54.200 19.595 64.720 22.330 ;
        RECT 66.330 21.985 67.940 22.460 ;
        RECT 69.520 28.720 71.130 28.865 ;
        RECT 72.740 28.850 83.260 31.590 ;
        RECT 86.340 28.850 96.860 31.590 ;
        RECT 72.740 28.720 96.860 28.850 ;
        RECT 98.470 28.720 100.080 31.590 ;
        RECT 69.520 27.250 100.080 28.720 ;
        RECT 69.520 27.130 83.270 27.250 ;
        RECT 69.520 27.120 74.460 27.130 ;
        RECT 69.520 24.060 71.130 27.120 ;
        RECT 72.860 24.060 74.460 27.120 ;
        RECT 69.520 24.050 74.460 24.060 ;
        RECT 77.200 24.050 78.800 27.130 ;
        RECT 81.540 27.120 83.270 27.130 ;
        RECT 86.330 27.130 100.080 27.250 ;
        RECT 86.330 27.120 88.060 27.130 ;
        RECT 81.540 24.060 83.140 27.120 ;
        RECT 86.460 24.060 88.060 27.120 ;
        RECT 81.540 24.050 83.270 24.060 ;
        RECT 69.520 23.930 83.270 24.050 ;
        RECT 86.330 24.050 88.060 24.060 ;
        RECT 90.800 24.050 92.400 27.130 ;
        RECT 95.140 27.120 100.080 27.130 ;
        RECT 95.140 24.060 96.740 27.120 ;
        RECT 98.470 24.060 100.080 27.120 ;
        RECT 95.140 24.050 100.080 24.060 ;
        RECT 86.330 23.930 100.080 24.050 ;
        RECT 69.520 22.460 100.080 23.930 ;
        RECT 69.520 21.985 71.130 22.460 ;
        RECT 66.330 20.385 71.130 21.985 ;
        RECT 66.330 19.595 67.940 20.385 ;
        RECT 54.200 19.590 67.940 19.595 ;
        RECT 0.560 16.850 3.460 18.450 ;
        RECT 5.060 16.850 7.960 18.450 ;
        RECT 10.180 18.195 67.940 19.590 ;
        RECT 1.860 15.250 6.660 16.850 ;
        RECT 10.180 15.530 11.790 18.195 ;
        RECT 13.400 17.995 67.940 18.195 ;
        RECT 13.400 17.990 64.720 17.995 ;
        RECT 13.400 15.530 23.920 17.990 ;
        RECT 10.180 15.250 23.920 15.530 ;
        RECT 27.000 15.250 37.520 17.990 ;
        RECT 40.600 15.250 51.120 17.990 ;
        RECT 54.200 15.250 64.720 17.990 ;
        RECT 0.560 13.650 3.460 15.250 ;
        RECT 1.860 10.850 3.460 13.650 ;
        RECT 5.060 15.130 64.720 15.250 ;
        RECT 66.330 17.515 67.940 17.995 ;
        RECT 69.520 19.800 71.130 20.385 ;
        RECT 72.740 22.330 96.860 22.460 ;
        RECT 72.740 19.800 83.260 22.330 ;
        RECT 69.520 19.590 83.260 19.800 ;
        RECT 86.340 19.595 96.860 22.330 ;
        RECT 98.470 19.595 100.080 22.460 ;
        RECT 86.340 19.590 100.080 19.595 ;
        RECT 69.520 18.195 100.080 19.590 ;
        RECT 69.520 17.515 71.130 18.195 ;
        RECT 66.330 15.915 71.130 17.515 ;
        RECT 66.330 15.130 67.940 15.915 ;
        RECT 5.060 13.930 67.940 15.130 ;
        RECT 5.060 13.650 11.790 13.930 ;
        RECT 5.060 10.850 6.660 13.650 ;
        RECT 10.180 11.920 11.790 13.650 ;
        RECT 13.400 13.650 67.940 13.930 ;
        RECT 13.400 13.530 23.930 13.650 ;
        RECT 13.400 11.920 15.000 13.530 ;
        RECT 17.865 11.920 19.465 13.530 ;
        RECT 22.330 11.920 23.930 13.530 ;
        RECT 26.990 13.530 37.530 13.650 ;
        RECT 26.990 11.920 28.590 13.530 ;
        RECT 31.460 11.920 33.060 13.530 ;
        RECT 35.930 11.920 37.530 13.530 ;
        RECT 40.590 13.530 51.130 13.650 ;
        RECT 40.590 11.920 42.190 13.530 ;
        RECT 45.060 11.920 46.660 13.530 ;
        RECT 49.530 11.920 51.130 13.530 ;
        RECT 54.190 13.530 67.940 13.650 ;
        RECT 54.190 11.920 55.790 13.530 ;
        RECT 58.450 11.920 60.055 13.530 ;
        RECT 62.720 11.920 64.320 13.530 ;
        RECT 66.330 13.045 67.940 13.530 ;
        RECT 69.520 15.530 71.130 15.915 ;
        RECT 72.740 17.995 100.080 18.195 ;
        RECT 72.740 17.990 96.860 17.995 ;
        RECT 72.740 15.530 83.260 17.990 ;
        RECT 69.520 15.250 83.260 15.530 ;
        RECT 86.340 15.250 96.860 17.990 ;
        RECT 69.520 15.130 96.860 15.250 ;
        RECT 98.470 15.130 100.080 17.995 ;
        RECT 69.520 13.930 100.080 15.130 ;
        RECT 69.520 13.045 71.130 13.930 ;
        RECT 66.330 11.920 71.130 13.045 ;
        RECT 72.740 13.650 100.080 13.930 ;
        RECT 72.740 13.530 83.270 13.650 ;
        RECT 72.740 11.920 74.340 13.530 ;
        RECT 77.205 11.920 78.805 13.530 ;
        RECT 81.670 11.920 83.270 13.530 ;
        RECT 86.330 13.530 100.080 13.650 ;
        RECT 86.330 11.920 87.930 13.530 ;
        RECT 90.590 11.920 92.195 13.530 ;
        RECT 94.860 11.920 96.460 13.530 ;
        RECT 98.470 11.920 100.080 13.530 ;
        RECT 10.180 11.445 100.080 11.920 ;
        RECT 10.180 10.310 67.940 11.445 ;
        RECT 69.520 10.310 100.080 11.445 ;
        RECT 140.300 121.790 170.860 122.470 ;
        RECT 172.440 121.790 230.200 122.470 ;
        RECT 232.420 122.450 235.320 124.050 ;
        RECT 236.920 122.450 239.820 124.050 ;
        RECT 140.300 120.860 230.200 121.790 ;
        RECT 140.300 118.850 141.910 120.860 ;
        RECT 143.520 119.250 145.120 120.860 ;
        RECT 147.985 119.250 149.585 120.860 ;
        RECT 152.450 119.250 154.050 120.860 ;
        RECT 143.520 119.130 154.050 119.250 ;
        RECT 157.110 119.250 158.710 120.860 ;
        RECT 161.370 119.250 162.975 120.860 ;
        RECT 165.640 119.250 167.240 120.860 ;
        RECT 169.250 120.190 174.050 120.860 ;
        RECT 169.250 119.250 170.860 120.190 ;
        RECT 157.110 119.130 170.860 119.250 ;
        RECT 143.520 118.850 170.860 119.130 ;
        RECT 140.300 117.650 170.860 118.850 ;
        RECT 140.300 117.530 167.640 117.650 ;
        RECT 140.300 117.250 154.040 117.530 ;
        RECT 140.300 114.585 141.910 117.250 ;
        RECT 143.520 114.790 154.040 117.250 ;
        RECT 157.120 114.790 167.640 117.530 ;
        RECT 143.520 114.785 167.640 114.790 ;
        RECT 169.250 114.785 170.860 117.650 ;
        RECT 143.520 114.635 170.860 114.785 ;
        RECT 172.440 118.850 174.050 120.190 ;
        RECT 175.660 119.250 177.260 120.860 ;
        RECT 180.125 119.250 181.725 120.860 ;
        RECT 184.590 119.250 186.190 120.860 ;
        RECT 175.660 119.130 186.190 119.250 ;
        RECT 189.250 119.250 190.850 120.860 ;
        RECT 193.720 119.250 195.320 120.860 ;
        RECT 198.190 119.250 199.790 120.860 ;
        RECT 189.250 119.130 199.790 119.250 ;
        RECT 202.850 119.250 204.450 120.860 ;
        RECT 207.320 119.250 208.920 120.860 ;
        RECT 211.790 119.250 213.390 120.860 ;
        RECT 202.850 119.130 213.390 119.250 ;
        RECT 216.450 119.250 218.050 120.860 ;
        RECT 220.710 119.250 222.315 120.860 ;
        RECT 224.980 119.250 226.580 120.860 ;
        RECT 228.590 119.250 230.200 120.860 ;
        RECT 233.720 120.850 238.520 122.450 ;
        RECT 232.420 119.250 235.320 120.850 ;
        RECT 236.920 119.250 239.820 120.850 ;
        RECT 216.450 119.130 230.200 119.250 ;
        RECT 175.660 118.850 230.200 119.130 ;
        RECT 172.440 117.650 230.200 118.850 ;
        RECT 233.720 117.650 238.520 119.250 ;
        RECT 172.440 117.530 226.980 117.650 ;
        RECT 172.440 117.250 186.180 117.530 ;
        RECT 172.440 114.635 174.050 117.250 ;
        RECT 143.520 114.585 174.050 114.635 ;
        RECT 175.660 114.790 186.180 117.250 ;
        RECT 189.260 114.790 199.780 117.530 ;
        RECT 202.860 114.790 213.380 117.530 ;
        RECT 216.460 114.790 226.980 117.530 ;
        RECT 175.660 114.785 226.980 114.790 ;
        RECT 228.590 116.050 235.320 117.650 ;
        RECT 236.920 116.050 239.820 117.650 ;
        RECT 228.590 114.785 230.200 116.050 ;
        RECT 175.660 114.585 230.200 114.785 ;
        RECT 140.300 113.190 230.200 114.585 ;
        RECT 233.720 114.450 238.520 116.050 ;
        RECT 140.300 112.980 154.040 113.190 ;
        RECT 140.300 110.320 141.910 112.980 ;
        RECT 143.520 110.450 154.040 112.980 ;
        RECT 157.120 113.185 186.180 113.190 ;
        RECT 157.120 110.450 167.640 113.185 ;
        RECT 143.520 110.320 167.640 110.450 ;
        RECT 169.250 113.035 186.180 113.185 ;
        RECT 169.250 110.320 170.860 113.035 ;
        RECT 140.300 109.025 170.860 110.320 ;
        RECT 172.440 112.980 186.180 113.035 ;
        RECT 172.440 110.320 174.050 112.980 ;
        RECT 175.660 110.450 186.180 112.980 ;
        RECT 189.260 110.450 199.780 113.190 ;
        RECT 202.860 110.450 213.380 113.190 ;
        RECT 216.460 113.185 230.200 113.190 ;
        RECT 216.460 110.450 226.980 113.185 ;
        RECT 175.660 110.320 226.980 110.450 ;
        RECT 228.590 111.250 230.200 113.185 ;
        RECT 232.420 112.850 235.320 114.450 ;
        RECT 236.920 112.850 239.820 114.450 ;
        RECT 233.720 111.250 238.520 112.850 ;
        RECT 228.590 110.320 235.320 111.250 ;
        RECT 172.440 109.650 235.320 110.320 ;
        RECT 236.920 109.650 239.820 111.250 ;
        RECT 172.440 109.025 230.200 109.650 ;
        RECT 140.300 108.850 230.200 109.025 ;
        RECT 140.300 108.730 154.050 108.850 ;
        RECT 140.300 108.720 145.240 108.730 ;
        RECT 140.300 105.660 141.910 108.720 ;
        RECT 143.640 105.660 145.240 108.720 ;
        RECT 140.300 105.650 145.240 105.660 ;
        RECT 147.980 105.650 149.580 108.730 ;
        RECT 152.320 108.720 154.050 108.730 ;
        RECT 157.110 108.730 186.190 108.850 ;
        RECT 157.110 108.720 158.840 108.730 ;
        RECT 152.320 105.660 153.920 108.720 ;
        RECT 157.240 105.660 158.840 108.720 ;
        RECT 152.320 105.650 154.050 105.660 ;
        RECT 140.300 105.530 154.050 105.650 ;
        RECT 157.110 105.650 158.840 105.660 ;
        RECT 161.580 105.650 163.180 108.730 ;
        RECT 165.920 108.720 177.380 108.730 ;
        RECT 165.920 105.660 167.520 108.720 ;
        RECT 169.250 107.425 174.050 108.720 ;
        RECT 169.250 105.660 170.860 107.425 ;
        RECT 165.920 105.650 170.860 105.660 ;
        RECT 157.110 105.530 170.860 105.650 ;
        RECT 140.300 104.550 170.860 105.530 ;
        RECT 172.440 105.660 174.050 107.425 ;
        RECT 175.780 105.660 177.380 108.720 ;
        RECT 172.440 105.650 177.380 105.660 ;
        RECT 180.120 105.650 181.720 108.730 ;
        RECT 184.460 108.720 186.190 108.730 ;
        RECT 189.250 108.730 199.790 108.850 ;
        RECT 189.250 108.720 190.980 108.730 ;
        RECT 184.460 105.660 186.060 108.720 ;
        RECT 189.380 105.660 190.980 108.720 ;
        RECT 184.460 105.650 186.190 105.660 ;
        RECT 172.440 105.530 186.190 105.650 ;
        RECT 189.250 105.650 190.980 105.660 ;
        RECT 193.720 105.650 195.320 108.730 ;
        RECT 198.060 108.720 199.790 108.730 ;
        RECT 202.850 108.730 213.390 108.850 ;
        RECT 202.850 108.720 204.580 108.730 ;
        RECT 198.060 105.660 199.660 108.720 ;
        RECT 202.980 105.660 204.580 108.720 ;
        RECT 198.060 105.650 199.790 105.660 ;
        RECT 189.250 105.530 199.790 105.650 ;
        RECT 202.850 105.650 204.580 105.660 ;
        RECT 207.320 105.650 208.920 108.730 ;
        RECT 211.660 108.720 213.390 108.730 ;
        RECT 216.450 108.730 230.200 108.850 ;
        RECT 216.450 108.720 218.180 108.730 ;
        RECT 211.660 105.660 213.260 108.720 ;
        RECT 216.580 105.660 218.180 108.720 ;
        RECT 211.660 105.650 213.390 105.660 ;
        RECT 202.850 105.530 213.390 105.650 ;
        RECT 216.450 105.650 218.180 105.660 ;
        RECT 220.920 105.650 222.520 108.730 ;
        RECT 225.260 108.720 230.200 108.730 ;
        RECT 225.260 105.660 226.860 108.720 ;
        RECT 228.590 105.660 230.200 108.720 ;
        RECT 233.720 108.050 238.520 109.650 ;
        RECT 232.420 106.450 235.320 108.050 ;
        RECT 236.920 106.450 239.820 108.050 ;
        RECT 225.260 105.650 230.200 105.660 ;
        RECT 216.450 105.530 230.200 105.650 ;
        RECT 172.440 104.850 230.200 105.530 ;
        RECT 233.720 104.850 238.520 106.450 ;
        RECT 172.440 104.550 235.320 104.850 ;
        RECT 140.300 104.060 235.320 104.550 ;
        RECT 140.300 101.190 141.910 104.060 ;
        RECT 143.520 103.930 167.640 104.060 ;
        RECT 143.520 101.190 154.040 103.930 ;
        RECT 157.120 101.190 167.640 103.930 ;
        RECT 169.250 102.950 174.050 104.060 ;
        RECT 169.250 101.190 170.860 102.950 ;
        RECT 140.300 100.135 170.860 101.190 ;
        RECT 172.440 101.190 174.050 102.950 ;
        RECT 175.660 103.930 226.980 104.060 ;
        RECT 175.660 101.190 186.180 103.930 ;
        RECT 189.260 101.190 199.780 103.930 ;
        RECT 202.860 101.190 213.380 103.930 ;
        RECT 216.460 101.190 226.980 103.930 ;
        RECT 228.590 103.250 235.320 104.060 ;
        RECT 236.920 103.250 239.820 104.850 ;
        RECT 228.590 101.190 230.200 103.250 ;
        RECT 233.720 101.650 238.520 103.250 ;
        RECT 172.440 100.135 230.200 101.190 ;
        RECT 140.300 99.590 230.200 100.135 ;
        RECT 232.420 100.050 235.320 101.650 ;
        RECT 236.920 100.050 239.820 101.650 ;
        RECT 140.300 96.720 141.910 99.590 ;
        RECT 143.520 96.850 154.040 99.590 ;
        RECT 157.120 96.850 167.640 99.590 ;
        RECT 143.520 96.720 167.640 96.850 ;
        RECT 169.250 98.535 174.050 99.590 ;
        RECT 169.250 96.720 170.860 98.535 ;
        RECT 140.300 95.250 170.860 96.720 ;
        RECT 140.300 95.130 154.050 95.250 ;
        RECT 140.300 95.120 145.240 95.130 ;
        RECT 140.300 92.060 141.910 95.120 ;
        RECT 143.640 92.060 145.240 95.120 ;
        RECT 140.300 92.050 145.240 92.060 ;
        RECT 147.980 92.050 149.580 95.130 ;
        RECT 152.320 95.120 154.050 95.130 ;
        RECT 157.110 95.130 170.860 95.250 ;
        RECT 157.110 95.120 158.840 95.130 ;
        RECT 152.320 92.060 153.920 95.120 ;
        RECT 157.240 92.060 158.840 95.120 ;
        RECT 152.320 92.050 154.050 92.060 ;
        RECT 140.300 91.930 154.050 92.050 ;
        RECT 157.110 92.050 158.840 92.060 ;
        RECT 161.580 92.050 163.180 95.130 ;
        RECT 165.920 95.120 170.860 95.130 ;
        RECT 165.920 92.060 167.520 95.120 ;
        RECT 169.250 92.060 170.860 95.120 ;
        RECT 165.920 92.050 170.860 92.060 ;
        RECT 157.110 91.930 170.860 92.050 ;
        RECT 140.300 91.615 170.860 91.930 ;
        RECT 172.440 96.720 174.050 98.535 ;
        RECT 175.660 96.850 186.180 99.590 ;
        RECT 189.260 96.850 199.780 99.590 ;
        RECT 202.860 96.850 213.380 99.590 ;
        RECT 216.460 96.850 226.980 99.590 ;
        RECT 175.660 96.720 226.980 96.850 ;
        RECT 228.590 98.450 230.200 99.590 ;
        RECT 233.720 98.450 238.520 100.050 ;
        RECT 228.590 96.850 235.320 98.450 ;
        RECT 236.920 96.850 239.820 98.450 ;
        RECT 228.590 96.720 230.200 96.850 ;
        RECT 172.440 95.250 230.200 96.720 ;
        RECT 233.720 95.250 238.520 96.850 ;
        RECT 172.440 95.130 186.190 95.250 ;
        RECT 172.440 95.120 177.380 95.130 ;
        RECT 172.440 92.060 174.050 95.120 ;
        RECT 175.780 92.060 177.380 95.120 ;
        RECT 172.440 92.050 177.380 92.060 ;
        RECT 180.120 92.050 181.720 95.130 ;
        RECT 184.460 95.120 186.190 95.130 ;
        RECT 189.250 95.130 199.790 95.250 ;
        RECT 189.250 95.120 190.980 95.130 ;
        RECT 184.460 92.060 186.060 95.120 ;
        RECT 189.380 92.060 190.980 95.120 ;
        RECT 184.460 92.050 186.190 92.060 ;
        RECT 172.440 91.930 186.190 92.050 ;
        RECT 189.250 92.050 190.980 92.060 ;
        RECT 193.720 92.050 195.320 95.130 ;
        RECT 198.060 95.120 199.790 95.130 ;
        RECT 202.850 95.130 213.390 95.250 ;
        RECT 202.850 95.120 204.580 95.130 ;
        RECT 198.060 92.060 199.660 95.120 ;
        RECT 202.980 92.060 204.580 95.120 ;
        RECT 198.060 92.050 199.790 92.060 ;
        RECT 189.250 91.930 199.790 92.050 ;
        RECT 202.850 92.050 204.580 92.060 ;
        RECT 207.320 92.050 208.920 95.130 ;
        RECT 211.660 95.120 213.390 95.130 ;
        RECT 216.450 95.130 230.200 95.250 ;
        RECT 216.450 95.120 218.180 95.130 ;
        RECT 211.660 92.060 213.260 95.120 ;
        RECT 216.580 92.060 218.180 95.120 ;
        RECT 211.660 92.050 213.390 92.060 ;
        RECT 202.850 91.930 213.390 92.050 ;
        RECT 216.450 92.050 218.180 92.060 ;
        RECT 220.920 92.050 222.520 95.130 ;
        RECT 225.260 95.120 230.200 95.130 ;
        RECT 225.260 92.060 226.860 95.120 ;
        RECT 228.590 92.060 230.200 95.120 ;
        RECT 232.420 93.650 235.320 95.250 ;
        RECT 236.920 93.650 239.820 95.250 ;
        RECT 225.260 92.050 230.200 92.060 ;
        RECT 233.720 92.050 238.520 93.650 ;
        RECT 216.450 91.930 235.320 92.050 ;
        RECT 172.440 91.615 235.320 91.930 ;
        RECT 140.300 90.460 235.320 91.615 ;
        RECT 140.300 87.590 141.910 90.460 ;
        RECT 143.520 90.330 167.640 90.460 ;
        RECT 143.520 87.590 154.040 90.330 ;
        RECT 157.120 87.590 167.640 90.330 ;
        RECT 169.250 90.015 174.050 90.460 ;
        RECT 169.250 87.590 170.860 90.015 ;
        RECT 140.300 87.205 170.860 87.590 ;
        RECT 172.440 87.590 174.050 90.015 ;
        RECT 175.660 90.330 226.980 90.460 ;
        RECT 175.660 87.590 186.180 90.330 ;
        RECT 189.260 87.590 199.780 90.330 ;
        RECT 202.860 87.590 213.380 90.330 ;
        RECT 216.460 87.590 226.980 90.330 ;
        RECT 228.590 90.450 235.320 90.460 ;
        RECT 236.920 90.450 239.820 92.050 ;
        RECT 228.590 87.590 230.200 90.450 ;
        RECT 233.720 88.850 238.520 90.450 ;
        RECT 172.440 87.205 230.200 87.590 ;
        RECT 232.420 87.250 235.320 88.850 ;
        RECT 236.920 87.250 239.820 88.850 ;
        RECT 140.300 85.990 230.200 87.205 ;
        RECT 140.300 83.120 141.910 85.990 ;
        RECT 143.520 83.250 154.040 85.990 ;
        RECT 157.120 83.250 167.640 85.990 ;
        RECT 143.520 83.120 167.640 83.250 ;
        RECT 169.250 85.605 174.050 85.990 ;
        RECT 169.250 83.120 170.860 85.605 ;
        RECT 140.300 82.720 170.860 83.120 ;
        RECT 172.440 83.120 174.050 85.605 ;
        RECT 175.660 83.250 186.180 85.990 ;
        RECT 189.260 83.250 199.780 85.990 ;
        RECT 202.860 83.250 213.380 85.990 ;
        RECT 216.460 83.250 226.980 85.990 ;
        RECT 175.660 83.120 226.980 83.250 ;
        RECT 228.590 85.650 230.200 85.990 ;
        RECT 233.720 85.650 238.520 87.250 ;
        RECT 228.590 84.050 235.320 85.650 ;
        RECT 236.920 84.050 239.820 85.650 ;
        RECT 228.590 83.120 230.200 84.050 ;
        RECT 172.440 82.720 230.200 83.120 ;
        RECT 140.300 81.650 230.200 82.720 ;
        RECT 233.720 82.450 238.520 84.050 ;
        RECT 140.300 81.530 154.050 81.650 ;
        RECT 140.300 81.520 145.240 81.530 ;
        RECT 140.300 78.460 141.910 81.520 ;
        RECT 143.640 78.460 145.240 81.520 ;
        RECT 140.300 78.450 145.240 78.460 ;
        RECT 147.980 78.450 149.580 81.530 ;
        RECT 152.320 81.520 154.050 81.530 ;
        RECT 157.110 81.530 186.190 81.650 ;
        RECT 157.110 81.520 158.840 81.530 ;
        RECT 152.320 78.460 153.920 81.520 ;
        RECT 157.240 78.460 158.840 81.520 ;
        RECT 152.320 78.450 154.050 78.460 ;
        RECT 140.300 78.330 154.050 78.450 ;
        RECT 157.110 78.450 158.840 78.460 ;
        RECT 161.580 78.450 163.180 81.530 ;
        RECT 165.920 81.520 177.380 81.530 ;
        RECT 165.920 78.460 167.520 81.520 ;
        RECT 169.250 81.120 174.050 81.520 ;
        RECT 169.250 78.460 170.860 81.120 ;
        RECT 165.920 78.450 170.860 78.460 ;
        RECT 157.110 78.330 170.860 78.450 ;
        RECT 140.300 76.860 170.860 78.330 ;
        RECT 140.300 73.990 141.910 76.860 ;
        RECT 143.520 76.730 167.640 76.860 ;
        RECT 143.520 73.990 154.040 76.730 ;
        RECT 157.120 73.990 167.640 76.730 ;
        RECT 169.250 74.255 170.860 76.860 ;
        RECT 172.440 78.460 174.050 81.120 ;
        RECT 175.780 78.460 177.380 81.520 ;
        RECT 172.440 78.450 177.380 78.460 ;
        RECT 180.120 78.450 181.720 81.530 ;
        RECT 184.460 81.520 186.190 81.530 ;
        RECT 189.250 81.530 199.790 81.650 ;
        RECT 189.250 81.520 190.980 81.530 ;
        RECT 184.460 78.460 186.060 81.520 ;
        RECT 189.380 78.460 190.980 81.520 ;
        RECT 184.460 78.450 186.190 78.460 ;
        RECT 172.440 78.330 186.190 78.450 ;
        RECT 189.250 78.450 190.980 78.460 ;
        RECT 193.720 78.450 195.320 81.530 ;
        RECT 198.060 81.520 199.790 81.530 ;
        RECT 202.850 81.530 213.390 81.650 ;
        RECT 202.850 81.520 204.580 81.530 ;
        RECT 198.060 78.460 199.660 81.520 ;
        RECT 202.980 78.460 204.580 81.520 ;
        RECT 198.060 78.450 199.790 78.460 ;
        RECT 189.250 78.330 199.790 78.450 ;
        RECT 202.850 78.450 204.580 78.460 ;
        RECT 207.320 78.450 208.920 81.530 ;
        RECT 211.660 81.520 213.390 81.530 ;
        RECT 216.450 81.530 230.200 81.650 ;
        RECT 216.450 81.520 218.180 81.530 ;
        RECT 211.660 78.460 213.260 81.520 ;
        RECT 216.580 78.460 218.180 81.520 ;
        RECT 211.660 78.450 213.390 78.460 ;
        RECT 202.850 78.330 213.390 78.450 ;
        RECT 216.450 78.450 218.180 78.460 ;
        RECT 220.920 78.450 222.520 81.530 ;
        RECT 225.260 81.520 230.200 81.530 ;
        RECT 225.260 78.460 226.860 81.520 ;
        RECT 228.590 79.250 230.200 81.520 ;
        RECT 232.420 80.850 235.320 82.450 ;
        RECT 236.920 80.850 239.820 82.450 ;
        RECT 233.720 79.250 238.520 80.850 ;
        RECT 228.590 78.460 235.320 79.250 ;
        RECT 225.260 78.450 235.320 78.460 ;
        RECT 216.450 78.330 235.320 78.450 ;
        RECT 172.440 77.650 235.320 78.330 ;
        RECT 236.920 77.650 239.820 79.250 ;
        RECT 172.440 76.860 230.200 77.650 ;
        RECT 172.440 74.255 174.050 76.860 ;
        RECT 169.250 73.990 174.050 74.255 ;
        RECT 175.660 76.730 226.980 76.860 ;
        RECT 175.660 73.990 186.180 76.730 ;
        RECT 189.260 73.990 199.780 76.730 ;
        RECT 202.860 73.990 213.380 76.730 ;
        RECT 216.460 73.990 226.980 76.730 ;
        RECT 228.590 73.990 230.200 76.860 ;
        RECT 233.720 76.050 238.520 77.650 ;
        RECT 232.420 74.450 235.320 76.050 ;
        RECT 236.920 74.450 239.820 76.050 ;
        RECT 140.300 72.850 230.200 73.990 ;
        RECT 233.720 72.850 238.520 74.450 ;
        RECT 140.300 72.655 235.320 72.850 ;
        RECT 140.300 72.390 170.860 72.655 ;
        RECT 140.300 69.520 141.910 72.390 ;
        RECT 143.520 69.650 154.040 72.390 ;
        RECT 157.120 69.650 167.640 72.390 ;
        RECT 143.520 69.520 167.640 69.650 ;
        RECT 169.250 69.765 170.860 72.390 ;
        RECT 172.440 72.390 235.320 72.655 ;
        RECT 172.440 69.765 174.050 72.390 ;
        RECT 169.250 69.520 174.050 69.765 ;
        RECT 175.660 69.650 186.180 72.390 ;
        RECT 189.260 69.650 199.780 72.390 ;
        RECT 202.860 69.650 213.380 72.390 ;
        RECT 216.460 69.650 226.980 72.390 ;
        RECT 175.660 69.520 226.980 69.650 ;
        RECT 228.590 71.250 235.320 72.390 ;
        RECT 236.920 71.250 239.820 72.850 ;
        RECT 228.590 69.520 230.200 71.250 ;
        RECT 233.720 69.650 238.520 71.250 ;
        RECT 140.300 68.165 230.200 69.520 ;
        RECT 140.300 68.050 170.860 68.165 ;
        RECT 140.300 67.930 154.050 68.050 ;
        RECT 140.300 67.920 145.240 67.930 ;
        RECT 140.300 64.860 141.910 67.920 ;
        RECT 143.640 64.860 145.240 67.920 ;
        RECT 140.300 64.850 145.240 64.860 ;
        RECT 147.980 64.850 149.580 67.930 ;
        RECT 152.320 67.920 154.050 67.930 ;
        RECT 157.110 67.930 170.860 68.050 ;
        RECT 157.110 67.920 158.840 67.930 ;
        RECT 152.320 64.860 153.920 67.920 ;
        RECT 157.240 64.860 158.840 67.920 ;
        RECT 152.320 64.850 154.050 64.860 ;
        RECT 140.300 64.730 154.050 64.850 ;
        RECT 157.110 64.850 158.840 64.860 ;
        RECT 161.580 64.850 163.180 67.930 ;
        RECT 165.920 67.920 170.860 67.930 ;
        RECT 165.920 64.860 167.520 67.920 ;
        RECT 169.250 65.300 170.860 67.920 ;
        RECT 172.440 68.050 230.200 68.165 ;
        RECT 232.420 68.050 235.320 69.650 ;
        RECT 236.920 68.050 239.820 69.650 ;
        RECT 172.440 67.930 186.190 68.050 ;
        RECT 172.440 67.920 177.380 67.930 ;
        RECT 172.440 65.300 174.050 67.920 ;
        RECT 169.250 64.860 174.050 65.300 ;
        RECT 175.780 64.860 177.380 67.920 ;
        RECT 165.920 64.850 177.380 64.860 ;
        RECT 180.120 64.850 181.720 67.930 ;
        RECT 184.460 67.920 186.190 67.930 ;
        RECT 189.250 67.930 199.790 68.050 ;
        RECT 189.250 67.920 190.980 67.930 ;
        RECT 184.460 64.860 186.060 67.920 ;
        RECT 189.380 64.860 190.980 67.920 ;
        RECT 184.460 64.850 186.190 64.860 ;
        RECT 157.110 64.730 186.190 64.850 ;
        RECT 189.250 64.850 190.980 64.860 ;
        RECT 193.720 64.850 195.320 67.930 ;
        RECT 198.060 67.920 199.790 67.930 ;
        RECT 202.850 67.930 213.390 68.050 ;
        RECT 202.850 67.920 204.580 67.930 ;
        RECT 198.060 64.860 199.660 67.920 ;
        RECT 202.980 64.860 204.580 67.920 ;
        RECT 198.060 64.850 199.790 64.860 ;
        RECT 189.250 64.730 199.790 64.850 ;
        RECT 202.850 64.850 204.580 64.860 ;
        RECT 207.320 64.850 208.920 67.930 ;
        RECT 211.660 67.920 213.390 67.930 ;
        RECT 216.450 67.930 230.200 68.050 ;
        RECT 216.450 67.920 218.180 67.930 ;
        RECT 211.660 64.860 213.260 67.920 ;
        RECT 216.580 64.860 218.180 67.920 ;
        RECT 211.660 64.850 213.390 64.860 ;
        RECT 202.850 64.730 213.390 64.850 ;
        RECT 216.450 64.850 218.180 64.860 ;
        RECT 220.920 64.850 222.520 67.930 ;
        RECT 225.260 67.920 230.200 67.930 ;
        RECT 225.260 64.860 226.860 67.920 ;
        RECT 228.590 66.450 230.200 67.920 ;
        RECT 233.720 66.450 238.520 68.050 ;
        RECT 228.590 64.860 235.320 66.450 ;
        RECT 225.260 64.850 235.320 64.860 ;
        RECT 236.920 64.850 239.820 66.450 ;
        RECT 216.450 64.730 230.200 64.850 ;
        RECT 140.300 63.700 230.200 64.730 ;
        RECT 140.300 63.260 170.860 63.700 ;
        RECT 140.300 60.390 141.910 63.260 ;
        RECT 143.520 63.130 167.640 63.260 ;
        RECT 143.520 60.390 154.040 63.130 ;
        RECT 157.120 60.390 167.640 63.130 ;
        RECT 169.250 60.390 170.860 63.260 ;
        RECT 140.300 58.790 170.860 60.390 ;
        RECT 140.300 55.920 141.910 58.790 ;
        RECT 143.520 56.050 154.040 58.790 ;
        RECT 157.120 56.050 167.640 58.790 ;
        RECT 143.520 55.920 167.640 56.050 ;
        RECT 169.250 56.820 170.860 58.790 ;
        RECT 172.440 63.260 230.200 63.700 ;
        RECT 172.440 60.390 174.050 63.260 ;
        RECT 175.660 63.130 226.980 63.260 ;
        RECT 175.660 60.390 186.180 63.130 ;
        RECT 189.260 60.390 199.780 63.130 ;
        RECT 202.860 60.390 213.380 63.130 ;
        RECT 216.460 60.390 226.980 63.130 ;
        RECT 228.590 60.390 230.200 63.260 ;
        RECT 233.720 63.250 238.520 64.850 ;
        RECT 232.420 61.650 235.320 63.250 ;
        RECT 236.920 61.650 239.820 63.250 ;
        RECT 172.440 60.050 230.200 60.390 ;
        RECT 233.720 60.050 238.520 61.650 ;
        RECT 172.440 58.790 235.320 60.050 ;
        RECT 172.440 56.820 174.050 58.790 ;
        RECT 169.250 55.920 174.050 56.820 ;
        RECT 175.660 56.050 186.180 58.790 ;
        RECT 189.260 56.050 199.780 58.790 ;
        RECT 202.860 56.050 213.380 58.790 ;
        RECT 216.460 56.050 226.980 58.790 ;
        RECT 175.660 55.920 226.980 56.050 ;
        RECT 228.590 58.450 235.320 58.790 ;
        RECT 236.920 58.450 239.820 60.050 ;
        RECT 228.590 55.920 230.200 58.450 ;
        RECT 233.720 56.850 238.520 58.450 ;
        RECT 140.300 55.220 230.200 55.920 ;
        RECT 232.420 55.250 235.320 56.850 ;
        RECT 236.920 55.250 239.820 56.850 ;
        RECT 140.300 54.450 170.860 55.220 ;
        RECT 140.300 54.330 154.050 54.450 ;
        RECT 140.300 54.320 145.240 54.330 ;
        RECT 140.300 51.260 141.910 54.320 ;
        RECT 143.640 51.260 145.240 54.320 ;
        RECT 140.300 51.250 145.240 51.260 ;
        RECT 147.980 51.250 149.580 54.330 ;
        RECT 152.320 54.320 154.050 54.330 ;
        RECT 157.110 54.330 170.860 54.450 ;
        RECT 157.110 54.320 158.840 54.330 ;
        RECT 152.320 51.260 153.920 54.320 ;
        RECT 157.240 51.260 158.840 54.320 ;
        RECT 152.320 51.250 154.050 51.260 ;
        RECT 140.300 51.130 154.050 51.250 ;
        RECT 157.110 51.250 158.840 51.260 ;
        RECT 161.580 51.250 163.180 54.330 ;
        RECT 165.920 54.320 170.860 54.330 ;
        RECT 165.920 51.260 167.520 54.320 ;
        RECT 169.250 52.355 170.860 54.320 ;
        RECT 172.440 54.450 230.200 55.220 ;
        RECT 172.440 54.330 186.190 54.450 ;
        RECT 172.440 54.320 177.380 54.330 ;
        RECT 172.440 52.355 174.050 54.320 ;
        RECT 169.250 51.260 174.050 52.355 ;
        RECT 175.780 51.260 177.380 54.320 ;
        RECT 165.920 51.250 177.380 51.260 ;
        RECT 180.120 51.250 181.720 54.330 ;
        RECT 184.460 54.320 186.190 54.330 ;
        RECT 189.250 54.330 199.790 54.450 ;
        RECT 189.250 54.320 190.980 54.330 ;
        RECT 184.460 51.260 186.060 54.320 ;
        RECT 189.380 51.260 190.980 54.320 ;
        RECT 184.460 51.250 186.190 51.260 ;
        RECT 157.110 51.130 186.190 51.250 ;
        RECT 189.250 51.250 190.980 51.260 ;
        RECT 193.720 51.250 195.320 54.330 ;
        RECT 198.060 54.320 199.790 54.330 ;
        RECT 202.850 54.330 213.390 54.450 ;
        RECT 202.850 54.320 204.580 54.330 ;
        RECT 198.060 51.260 199.660 54.320 ;
        RECT 202.980 51.260 204.580 54.320 ;
        RECT 198.060 51.250 199.790 51.260 ;
        RECT 189.250 51.130 199.790 51.250 ;
        RECT 202.850 51.250 204.580 51.260 ;
        RECT 207.320 51.250 208.920 54.330 ;
        RECT 211.660 54.320 213.390 54.330 ;
        RECT 216.450 54.330 230.200 54.450 ;
        RECT 216.450 54.320 218.180 54.330 ;
        RECT 211.660 51.260 213.260 54.320 ;
        RECT 216.580 51.260 218.180 54.320 ;
        RECT 211.660 51.250 213.390 51.260 ;
        RECT 202.850 51.130 213.390 51.250 ;
        RECT 216.450 51.250 218.180 51.260 ;
        RECT 220.920 51.250 222.520 54.330 ;
        RECT 225.260 54.320 230.200 54.330 ;
        RECT 225.260 51.260 226.860 54.320 ;
        RECT 228.590 53.650 230.200 54.320 ;
        RECT 233.720 53.650 238.520 55.250 ;
        RECT 228.590 52.050 235.320 53.650 ;
        RECT 236.920 52.050 239.820 53.650 ;
        RECT 228.590 51.260 230.200 52.050 ;
        RECT 225.260 51.250 230.200 51.260 ;
        RECT 216.450 51.130 230.200 51.250 ;
        RECT 140.300 50.755 230.200 51.130 ;
        RECT 140.300 49.660 170.860 50.755 ;
        RECT 140.300 46.790 141.910 49.660 ;
        RECT 143.520 49.530 167.640 49.660 ;
        RECT 143.520 46.790 154.040 49.530 ;
        RECT 157.120 46.790 167.640 49.530 ;
        RECT 169.250 47.880 170.860 49.660 ;
        RECT 172.440 49.660 230.200 50.755 ;
        RECT 233.720 50.450 238.520 52.050 ;
        RECT 172.440 47.880 174.050 49.660 ;
        RECT 169.250 46.790 174.050 47.880 ;
        RECT 175.660 49.530 226.980 49.660 ;
        RECT 175.660 46.790 186.180 49.530 ;
        RECT 189.260 46.790 199.780 49.530 ;
        RECT 202.860 46.790 213.380 49.530 ;
        RECT 216.460 46.790 226.980 49.530 ;
        RECT 228.590 47.250 230.200 49.660 ;
        RECT 232.420 48.850 235.320 50.450 ;
        RECT 236.920 48.850 239.820 50.450 ;
        RECT 233.720 47.250 238.520 48.850 ;
        RECT 228.590 46.790 235.320 47.250 ;
        RECT 140.300 46.280 235.320 46.790 ;
        RECT 140.300 45.190 170.860 46.280 ;
        RECT 140.300 42.320 141.910 45.190 ;
        RECT 143.520 42.450 154.040 45.190 ;
        RECT 157.120 42.450 167.640 45.190 ;
        RECT 143.520 42.320 167.640 42.450 ;
        RECT 169.250 42.320 170.860 45.190 ;
        RECT 140.300 40.850 170.860 42.320 ;
        RECT 140.300 40.730 154.050 40.850 ;
        RECT 140.300 40.720 145.240 40.730 ;
        RECT 140.300 37.660 141.910 40.720 ;
        RECT 143.640 37.660 145.240 40.720 ;
        RECT 140.300 37.650 145.240 37.660 ;
        RECT 147.980 37.650 149.580 40.730 ;
        RECT 152.320 40.720 154.050 40.730 ;
        RECT 157.110 40.730 170.860 40.850 ;
        RECT 157.110 40.720 158.840 40.730 ;
        RECT 152.320 37.660 153.920 40.720 ;
        RECT 157.240 37.660 158.840 40.720 ;
        RECT 152.320 37.650 154.050 37.660 ;
        RECT 140.300 37.530 154.050 37.650 ;
        RECT 157.110 37.650 158.840 37.660 ;
        RECT 161.580 37.650 163.180 40.730 ;
        RECT 165.920 40.720 170.860 40.730 ;
        RECT 165.920 37.660 167.520 40.720 ;
        RECT 169.250 39.390 170.860 40.720 ;
        RECT 172.440 45.650 235.320 46.280 ;
        RECT 236.920 45.650 239.820 47.250 ;
        RECT 172.440 45.190 230.200 45.650 ;
        RECT 172.440 42.320 174.050 45.190 ;
        RECT 175.660 42.450 186.180 45.190 ;
        RECT 189.260 42.450 199.780 45.190 ;
        RECT 202.860 42.450 213.380 45.190 ;
        RECT 216.460 42.450 226.980 45.190 ;
        RECT 175.660 42.320 226.980 42.450 ;
        RECT 228.590 42.320 230.200 45.190 ;
        RECT 233.720 44.050 238.520 45.650 ;
        RECT 232.420 42.450 235.320 44.050 ;
        RECT 236.920 42.450 239.820 44.050 ;
        RECT 172.440 40.850 230.200 42.320 ;
        RECT 233.720 40.850 238.520 42.450 ;
        RECT 172.440 40.730 186.190 40.850 ;
        RECT 172.440 40.720 177.380 40.730 ;
        RECT 172.440 39.390 174.050 40.720 ;
        RECT 169.250 37.790 174.050 39.390 ;
        RECT 169.250 37.660 170.860 37.790 ;
        RECT 165.920 37.650 170.860 37.660 ;
        RECT 157.110 37.530 170.860 37.650 ;
        RECT 140.300 36.060 170.860 37.530 ;
        RECT 140.300 33.190 141.910 36.060 ;
        RECT 143.520 35.930 167.640 36.060 ;
        RECT 143.520 33.190 154.040 35.930 ;
        RECT 157.120 33.190 167.640 35.930 ;
        RECT 169.250 34.925 170.860 36.060 ;
        RECT 172.440 37.660 174.050 37.790 ;
        RECT 175.780 37.660 177.380 40.720 ;
        RECT 172.440 37.650 177.380 37.660 ;
        RECT 180.120 37.650 181.720 40.730 ;
        RECT 184.460 40.720 186.190 40.730 ;
        RECT 189.250 40.730 199.790 40.850 ;
        RECT 189.250 40.720 190.980 40.730 ;
        RECT 184.460 37.660 186.060 40.720 ;
        RECT 189.380 37.660 190.980 40.720 ;
        RECT 184.460 37.650 186.190 37.660 ;
        RECT 172.440 37.530 186.190 37.650 ;
        RECT 189.250 37.650 190.980 37.660 ;
        RECT 193.720 37.650 195.320 40.730 ;
        RECT 198.060 40.720 199.790 40.730 ;
        RECT 202.850 40.730 213.390 40.850 ;
        RECT 202.850 40.720 204.580 40.730 ;
        RECT 198.060 37.660 199.660 40.720 ;
        RECT 202.980 37.660 204.580 40.720 ;
        RECT 198.060 37.650 199.790 37.660 ;
        RECT 189.250 37.530 199.790 37.650 ;
        RECT 202.850 37.650 204.580 37.660 ;
        RECT 207.320 37.650 208.920 40.730 ;
        RECT 211.660 40.720 213.390 40.730 ;
        RECT 216.450 40.730 235.320 40.850 ;
        RECT 216.450 40.720 218.180 40.730 ;
        RECT 211.660 37.660 213.260 40.720 ;
        RECT 216.580 37.660 218.180 40.720 ;
        RECT 211.660 37.650 213.390 37.660 ;
        RECT 202.850 37.530 213.390 37.650 ;
        RECT 216.450 37.650 218.180 37.660 ;
        RECT 220.920 37.650 222.520 40.730 ;
        RECT 225.260 40.720 235.320 40.730 ;
        RECT 225.260 37.660 226.860 40.720 ;
        RECT 228.590 39.250 235.320 40.720 ;
        RECT 236.920 39.250 239.820 40.850 ;
        RECT 228.590 37.660 230.200 39.250 ;
        RECT 225.260 37.650 230.200 37.660 ;
        RECT 233.720 37.650 238.520 39.250 ;
        RECT 216.450 37.530 230.200 37.650 ;
        RECT 172.440 36.060 230.200 37.530 ;
        RECT 172.440 34.925 174.050 36.060 ;
        RECT 169.250 33.325 174.050 34.925 ;
        RECT 169.250 33.190 170.860 33.325 ;
        RECT 140.300 31.590 170.860 33.190 ;
        RECT 140.300 28.720 141.910 31.590 ;
        RECT 143.520 28.850 154.040 31.590 ;
        RECT 157.120 28.850 167.640 31.590 ;
        RECT 143.520 28.720 167.640 28.850 ;
        RECT 169.250 30.465 170.860 31.590 ;
        RECT 172.440 33.190 174.050 33.325 ;
        RECT 175.660 35.930 226.980 36.060 ;
        RECT 175.660 33.190 186.180 35.930 ;
        RECT 189.260 33.190 199.780 35.930 ;
        RECT 202.860 33.190 213.380 35.930 ;
        RECT 216.460 33.190 226.980 35.930 ;
        RECT 228.590 34.450 230.200 36.060 ;
        RECT 232.420 36.050 235.320 37.650 ;
        RECT 236.920 36.050 239.820 37.650 ;
        RECT 233.720 34.450 238.520 36.050 ;
        RECT 228.590 33.190 235.320 34.450 ;
        RECT 172.440 32.850 235.320 33.190 ;
        RECT 236.920 32.850 239.820 34.450 ;
        RECT 172.440 31.590 230.200 32.850 ;
        RECT 172.440 30.465 174.050 31.590 ;
        RECT 169.250 28.865 174.050 30.465 ;
        RECT 169.250 28.720 170.860 28.865 ;
        RECT 140.300 27.250 170.860 28.720 ;
        RECT 140.300 27.130 154.050 27.250 ;
        RECT 140.300 27.120 145.240 27.130 ;
        RECT 140.300 24.060 141.910 27.120 ;
        RECT 143.640 24.060 145.240 27.120 ;
        RECT 140.300 24.050 145.240 24.060 ;
        RECT 147.980 24.050 149.580 27.130 ;
        RECT 152.320 27.120 154.050 27.130 ;
        RECT 157.110 27.130 170.860 27.250 ;
        RECT 157.110 27.120 158.840 27.130 ;
        RECT 152.320 24.060 153.920 27.120 ;
        RECT 157.240 24.060 158.840 27.120 ;
        RECT 152.320 24.050 154.050 24.060 ;
        RECT 140.300 23.930 154.050 24.050 ;
        RECT 157.110 24.050 158.840 24.060 ;
        RECT 161.580 24.050 163.180 27.130 ;
        RECT 165.920 27.120 170.860 27.130 ;
        RECT 165.920 24.060 167.520 27.120 ;
        RECT 169.250 24.060 170.860 27.120 ;
        RECT 165.920 24.050 170.860 24.060 ;
        RECT 157.110 23.930 170.860 24.050 ;
        RECT 140.300 22.460 170.860 23.930 ;
        RECT 140.300 19.595 141.910 22.460 ;
        RECT 143.520 22.330 167.640 22.460 ;
        RECT 143.520 19.595 154.040 22.330 ;
        RECT 140.300 19.590 154.040 19.595 ;
        RECT 157.120 19.800 167.640 22.330 ;
        RECT 169.250 21.985 170.860 22.460 ;
        RECT 172.440 28.720 174.050 28.865 ;
        RECT 175.660 28.850 186.180 31.590 ;
        RECT 189.260 28.850 199.780 31.590 ;
        RECT 202.860 28.850 213.380 31.590 ;
        RECT 216.460 28.850 226.980 31.590 ;
        RECT 175.660 28.720 226.980 28.850 ;
        RECT 228.590 28.720 230.200 31.590 ;
        RECT 233.720 31.250 238.520 32.850 ;
        RECT 232.420 29.650 235.320 31.250 ;
        RECT 236.920 29.650 239.820 31.250 ;
        RECT 172.440 28.050 230.200 28.720 ;
        RECT 233.720 28.050 238.520 29.650 ;
        RECT 172.440 27.250 235.320 28.050 ;
        RECT 172.440 27.130 186.190 27.250 ;
        RECT 172.440 27.120 177.380 27.130 ;
        RECT 172.440 24.060 174.050 27.120 ;
        RECT 175.780 24.060 177.380 27.120 ;
        RECT 172.440 24.050 177.380 24.060 ;
        RECT 180.120 24.050 181.720 27.130 ;
        RECT 184.460 27.120 186.190 27.130 ;
        RECT 189.250 27.130 199.790 27.250 ;
        RECT 189.250 27.120 190.980 27.130 ;
        RECT 184.460 24.060 186.060 27.120 ;
        RECT 189.380 24.060 190.980 27.120 ;
        RECT 184.460 24.050 186.190 24.060 ;
        RECT 172.440 23.930 186.190 24.050 ;
        RECT 189.250 24.050 190.980 24.060 ;
        RECT 193.720 24.050 195.320 27.130 ;
        RECT 198.060 27.120 199.790 27.130 ;
        RECT 202.850 27.130 213.390 27.250 ;
        RECT 202.850 27.120 204.580 27.130 ;
        RECT 198.060 24.060 199.660 27.120 ;
        RECT 202.980 24.060 204.580 27.120 ;
        RECT 198.060 24.050 199.790 24.060 ;
        RECT 189.250 23.930 199.790 24.050 ;
        RECT 202.850 24.050 204.580 24.060 ;
        RECT 207.320 24.050 208.920 27.130 ;
        RECT 211.660 27.120 213.390 27.130 ;
        RECT 216.450 27.130 235.320 27.250 ;
        RECT 216.450 27.120 218.180 27.130 ;
        RECT 211.660 24.060 213.260 27.120 ;
        RECT 216.580 24.060 218.180 27.120 ;
        RECT 211.660 24.050 213.390 24.060 ;
        RECT 202.850 23.930 213.390 24.050 ;
        RECT 216.450 24.050 218.180 24.060 ;
        RECT 220.920 24.050 222.520 27.130 ;
        RECT 225.260 27.120 235.320 27.130 ;
        RECT 225.260 24.060 226.860 27.120 ;
        RECT 228.590 26.450 235.320 27.120 ;
        RECT 236.920 26.450 239.820 28.050 ;
        RECT 228.590 24.060 230.200 26.450 ;
        RECT 233.720 24.850 238.520 26.450 ;
        RECT 225.260 24.050 230.200 24.060 ;
        RECT 216.450 23.930 230.200 24.050 ;
        RECT 172.440 22.460 230.200 23.930 ;
        RECT 232.420 23.250 235.320 24.850 ;
        RECT 236.920 23.250 239.820 24.850 ;
        RECT 172.440 21.985 174.050 22.460 ;
        RECT 169.250 20.385 174.050 21.985 ;
        RECT 169.250 19.800 170.860 20.385 ;
        RECT 157.120 19.590 170.860 19.800 ;
        RECT 140.300 18.195 170.860 19.590 ;
        RECT 140.300 17.995 167.640 18.195 ;
        RECT 140.300 15.130 141.910 17.995 ;
        RECT 143.520 17.990 167.640 17.995 ;
        RECT 143.520 15.250 154.040 17.990 ;
        RECT 157.120 15.530 167.640 17.990 ;
        RECT 169.250 17.515 170.860 18.195 ;
        RECT 172.440 19.595 174.050 20.385 ;
        RECT 175.660 22.330 226.980 22.460 ;
        RECT 175.660 19.595 186.180 22.330 ;
        RECT 172.440 19.590 186.180 19.595 ;
        RECT 189.260 19.590 199.780 22.330 ;
        RECT 202.860 19.590 213.380 22.330 ;
        RECT 216.460 19.800 226.980 22.330 ;
        RECT 228.590 21.650 230.200 22.460 ;
        RECT 233.720 21.650 238.520 23.250 ;
        RECT 228.590 20.050 235.320 21.650 ;
        RECT 236.920 20.050 239.820 21.650 ;
        RECT 228.590 19.800 230.200 20.050 ;
        RECT 216.460 19.590 230.200 19.800 ;
        RECT 172.440 18.195 230.200 19.590 ;
        RECT 233.720 18.450 238.520 20.050 ;
        RECT 172.440 17.995 226.980 18.195 ;
        RECT 172.440 17.515 174.050 17.995 ;
        RECT 169.250 15.915 174.050 17.515 ;
        RECT 169.250 15.530 170.860 15.915 ;
        RECT 157.120 15.250 170.860 15.530 ;
        RECT 143.520 15.130 170.860 15.250 ;
        RECT 140.300 13.930 170.860 15.130 ;
        RECT 140.300 13.650 167.640 13.930 ;
        RECT 140.300 13.530 154.050 13.650 ;
        RECT 140.300 11.920 141.910 13.530 ;
        RECT 143.920 11.920 145.520 13.530 ;
        RECT 148.185 11.920 149.790 13.530 ;
        RECT 152.450 11.920 154.050 13.530 ;
        RECT 157.110 13.530 167.640 13.650 ;
        RECT 157.110 11.920 158.710 13.530 ;
        RECT 161.575 11.920 163.175 13.530 ;
        RECT 166.040 11.920 167.640 13.530 ;
        RECT 169.250 13.045 170.860 13.930 ;
        RECT 172.440 15.130 174.050 15.915 ;
        RECT 175.660 17.990 226.980 17.995 ;
        RECT 175.660 15.250 186.180 17.990 ;
        RECT 189.260 15.250 199.780 17.990 ;
        RECT 202.860 15.250 213.380 17.990 ;
        RECT 216.460 15.530 226.980 17.990 ;
        RECT 228.590 15.530 230.200 18.195 ;
        RECT 232.420 16.850 235.320 18.450 ;
        RECT 236.920 16.850 239.820 18.450 ;
        RECT 216.460 15.250 230.200 15.530 ;
        RECT 233.720 15.250 238.520 16.850 ;
        RECT 175.660 15.130 235.320 15.250 ;
        RECT 172.440 13.930 235.320 15.130 ;
        RECT 172.440 13.650 226.980 13.930 ;
        RECT 172.440 13.530 186.190 13.650 ;
        RECT 172.440 13.045 174.050 13.530 ;
        RECT 169.250 11.920 174.050 13.045 ;
        RECT 176.060 11.920 177.660 13.530 ;
        RECT 180.325 11.920 181.930 13.530 ;
        RECT 184.590 11.920 186.190 13.530 ;
        RECT 189.250 13.530 199.790 13.650 ;
        RECT 189.250 11.920 190.850 13.530 ;
        RECT 193.720 11.920 195.320 13.530 ;
        RECT 198.190 11.920 199.790 13.530 ;
        RECT 202.850 13.530 213.390 13.650 ;
        RECT 202.850 11.920 204.450 13.530 ;
        RECT 207.320 11.920 208.920 13.530 ;
        RECT 211.790 11.920 213.390 13.530 ;
        RECT 216.450 13.530 226.980 13.650 ;
        RECT 216.450 11.920 218.050 13.530 ;
        RECT 220.915 11.920 222.515 13.530 ;
        RECT 225.380 11.920 226.980 13.530 ;
        RECT 228.590 13.650 235.320 13.930 ;
        RECT 228.590 11.920 230.200 13.650 ;
        RECT 140.300 11.445 230.200 11.920 ;
        RECT 140.300 10.310 170.860 11.445 ;
        RECT 172.440 10.310 230.200 11.445 ;
        RECT 233.720 10.850 235.320 13.650 ;
        RECT 236.920 13.650 239.820 15.250 ;
        RECT 236.920 10.850 238.520 13.650 ;
        RECT 9.570 6.100 11.170 7.400 ;
        RECT 12.770 6.100 14.370 10.310 ;
        RECT 15.970 6.100 17.570 7.400 ;
        RECT 19.170 6.100 20.770 10.310 ;
        RECT 22.370 6.100 23.970 7.400 ;
        RECT 25.570 6.100 27.170 10.310 ;
        RECT 28.770 6.100 30.370 7.400 ;
        RECT 31.970 6.100 33.570 10.310 ;
        RECT 35.170 6.100 36.770 7.400 ;
        RECT 38.370 6.100 39.970 10.310 ;
        RECT 41.570 6.100 43.170 7.400 ;
        RECT 44.770 6.100 46.370 10.310 ;
        RECT 47.970 6.100 49.570 7.400 ;
        RECT 51.170 6.100 52.770 10.310 ;
        RECT 54.370 6.100 55.970 7.400 ;
        RECT 57.570 6.100 59.170 10.310 ;
        RECT 60.770 6.100 62.370 7.400 ;
        RECT 63.970 6.100 65.570 10.310 ;
        RECT 67.170 6.100 68.770 7.400 ;
        RECT 70.370 6.100 71.970 10.310 ;
        RECT 73.570 6.100 75.170 7.400 ;
        RECT 76.770 6.100 78.370 7.400 ;
        RECT 79.970 6.100 81.570 7.400 ;
        RECT 83.170 6.100 84.770 10.310 ;
        RECT 86.370 6.100 87.970 7.400 ;
        RECT 89.570 6.100 91.170 10.310 ;
        RECT 92.770 6.100 94.370 7.400 ;
        RECT 95.970 6.100 97.570 10.310 ;
        RECT 99.170 6.100 100.770 7.400 ;
        RECT 102.370 6.100 103.970 7.400 ;
        RECT 105.570 6.100 107.170 7.400 ;
        RECT 108.770 6.100 110.370 7.400 ;
        RECT 111.970 6.100 113.570 7.400 ;
        RECT 115.170 6.100 116.770 7.400 ;
        RECT 123.610 6.100 125.210 7.400 ;
        RECT 126.810 6.100 128.410 7.400 ;
        RECT 130.010 6.100 131.610 7.400 ;
        RECT 133.210 6.100 134.810 7.400 ;
        RECT 136.410 6.100 138.010 7.400 ;
        RECT 139.610 6.100 141.210 7.400 ;
        RECT 142.810 6.100 144.410 10.310 ;
        RECT 146.010 6.100 147.610 7.400 ;
        RECT 149.210 6.100 150.810 10.310 ;
        RECT 152.410 6.100 154.010 7.400 ;
        RECT 155.610 6.100 157.210 10.310 ;
        RECT 158.810 6.100 160.410 7.400 ;
        RECT 162.010 6.100 163.610 7.400 ;
        RECT 165.210 6.100 166.810 7.400 ;
        RECT 168.410 6.100 170.010 10.310 ;
        RECT 171.610 6.100 173.210 7.400 ;
        RECT 174.810 6.100 176.410 10.310 ;
        RECT 178.010 6.100 179.610 7.400 ;
        RECT 181.210 6.100 182.810 10.310 ;
        RECT 184.410 6.100 186.010 7.400 ;
        RECT 187.610 6.100 189.210 10.310 ;
        RECT 190.810 6.100 192.410 7.400 ;
        RECT 194.010 6.100 195.610 10.310 ;
        RECT 197.210 6.100 198.810 7.400 ;
        RECT 200.410 6.100 202.010 10.310 ;
        RECT 203.610 6.100 205.210 7.400 ;
        RECT 206.810 6.100 208.410 10.310 ;
        RECT 210.010 6.100 211.610 7.400 ;
        RECT 213.210 6.100 214.810 10.310 ;
        RECT 216.410 6.100 218.010 7.400 ;
        RECT 219.610 6.100 221.210 10.310 ;
        RECT 222.810 6.100 224.410 7.400 ;
        RECT 226.010 6.100 227.610 10.310 ;
        RECT 229.210 6.100 230.810 7.400 ;
        RECT 6.710 4.500 233.670 6.100 ;
        RECT 7.970 2.900 9.570 4.500 ;
        RECT 11.170 2.900 12.770 4.500 ;
        RECT 14.370 2.900 15.970 4.500 ;
        RECT 17.570 2.900 19.170 4.500 ;
        RECT 20.770 2.900 22.370 4.500 ;
        RECT 23.970 2.900 25.570 4.500 ;
        RECT 27.170 2.900 28.770 4.500 ;
        RECT 30.370 2.900 31.970 4.500 ;
        RECT 33.570 2.900 35.170 4.500 ;
        RECT 36.770 2.900 38.370 4.500 ;
        RECT 39.970 2.900 41.570 4.500 ;
        RECT 43.170 2.900 44.770 4.500 ;
        RECT 46.370 2.900 47.970 4.500 ;
        RECT 49.570 2.900 51.170 4.500 ;
        RECT 52.770 2.900 54.370 4.500 ;
        RECT 55.970 2.900 57.570 4.500 ;
        RECT 59.170 2.900 60.770 4.500 ;
        RECT 62.370 2.900 63.970 4.500 ;
        RECT 65.570 2.900 67.170 4.500 ;
        RECT 68.770 2.900 70.370 4.500 ;
        RECT 71.970 2.900 73.570 4.500 ;
        RECT 75.170 2.900 76.770 4.500 ;
        RECT 78.370 2.900 79.970 4.500 ;
        RECT 81.570 2.900 83.170 4.500 ;
        RECT 84.770 2.900 86.370 4.500 ;
        RECT 87.970 2.900 89.570 4.500 ;
        RECT 91.170 2.900 92.770 4.500 ;
        RECT 94.370 2.900 95.970 4.500 ;
        RECT 97.570 2.900 99.170 4.500 ;
        RECT 100.770 2.900 102.370 4.500 ;
        RECT 103.970 2.900 105.570 4.500 ;
        RECT 107.170 2.900 108.770 4.500 ;
        RECT 110.370 2.900 111.970 4.500 ;
        RECT 113.570 2.900 115.170 4.500 ;
        RECT 116.770 2.900 118.370 4.500 ;
        RECT 122.010 2.900 123.610 4.500 ;
        RECT 125.210 2.900 126.810 4.500 ;
        RECT 128.410 2.900 130.010 4.500 ;
        RECT 131.610 2.900 133.210 4.500 ;
        RECT 134.810 2.900 136.410 4.500 ;
        RECT 138.010 2.900 139.610 4.500 ;
        RECT 141.210 2.900 142.810 4.500 ;
        RECT 144.410 2.900 146.010 4.500 ;
        RECT 147.610 2.900 149.210 4.500 ;
        RECT 150.810 2.900 152.410 4.500 ;
        RECT 154.010 2.900 155.610 4.500 ;
        RECT 157.210 2.900 158.810 4.500 ;
        RECT 160.410 2.900 162.010 4.500 ;
        RECT 163.610 2.900 165.210 4.500 ;
        RECT 166.810 2.900 168.410 4.500 ;
        RECT 170.010 2.900 171.610 4.500 ;
        RECT 173.210 2.900 174.810 4.500 ;
        RECT 176.410 2.900 178.010 4.500 ;
        RECT 179.610 2.900 181.210 4.500 ;
        RECT 182.810 2.900 184.410 4.500 ;
        RECT 186.010 2.900 187.610 4.500 ;
        RECT 189.210 2.900 190.810 4.500 ;
        RECT 192.410 2.900 194.010 4.500 ;
        RECT 195.610 2.900 197.210 4.500 ;
        RECT 198.810 2.900 200.410 4.500 ;
        RECT 202.010 2.900 203.610 4.500 ;
        RECT 205.210 2.900 206.810 4.500 ;
        RECT 208.410 2.900 210.010 4.500 ;
        RECT 211.610 2.900 213.210 4.500 ;
        RECT 214.810 2.900 216.410 4.500 ;
        RECT 218.010 2.900 219.610 4.500 ;
        RECT 221.210 2.900 222.810 4.500 ;
        RECT 224.410 2.900 226.010 4.500 ;
        RECT 227.610 2.900 229.210 4.500 ;
        RECT 230.810 2.900 232.410 4.500 ;
        RECT 3.505 1.300 236.875 2.900 ;
        RECT 9.570 0.000 11.170 1.300 ;
        RECT 12.770 0.000 14.370 1.300 ;
        RECT 15.970 0.000 17.570 1.300 ;
        RECT 19.170 0.000 20.770 1.300 ;
        RECT 22.370 0.000 23.970 1.300 ;
        RECT 25.570 0.000 27.170 1.300 ;
        RECT 28.770 0.000 30.370 1.300 ;
        RECT 31.970 0.000 33.570 1.300 ;
        RECT 35.170 0.000 36.770 1.300 ;
        RECT 38.370 0.000 39.970 1.300 ;
        RECT 41.570 0.000 43.170 1.300 ;
        RECT 44.770 0.000 46.370 1.300 ;
        RECT 47.970 0.000 49.570 1.300 ;
        RECT 51.170 0.000 52.770 1.300 ;
        RECT 54.370 0.000 55.970 1.300 ;
        RECT 57.570 0.000 59.170 1.300 ;
        RECT 60.770 0.000 62.370 1.300 ;
        RECT 63.970 0.000 65.570 1.300 ;
        RECT 67.170 0.000 68.770 1.300 ;
        RECT 70.370 0.000 71.970 1.300 ;
        RECT 73.570 0.000 75.170 1.300 ;
        RECT 76.770 0.000 78.370 1.300 ;
        RECT 79.970 0.000 81.570 1.300 ;
        RECT 83.170 0.000 84.770 1.300 ;
        RECT 86.370 0.000 87.970 1.300 ;
        RECT 89.570 0.000 91.170 1.300 ;
        RECT 92.770 0.000 94.370 1.300 ;
        RECT 95.970 0.000 97.570 1.300 ;
        RECT 99.170 0.000 100.770 1.300 ;
        RECT 102.370 0.000 103.970 1.300 ;
        RECT 105.570 0.000 107.170 1.300 ;
        RECT 108.770 0.000 110.370 1.300 ;
        RECT 111.970 0.000 113.570 1.300 ;
        RECT 115.170 0.000 116.770 1.300 ;
        RECT 123.610 0.000 125.210 1.300 ;
        RECT 126.810 0.000 128.410 1.300 ;
        RECT 130.010 0.000 131.610 1.300 ;
        RECT 133.210 0.000 134.810 1.300 ;
        RECT 136.410 0.000 138.010 1.300 ;
        RECT 139.610 0.000 141.210 1.300 ;
        RECT 142.810 0.000 144.410 1.300 ;
        RECT 146.010 0.000 147.610 1.300 ;
        RECT 149.210 0.000 150.810 1.300 ;
        RECT 152.410 0.000 154.010 1.300 ;
        RECT 155.610 0.000 157.210 1.300 ;
        RECT 158.810 0.000 160.410 1.300 ;
        RECT 162.010 0.000 163.610 1.300 ;
        RECT 165.210 0.000 166.810 1.300 ;
        RECT 168.410 0.000 170.010 1.300 ;
        RECT 171.610 0.000 173.210 1.300 ;
        RECT 174.810 0.000 176.410 1.300 ;
        RECT 178.010 0.000 179.610 1.300 ;
        RECT 181.210 0.000 182.810 1.300 ;
        RECT 184.410 0.000 186.010 1.300 ;
        RECT 187.610 0.000 189.210 1.300 ;
        RECT 190.810 0.000 192.410 1.300 ;
        RECT 194.010 0.000 195.610 1.300 ;
        RECT 197.210 0.000 198.810 1.300 ;
        RECT 200.410 0.000 202.010 1.300 ;
        RECT 203.610 0.000 205.210 1.300 ;
        RECT 206.810 0.000 208.410 1.300 ;
        RECT 210.010 0.000 211.610 1.300 ;
        RECT 213.210 0.000 214.810 1.300 ;
        RECT 216.410 0.000 218.010 1.300 ;
        RECT 219.610 0.000 221.210 1.300 ;
        RECT 222.810 0.000 224.410 1.300 ;
        RECT 226.010 0.000 227.610 1.300 ;
        RECT 229.210 0.000 230.810 1.300 ;
      LAYER via3 ;
        RECT 105.480 173.120 105.800 173.440 ;
        RECT 110.015 172.900 110.335 173.220 ;
        RECT 114.745 172.895 115.065 173.215 ;
        RECT 95.490 169.095 95.810 169.415 ;
        RECT 105.510 167.605 105.830 167.925 ;
        RECT 110.150 167.455 110.470 167.775 ;
        RECT 114.755 167.455 115.075 167.775 ;
        RECT 97.540 166.355 98.200 166.725 ;
        RECT 95.505 163.680 95.825 164.000 ;
        RECT 105.535 162.200 105.855 162.520 ;
        RECT 110.135 162.010 110.455 162.330 ;
        RECT 114.745 162.010 115.065 162.330 ;
        RECT 114.700 147.825 115.070 148.180 ;
        RECT 0.685 125.865 1.855 127.035 ;
        RECT 6.665 125.865 7.835 127.035 ;
        RECT 3.465 124.265 5.055 125.435 ;
        RECT 0.685 122.665 1.855 123.835 ;
        RECT 6.665 122.665 7.835 123.835 ;
        RECT 232.545 125.865 233.715 127.035 ;
        RECT 238.525 125.865 239.695 127.035 ;
        RECT 235.325 124.265 236.915 125.435 ;
        RECT 232.545 122.665 233.715 123.835 ;
        RECT 3.465 121.065 5.055 122.235 ;
        RECT 0.685 119.465 1.855 120.635 ;
        RECT 6.665 119.465 7.835 120.635 ;
        RECT 3.465 117.865 5.055 119.035 ;
        RECT 10.345 121.015 19.670 122.305 ;
        RECT 22.330 121.015 24.530 122.305 ;
        RECT 26.390 121.015 38.120 122.305 ;
        RECT 39.990 121.015 51.720 122.305 ;
        RECT 53.590 121.015 60.255 122.305 ;
        RECT 63.120 121.015 67.775 122.305 ;
        RECT 10.345 117.650 11.635 121.015 ;
        RECT 0.685 116.265 1.855 117.435 ;
        RECT 6.665 116.265 7.835 117.435 ;
        RECT 3.465 114.665 5.055 115.835 ;
        RECT 0.685 113.065 1.855 114.235 ;
        RECT 6.665 113.065 7.835 114.235 ;
        RECT 3.465 111.465 5.055 112.635 ;
        RECT 0.685 109.865 1.855 111.035 ;
        RECT 6.665 109.865 7.835 111.035 ;
        RECT 3.465 108.265 5.055 109.435 ;
        RECT 10.345 108.120 11.635 114.785 ;
        RECT 66.485 112.980 67.775 121.015 ;
        RECT 69.685 121.015 79.010 122.305 ;
        RECT 81.670 121.015 83.870 122.305 ;
        RECT 85.730 121.015 92.395 122.305 ;
        RECT 95.260 121.015 99.915 122.305 ;
        RECT 69.685 117.650 70.975 121.015 ;
        RECT 0.685 106.665 1.855 107.835 ;
        RECT 6.665 106.665 7.835 107.835 ;
        RECT 3.465 105.065 5.055 106.235 ;
        RECT 0.685 103.465 1.855 104.635 ;
        RECT 6.665 103.465 7.835 104.635 ;
        RECT 3.465 101.865 5.055 103.035 ;
        RECT 0.685 100.265 1.855 101.435 ;
        RECT 6.665 100.265 7.835 101.435 ;
        RECT 3.465 98.665 5.055 99.835 ;
        RECT 0.685 97.065 1.855 98.235 ;
        RECT 6.665 97.065 7.835 98.235 ;
        RECT 3.465 95.465 5.055 96.635 ;
        RECT 0.685 93.865 1.855 95.035 ;
        RECT 6.665 93.865 7.835 95.035 ;
        RECT 10.345 94.520 11.635 106.250 ;
        RECT 66.485 108.120 67.775 110.320 ;
        RECT 69.685 108.120 70.975 114.785 ;
        RECT 98.625 112.980 99.915 121.015 ;
        RECT 3.465 92.265 5.055 93.435 ;
        RECT 0.685 90.665 1.855 91.835 ;
        RECT 6.665 90.665 7.835 91.835 ;
        RECT 3.465 89.065 5.055 90.235 ;
        RECT 0.685 87.465 1.855 88.635 ;
        RECT 6.665 87.465 7.835 88.635 ;
        RECT 3.465 85.865 5.055 87.035 ;
        RECT 0.685 84.265 1.855 85.435 ;
        RECT 6.665 84.265 7.835 85.435 ;
        RECT 3.465 82.665 5.055 83.835 ;
        RECT 0.685 81.065 1.855 82.235 ;
        RECT 6.665 81.065 7.835 82.235 ;
        RECT 10.345 80.920 11.635 92.650 ;
        RECT 66.485 94.530 67.775 106.260 ;
        RECT 3.465 79.465 5.055 80.635 ;
        RECT 0.685 77.865 1.855 79.035 ;
        RECT 6.665 77.865 7.835 79.035 ;
        RECT 3.465 76.265 5.055 77.435 ;
        RECT 0.685 74.665 1.855 75.835 ;
        RECT 6.665 74.665 7.835 75.835 ;
        RECT 3.465 73.065 5.055 74.235 ;
        RECT 0.685 71.465 1.855 72.635 ;
        RECT 6.665 71.465 7.835 72.635 ;
        RECT 3.465 69.865 5.055 71.035 ;
        RECT 0.685 68.265 1.855 69.435 ;
        RECT 6.665 68.265 7.835 69.435 ;
        RECT 3.465 66.665 5.055 67.835 ;
        RECT 10.345 67.320 11.635 79.050 ;
        RECT 66.485 80.930 67.775 92.660 ;
        RECT 69.685 94.520 70.975 106.250 ;
        RECT 98.625 108.120 99.915 110.320 ;
        RECT 0.685 65.065 1.855 66.235 ;
        RECT 6.665 65.065 7.835 66.235 ;
        RECT 3.465 63.465 5.055 64.635 ;
        RECT 0.685 61.865 1.855 63.035 ;
        RECT 6.665 61.865 7.835 63.035 ;
        RECT 3.465 60.265 5.055 61.435 ;
        RECT 0.685 58.665 1.855 59.835 ;
        RECT 6.665 58.665 7.835 59.835 ;
        RECT 3.465 57.065 5.055 58.235 ;
        RECT 0.685 55.465 1.855 56.635 ;
        RECT 6.665 55.465 7.835 56.635 ;
        RECT 3.465 53.865 5.055 55.035 ;
        RECT 10.345 53.720 11.635 65.450 ;
        RECT 66.485 67.330 67.775 79.060 ;
        RECT 69.685 80.920 70.975 92.650 ;
        RECT 98.625 94.530 99.915 106.260 ;
        RECT 0.685 52.265 1.855 53.435 ;
        RECT 6.665 52.265 7.835 53.435 ;
        RECT 3.465 50.665 5.055 51.835 ;
        RECT 0.685 49.065 1.855 50.235 ;
        RECT 6.665 49.065 7.835 50.235 ;
        RECT 3.465 47.465 5.055 48.635 ;
        RECT 0.685 45.865 1.855 47.035 ;
        RECT 6.665 45.865 7.835 47.035 ;
        RECT 3.465 44.265 5.055 45.435 ;
        RECT 0.685 42.665 1.855 43.835 ;
        RECT 6.665 42.665 7.835 43.835 ;
        RECT 3.465 41.065 5.055 42.235 ;
        RECT 0.685 39.465 1.855 40.635 ;
        RECT 6.665 39.465 7.835 40.635 ;
        RECT 10.345 40.120 11.635 51.850 ;
        RECT 66.485 53.730 67.775 65.460 ;
        RECT 69.685 67.320 70.975 79.050 ;
        RECT 98.625 80.930 99.915 92.660 ;
        RECT 69.685 53.720 70.975 65.450 ;
        RECT 98.625 67.330 99.915 79.060 ;
        RECT 3.465 37.865 5.055 39.035 ;
        RECT 0.685 36.265 1.855 37.435 ;
        RECT 6.665 36.265 7.835 37.435 ;
        RECT 3.465 34.665 5.055 35.835 ;
        RECT 0.685 33.065 1.855 34.235 ;
        RECT 6.665 33.065 7.835 34.235 ;
        RECT 3.465 31.465 5.055 32.635 ;
        RECT 0.685 29.865 1.855 31.035 ;
        RECT 6.665 29.865 7.835 31.035 ;
        RECT 3.465 28.265 5.055 29.435 ;
        RECT 0.685 26.665 1.855 27.835 ;
        RECT 6.665 26.665 7.835 27.835 ;
        RECT 10.345 26.520 11.635 38.250 ;
        RECT 66.485 40.130 67.775 51.860 ;
        RECT 69.685 40.120 70.975 51.850 ;
        RECT 98.625 53.730 99.915 65.460 ;
        RECT 3.465 25.065 5.055 26.235 ;
        RECT 0.685 23.465 1.855 24.635 ;
        RECT 6.665 23.465 7.835 24.635 ;
        RECT 3.465 21.865 5.055 23.035 ;
        RECT 10.345 22.460 11.635 24.660 ;
        RECT 66.485 26.530 67.775 38.260 ;
        RECT 0.685 20.265 1.855 21.435 ;
        RECT 6.665 20.265 7.835 21.435 ;
        RECT 3.465 18.665 5.055 19.835 ;
        RECT 0.685 17.065 1.855 18.235 ;
        RECT 6.665 17.065 7.835 18.235 ;
        RECT 3.465 15.465 5.055 16.635 ;
        RECT 0.685 13.865 1.855 15.035 ;
        RECT 6.665 13.865 7.835 15.035 ;
        RECT 10.345 11.765 11.635 19.800 ;
        RECT 66.485 17.995 67.775 24.660 ;
        RECT 69.685 26.520 70.975 38.250 ;
        RECT 98.625 40.130 99.915 51.860 ;
        RECT 69.685 22.460 70.975 24.660 ;
        RECT 98.625 26.530 99.915 38.260 ;
        RECT 66.485 11.765 67.775 15.130 ;
        RECT 10.345 10.475 15.000 11.765 ;
        RECT 17.865 10.475 24.530 11.765 ;
        RECT 26.400 10.475 38.130 11.765 ;
        RECT 40.000 10.475 51.730 11.765 ;
        RECT 53.590 10.475 55.790 11.765 ;
        RECT 58.450 10.475 67.775 11.765 ;
        RECT 69.685 11.765 70.975 19.800 ;
        RECT 98.625 17.995 99.915 24.660 ;
        RECT 98.625 11.765 99.915 15.130 ;
        RECT 69.685 10.475 74.340 11.765 ;
        RECT 77.205 10.475 83.870 11.765 ;
        RECT 85.730 10.475 87.930 11.765 ;
        RECT 90.590 10.475 99.915 11.765 ;
        RECT 140.465 121.015 145.120 122.305 ;
        RECT 147.985 121.015 154.650 122.305 ;
        RECT 156.510 121.015 158.710 122.305 ;
        RECT 161.370 121.015 170.695 122.305 ;
        RECT 238.525 122.665 239.695 123.835 ;
        RECT 140.465 112.980 141.755 121.015 ;
        RECT 169.405 117.650 170.695 121.015 ;
        RECT 172.605 121.015 177.260 122.305 ;
        RECT 180.125 121.015 186.790 122.305 ;
        RECT 188.660 121.015 200.390 122.305 ;
        RECT 202.260 121.015 213.990 122.305 ;
        RECT 215.850 121.015 218.050 122.305 ;
        RECT 220.710 121.015 230.035 122.305 ;
        RECT 140.465 108.120 141.755 110.320 ;
        RECT 140.465 94.530 141.755 106.260 ;
        RECT 169.405 108.120 170.695 114.785 ;
        RECT 172.605 112.980 173.895 121.015 ;
        RECT 228.745 117.650 230.035 121.015 ;
        RECT 235.325 121.065 236.915 122.235 ;
        RECT 232.545 119.465 233.715 120.635 ;
        RECT 238.525 119.465 239.695 120.635 ;
        RECT 235.325 117.865 236.915 119.035 ;
        RECT 232.545 116.265 233.715 117.435 ;
        RECT 238.525 116.265 239.695 117.435 ;
        RECT 172.605 108.120 173.895 110.320 ;
        RECT 140.465 80.930 141.755 92.660 ;
        RECT 169.405 94.520 170.695 106.250 ;
        RECT 140.465 67.330 141.755 79.060 ;
        RECT 169.405 80.920 170.695 92.650 ;
        RECT 172.605 94.530 173.895 106.260 ;
        RECT 228.745 108.120 230.035 114.785 ;
        RECT 235.325 114.665 236.915 115.835 ;
        RECT 232.545 113.065 233.715 114.235 ;
        RECT 238.525 113.065 239.695 114.235 ;
        RECT 235.325 111.465 236.915 112.635 ;
        RECT 232.545 109.865 233.715 111.035 ;
        RECT 238.525 109.865 239.695 111.035 ;
        RECT 235.325 108.265 236.915 109.435 ;
        RECT 232.545 106.665 233.715 107.835 ;
        RECT 238.525 106.665 239.695 107.835 ;
        RECT 140.465 53.730 141.755 65.460 ;
        RECT 169.405 67.320 170.695 79.050 ;
        RECT 172.605 80.930 173.895 92.660 ;
        RECT 228.745 94.520 230.035 106.250 ;
        RECT 235.325 105.065 236.915 106.235 ;
        RECT 232.545 103.465 233.715 104.635 ;
        RECT 238.525 103.465 239.695 104.635 ;
        RECT 235.325 101.865 236.915 103.035 ;
        RECT 232.545 100.265 233.715 101.435 ;
        RECT 238.525 100.265 239.695 101.435 ;
        RECT 235.325 98.665 236.915 99.835 ;
        RECT 232.545 97.065 233.715 98.235 ;
        RECT 238.525 97.065 239.695 98.235 ;
        RECT 235.325 95.465 236.915 96.635 ;
        RECT 232.545 93.865 233.715 95.035 ;
        RECT 238.525 93.865 239.695 95.035 ;
        RECT 140.465 40.130 141.755 51.860 ;
        RECT 169.405 53.720 170.695 65.450 ;
        RECT 172.605 67.330 173.895 79.060 ;
        RECT 228.745 80.920 230.035 92.650 ;
        RECT 235.325 92.265 236.915 93.435 ;
        RECT 232.545 90.665 233.715 91.835 ;
        RECT 238.525 90.665 239.695 91.835 ;
        RECT 235.325 89.065 236.915 90.235 ;
        RECT 232.545 87.465 233.715 88.635 ;
        RECT 238.525 87.465 239.695 88.635 ;
        RECT 235.325 85.865 236.915 87.035 ;
        RECT 232.545 84.265 233.715 85.435 ;
        RECT 238.525 84.265 239.695 85.435 ;
        RECT 235.325 82.665 236.915 83.835 ;
        RECT 232.545 81.065 233.715 82.235 ;
        RECT 238.525 81.065 239.695 82.235 ;
        RECT 235.325 79.465 236.915 80.635 ;
        RECT 172.605 53.730 173.895 65.460 ;
        RECT 228.745 67.320 230.035 79.050 ;
        RECT 232.545 77.865 233.715 79.035 ;
        RECT 238.525 77.865 239.695 79.035 ;
        RECT 235.325 76.265 236.915 77.435 ;
        RECT 232.545 74.665 233.715 75.835 ;
        RECT 238.525 74.665 239.695 75.835 ;
        RECT 235.325 73.065 236.915 74.235 ;
        RECT 232.545 71.465 233.715 72.635 ;
        RECT 238.525 71.465 239.695 72.635 ;
        RECT 235.325 69.865 236.915 71.035 ;
        RECT 232.545 68.265 233.715 69.435 ;
        RECT 238.525 68.265 239.695 69.435 ;
        RECT 235.325 66.665 236.915 67.835 ;
        RECT 140.465 26.530 141.755 38.260 ;
        RECT 169.405 40.120 170.695 51.850 ;
        RECT 172.605 40.130 173.895 51.860 ;
        RECT 228.745 53.720 230.035 65.450 ;
        RECT 232.545 65.065 233.715 66.235 ;
        RECT 238.525 65.065 239.695 66.235 ;
        RECT 235.325 63.465 236.915 64.635 ;
        RECT 232.545 61.865 233.715 63.035 ;
        RECT 238.525 61.865 239.695 63.035 ;
        RECT 235.325 60.265 236.915 61.435 ;
        RECT 232.545 58.665 233.715 59.835 ;
        RECT 238.525 58.665 239.695 59.835 ;
        RECT 235.325 57.065 236.915 58.235 ;
        RECT 232.545 55.465 233.715 56.635 ;
        RECT 238.525 55.465 239.695 56.635 ;
        RECT 235.325 53.865 236.915 55.035 ;
        RECT 232.545 52.265 233.715 53.435 ;
        RECT 238.525 52.265 239.695 53.435 ;
        RECT 140.465 17.995 141.755 24.660 ;
        RECT 169.405 26.520 170.695 38.250 ;
        RECT 169.405 22.460 170.695 24.660 ;
        RECT 172.605 26.530 173.895 38.260 ;
        RECT 228.745 40.120 230.035 51.850 ;
        RECT 235.325 50.665 236.915 51.835 ;
        RECT 232.545 49.065 233.715 50.235 ;
        RECT 238.525 49.065 239.695 50.235 ;
        RECT 235.325 47.465 236.915 48.635 ;
        RECT 232.545 45.865 233.715 47.035 ;
        RECT 238.525 45.865 239.695 47.035 ;
        RECT 235.325 44.265 236.915 45.435 ;
        RECT 232.545 42.665 233.715 43.835 ;
        RECT 238.525 42.665 239.695 43.835 ;
        RECT 235.325 41.065 236.915 42.235 ;
        RECT 232.545 39.465 233.715 40.635 ;
        RECT 238.525 39.465 239.695 40.635 ;
        RECT 140.465 11.765 141.755 15.130 ;
        RECT 169.405 11.765 170.695 19.800 ;
        RECT 172.605 17.995 173.895 24.660 ;
        RECT 228.745 26.520 230.035 38.250 ;
        RECT 235.325 37.865 236.915 39.035 ;
        RECT 232.545 36.265 233.715 37.435 ;
        RECT 238.525 36.265 239.695 37.435 ;
        RECT 235.325 34.665 236.915 35.835 ;
        RECT 232.545 33.065 233.715 34.235 ;
        RECT 238.525 33.065 239.695 34.235 ;
        RECT 235.325 31.465 236.915 32.635 ;
        RECT 232.545 29.865 233.715 31.035 ;
        RECT 238.525 29.865 239.695 31.035 ;
        RECT 235.325 28.265 236.915 29.435 ;
        RECT 232.545 26.665 233.715 27.835 ;
        RECT 238.525 26.665 239.695 27.835 ;
        RECT 235.325 25.065 236.915 26.235 ;
        RECT 228.745 22.460 230.035 24.660 ;
        RECT 232.545 23.465 233.715 24.635 ;
        RECT 238.525 23.465 239.695 24.635 ;
        RECT 235.325 21.865 236.915 23.035 ;
        RECT 232.545 20.265 233.715 21.435 ;
        RECT 238.525 20.265 239.695 21.435 ;
        RECT 140.465 10.475 149.790 11.765 ;
        RECT 152.450 10.475 154.650 11.765 ;
        RECT 156.510 10.475 163.175 11.765 ;
        RECT 166.040 10.475 170.695 11.765 ;
        RECT 172.605 11.765 173.895 15.130 ;
        RECT 228.745 11.765 230.035 19.800 ;
        RECT 235.325 18.665 236.915 19.835 ;
        RECT 232.545 17.065 233.715 18.235 ;
        RECT 238.525 17.065 239.695 18.235 ;
        RECT 235.325 15.465 236.915 16.635 ;
        RECT 232.545 13.865 233.715 15.035 ;
        RECT 172.605 10.475 181.930 11.765 ;
        RECT 184.590 10.475 186.790 11.765 ;
        RECT 188.650 10.475 200.380 11.765 ;
        RECT 202.250 10.475 213.980 11.765 ;
        RECT 215.850 10.475 222.515 11.765 ;
        RECT 225.380 10.475 230.035 11.765 ;
        RECT 238.525 13.865 239.695 15.035 ;
        RECT 9.785 6.105 10.955 7.275 ;
        RECT 12.985 6.105 14.155 7.275 ;
        RECT 16.185 6.105 17.355 7.275 ;
        RECT 19.385 6.105 20.555 7.275 ;
        RECT 22.585 6.105 23.755 7.275 ;
        RECT 25.785 6.105 26.955 7.275 ;
        RECT 28.985 6.105 30.155 7.275 ;
        RECT 32.185 6.105 33.355 7.275 ;
        RECT 35.385 6.105 36.555 7.275 ;
        RECT 38.585 6.105 39.755 7.275 ;
        RECT 41.785 6.105 42.955 7.275 ;
        RECT 44.985 6.105 46.155 7.275 ;
        RECT 48.185 6.105 49.355 7.275 ;
        RECT 51.385 6.105 52.555 7.275 ;
        RECT 54.585 6.105 55.755 7.275 ;
        RECT 57.785 6.105 58.955 7.275 ;
        RECT 60.985 6.105 62.155 7.275 ;
        RECT 64.185 6.105 65.355 7.275 ;
        RECT 67.385 6.105 68.555 7.275 ;
        RECT 70.585 6.105 71.755 7.275 ;
        RECT 73.785 6.105 74.955 7.275 ;
        RECT 76.985 6.105 78.155 7.275 ;
        RECT 80.185 6.105 81.355 7.275 ;
        RECT 83.385 6.105 84.555 7.275 ;
        RECT 86.585 6.105 87.755 7.275 ;
        RECT 89.785 6.105 90.955 7.275 ;
        RECT 92.985 6.105 94.155 7.275 ;
        RECT 96.185 6.105 97.355 7.275 ;
        RECT 99.385 6.105 100.555 7.275 ;
        RECT 102.585 6.105 103.755 7.275 ;
        RECT 105.785 6.105 106.955 7.275 ;
        RECT 108.985 6.105 110.155 7.275 ;
        RECT 112.185 6.105 113.355 7.275 ;
        RECT 115.385 6.105 116.555 7.275 ;
        RECT 123.825 6.105 124.995 7.275 ;
        RECT 127.025 6.105 128.195 7.275 ;
        RECT 130.225 6.105 131.395 7.275 ;
        RECT 133.425 6.105 134.595 7.275 ;
        RECT 136.625 6.105 137.795 7.275 ;
        RECT 139.825 6.105 140.995 7.275 ;
        RECT 143.025 6.105 144.195 7.275 ;
        RECT 146.225 6.105 147.395 7.275 ;
        RECT 149.425 6.105 150.595 7.275 ;
        RECT 152.625 6.105 153.795 7.275 ;
        RECT 155.825 6.105 156.995 7.275 ;
        RECT 159.025 6.105 160.195 7.275 ;
        RECT 162.225 6.105 163.395 7.275 ;
        RECT 165.425 6.105 166.595 7.275 ;
        RECT 168.625 6.105 169.795 7.275 ;
        RECT 171.825 6.105 172.995 7.275 ;
        RECT 175.025 6.105 176.195 7.275 ;
        RECT 178.225 6.105 179.395 7.275 ;
        RECT 181.425 6.105 182.595 7.275 ;
        RECT 184.625 6.105 185.795 7.275 ;
        RECT 187.825 6.105 188.995 7.275 ;
        RECT 191.025 6.105 192.195 7.275 ;
        RECT 194.225 6.105 195.395 7.275 ;
        RECT 197.425 6.105 198.595 7.275 ;
        RECT 200.625 6.105 201.795 7.275 ;
        RECT 203.825 6.105 204.995 7.275 ;
        RECT 207.025 6.105 208.195 7.275 ;
        RECT 210.225 6.105 211.395 7.275 ;
        RECT 213.425 6.105 214.595 7.275 ;
        RECT 216.625 6.105 217.795 7.275 ;
        RECT 219.825 6.105 220.995 7.275 ;
        RECT 223.025 6.105 224.195 7.275 ;
        RECT 226.225 6.105 227.395 7.275 ;
        RECT 229.425 6.105 230.595 7.275 ;
        RECT 8.185 2.905 9.355 4.495 ;
        RECT 11.385 2.905 12.555 4.495 ;
        RECT 14.585 2.905 15.755 4.495 ;
        RECT 17.785 2.905 18.955 4.495 ;
        RECT 20.985 2.905 22.155 4.495 ;
        RECT 24.185 2.905 25.355 4.495 ;
        RECT 27.385 2.905 28.555 4.495 ;
        RECT 30.585 2.905 31.755 4.495 ;
        RECT 33.785 2.905 34.955 4.495 ;
        RECT 36.985 2.905 38.155 4.495 ;
        RECT 40.185 2.905 41.355 4.495 ;
        RECT 43.385 2.905 44.555 4.495 ;
        RECT 46.585 2.905 47.755 4.495 ;
        RECT 49.785 2.905 50.955 4.495 ;
        RECT 52.985 2.905 54.155 4.495 ;
        RECT 56.185 2.905 57.355 4.495 ;
        RECT 59.385 2.905 60.555 4.495 ;
        RECT 62.585 2.905 63.755 4.495 ;
        RECT 65.785 2.905 66.955 4.495 ;
        RECT 68.985 2.905 70.155 4.495 ;
        RECT 72.185 2.905 73.355 4.495 ;
        RECT 75.385 2.905 76.555 4.495 ;
        RECT 78.585 2.905 79.755 4.495 ;
        RECT 81.785 2.905 82.955 4.495 ;
        RECT 84.985 2.905 86.155 4.495 ;
        RECT 88.185 2.905 89.355 4.495 ;
        RECT 91.385 2.905 92.555 4.495 ;
        RECT 94.585 2.905 95.755 4.495 ;
        RECT 97.785 2.905 98.955 4.495 ;
        RECT 100.985 2.905 102.155 4.495 ;
        RECT 104.185 2.905 105.355 4.495 ;
        RECT 107.385 2.905 108.555 4.495 ;
        RECT 110.585 2.905 111.755 4.495 ;
        RECT 113.785 2.905 114.955 4.495 ;
        RECT 116.985 2.905 118.155 4.495 ;
        RECT 122.225 2.905 123.395 4.495 ;
        RECT 125.425 2.905 126.595 4.495 ;
        RECT 128.625 2.905 129.795 4.495 ;
        RECT 131.825 2.905 132.995 4.495 ;
        RECT 135.025 2.905 136.195 4.495 ;
        RECT 138.225 2.905 139.395 4.495 ;
        RECT 141.425 2.905 142.595 4.495 ;
        RECT 144.625 2.905 145.795 4.495 ;
        RECT 147.825 2.905 148.995 4.495 ;
        RECT 151.025 2.905 152.195 4.495 ;
        RECT 154.225 2.905 155.395 4.495 ;
        RECT 157.425 2.905 158.595 4.495 ;
        RECT 160.625 2.905 161.795 4.495 ;
        RECT 163.825 2.905 164.995 4.495 ;
        RECT 167.025 2.905 168.195 4.495 ;
        RECT 170.225 2.905 171.395 4.495 ;
        RECT 173.425 2.905 174.595 4.495 ;
        RECT 176.625 2.905 177.795 4.495 ;
        RECT 179.825 2.905 180.995 4.495 ;
        RECT 183.025 2.905 184.195 4.495 ;
        RECT 186.225 2.905 187.395 4.495 ;
        RECT 189.425 2.905 190.595 4.495 ;
        RECT 192.625 2.905 193.795 4.495 ;
        RECT 195.825 2.905 196.995 4.495 ;
        RECT 199.025 2.905 200.195 4.495 ;
        RECT 202.225 2.905 203.395 4.495 ;
        RECT 205.425 2.905 206.595 4.495 ;
        RECT 208.625 2.905 209.795 4.495 ;
        RECT 211.825 2.905 212.995 4.495 ;
        RECT 215.025 2.905 216.195 4.495 ;
        RECT 218.225 2.905 219.395 4.495 ;
        RECT 221.425 2.905 222.595 4.495 ;
        RECT 224.625 2.905 225.795 4.495 ;
        RECT 227.825 2.905 228.995 4.495 ;
        RECT 231.025 2.905 232.195 4.495 ;
        RECT 9.785 0.125 10.955 1.295 ;
        RECT 12.985 0.125 14.155 1.295 ;
        RECT 16.185 0.125 17.355 1.295 ;
        RECT 19.385 0.125 20.555 1.295 ;
        RECT 22.585 0.125 23.755 1.295 ;
        RECT 25.785 0.125 26.955 1.295 ;
        RECT 28.985 0.125 30.155 1.295 ;
        RECT 32.185 0.125 33.355 1.295 ;
        RECT 35.385 0.125 36.555 1.295 ;
        RECT 38.585 0.125 39.755 1.295 ;
        RECT 41.785 0.125 42.955 1.295 ;
        RECT 44.985 0.125 46.155 1.295 ;
        RECT 48.185 0.125 49.355 1.295 ;
        RECT 51.385 0.125 52.555 1.295 ;
        RECT 54.585 0.125 55.755 1.295 ;
        RECT 57.785 0.125 58.955 1.295 ;
        RECT 60.985 0.125 62.155 1.295 ;
        RECT 64.185 0.125 65.355 1.295 ;
        RECT 67.385 0.125 68.555 1.295 ;
        RECT 70.585 0.125 71.755 1.295 ;
        RECT 73.785 0.125 74.955 1.295 ;
        RECT 76.985 0.125 78.155 1.295 ;
        RECT 80.185 0.125 81.355 1.295 ;
        RECT 83.385 0.125 84.555 1.295 ;
        RECT 86.585 0.125 87.755 1.295 ;
        RECT 89.785 0.125 90.955 1.295 ;
        RECT 92.985 0.125 94.155 1.295 ;
        RECT 96.185 0.125 97.355 1.295 ;
        RECT 99.385 0.125 100.555 1.295 ;
        RECT 102.585 0.125 103.755 1.295 ;
        RECT 105.785 0.125 106.955 1.295 ;
        RECT 108.985 0.125 110.155 1.295 ;
        RECT 112.185 0.125 113.355 1.295 ;
        RECT 115.385 0.125 116.555 1.295 ;
        RECT 123.825 0.125 124.995 1.295 ;
        RECT 127.025 0.125 128.195 1.295 ;
        RECT 130.225 0.125 131.395 1.295 ;
        RECT 133.425 0.125 134.595 1.295 ;
        RECT 136.625 0.125 137.795 1.295 ;
        RECT 139.825 0.125 140.995 1.295 ;
        RECT 143.025 0.125 144.195 1.295 ;
        RECT 146.225 0.125 147.395 1.295 ;
        RECT 149.425 0.125 150.595 1.295 ;
        RECT 152.625 0.125 153.795 1.295 ;
        RECT 155.825 0.125 156.995 1.295 ;
        RECT 159.025 0.125 160.195 1.295 ;
        RECT 162.225 0.125 163.395 1.295 ;
        RECT 165.425 0.125 166.595 1.295 ;
        RECT 168.625 0.125 169.795 1.295 ;
        RECT 171.825 0.125 172.995 1.295 ;
        RECT 175.025 0.125 176.195 1.295 ;
        RECT 178.225 0.125 179.395 1.295 ;
        RECT 181.425 0.125 182.595 1.295 ;
        RECT 184.625 0.125 185.795 1.295 ;
        RECT 187.825 0.125 188.995 1.295 ;
        RECT 191.025 0.125 192.195 1.295 ;
        RECT 194.225 0.125 195.395 1.295 ;
        RECT 197.425 0.125 198.595 1.295 ;
        RECT 200.625 0.125 201.795 1.295 ;
        RECT 203.825 0.125 204.995 1.295 ;
        RECT 207.025 0.125 208.195 1.295 ;
        RECT 210.225 0.125 211.395 1.295 ;
        RECT 213.425 0.125 214.595 1.295 ;
        RECT 216.625 0.125 217.795 1.295 ;
        RECT 219.825 0.125 220.995 1.295 ;
        RECT 223.025 0.125 224.195 1.295 ;
        RECT 226.225 0.125 227.395 1.295 ;
        RECT 229.425 0.125 230.595 1.295 ;
      LAYER met4 ;
        RECT 95.390 166.780 95.860 169.545 ;
        RECT 95.390 166.300 98.250 166.780 ;
        RECT 95.390 163.550 95.860 166.300 ;
        RECT 105.460 159.205 105.890 176.005 ;
        RECT 110.060 173.225 110.490 176.005 ;
        RECT 110.010 172.895 110.490 173.225 ;
        RECT 110.060 159.205 110.490 172.895 ;
        RECT 114.665 147.660 115.095 176.005 ;
        RECT 0.680 125.860 1.860 127.040 ;
        RECT 6.660 125.860 7.840 127.040 ;
        RECT 232.540 125.860 233.720 127.040 ;
        RECT 238.520 125.860 239.700 127.040 ;
        RECT 3.460 124.260 5.060 125.440 ;
        RECT 235.320 124.260 236.920 125.440 ;
        RECT 0.680 122.660 1.860 123.840 ;
        RECT 6.660 122.660 7.840 123.840 ;
        RECT 232.540 122.660 233.720 123.840 ;
        RECT 238.520 122.660 239.700 123.840 ;
        RECT 3.460 121.060 5.060 122.240 ;
        RECT 10.310 120.980 19.675 122.340 ;
        RECT 22.325 120.980 24.535 122.340 ;
        RECT 26.385 120.980 38.125 122.340 ;
        RECT 39.985 120.980 51.725 122.340 ;
        RECT 52.660 120.980 60.260 122.340 ;
        RECT 63.115 121.790 67.810 122.340 ;
        RECT 69.650 121.790 79.015 122.340 ;
        RECT 63.115 120.980 79.015 121.790 ;
        RECT 81.665 120.980 83.875 122.340 ;
        RECT 84.800 120.980 92.400 122.340 ;
        RECT 95.255 120.980 99.950 122.340 ;
        RECT 0.680 119.460 1.860 120.640 ;
        RECT 6.660 119.460 7.840 120.640 ;
        RECT 3.460 117.860 5.060 119.040 ;
        RECT 10.310 117.645 11.670 120.980 ;
        RECT 66.450 120.190 71.010 120.980 ;
        RECT 0.680 116.260 1.860 117.440 ;
        RECT 6.660 116.260 7.840 117.440 ;
        RECT 3.460 114.660 5.060 115.840 ;
        RECT 0.680 113.060 1.860 114.240 ;
        RECT 6.660 113.060 7.840 114.240 ;
        RECT 3.460 111.460 5.060 112.640 ;
        RECT 0.680 109.860 1.860 111.040 ;
        RECT 6.660 109.860 7.840 111.040 ;
        RECT 3.460 108.260 5.060 109.440 ;
        RECT 0.680 106.660 1.860 107.840 ;
        RECT 6.660 106.660 7.840 107.840 ;
        RECT 10.310 107.190 11.670 114.790 ;
        RECT 66.450 114.635 67.810 120.190 ;
        RECT 69.650 117.645 71.010 120.190 ;
        RECT 69.650 114.635 71.010 114.790 ;
        RECT 66.450 113.035 71.010 114.635 ;
        RECT 66.450 112.975 67.810 113.035 ;
        RECT 66.450 109.025 67.810 110.325 ;
        RECT 69.650 109.025 71.010 113.035 ;
        RECT 98.590 112.975 99.950 120.980 ;
        RECT 140.430 120.980 145.125 122.340 ;
        RECT 147.980 120.980 155.580 122.340 ;
        RECT 156.505 120.980 158.715 122.340 ;
        RECT 161.365 121.790 170.730 122.340 ;
        RECT 172.570 121.790 177.265 122.340 ;
        RECT 161.365 120.980 177.265 121.790 ;
        RECT 180.120 120.980 187.720 122.340 ;
        RECT 188.655 120.980 200.395 122.340 ;
        RECT 202.255 120.980 213.995 122.340 ;
        RECT 215.845 120.980 218.055 122.340 ;
        RECT 220.705 120.980 230.070 122.340 ;
        RECT 235.320 121.060 236.920 122.240 ;
        RECT 140.430 112.975 141.790 120.980 ;
        RECT 169.370 120.190 173.930 120.980 ;
        RECT 169.370 117.645 170.730 120.190 ;
        RECT 169.370 114.635 170.730 114.790 ;
        RECT 172.570 114.635 173.930 120.190 ;
        RECT 228.710 117.645 230.070 120.980 ;
        RECT 232.540 119.460 233.720 120.640 ;
        RECT 238.520 119.460 239.700 120.640 ;
        RECT 235.320 117.860 236.920 119.040 ;
        RECT 232.540 116.260 233.720 117.440 ;
        RECT 238.520 116.260 239.700 117.440 ;
        RECT 169.370 113.035 173.930 114.635 ;
        RECT 66.450 108.115 71.010 109.025 ;
        RECT 98.590 108.115 99.950 110.325 ;
        RECT 140.430 108.115 141.790 110.325 ;
        RECT 169.370 109.025 170.730 113.035 ;
        RECT 172.570 112.975 173.930 113.035 ;
        RECT 172.570 109.025 173.930 110.325 ;
        RECT 169.370 108.115 173.930 109.025 ;
        RECT 67.600 107.425 71.010 108.115 ;
        RECT 69.650 107.190 71.010 107.425 ;
        RECT 169.370 107.425 172.780 108.115 ;
        RECT 169.370 107.190 170.730 107.425 ;
        RECT 228.710 107.190 230.070 114.790 ;
        RECT 235.320 114.660 236.920 115.840 ;
        RECT 232.540 113.060 233.720 114.240 ;
        RECT 238.520 113.060 239.700 114.240 ;
        RECT 235.320 111.460 236.920 112.640 ;
        RECT 232.540 109.860 233.720 111.040 ;
        RECT 238.520 109.860 239.700 111.040 ;
        RECT 235.320 108.260 236.920 109.440 ;
        RECT 232.540 106.660 233.720 107.840 ;
        RECT 238.520 106.660 239.700 107.840 ;
        RECT 3.460 105.060 5.060 106.240 ;
        RECT 0.680 103.460 1.860 104.640 ;
        RECT 6.660 103.460 7.840 104.640 ;
        RECT 3.460 101.860 5.060 103.040 ;
        RECT 0.680 100.260 1.860 101.440 ;
        RECT 6.660 100.260 7.840 101.440 ;
        RECT 3.460 98.660 5.060 99.840 ;
        RECT 0.680 97.060 1.860 98.240 ;
        RECT 6.660 97.060 7.840 98.240 ;
        RECT 3.460 95.460 5.060 96.640 ;
        RECT 0.680 93.860 1.860 95.040 ;
        RECT 6.660 93.860 7.840 95.040 ;
        RECT 10.310 94.515 11.670 106.255 ;
        RECT 66.450 104.550 67.810 106.265 ;
        RECT 69.650 104.550 71.010 106.255 ;
        RECT 66.450 102.950 71.010 104.550 ;
        RECT 66.450 100.135 67.810 102.950 ;
        RECT 69.650 100.135 71.010 102.950 ;
        RECT 66.450 98.535 71.010 100.135 ;
        RECT 66.450 94.525 67.810 98.535 ;
        RECT 69.650 94.515 71.010 98.535 ;
        RECT 98.590 94.525 99.950 106.265 ;
        RECT 140.430 94.525 141.790 106.265 ;
        RECT 169.370 104.550 170.730 106.255 ;
        RECT 172.570 104.550 173.930 106.265 ;
        RECT 169.370 102.950 173.930 104.550 ;
        RECT 169.370 100.135 170.730 102.950 ;
        RECT 172.570 100.135 173.930 102.950 ;
        RECT 169.370 98.535 173.930 100.135 ;
        RECT 169.370 94.515 170.730 98.535 ;
        RECT 172.570 94.525 173.930 98.535 ;
        RECT 228.710 94.515 230.070 106.255 ;
        RECT 235.320 105.060 236.920 106.240 ;
        RECT 232.540 103.460 233.720 104.640 ;
        RECT 238.520 103.460 239.700 104.640 ;
        RECT 235.320 101.860 236.920 103.040 ;
        RECT 232.540 100.260 233.720 101.440 ;
        RECT 238.520 100.260 239.700 101.440 ;
        RECT 235.320 98.660 236.920 99.840 ;
        RECT 232.540 97.060 233.720 98.240 ;
        RECT 238.520 97.060 239.700 98.240 ;
        RECT 235.320 95.460 236.920 96.640 ;
        RECT 232.540 93.860 233.720 95.040 ;
        RECT 238.520 93.860 239.700 95.040 ;
        RECT 3.460 92.260 5.060 93.440 ;
        RECT 0.680 90.660 1.860 91.840 ;
        RECT 6.660 90.660 7.840 91.840 ;
        RECT 3.460 89.060 5.060 90.240 ;
        RECT 0.680 87.460 1.860 88.640 ;
        RECT 6.660 87.460 7.840 88.640 ;
        RECT 3.460 85.860 5.060 87.040 ;
        RECT 0.680 84.260 1.860 85.440 ;
        RECT 6.660 84.260 7.840 85.440 ;
        RECT 3.460 82.660 5.060 83.840 ;
        RECT 0.680 81.060 1.860 82.240 ;
        RECT 6.660 81.060 7.840 82.240 ;
        RECT 10.310 80.915 11.670 92.655 ;
        RECT 66.450 91.615 67.810 92.665 ;
        RECT 69.650 91.615 71.010 92.655 ;
        RECT 66.450 90.015 71.010 91.615 ;
        RECT 66.450 87.205 67.810 90.015 ;
        RECT 69.650 87.205 71.010 90.015 ;
        RECT 66.450 85.605 71.010 87.205 ;
        RECT 66.450 82.720 67.810 85.605 ;
        RECT 69.650 82.720 71.010 85.605 ;
        RECT 66.450 81.120 71.010 82.720 ;
        RECT 66.450 80.925 67.810 81.120 ;
        RECT 69.650 80.915 71.010 81.120 ;
        RECT 98.590 80.925 99.950 92.665 ;
        RECT 140.430 80.925 141.790 92.665 ;
        RECT 169.370 91.615 170.730 92.655 ;
        RECT 172.570 91.615 173.930 92.665 ;
        RECT 169.370 90.015 173.930 91.615 ;
        RECT 169.370 87.205 170.730 90.015 ;
        RECT 172.570 87.205 173.930 90.015 ;
        RECT 169.370 85.605 173.930 87.205 ;
        RECT 169.370 82.720 170.730 85.605 ;
        RECT 172.570 82.720 173.930 85.605 ;
        RECT 169.370 81.120 173.930 82.720 ;
        RECT 169.370 80.915 170.730 81.120 ;
        RECT 172.570 80.925 173.930 81.120 ;
        RECT 228.710 80.915 230.070 92.655 ;
        RECT 235.320 92.260 236.920 93.440 ;
        RECT 232.540 90.660 233.720 91.840 ;
        RECT 238.520 90.660 239.700 91.840 ;
        RECT 235.320 89.060 236.920 90.240 ;
        RECT 232.540 87.460 233.720 88.640 ;
        RECT 238.520 87.460 239.700 88.640 ;
        RECT 235.320 85.860 236.920 87.040 ;
        RECT 232.540 84.260 233.720 85.440 ;
        RECT 238.520 84.260 239.700 85.440 ;
        RECT 235.320 82.660 236.920 83.840 ;
        RECT 232.540 81.060 233.720 82.240 ;
        RECT 238.520 81.060 239.700 82.240 ;
        RECT 3.460 79.460 5.060 80.640 ;
        RECT 235.320 79.460 236.920 80.640 ;
        RECT 0.680 77.860 1.860 79.040 ;
        RECT 6.660 77.860 7.840 79.040 ;
        RECT 3.460 76.260 5.060 77.440 ;
        RECT 0.680 74.660 1.860 75.840 ;
        RECT 6.660 74.660 7.840 75.840 ;
        RECT 3.460 73.060 5.060 74.240 ;
        RECT 0.680 71.460 1.860 72.640 ;
        RECT 6.660 71.460 7.840 72.640 ;
        RECT 3.460 69.860 5.060 71.040 ;
        RECT 0.680 68.260 1.860 69.440 ;
        RECT 6.660 68.260 7.840 69.440 ;
        RECT 3.460 66.660 5.060 67.840 ;
        RECT 10.310 67.315 11.670 79.055 ;
        RECT 66.450 74.255 67.810 79.065 ;
        RECT 69.650 74.255 71.010 79.055 ;
        RECT 66.450 72.655 71.010 74.255 ;
        RECT 66.450 69.765 67.810 72.655 ;
        RECT 69.650 69.765 71.010 72.655 ;
        RECT 66.450 68.165 71.010 69.765 ;
        RECT 66.450 67.325 67.810 68.165 ;
        RECT 69.650 67.315 71.010 68.165 ;
        RECT 98.590 67.325 99.950 79.065 ;
        RECT 140.430 67.325 141.790 79.065 ;
        RECT 169.370 74.255 170.730 79.055 ;
        RECT 172.570 74.255 173.930 79.065 ;
        RECT 169.370 72.655 173.930 74.255 ;
        RECT 169.370 69.765 170.730 72.655 ;
        RECT 172.570 69.765 173.930 72.655 ;
        RECT 169.370 68.165 173.930 69.765 ;
        RECT 169.370 67.315 170.730 68.165 ;
        RECT 172.570 67.325 173.930 68.165 ;
        RECT 228.710 67.315 230.070 79.055 ;
        RECT 232.540 77.860 233.720 79.040 ;
        RECT 238.520 77.860 239.700 79.040 ;
        RECT 235.320 76.260 236.920 77.440 ;
        RECT 232.540 74.660 233.720 75.840 ;
        RECT 238.520 74.660 239.700 75.840 ;
        RECT 235.320 73.060 236.920 74.240 ;
        RECT 232.540 71.460 233.720 72.640 ;
        RECT 238.520 71.460 239.700 72.640 ;
        RECT 235.320 69.860 236.920 71.040 ;
        RECT 232.540 68.260 233.720 69.440 ;
        RECT 238.520 68.260 239.700 69.440 ;
        RECT 235.320 66.660 236.920 67.840 ;
        RECT 0.680 65.060 1.860 66.240 ;
        RECT 6.660 65.060 7.840 66.240 ;
        RECT 3.460 63.460 5.060 64.640 ;
        RECT 0.680 61.860 1.860 63.040 ;
        RECT 6.660 61.860 7.840 63.040 ;
        RECT 3.460 60.260 5.060 61.440 ;
        RECT 0.680 58.660 1.860 59.840 ;
        RECT 6.660 58.660 7.840 59.840 ;
        RECT 3.460 57.060 5.060 58.240 ;
        RECT 0.680 55.460 1.860 56.640 ;
        RECT 6.660 55.460 7.840 56.640 ;
        RECT 3.460 53.860 5.060 55.040 ;
        RECT 10.310 53.715 11.670 65.455 ;
        RECT 66.450 65.300 67.810 65.465 ;
        RECT 69.650 65.300 71.010 65.455 ;
        RECT 66.450 63.700 71.010 65.300 ;
        RECT 66.450 56.820 67.810 63.700 ;
        RECT 69.650 56.820 71.010 63.700 ;
        RECT 66.450 55.220 71.010 56.820 ;
        RECT 66.450 53.725 67.810 55.220 ;
        RECT 69.650 53.715 71.010 55.220 ;
        RECT 98.590 53.725 99.950 65.465 ;
        RECT 140.430 53.725 141.790 65.465 ;
        RECT 169.370 65.300 170.730 65.455 ;
        RECT 172.570 65.300 173.930 65.465 ;
        RECT 169.370 63.700 173.930 65.300 ;
        RECT 169.370 56.820 170.730 63.700 ;
        RECT 172.570 56.820 173.930 63.700 ;
        RECT 169.370 55.220 173.930 56.820 ;
        RECT 169.370 53.715 170.730 55.220 ;
        RECT 172.570 53.725 173.930 55.220 ;
        RECT 228.710 53.715 230.070 65.455 ;
        RECT 232.540 65.060 233.720 66.240 ;
        RECT 238.520 65.060 239.700 66.240 ;
        RECT 235.320 63.460 236.920 64.640 ;
        RECT 232.540 61.860 233.720 63.040 ;
        RECT 238.520 61.860 239.700 63.040 ;
        RECT 235.320 60.260 236.920 61.440 ;
        RECT 232.540 58.660 233.720 59.840 ;
        RECT 238.520 58.660 239.700 59.840 ;
        RECT 235.320 57.060 236.920 58.240 ;
        RECT 232.540 55.460 233.720 56.640 ;
        RECT 238.520 55.460 239.700 56.640 ;
        RECT 235.320 53.860 236.920 55.040 ;
        RECT 0.680 52.260 1.860 53.440 ;
        RECT 6.660 52.260 7.840 53.440 ;
        RECT 67.720 51.865 69.765 52.355 ;
        RECT 170.615 51.865 172.660 52.355 ;
        RECT 232.540 52.260 233.720 53.440 ;
        RECT 238.520 52.260 239.700 53.440 ;
        RECT 66.450 51.855 69.765 51.865 ;
        RECT 3.460 50.660 5.060 51.840 ;
        RECT 0.680 49.060 1.860 50.240 ;
        RECT 6.660 49.060 7.840 50.240 ;
        RECT 3.460 47.460 5.060 48.640 ;
        RECT 0.680 45.860 1.860 47.040 ;
        RECT 6.660 45.860 7.840 47.040 ;
        RECT 3.460 44.260 5.060 45.440 ;
        RECT 0.680 42.660 1.860 43.840 ;
        RECT 6.660 42.660 7.840 43.840 ;
        RECT 3.460 41.060 5.060 42.240 ;
        RECT 0.680 39.460 1.860 40.640 ;
        RECT 6.660 39.460 7.840 40.640 ;
        RECT 10.310 40.115 11.670 51.855 ;
        RECT 66.450 50.755 71.010 51.855 ;
        RECT 66.450 47.880 67.810 50.755 ;
        RECT 69.650 47.880 71.010 50.755 ;
        RECT 66.450 46.280 71.010 47.880 ;
        RECT 66.450 40.125 67.810 46.280 ;
        RECT 69.650 40.115 71.010 46.280 ;
        RECT 98.590 40.125 99.950 51.865 ;
        RECT 140.430 40.125 141.790 51.865 ;
        RECT 170.615 51.855 173.930 51.865 ;
        RECT 169.370 50.755 173.930 51.855 ;
        RECT 169.370 47.880 170.730 50.755 ;
        RECT 172.570 47.880 173.930 50.755 ;
        RECT 169.370 46.280 173.930 47.880 ;
        RECT 169.370 40.115 170.730 46.280 ;
        RECT 172.570 40.125 173.930 46.280 ;
        RECT 228.710 40.115 230.070 51.855 ;
        RECT 235.320 50.660 236.920 51.840 ;
        RECT 232.540 49.060 233.720 50.240 ;
        RECT 238.520 49.060 239.700 50.240 ;
        RECT 235.320 47.460 236.920 48.640 ;
        RECT 232.540 45.860 233.720 47.040 ;
        RECT 238.520 45.860 239.700 47.040 ;
        RECT 235.320 44.260 236.920 45.440 ;
        RECT 232.540 42.660 233.720 43.840 ;
        RECT 238.520 42.660 239.700 43.840 ;
        RECT 235.320 41.060 236.920 42.240 ;
        RECT 232.540 39.460 233.720 40.640 ;
        RECT 238.520 39.460 239.700 40.640 ;
        RECT 3.460 37.860 5.060 39.040 ;
        RECT 67.740 38.265 69.785 39.390 ;
        RECT 170.595 38.265 172.640 39.390 ;
        RECT 66.450 38.255 69.785 38.265 ;
        RECT 0.680 36.260 1.860 37.440 ;
        RECT 6.660 36.260 7.840 37.440 ;
        RECT 3.460 34.660 5.060 35.840 ;
        RECT 0.680 33.060 1.860 34.240 ;
        RECT 6.660 33.060 7.840 34.240 ;
        RECT 3.460 31.460 5.060 32.640 ;
        RECT 0.680 29.860 1.860 31.040 ;
        RECT 6.660 29.860 7.840 31.040 ;
        RECT 3.460 28.260 5.060 29.440 ;
        RECT 0.680 26.660 1.860 27.840 ;
        RECT 6.660 26.660 7.840 27.840 ;
        RECT 10.310 26.515 11.670 38.255 ;
        RECT 66.450 37.790 71.010 38.255 ;
        RECT 66.450 34.925 67.810 37.790 ;
        RECT 69.650 34.925 71.010 37.790 ;
        RECT 66.450 33.325 71.010 34.925 ;
        RECT 66.450 30.465 67.810 33.325 ;
        RECT 69.650 30.465 71.010 33.325 ;
        RECT 66.450 28.865 71.010 30.465 ;
        RECT 66.450 26.525 67.810 28.865 ;
        RECT 69.650 26.515 71.010 28.865 ;
        RECT 98.590 26.525 99.950 38.265 ;
        RECT 140.430 26.525 141.790 38.265 ;
        RECT 170.595 38.255 173.930 38.265 ;
        RECT 169.370 37.790 173.930 38.255 ;
        RECT 169.370 34.925 170.730 37.790 ;
        RECT 172.570 34.925 173.930 37.790 ;
        RECT 169.370 33.325 173.930 34.925 ;
        RECT 169.370 30.465 170.730 33.325 ;
        RECT 172.570 30.465 173.930 33.325 ;
        RECT 169.370 28.865 173.930 30.465 ;
        RECT 169.370 26.515 170.730 28.865 ;
        RECT 172.570 26.525 173.930 28.865 ;
        RECT 228.710 26.515 230.070 38.255 ;
        RECT 235.320 37.860 236.920 39.040 ;
        RECT 232.540 36.260 233.720 37.440 ;
        RECT 238.520 36.260 239.700 37.440 ;
        RECT 235.320 34.660 236.920 35.840 ;
        RECT 232.540 33.060 233.720 34.240 ;
        RECT 238.520 33.060 239.700 34.240 ;
        RECT 235.320 31.460 236.920 32.640 ;
        RECT 232.540 29.860 233.720 31.040 ;
        RECT 238.520 29.860 239.700 31.040 ;
        RECT 235.320 28.260 236.920 29.440 ;
        RECT 232.540 26.660 233.720 27.840 ;
        RECT 238.520 26.660 239.700 27.840 ;
        RECT 3.460 25.060 5.060 26.240 ;
        RECT 0.680 23.460 1.860 24.640 ;
        RECT 6.660 23.460 7.840 24.640 ;
        RECT 3.460 21.860 5.060 23.040 ;
        RECT 10.310 22.455 11.670 24.665 ;
        RECT 66.450 21.985 67.810 25.590 ;
        RECT 69.650 22.455 71.010 24.665 ;
        RECT 0.680 20.260 1.860 21.440 ;
        RECT 6.660 20.260 7.840 21.440 ;
        RECT 66.450 20.385 69.725 21.985 ;
        RECT 3.460 18.660 5.060 19.840 ;
        RECT 0.680 17.060 1.860 18.240 ;
        RECT 6.660 17.060 7.840 18.240 ;
        RECT 3.460 15.460 5.060 16.640 ;
        RECT 0.680 13.860 1.860 15.040 ;
        RECT 6.660 13.860 7.840 15.040 ;
        RECT 10.310 11.800 11.670 19.805 ;
        RECT 66.450 17.990 67.810 20.385 ;
        RECT 69.650 17.515 71.010 19.805 ;
        RECT 98.590 17.990 99.950 25.590 ;
        RECT 140.430 17.990 141.790 25.590 ;
        RECT 169.370 22.455 170.730 24.665 ;
        RECT 172.570 21.985 173.930 25.590 ;
        RECT 235.320 25.060 236.920 26.240 ;
        RECT 228.710 22.455 230.070 24.665 ;
        RECT 232.540 23.460 233.720 24.640 ;
        RECT 238.520 23.460 239.700 24.640 ;
        RECT 170.655 20.385 173.930 21.985 ;
        RECT 235.320 21.860 236.920 23.040 ;
        RECT 67.735 15.915 71.010 17.515 ;
        RECT 66.450 13.045 67.810 15.135 ;
        RECT 69.650 13.045 71.010 15.915 ;
        RECT 169.370 17.515 170.730 19.805 ;
        RECT 172.570 17.990 173.930 20.385 ;
        RECT 232.540 20.260 233.720 21.440 ;
        RECT 238.520 20.260 239.700 21.440 ;
        RECT 169.370 15.915 172.645 17.515 ;
        RECT 66.450 11.800 71.010 13.045 ;
        RECT 98.590 11.800 99.950 15.135 ;
        RECT 10.310 10.440 15.005 11.800 ;
        RECT 17.860 10.440 25.460 11.800 ;
        RECT 26.395 10.440 38.135 11.800 ;
        RECT 39.995 10.440 51.735 11.800 ;
        RECT 53.585 10.440 55.795 11.800 ;
        RECT 58.445 11.445 74.345 11.800 ;
        RECT 58.445 10.440 67.810 11.445 ;
        RECT 69.650 10.440 74.345 11.445 ;
        RECT 77.200 10.440 84.800 11.800 ;
        RECT 85.725 10.440 87.935 11.800 ;
        RECT 90.585 10.440 99.950 11.800 ;
        RECT 140.430 11.800 141.790 15.135 ;
        RECT 169.370 13.045 170.730 15.915 ;
        RECT 172.570 13.045 173.930 15.135 ;
        RECT 169.370 11.800 173.930 13.045 ;
        RECT 228.710 11.800 230.070 19.805 ;
        RECT 235.320 18.660 236.920 19.840 ;
        RECT 232.540 17.060 233.720 18.240 ;
        RECT 238.520 17.060 239.700 18.240 ;
        RECT 235.320 15.460 236.920 16.640 ;
        RECT 232.540 13.860 233.720 15.040 ;
        RECT 238.520 13.860 239.700 15.040 ;
        RECT 140.430 10.440 149.795 11.800 ;
        RECT 152.445 10.440 154.655 11.800 ;
        RECT 155.580 10.440 163.180 11.800 ;
        RECT 166.035 11.445 181.935 11.800 ;
        RECT 166.035 10.440 170.730 11.445 ;
        RECT 172.570 10.440 181.935 11.445 ;
        RECT 184.585 10.440 186.795 11.800 ;
        RECT 188.645 10.440 200.385 11.800 ;
        RECT 202.245 10.440 213.985 11.800 ;
        RECT 214.920 10.440 222.520 11.800 ;
        RECT 225.375 10.440 230.070 11.800 ;
        RECT 9.780 6.100 10.960 7.280 ;
        RECT 12.980 6.100 14.160 7.280 ;
        RECT 16.180 6.100 17.360 7.280 ;
        RECT 19.380 6.100 20.560 7.280 ;
        RECT 22.580 6.100 23.760 7.280 ;
        RECT 25.780 6.100 26.960 7.280 ;
        RECT 28.980 6.100 30.160 7.280 ;
        RECT 32.180 6.100 33.360 7.280 ;
        RECT 35.380 6.100 36.560 7.280 ;
        RECT 38.580 6.100 39.760 7.280 ;
        RECT 41.780 6.100 42.960 7.280 ;
        RECT 44.980 6.100 46.160 7.280 ;
        RECT 48.180 6.100 49.360 7.280 ;
        RECT 51.380 6.100 52.560 7.280 ;
        RECT 54.580 6.100 55.760 7.280 ;
        RECT 57.780 6.100 58.960 7.280 ;
        RECT 60.980 6.100 62.160 7.280 ;
        RECT 64.180 6.100 65.360 7.280 ;
        RECT 67.380 6.100 68.560 7.280 ;
        RECT 70.580 6.100 71.760 7.280 ;
        RECT 73.780 6.100 74.960 7.280 ;
        RECT 76.980 6.100 78.160 7.280 ;
        RECT 80.180 6.100 81.360 7.280 ;
        RECT 83.380 6.100 84.560 7.280 ;
        RECT 86.580 6.100 87.760 7.280 ;
        RECT 89.780 6.100 90.960 7.280 ;
        RECT 92.980 6.100 94.160 7.280 ;
        RECT 96.180 6.100 97.360 7.280 ;
        RECT 99.380 6.100 100.560 7.280 ;
        RECT 102.580 6.100 103.760 7.280 ;
        RECT 105.780 6.100 106.960 7.280 ;
        RECT 108.980 6.100 110.160 7.280 ;
        RECT 112.180 6.100 113.360 7.280 ;
        RECT 115.380 6.100 116.560 7.280 ;
        RECT 123.820 6.100 125.000 7.280 ;
        RECT 127.020 6.100 128.200 7.280 ;
        RECT 130.220 6.100 131.400 7.280 ;
        RECT 133.420 6.100 134.600 7.280 ;
        RECT 136.620 6.100 137.800 7.280 ;
        RECT 139.820 6.100 141.000 7.280 ;
        RECT 143.020 6.100 144.200 7.280 ;
        RECT 146.220 6.100 147.400 7.280 ;
        RECT 149.420 6.100 150.600 7.280 ;
        RECT 152.620 6.100 153.800 7.280 ;
        RECT 155.820 6.100 157.000 7.280 ;
        RECT 159.020 6.100 160.200 7.280 ;
        RECT 162.220 6.100 163.400 7.280 ;
        RECT 165.420 6.100 166.600 7.280 ;
        RECT 168.620 6.100 169.800 7.280 ;
        RECT 171.820 6.100 173.000 7.280 ;
        RECT 175.020 6.100 176.200 7.280 ;
        RECT 178.220 6.100 179.400 7.280 ;
        RECT 181.420 6.100 182.600 7.280 ;
        RECT 184.620 6.100 185.800 7.280 ;
        RECT 187.820 6.100 189.000 7.280 ;
        RECT 191.020 6.100 192.200 7.280 ;
        RECT 194.220 6.100 195.400 7.280 ;
        RECT 197.420 6.100 198.600 7.280 ;
        RECT 200.620 6.100 201.800 7.280 ;
        RECT 203.820 6.100 205.000 7.280 ;
        RECT 207.020 6.100 208.200 7.280 ;
        RECT 210.220 6.100 211.400 7.280 ;
        RECT 213.420 6.100 214.600 7.280 ;
        RECT 216.620 6.100 217.800 7.280 ;
        RECT 219.820 6.100 221.000 7.280 ;
        RECT 223.020 6.100 224.200 7.280 ;
        RECT 226.220 6.100 227.400 7.280 ;
        RECT 229.420 6.100 230.600 7.280 ;
        RECT 8.180 2.900 9.360 4.500 ;
        RECT 11.380 2.900 12.560 4.500 ;
        RECT 14.580 2.900 15.760 4.500 ;
        RECT 17.780 2.900 18.960 4.500 ;
        RECT 20.980 2.900 22.160 4.500 ;
        RECT 24.180 2.900 25.360 4.500 ;
        RECT 27.380 2.900 28.560 4.500 ;
        RECT 30.580 2.900 31.760 4.500 ;
        RECT 33.780 2.900 34.960 4.500 ;
        RECT 36.980 2.900 38.160 4.500 ;
        RECT 40.180 2.900 41.360 4.500 ;
        RECT 43.380 2.900 44.560 4.500 ;
        RECT 46.580 2.900 47.760 4.500 ;
        RECT 49.780 2.900 50.960 4.500 ;
        RECT 52.980 2.900 54.160 4.500 ;
        RECT 56.180 2.900 57.360 4.500 ;
        RECT 59.380 2.900 60.560 4.500 ;
        RECT 62.580 2.900 63.760 4.500 ;
        RECT 65.780 2.900 66.960 4.500 ;
        RECT 68.980 2.900 70.160 4.500 ;
        RECT 72.180 2.900 73.360 4.500 ;
        RECT 75.380 2.900 76.560 4.500 ;
        RECT 78.580 2.900 79.760 4.500 ;
        RECT 81.780 2.900 82.960 4.500 ;
        RECT 84.980 2.900 86.160 4.500 ;
        RECT 88.180 2.900 89.360 4.500 ;
        RECT 91.380 2.900 92.560 4.500 ;
        RECT 94.580 2.900 95.760 4.500 ;
        RECT 97.780 2.900 98.960 4.500 ;
        RECT 100.980 2.900 102.160 4.500 ;
        RECT 104.180 2.900 105.360 4.500 ;
        RECT 107.380 2.900 108.560 4.500 ;
        RECT 110.580 2.900 111.760 4.500 ;
        RECT 113.780 2.900 114.960 4.500 ;
        RECT 116.980 2.900 118.160 4.500 ;
        RECT 122.220 2.900 123.400 4.500 ;
        RECT 125.420 2.900 126.600 4.500 ;
        RECT 128.620 2.900 129.800 4.500 ;
        RECT 131.820 2.900 133.000 4.500 ;
        RECT 135.020 2.900 136.200 4.500 ;
        RECT 138.220 2.900 139.400 4.500 ;
        RECT 141.420 2.900 142.600 4.500 ;
        RECT 144.620 2.900 145.800 4.500 ;
        RECT 147.820 2.900 149.000 4.500 ;
        RECT 151.020 2.900 152.200 4.500 ;
        RECT 154.220 2.900 155.400 4.500 ;
        RECT 157.420 2.900 158.600 4.500 ;
        RECT 160.620 2.900 161.800 4.500 ;
        RECT 163.820 2.900 165.000 4.500 ;
        RECT 167.020 2.900 168.200 4.500 ;
        RECT 170.220 2.900 171.400 4.500 ;
        RECT 173.420 2.900 174.600 4.500 ;
        RECT 176.620 2.900 177.800 4.500 ;
        RECT 179.820 2.900 181.000 4.500 ;
        RECT 183.020 2.900 184.200 4.500 ;
        RECT 186.220 2.900 187.400 4.500 ;
        RECT 189.420 2.900 190.600 4.500 ;
        RECT 192.620 2.900 193.800 4.500 ;
        RECT 195.820 2.900 197.000 4.500 ;
        RECT 199.020 2.900 200.200 4.500 ;
        RECT 202.220 2.900 203.400 4.500 ;
        RECT 205.420 2.900 206.600 4.500 ;
        RECT 208.620 2.900 209.800 4.500 ;
        RECT 211.820 2.900 213.000 4.500 ;
        RECT 215.020 2.900 216.200 4.500 ;
        RECT 218.220 2.900 219.400 4.500 ;
        RECT 221.420 2.900 222.600 4.500 ;
        RECT 224.620 2.900 225.800 4.500 ;
        RECT 227.820 2.900 229.000 4.500 ;
        RECT 231.020 2.900 232.200 4.500 ;
        RECT 9.780 0.120 10.960 1.300 ;
        RECT 12.980 0.120 14.160 1.300 ;
        RECT 16.180 0.120 17.360 1.300 ;
        RECT 19.380 0.120 20.560 1.300 ;
        RECT 22.580 0.120 23.760 1.300 ;
        RECT 25.780 0.120 26.960 1.300 ;
        RECT 28.980 0.120 30.160 1.300 ;
        RECT 32.180 0.120 33.360 1.300 ;
        RECT 35.380 0.120 36.560 1.300 ;
        RECT 38.580 0.120 39.760 1.300 ;
        RECT 41.780 0.120 42.960 1.300 ;
        RECT 44.980 0.120 46.160 1.300 ;
        RECT 48.180 0.120 49.360 1.300 ;
        RECT 51.380 0.120 52.560 1.300 ;
        RECT 54.580 0.120 55.760 1.300 ;
        RECT 57.780 0.120 58.960 1.300 ;
        RECT 60.980 0.120 62.160 1.300 ;
        RECT 64.180 0.120 65.360 1.300 ;
        RECT 67.380 0.120 68.560 1.300 ;
        RECT 70.580 0.120 71.760 1.300 ;
        RECT 73.780 0.120 74.960 1.300 ;
        RECT 76.980 0.120 78.160 1.300 ;
        RECT 80.180 0.120 81.360 1.300 ;
        RECT 83.380 0.120 84.560 1.300 ;
        RECT 86.580 0.120 87.760 1.300 ;
        RECT 89.780 0.120 90.960 1.300 ;
        RECT 92.980 0.120 94.160 1.300 ;
        RECT 96.180 0.120 97.360 1.300 ;
        RECT 99.380 0.120 100.560 1.300 ;
        RECT 102.580 0.120 103.760 1.300 ;
        RECT 105.780 0.120 106.960 1.300 ;
        RECT 108.980 0.120 110.160 1.300 ;
        RECT 112.180 0.120 113.360 1.300 ;
        RECT 115.380 0.120 116.560 1.300 ;
        RECT 123.820 0.120 125.000 1.300 ;
        RECT 127.020 0.120 128.200 1.300 ;
        RECT 130.220 0.120 131.400 1.300 ;
        RECT 133.420 0.120 134.600 1.300 ;
        RECT 136.620 0.120 137.800 1.300 ;
        RECT 139.820 0.120 141.000 1.300 ;
        RECT 143.020 0.120 144.200 1.300 ;
        RECT 146.220 0.120 147.400 1.300 ;
        RECT 149.420 0.120 150.600 1.300 ;
        RECT 152.620 0.120 153.800 1.300 ;
        RECT 155.820 0.120 157.000 1.300 ;
        RECT 159.020 0.120 160.200 1.300 ;
        RECT 162.220 0.120 163.400 1.300 ;
        RECT 165.420 0.120 166.600 1.300 ;
        RECT 168.620 0.120 169.800 1.300 ;
        RECT 171.820 0.120 173.000 1.300 ;
        RECT 175.020 0.120 176.200 1.300 ;
        RECT 178.220 0.120 179.400 1.300 ;
        RECT 181.420 0.120 182.600 1.300 ;
        RECT 184.620 0.120 185.800 1.300 ;
        RECT 187.820 0.120 189.000 1.300 ;
        RECT 191.020 0.120 192.200 1.300 ;
        RECT 194.220 0.120 195.400 1.300 ;
        RECT 197.420 0.120 198.600 1.300 ;
        RECT 200.620 0.120 201.800 1.300 ;
        RECT 203.820 0.120 205.000 1.300 ;
        RECT 207.020 0.120 208.200 1.300 ;
        RECT 210.220 0.120 211.400 1.300 ;
        RECT 213.420 0.120 214.600 1.300 ;
        RECT 216.620 0.120 217.800 1.300 ;
        RECT 219.820 0.120 221.000 1.300 ;
        RECT 223.020 0.120 224.200 1.300 ;
        RECT 226.220 0.120 227.400 1.300 ;
        RECT 229.420 0.120 230.600 1.300 ;
      LAYER via4 ;
        RECT 10.310 120.980 19.670 122.340 ;
        RECT 22.330 120.980 24.530 122.340 ;
        RECT 26.390 120.980 38.120 122.340 ;
        RECT 39.990 120.980 51.720 122.340 ;
        RECT 53.590 120.980 60.255 122.340 ;
        RECT 63.120 120.980 67.810 122.340 ;
        RECT 10.310 117.650 11.670 120.980 ;
        RECT 10.310 108.120 11.670 114.785 ;
        RECT 66.450 112.980 67.810 120.980 ;
        RECT 69.650 120.980 79.010 122.340 ;
        RECT 81.670 120.980 83.870 122.340 ;
        RECT 85.730 120.980 92.395 122.340 ;
        RECT 95.260 120.980 99.950 122.340 ;
        RECT 69.650 117.650 71.010 120.980 ;
        RECT 66.450 108.120 67.810 110.320 ;
        RECT 69.650 108.120 71.010 114.785 ;
        RECT 98.590 112.980 99.950 120.980 ;
        RECT 140.430 120.980 145.120 122.340 ;
        RECT 147.985 120.980 154.650 122.340 ;
        RECT 156.510 120.980 158.710 122.340 ;
        RECT 161.370 120.980 170.730 122.340 ;
        RECT 140.430 112.980 141.790 120.980 ;
        RECT 169.370 117.650 170.730 120.980 ;
        RECT 172.570 120.980 177.260 122.340 ;
        RECT 180.125 120.980 186.790 122.340 ;
        RECT 188.660 120.980 200.390 122.340 ;
        RECT 202.260 120.980 213.990 122.340 ;
        RECT 215.850 120.980 218.050 122.340 ;
        RECT 220.710 120.980 230.070 122.340 ;
        RECT 98.590 108.120 99.950 110.320 ;
        RECT 140.430 108.120 141.790 110.320 ;
        RECT 169.370 108.120 170.730 114.785 ;
        RECT 172.570 112.980 173.930 120.980 ;
        RECT 228.710 117.650 230.070 120.980 ;
        RECT 172.570 108.120 173.930 110.320 ;
        RECT 228.710 108.120 230.070 114.785 ;
        RECT 10.310 94.520 11.670 106.250 ;
        RECT 66.450 94.530 67.810 106.260 ;
        RECT 69.650 94.520 71.010 106.250 ;
        RECT 98.590 94.530 99.950 106.260 ;
        RECT 140.430 94.530 141.790 106.260 ;
        RECT 169.370 94.520 170.730 106.250 ;
        RECT 172.570 94.530 173.930 106.260 ;
        RECT 228.710 94.520 230.070 106.250 ;
        RECT 10.310 80.920 11.670 92.650 ;
        RECT 66.450 80.930 67.810 92.660 ;
        RECT 69.650 80.920 71.010 92.650 ;
        RECT 98.590 80.930 99.950 92.660 ;
        RECT 140.430 80.930 141.790 92.660 ;
        RECT 169.370 80.920 170.730 92.650 ;
        RECT 172.570 80.930 173.930 92.660 ;
        RECT 228.710 80.920 230.070 92.650 ;
        RECT 10.310 67.320 11.670 79.050 ;
        RECT 66.450 67.330 67.810 79.060 ;
        RECT 69.650 67.320 71.010 79.050 ;
        RECT 98.590 67.330 99.950 79.060 ;
        RECT 140.430 67.330 141.790 79.060 ;
        RECT 169.370 67.320 170.730 79.050 ;
        RECT 172.570 67.330 173.930 79.060 ;
        RECT 228.710 67.320 230.070 79.050 ;
        RECT 10.310 53.720 11.670 65.450 ;
        RECT 66.450 53.730 67.810 65.460 ;
        RECT 69.650 53.720 71.010 65.450 ;
        RECT 98.590 53.730 99.950 65.460 ;
        RECT 140.430 53.730 141.790 65.460 ;
        RECT 169.370 53.720 170.730 65.450 ;
        RECT 172.570 53.730 173.930 65.460 ;
        RECT 228.710 53.720 230.070 65.450 ;
        RECT 10.310 40.120 11.670 51.850 ;
        RECT 66.450 40.130 67.810 51.860 ;
        RECT 69.650 40.120 71.010 51.850 ;
        RECT 98.590 40.130 99.950 51.860 ;
        RECT 140.430 40.130 141.790 51.860 ;
        RECT 169.370 40.120 170.730 51.850 ;
        RECT 172.570 40.130 173.930 51.860 ;
        RECT 228.710 40.120 230.070 51.850 ;
        RECT 10.310 26.520 11.670 38.250 ;
        RECT 66.450 26.530 67.810 38.260 ;
        RECT 69.650 26.520 71.010 38.250 ;
        RECT 98.590 26.530 99.950 38.260 ;
        RECT 140.430 26.530 141.790 38.260 ;
        RECT 169.370 26.520 170.730 38.250 ;
        RECT 172.570 26.530 173.930 38.260 ;
        RECT 228.710 26.520 230.070 38.250 ;
        RECT 10.310 22.460 11.670 24.660 ;
        RECT 10.310 11.800 11.670 19.800 ;
        RECT 66.450 17.995 67.810 24.660 ;
        RECT 69.650 22.460 71.010 24.660 ;
        RECT 66.450 11.800 67.810 15.130 ;
        RECT 17.865 10.440 24.530 11.800 ;
        RECT 26.400 10.440 38.130 11.800 ;
        RECT 40.000 10.440 51.730 11.800 ;
        RECT 53.590 10.440 55.790 11.800 ;
        RECT 58.450 10.440 67.810 11.800 ;
        RECT 69.650 11.800 71.010 19.800 ;
        RECT 98.590 17.995 99.950 24.660 ;
        RECT 140.430 17.995 141.790 24.660 ;
        RECT 169.370 22.460 170.730 24.660 ;
        RECT 98.590 11.800 99.950 15.130 ;
        RECT 77.205 10.440 83.870 11.800 ;
        RECT 85.730 10.440 87.930 11.800 ;
        RECT 90.590 10.440 99.950 11.800 ;
        RECT 140.430 11.800 141.790 15.130 ;
        RECT 169.370 11.800 170.730 19.800 ;
        RECT 172.570 17.995 173.930 24.660 ;
        RECT 228.710 22.460 230.070 24.660 ;
        RECT 152.450 10.440 154.650 11.800 ;
        RECT 156.510 10.440 163.175 11.800 ;
        RECT 166.040 10.440 170.730 11.800 ;
        RECT 172.570 11.800 173.930 15.130 ;
        RECT 228.710 11.800 230.070 19.800 ;
        RECT 184.590 10.440 186.790 11.800 ;
        RECT 188.650 10.440 200.380 11.800 ;
        RECT 202.250 10.440 213.980 11.800 ;
        RECT 215.850 10.440 222.515 11.800 ;
        RECT 225.380 10.440 230.070 11.800 ;
      LAYER met5 ;
        RECT 1.860 127.250 3.460 128.375 ;
        RECT 0.560 125.650 3.460 127.250 ;
        RECT 5.060 127.250 6.660 128.410 ;
        RECT 233.720 127.250 235.320 128.410 ;
        RECT 5.060 125.650 7.960 127.250 ;
        RECT 232.420 125.650 235.320 127.250 ;
        RECT 236.920 127.250 238.520 128.375 ;
        RECT 236.920 125.650 239.820 127.250 ;
        RECT 1.860 124.050 6.660 125.650 ;
        RECT 233.720 124.050 238.520 125.650 ;
        RECT 0.560 122.450 3.460 124.050 ;
        RECT 5.060 122.450 7.960 124.050 ;
        RECT 1.860 120.850 6.660 122.450 ;
        RECT 10.190 121.790 67.930 122.460 ;
        RECT 69.530 121.790 100.070 122.460 ;
        RECT 10.190 120.860 100.070 121.790 ;
        RECT 0.560 119.250 3.460 120.850 ;
        RECT 5.060 119.250 7.960 120.850 ;
        RECT 10.190 119.250 11.790 120.860 ;
        RECT 13.800 119.250 15.400 120.860 ;
        RECT 18.065 119.250 19.670 120.860 ;
        RECT 22.330 119.250 23.930 120.860 ;
        RECT 1.860 117.650 6.660 119.250 ;
        RECT 10.190 119.130 23.930 119.250 ;
        RECT 26.990 119.250 28.590 120.860 ;
        RECT 31.460 119.250 33.060 120.860 ;
        RECT 35.930 119.250 37.530 120.860 ;
        RECT 26.990 119.130 37.530 119.250 ;
        RECT 40.590 119.250 42.190 120.860 ;
        RECT 45.060 119.250 46.660 120.860 ;
        RECT 49.530 119.250 51.130 120.860 ;
        RECT 40.590 119.130 51.130 119.250 ;
        RECT 54.190 119.250 55.790 120.860 ;
        RECT 58.655 119.250 60.255 120.860 ;
        RECT 63.120 119.250 64.720 120.860 ;
        RECT 54.190 119.130 64.720 119.250 ;
        RECT 10.190 118.850 64.720 119.130 ;
        RECT 66.330 120.190 71.130 120.860 ;
        RECT 66.330 118.850 67.930 120.190 ;
        RECT 10.190 117.650 67.930 118.850 ;
        RECT 0.560 116.050 3.460 117.650 ;
        RECT 5.060 116.050 11.790 117.650 ;
        RECT 1.860 114.450 6.660 116.050 ;
        RECT 10.190 114.785 11.790 116.050 ;
        RECT 13.400 117.530 67.930 117.650 ;
        RECT 13.400 114.790 23.920 117.530 ;
        RECT 27.000 114.790 37.520 117.530 ;
        RECT 40.600 114.790 51.120 117.530 ;
        RECT 54.200 117.250 67.930 117.530 ;
        RECT 54.200 114.790 64.720 117.250 ;
        RECT 13.400 114.785 64.720 114.790 ;
        RECT 10.190 114.585 64.720 114.785 ;
        RECT 66.330 114.635 67.930 117.250 ;
        RECT 69.530 119.250 71.130 120.190 ;
        RECT 73.140 119.250 74.740 120.860 ;
        RECT 77.405 119.250 79.010 120.860 ;
        RECT 81.670 119.250 83.270 120.860 ;
        RECT 69.530 119.130 83.270 119.250 ;
        RECT 86.330 119.250 87.930 120.860 ;
        RECT 90.795 119.250 92.395 120.860 ;
        RECT 95.260 119.250 96.860 120.860 ;
        RECT 86.330 119.130 96.860 119.250 ;
        RECT 69.530 118.850 96.860 119.130 ;
        RECT 98.470 118.850 100.070 120.860 ;
        RECT 69.530 117.650 100.070 118.850 ;
        RECT 69.530 114.785 71.130 117.650 ;
        RECT 72.740 117.530 100.070 117.650 ;
        RECT 72.740 114.790 83.260 117.530 ;
        RECT 86.340 117.250 100.070 117.530 ;
        RECT 86.340 114.790 96.860 117.250 ;
        RECT 72.740 114.785 96.860 114.790 ;
        RECT 69.530 114.635 96.860 114.785 ;
        RECT 66.330 114.585 96.860 114.635 ;
        RECT 98.470 114.585 100.070 117.250 ;
        RECT 0.560 112.850 3.460 114.450 ;
        RECT 5.060 112.850 7.960 114.450 ;
        RECT 10.190 113.190 100.070 114.585 ;
        RECT 10.190 113.185 23.920 113.190 ;
        RECT 1.860 111.250 6.660 112.850 ;
        RECT 10.190 111.250 11.790 113.185 ;
        RECT 0.560 109.650 3.460 111.250 ;
        RECT 5.060 110.320 11.790 111.250 ;
        RECT 13.400 110.450 23.920 113.185 ;
        RECT 27.000 110.450 37.520 113.190 ;
        RECT 40.600 110.450 51.120 113.190 ;
        RECT 54.200 113.185 83.260 113.190 ;
        RECT 54.200 113.035 71.130 113.185 ;
        RECT 54.200 112.980 67.930 113.035 ;
        RECT 54.200 110.450 64.720 112.980 ;
        RECT 13.400 110.320 64.720 110.450 ;
        RECT 66.330 110.320 67.930 112.980 ;
        RECT 5.060 109.650 67.930 110.320 ;
        RECT 1.860 108.050 6.660 109.650 ;
        RECT 10.190 109.025 67.930 109.650 ;
        RECT 69.530 110.320 71.130 113.035 ;
        RECT 72.740 110.450 83.260 113.185 ;
        RECT 86.340 112.980 100.070 113.190 ;
        RECT 86.340 110.450 96.860 112.980 ;
        RECT 72.740 110.320 96.860 110.450 ;
        RECT 98.470 110.320 100.070 112.980 ;
        RECT 69.530 109.025 100.070 110.320 ;
        RECT 10.190 108.850 100.070 109.025 ;
        RECT 10.190 108.730 23.930 108.850 ;
        RECT 10.190 108.720 15.120 108.730 ;
        RECT 0.560 106.450 3.460 108.050 ;
        RECT 5.060 106.450 7.960 108.050 ;
        RECT 1.860 104.850 6.660 106.450 ;
        RECT 10.190 105.660 11.790 108.720 ;
        RECT 13.520 105.660 15.120 108.720 ;
        RECT 10.190 105.650 15.120 105.660 ;
        RECT 17.860 105.650 19.460 108.730 ;
        RECT 22.200 108.720 23.930 108.730 ;
        RECT 26.990 108.730 37.530 108.850 ;
        RECT 26.990 108.720 28.720 108.730 ;
        RECT 22.200 105.660 23.800 108.720 ;
        RECT 27.120 105.660 28.720 108.720 ;
        RECT 22.200 105.650 23.930 105.660 ;
        RECT 10.190 105.530 23.930 105.650 ;
        RECT 26.990 105.650 28.720 105.660 ;
        RECT 31.460 105.650 33.060 108.730 ;
        RECT 35.800 108.720 37.530 108.730 ;
        RECT 40.590 108.730 51.130 108.850 ;
        RECT 40.590 108.720 42.320 108.730 ;
        RECT 35.800 105.660 37.400 108.720 ;
        RECT 40.720 105.660 42.320 108.720 ;
        RECT 35.800 105.650 37.530 105.660 ;
        RECT 26.990 105.530 37.530 105.650 ;
        RECT 40.590 105.650 42.320 105.660 ;
        RECT 45.060 105.650 46.660 108.730 ;
        RECT 49.400 108.720 51.130 108.730 ;
        RECT 54.190 108.730 83.270 108.850 ;
        RECT 54.190 108.720 55.920 108.730 ;
        RECT 49.400 105.660 51.000 108.720 ;
        RECT 54.320 105.660 55.920 108.720 ;
        RECT 49.400 105.650 51.130 105.660 ;
        RECT 40.590 105.530 51.130 105.650 ;
        RECT 54.190 105.650 55.920 105.660 ;
        RECT 58.660 105.650 60.260 108.730 ;
        RECT 63.000 108.720 74.460 108.730 ;
        RECT 63.000 105.660 64.600 108.720 ;
        RECT 66.330 107.425 71.130 108.720 ;
        RECT 66.330 105.660 67.930 107.425 ;
        RECT 63.000 105.650 67.930 105.660 ;
        RECT 54.190 105.530 67.930 105.650 ;
        RECT 10.190 104.850 67.930 105.530 ;
        RECT 0.560 103.250 3.460 104.850 ;
        RECT 5.060 104.550 67.930 104.850 ;
        RECT 69.530 105.660 71.130 107.425 ;
        RECT 72.860 105.660 74.460 108.720 ;
        RECT 69.530 105.650 74.460 105.660 ;
        RECT 77.200 105.650 78.800 108.730 ;
        RECT 81.540 108.720 83.270 108.730 ;
        RECT 86.330 108.730 100.070 108.850 ;
        RECT 86.330 108.720 88.060 108.730 ;
        RECT 81.540 105.660 83.140 108.720 ;
        RECT 86.460 105.660 88.060 108.720 ;
        RECT 81.540 105.650 83.270 105.660 ;
        RECT 69.530 105.530 83.270 105.650 ;
        RECT 86.330 105.650 88.060 105.660 ;
        RECT 90.800 105.650 92.400 108.730 ;
        RECT 95.140 108.720 100.070 108.730 ;
        RECT 95.140 105.660 96.740 108.720 ;
        RECT 98.470 105.660 100.070 108.720 ;
        RECT 95.140 105.650 100.070 105.660 ;
        RECT 86.330 105.530 100.070 105.650 ;
        RECT 69.530 104.550 100.070 105.530 ;
        RECT 5.060 104.060 100.070 104.550 ;
        RECT 5.060 103.250 11.790 104.060 ;
        RECT 1.860 101.650 6.660 103.250 ;
        RECT 0.560 100.050 3.460 101.650 ;
        RECT 5.060 100.050 7.960 101.650 ;
        RECT 10.190 101.190 11.790 103.250 ;
        RECT 13.400 103.930 64.720 104.060 ;
        RECT 13.400 101.190 23.920 103.930 ;
        RECT 27.000 101.190 37.520 103.930 ;
        RECT 40.600 101.190 51.120 103.930 ;
        RECT 54.200 101.190 64.720 103.930 ;
        RECT 66.330 102.950 71.130 104.060 ;
        RECT 66.330 101.190 67.930 102.950 ;
        RECT 10.190 100.135 67.930 101.190 ;
        RECT 69.530 101.190 71.130 102.950 ;
        RECT 72.740 103.930 96.860 104.060 ;
        RECT 72.740 101.190 83.260 103.930 ;
        RECT 86.340 101.190 96.860 103.930 ;
        RECT 98.470 101.190 100.070 104.060 ;
        RECT 69.530 100.135 100.070 101.190 ;
        RECT 1.860 98.450 6.660 100.050 ;
        RECT 10.190 99.590 100.070 100.135 ;
        RECT 10.190 98.450 11.790 99.590 ;
        RECT 0.560 96.850 3.460 98.450 ;
        RECT 5.060 96.850 11.790 98.450 ;
        RECT 1.860 95.250 6.660 96.850 ;
        RECT 10.190 96.720 11.790 96.850 ;
        RECT 13.400 96.850 23.920 99.590 ;
        RECT 27.000 96.850 37.520 99.590 ;
        RECT 40.600 96.850 51.120 99.590 ;
        RECT 54.200 96.850 64.720 99.590 ;
        RECT 13.400 96.720 64.720 96.850 ;
        RECT 66.330 98.535 71.130 99.590 ;
        RECT 66.330 96.720 67.930 98.535 ;
        RECT 10.190 95.250 67.930 96.720 ;
        RECT 0.560 93.650 3.460 95.250 ;
        RECT 5.060 93.650 7.960 95.250 ;
        RECT 10.190 95.130 23.930 95.250 ;
        RECT 10.190 95.120 15.120 95.130 ;
        RECT 1.860 92.050 6.660 93.650 ;
        RECT 10.190 92.060 11.790 95.120 ;
        RECT 13.520 92.060 15.120 95.120 ;
        RECT 10.190 92.050 15.120 92.060 ;
        RECT 17.860 92.050 19.460 95.130 ;
        RECT 22.200 95.120 23.930 95.130 ;
        RECT 26.990 95.130 37.530 95.250 ;
        RECT 26.990 95.120 28.720 95.130 ;
        RECT 22.200 92.060 23.800 95.120 ;
        RECT 27.120 92.060 28.720 95.120 ;
        RECT 22.200 92.050 23.930 92.060 ;
        RECT 0.560 90.450 3.460 92.050 ;
        RECT 5.060 91.930 23.930 92.050 ;
        RECT 26.990 92.050 28.720 92.060 ;
        RECT 31.460 92.050 33.060 95.130 ;
        RECT 35.800 95.120 37.530 95.130 ;
        RECT 40.590 95.130 51.130 95.250 ;
        RECT 40.590 95.120 42.320 95.130 ;
        RECT 35.800 92.060 37.400 95.120 ;
        RECT 40.720 92.060 42.320 95.120 ;
        RECT 35.800 92.050 37.530 92.060 ;
        RECT 26.990 91.930 37.530 92.050 ;
        RECT 40.590 92.050 42.320 92.060 ;
        RECT 45.060 92.050 46.660 95.130 ;
        RECT 49.400 95.120 51.130 95.130 ;
        RECT 54.190 95.130 67.930 95.250 ;
        RECT 54.190 95.120 55.920 95.130 ;
        RECT 49.400 92.060 51.000 95.120 ;
        RECT 54.320 92.060 55.920 95.120 ;
        RECT 49.400 92.050 51.130 92.060 ;
        RECT 40.590 91.930 51.130 92.050 ;
        RECT 54.190 92.050 55.920 92.060 ;
        RECT 58.660 92.050 60.260 95.130 ;
        RECT 63.000 95.120 67.930 95.130 ;
        RECT 63.000 92.060 64.600 95.120 ;
        RECT 66.330 92.060 67.930 95.120 ;
        RECT 63.000 92.050 67.930 92.060 ;
        RECT 54.190 91.930 67.930 92.050 ;
        RECT 5.060 91.615 67.930 91.930 ;
        RECT 69.530 96.720 71.130 98.535 ;
        RECT 72.740 96.850 83.260 99.590 ;
        RECT 86.340 96.850 96.860 99.590 ;
        RECT 72.740 96.720 96.860 96.850 ;
        RECT 98.470 96.720 100.070 99.590 ;
        RECT 69.530 95.250 100.070 96.720 ;
        RECT 69.530 95.130 83.270 95.250 ;
        RECT 69.530 95.120 74.460 95.130 ;
        RECT 69.530 92.060 71.130 95.120 ;
        RECT 72.860 92.060 74.460 95.120 ;
        RECT 69.530 92.050 74.460 92.060 ;
        RECT 77.200 92.050 78.800 95.130 ;
        RECT 81.540 95.120 83.270 95.130 ;
        RECT 86.330 95.130 100.070 95.250 ;
        RECT 86.330 95.120 88.060 95.130 ;
        RECT 81.540 92.060 83.140 95.120 ;
        RECT 86.460 92.060 88.060 95.120 ;
        RECT 81.540 92.050 83.270 92.060 ;
        RECT 69.530 91.930 83.270 92.050 ;
        RECT 86.330 92.050 88.060 92.060 ;
        RECT 90.800 92.050 92.400 95.130 ;
        RECT 95.140 95.120 100.070 95.130 ;
        RECT 95.140 92.060 96.740 95.120 ;
        RECT 98.470 92.060 100.070 95.120 ;
        RECT 95.140 92.050 100.070 92.060 ;
        RECT 86.330 91.930 100.070 92.050 ;
        RECT 69.530 91.615 100.070 91.930 ;
        RECT 5.060 90.460 100.070 91.615 ;
        RECT 5.060 90.450 11.790 90.460 ;
        RECT 1.860 88.850 6.660 90.450 ;
        RECT 0.560 87.250 3.460 88.850 ;
        RECT 5.060 87.250 7.960 88.850 ;
        RECT 10.190 87.590 11.790 90.450 ;
        RECT 13.400 90.330 64.720 90.460 ;
        RECT 13.400 87.590 23.920 90.330 ;
        RECT 27.000 87.590 37.520 90.330 ;
        RECT 40.600 87.590 51.120 90.330 ;
        RECT 54.200 87.590 64.720 90.330 ;
        RECT 66.330 90.015 71.130 90.460 ;
        RECT 66.330 87.590 67.930 90.015 ;
        RECT 1.860 85.650 6.660 87.250 ;
        RECT 10.190 87.205 67.930 87.590 ;
        RECT 69.530 87.590 71.130 90.015 ;
        RECT 72.740 90.330 96.860 90.460 ;
        RECT 72.740 87.590 83.260 90.330 ;
        RECT 86.340 87.590 96.860 90.330 ;
        RECT 98.470 87.590 100.070 90.460 ;
        RECT 69.530 87.205 100.070 87.590 ;
        RECT 10.190 85.990 100.070 87.205 ;
        RECT 10.190 85.650 11.790 85.990 ;
        RECT 0.560 84.050 3.460 85.650 ;
        RECT 5.060 84.050 11.790 85.650 ;
        RECT 1.860 82.450 6.660 84.050 ;
        RECT 10.190 83.120 11.790 84.050 ;
        RECT 13.400 83.250 23.920 85.990 ;
        RECT 27.000 83.250 37.520 85.990 ;
        RECT 40.600 83.250 51.120 85.990 ;
        RECT 54.200 83.250 64.720 85.990 ;
        RECT 13.400 83.120 64.720 83.250 ;
        RECT 66.330 85.605 71.130 85.990 ;
        RECT 66.330 83.120 67.930 85.605 ;
        RECT 10.190 82.720 67.930 83.120 ;
        RECT 69.530 83.120 71.130 85.605 ;
        RECT 72.740 83.250 83.260 85.990 ;
        RECT 86.340 83.250 96.860 85.990 ;
        RECT 72.740 83.120 96.860 83.250 ;
        RECT 98.470 83.120 100.070 85.990 ;
        RECT 69.530 82.720 100.070 83.120 ;
        RECT 0.560 80.850 3.460 82.450 ;
        RECT 5.060 80.850 7.960 82.450 ;
        RECT 10.190 81.650 100.070 82.720 ;
        RECT 10.190 81.530 23.930 81.650 ;
        RECT 10.190 81.520 15.120 81.530 ;
        RECT 1.860 79.250 6.660 80.850 ;
        RECT 10.190 79.250 11.790 81.520 ;
        RECT 0.560 77.650 3.460 79.250 ;
        RECT 5.060 78.460 11.790 79.250 ;
        RECT 13.520 78.460 15.120 81.520 ;
        RECT 5.060 78.450 15.120 78.460 ;
        RECT 17.860 78.450 19.460 81.530 ;
        RECT 22.200 81.520 23.930 81.530 ;
        RECT 26.990 81.530 37.530 81.650 ;
        RECT 26.990 81.520 28.720 81.530 ;
        RECT 22.200 78.460 23.800 81.520 ;
        RECT 27.120 78.460 28.720 81.520 ;
        RECT 22.200 78.450 23.930 78.460 ;
        RECT 5.060 78.330 23.930 78.450 ;
        RECT 26.990 78.450 28.720 78.460 ;
        RECT 31.460 78.450 33.060 81.530 ;
        RECT 35.800 81.520 37.530 81.530 ;
        RECT 40.590 81.530 51.130 81.650 ;
        RECT 40.590 81.520 42.320 81.530 ;
        RECT 35.800 78.460 37.400 81.520 ;
        RECT 40.720 78.460 42.320 81.520 ;
        RECT 35.800 78.450 37.530 78.460 ;
        RECT 26.990 78.330 37.530 78.450 ;
        RECT 40.590 78.450 42.320 78.460 ;
        RECT 45.060 78.450 46.660 81.530 ;
        RECT 49.400 81.520 51.130 81.530 ;
        RECT 54.190 81.530 83.270 81.650 ;
        RECT 54.190 81.520 55.920 81.530 ;
        RECT 49.400 78.460 51.000 81.520 ;
        RECT 54.320 78.460 55.920 81.520 ;
        RECT 49.400 78.450 51.130 78.460 ;
        RECT 40.590 78.330 51.130 78.450 ;
        RECT 54.190 78.450 55.920 78.460 ;
        RECT 58.660 78.450 60.260 81.530 ;
        RECT 63.000 81.520 74.460 81.530 ;
        RECT 63.000 78.460 64.600 81.520 ;
        RECT 66.330 81.120 71.130 81.520 ;
        RECT 66.330 78.460 67.930 81.120 ;
        RECT 63.000 78.450 67.930 78.460 ;
        RECT 54.190 78.330 67.930 78.450 ;
        RECT 5.060 77.650 67.930 78.330 ;
        RECT 1.860 76.050 6.660 77.650 ;
        RECT 10.190 76.860 67.930 77.650 ;
        RECT 0.560 74.450 3.460 76.050 ;
        RECT 5.060 74.450 7.960 76.050 ;
        RECT 1.860 72.850 6.660 74.450 ;
        RECT 10.190 73.990 11.790 76.860 ;
        RECT 13.400 76.730 64.720 76.860 ;
        RECT 13.400 73.990 23.920 76.730 ;
        RECT 27.000 73.990 37.520 76.730 ;
        RECT 40.600 73.990 51.120 76.730 ;
        RECT 54.200 73.990 64.720 76.730 ;
        RECT 66.330 74.255 67.930 76.860 ;
        RECT 69.530 78.460 71.130 81.120 ;
        RECT 72.860 78.460 74.460 81.520 ;
        RECT 69.530 78.450 74.460 78.460 ;
        RECT 77.200 78.450 78.800 81.530 ;
        RECT 81.540 81.520 83.270 81.530 ;
        RECT 86.330 81.530 100.070 81.650 ;
        RECT 86.330 81.520 88.060 81.530 ;
        RECT 81.540 78.460 83.140 81.520 ;
        RECT 86.460 78.460 88.060 81.520 ;
        RECT 81.540 78.450 83.270 78.460 ;
        RECT 69.530 78.330 83.270 78.450 ;
        RECT 86.330 78.450 88.060 78.460 ;
        RECT 90.800 78.450 92.400 81.530 ;
        RECT 95.140 81.520 100.070 81.530 ;
        RECT 95.140 78.460 96.740 81.520 ;
        RECT 98.470 78.460 100.070 81.520 ;
        RECT 95.140 78.450 100.070 78.460 ;
        RECT 86.330 78.330 100.070 78.450 ;
        RECT 69.530 76.860 100.070 78.330 ;
        RECT 69.530 74.255 71.130 76.860 ;
        RECT 66.330 73.990 71.130 74.255 ;
        RECT 72.740 76.730 96.860 76.860 ;
        RECT 72.740 73.990 83.260 76.730 ;
        RECT 86.340 73.990 96.860 76.730 ;
        RECT 98.470 73.990 100.070 76.860 ;
        RECT 10.190 72.850 100.070 73.990 ;
        RECT 0.560 71.250 3.460 72.850 ;
        RECT 5.060 72.655 100.070 72.850 ;
        RECT 5.060 72.390 67.930 72.655 ;
        RECT 5.060 71.250 11.790 72.390 ;
        RECT 1.860 69.650 6.660 71.250 ;
        RECT 0.560 68.050 3.460 69.650 ;
        RECT 5.060 68.050 7.960 69.650 ;
        RECT 10.190 69.520 11.790 71.250 ;
        RECT 13.400 69.650 23.920 72.390 ;
        RECT 27.000 69.650 37.520 72.390 ;
        RECT 40.600 69.650 51.120 72.390 ;
        RECT 54.200 69.650 64.720 72.390 ;
        RECT 13.400 69.520 64.720 69.650 ;
        RECT 66.330 69.765 67.930 72.390 ;
        RECT 69.530 72.390 100.070 72.655 ;
        RECT 69.530 69.765 71.130 72.390 ;
        RECT 66.330 69.520 71.130 69.765 ;
        RECT 72.740 69.650 83.260 72.390 ;
        RECT 86.340 69.650 96.860 72.390 ;
        RECT 72.740 69.520 96.860 69.650 ;
        RECT 98.470 69.520 100.070 72.390 ;
        RECT 10.190 68.165 100.070 69.520 ;
        RECT 10.190 68.050 67.930 68.165 ;
        RECT 1.860 66.450 6.660 68.050 ;
        RECT 10.190 67.930 23.930 68.050 ;
        RECT 10.190 67.920 15.120 67.930 ;
        RECT 10.190 66.450 11.790 67.920 ;
        RECT 0.560 64.850 3.460 66.450 ;
        RECT 5.060 64.860 11.790 66.450 ;
        RECT 13.520 64.860 15.120 67.920 ;
        RECT 5.060 64.850 15.120 64.860 ;
        RECT 17.860 64.850 19.460 67.930 ;
        RECT 22.200 67.920 23.930 67.930 ;
        RECT 26.990 67.930 37.530 68.050 ;
        RECT 26.990 67.920 28.720 67.930 ;
        RECT 22.200 64.860 23.800 67.920 ;
        RECT 27.120 64.860 28.720 67.920 ;
        RECT 22.200 64.850 23.930 64.860 ;
        RECT 1.860 63.250 6.660 64.850 ;
        RECT 10.190 64.730 23.930 64.850 ;
        RECT 26.990 64.850 28.720 64.860 ;
        RECT 31.460 64.850 33.060 67.930 ;
        RECT 35.800 67.920 37.530 67.930 ;
        RECT 40.590 67.930 51.130 68.050 ;
        RECT 40.590 67.920 42.320 67.930 ;
        RECT 35.800 64.860 37.400 67.920 ;
        RECT 40.720 64.860 42.320 67.920 ;
        RECT 35.800 64.850 37.530 64.860 ;
        RECT 26.990 64.730 37.530 64.850 ;
        RECT 40.590 64.850 42.320 64.860 ;
        RECT 45.060 64.850 46.660 67.930 ;
        RECT 49.400 67.920 51.130 67.930 ;
        RECT 54.190 67.930 67.930 68.050 ;
        RECT 54.190 67.920 55.920 67.930 ;
        RECT 49.400 64.860 51.000 67.920 ;
        RECT 54.320 64.860 55.920 67.920 ;
        RECT 49.400 64.850 51.130 64.860 ;
        RECT 40.590 64.730 51.130 64.850 ;
        RECT 54.190 64.850 55.920 64.860 ;
        RECT 58.660 64.850 60.260 67.930 ;
        RECT 63.000 67.920 67.930 67.930 ;
        RECT 63.000 64.860 64.600 67.920 ;
        RECT 66.330 65.300 67.930 67.920 ;
        RECT 69.530 68.050 100.070 68.165 ;
        RECT 69.530 67.930 83.270 68.050 ;
        RECT 69.530 67.920 74.460 67.930 ;
        RECT 69.530 65.300 71.130 67.920 ;
        RECT 66.330 64.860 71.130 65.300 ;
        RECT 72.860 64.860 74.460 67.920 ;
        RECT 63.000 64.850 74.460 64.860 ;
        RECT 77.200 64.850 78.800 67.930 ;
        RECT 81.540 67.920 83.270 67.930 ;
        RECT 86.330 67.930 100.070 68.050 ;
        RECT 86.330 67.920 88.060 67.930 ;
        RECT 81.540 64.860 83.140 67.920 ;
        RECT 86.460 64.860 88.060 67.920 ;
        RECT 81.540 64.850 83.270 64.860 ;
        RECT 54.190 64.730 83.270 64.850 ;
        RECT 86.330 64.850 88.060 64.860 ;
        RECT 90.800 64.850 92.400 67.930 ;
        RECT 95.140 67.920 100.070 67.930 ;
        RECT 95.140 64.860 96.740 67.920 ;
        RECT 98.470 64.860 100.070 67.920 ;
        RECT 95.140 64.850 100.070 64.860 ;
        RECT 86.330 64.730 100.070 64.850 ;
        RECT 10.190 63.700 100.070 64.730 ;
        RECT 10.190 63.260 67.930 63.700 ;
        RECT 0.560 61.650 3.460 63.250 ;
        RECT 5.060 61.650 7.960 63.250 ;
        RECT 1.860 60.050 6.660 61.650 ;
        RECT 10.190 60.390 11.790 63.260 ;
        RECT 13.400 63.130 64.720 63.260 ;
        RECT 13.400 60.390 23.920 63.130 ;
        RECT 27.000 60.390 37.520 63.130 ;
        RECT 40.600 60.390 51.120 63.130 ;
        RECT 54.200 60.390 64.720 63.130 ;
        RECT 66.330 60.390 67.930 63.260 ;
        RECT 10.190 60.050 67.930 60.390 ;
        RECT 0.560 58.450 3.460 60.050 ;
        RECT 5.060 58.790 67.930 60.050 ;
        RECT 5.060 58.450 11.790 58.790 ;
        RECT 1.860 56.850 6.660 58.450 ;
        RECT 0.560 55.250 3.460 56.850 ;
        RECT 5.060 55.250 7.960 56.850 ;
        RECT 10.190 55.920 11.790 58.450 ;
        RECT 13.400 56.050 23.920 58.790 ;
        RECT 27.000 56.050 37.520 58.790 ;
        RECT 40.600 56.050 51.120 58.790 ;
        RECT 54.200 56.050 64.720 58.790 ;
        RECT 13.400 55.920 64.720 56.050 ;
        RECT 66.330 56.820 67.930 58.790 ;
        RECT 69.530 63.260 100.070 63.700 ;
        RECT 69.530 60.390 71.130 63.260 ;
        RECT 72.740 63.130 96.860 63.260 ;
        RECT 72.740 60.390 83.260 63.130 ;
        RECT 86.340 60.390 96.860 63.130 ;
        RECT 98.470 60.390 100.070 63.260 ;
        RECT 69.530 58.790 100.070 60.390 ;
        RECT 69.530 56.820 71.130 58.790 ;
        RECT 66.330 55.920 71.130 56.820 ;
        RECT 72.740 56.050 83.260 58.790 ;
        RECT 86.340 56.050 96.860 58.790 ;
        RECT 72.740 55.920 96.860 56.050 ;
        RECT 98.470 55.920 100.070 58.790 ;
        RECT 1.860 53.650 6.660 55.250 ;
        RECT 10.190 55.220 100.070 55.920 ;
        RECT 10.190 54.450 67.930 55.220 ;
        RECT 10.190 54.330 23.930 54.450 ;
        RECT 10.190 54.320 15.120 54.330 ;
        RECT 10.190 53.650 11.790 54.320 ;
        RECT 0.560 52.050 3.460 53.650 ;
        RECT 5.060 52.050 11.790 53.650 ;
        RECT 1.860 50.450 6.660 52.050 ;
        RECT 10.190 51.260 11.790 52.050 ;
        RECT 13.520 51.260 15.120 54.320 ;
        RECT 10.190 51.250 15.120 51.260 ;
        RECT 17.860 51.250 19.460 54.330 ;
        RECT 22.200 54.320 23.930 54.330 ;
        RECT 26.990 54.330 37.530 54.450 ;
        RECT 26.990 54.320 28.720 54.330 ;
        RECT 22.200 51.260 23.800 54.320 ;
        RECT 27.120 51.260 28.720 54.320 ;
        RECT 22.200 51.250 23.930 51.260 ;
        RECT 10.190 51.130 23.930 51.250 ;
        RECT 26.990 51.250 28.720 51.260 ;
        RECT 31.460 51.250 33.060 54.330 ;
        RECT 35.800 54.320 37.530 54.330 ;
        RECT 40.590 54.330 51.130 54.450 ;
        RECT 40.590 54.320 42.320 54.330 ;
        RECT 35.800 51.260 37.400 54.320 ;
        RECT 40.720 51.260 42.320 54.320 ;
        RECT 35.800 51.250 37.530 51.260 ;
        RECT 26.990 51.130 37.530 51.250 ;
        RECT 40.590 51.250 42.320 51.260 ;
        RECT 45.060 51.250 46.660 54.330 ;
        RECT 49.400 54.320 51.130 54.330 ;
        RECT 54.190 54.330 67.930 54.450 ;
        RECT 54.190 54.320 55.920 54.330 ;
        RECT 49.400 51.260 51.000 54.320 ;
        RECT 54.320 51.260 55.920 54.320 ;
        RECT 49.400 51.250 51.130 51.260 ;
        RECT 40.590 51.130 51.130 51.250 ;
        RECT 54.190 51.250 55.920 51.260 ;
        RECT 58.660 51.250 60.260 54.330 ;
        RECT 63.000 54.320 67.930 54.330 ;
        RECT 63.000 51.260 64.600 54.320 ;
        RECT 66.330 52.355 67.930 54.320 ;
        RECT 69.530 54.450 100.070 55.220 ;
        RECT 69.530 54.330 83.270 54.450 ;
        RECT 69.530 54.320 74.460 54.330 ;
        RECT 69.530 52.355 71.130 54.320 ;
        RECT 66.330 51.260 71.130 52.355 ;
        RECT 72.860 51.260 74.460 54.320 ;
        RECT 63.000 51.250 74.460 51.260 ;
        RECT 77.200 51.250 78.800 54.330 ;
        RECT 81.540 54.320 83.270 54.330 ;
        RECT 86.330 54.330 100.070 54.450 ;
        RECT 86.330 54.320 88.060 54.330 ;
        RECT 81.540 51.260 83.140 54.320 ;
        RECT 86.460 51.260 88.060 54.320 ;
        RECT 81.540 51.250 83.270 51.260 ;
        RECT 54.190 51.130 83.270 51.250 ;
        RECT 86.330 51.250 88.060 51.260 ;
        RECT 90.800 51.250 92.400 54.330 ;
        RECT 95.140 54.320 100.070 54.330 ;
        RECT 95.140 51.260 96.740 54.320 ;
        RECT 98.470 51.260 100.070 54.320 ;
        RECT 95.140 51.250 100.070 51.260 ;
        RECT 86.330 51.130 100.070 51.250 ;
        RECT 10.190 50.755 100.070 51.130 ;
        RECT 0.560 48.850 3.460 50.450 ;
        RECT 5.060 48.850 7.960 50.450 ;
        RECT 10.190 49.660 67.930 50.755 ;
        RECT 1.860 47.250 6.660 48.850 ;
        RECT 10.190 47.250 11.790 49.660 ;
        RECT 0.560 45.650 3.460 47.250 ;
        RECT 5.060 46.790 11.790 47.250 ;
        RECT 13.400 49.530 64.720 49.660 ;
        RECT 13.400 46.790 23.920 49.530 ;
        RECT 27.000 46.790 37.520 49.530 ;
        RECT 40.600 46.790 51.120 49.530 ;
        RECT 54.200 46.790 64.720 49.530 ;
        RECT 66.330 47.880 67.930 49.660 ;
        RECT 69.530 49.660 100.070 50.755 ;
        RECT 69.530 47.880 71.130 49.660 ;
        RECT 66.330 46.790 71.130 47.880 ;
        RECT 72.740 49.530 96.860 49.660 ;
        RECT 72.740 46.790 83.260 49.530 ;
        RECT 86.340 46.790 96.860 49.530 ;
        RECT 98.470 46.790 100.070 49.660 ;
        RECT 5.060 46.280 100.070 46.790 ;
        RECT 5.060 45.650 67.930 46.280 ;
        RECT 1.860 44.050 6.660 45.650 ;
        RECT 10.190 45.190 67.930 45.650 ;
        RECT 0.560 42.450 3.460 44.050 ;
        RECT 5.060 42.450 7.960 44.050 ;
        RECT 1.860 40.850 6.660 42.450 ;
        RECT 10.190 42.320 11.790 45.190 ;
        RECT 13.400 42.450 23.920 45.190 ;
        RECT 27.000 42.450 37.520 45.190 ;
        RECT 40.600 42.450 51.120 45.190 ;
        RECT 54.200 42.450 64.720 45.190 ;
        RECT 13.400 42.320 64.720 42.450 ;
        RECT 66.330 42.320 67.930 45.190 ;
        RECT 10.190 40.850 67.930 42.320 ;
        RECT 0.560 39.250 3.460 40.850 ;
        RECT 5.060 40.730 23.930 40.850 ;
        RECT 5.060 40.720 15.120 40.730 ;
        RECT 5.060 39.250 11.790 40.720 ;
        RECT 1.860 37.650 6.660 39.250 ;
        RECT 10.190 37.660 11.790 39.250 ;
        RECT 13.520 37.660 15.120 40.720 ;
        RECT 10.190 37.650 15.120 37.660 ;
        RECT 17.860 37.650 19.460 40.730 ;
        RECT 22.200 40.720 23.930 40.730 ;
        RECT 26.990 40.730 37.530 40.850 ;
        RECT 26.990 40.720 28.720 40.730 ;
        RECT 22.200 37.660 23.800 40.720 ;
        RECT 27.120 37.660 28.720 40.720 ;
        RECT 22.200 37.650 23.930 37.660 ;
        RECT 0.560 36.050 3.460 37.650 ;
        RECT 5.060 36.050 7.960 37.650 ;
        RECT 10.190 37.530 23.930 37.650 ;
        RECT 26.990 37.650 28.720 37.660 ;
        RECT 31.460 37.650 33.060 40.730 ;
        RECT 35.800 40.720 37.530 40.730 ;
        RECT 40.590 40.730 51.130 40.850 ;
        RECT 40.590 40.720 42.320 40.730 ;
        RECT 35.800 37.660 37.400 40.720 ;
        RECT 40.720 37.660 42.320 40.720 ;
        RECT 35.800 37.650 37.530 37.660 ;
        RECT 26.990 37.530 37.530 37.650 ;
        RECT 40.590 37.650 42.320 37.660 ;
        RECT 45.060 37.650 46.660 40.730 ;
        RECT 49.400 40.720 51.130 40.730 ;
        RECT 54.190 40.730 67.930 40.850 ;
        RECT 54.190 40.720 55.920 40.730 ;
        RECT 49.400 37.660 51.000 40.720 ;
        RECT 54.320 37.660 55.920 40.720 ;
        RECT 49.400 37.650 51.130 37.660 ;
        RECT 40.590 37.530 51.130 37.650 ;
        RECT 54.190 37.650 55.920 37.660 ;
        RECT 58.660 37.650 60.260 40.730 ;
        RECT 63.000 40.720 67.930 40.730 ;
        RECT 63.000 37.660 64.600 40.720 ;
        RECT 66.330 39.390 67.930 40.720 ;
        RECT 69.530 45.190 100.070 46.280 ;
        RECT 69.530 42.320 71.130 45.190 ;
        RECT 72.740 42.450 83.260 45.190 ;
        RECT 86.340 42.450 96.860 45.190 ;
        RECT 72.740 42.320 96.860 42.450 ;
        RECT 98.470 42.320 100.070 45.190 ;
        RECT 69.530 40.850 100.070 42.320 ;
        RECT 69.530 40.730 83.270 40.850 ;
        RECT 69.530 40.720 74.460 40.730 ;
        RECT 69.530 39.390 71.130 40.720 ;
        RECT 66.330 37.790 71.130 39.390 ;
        RECT 66.330 37.660 67.930 37.790 ;
        RECT 63.000 37.650 67.930 37.660 ;
        RECT 54.190 37.530 67.930 37.650 ;
        RECT 10.190 36.060 67.930 37.530 ;
        RECT 1.860 34.450 6.660 36.050 ;
        RECT 10.190 34.450 11.790 36.060 ;
        RECT 0.560 32.850 3.460 34.450 ;
        RECT 5.060 33.190 11.790 34.450 ;
        RECT 13.400 35.930 64.720 36.060 ;
        RECT 13.400 33.190 23.920 35.930 ;
        RECT 27.000 33.190 37.520 35.930 ;
        RECT 40.600 33.190 51.120 35.930 ;
        RECT 54.200 33.190 64.720 35.930 ;
        RECT 66.330 34.925 67.930 36.060 ;
        RECT 69.530 37.660 71.130 37.790 ;
        RECT 72.860 37.660 74.460 40.720 ;
        RECT 69.530 37.650 74.460 37.660 ;
        RECT 77.200 37.650 78.800 40.730 ;
        RECT 81.540 40.720 83.270 40.730 ;
        RECT 86.330 40.730 100.070 40.850 ;
        RECT 86.330 40.720 88.060 40.730 ;
        RECT 81.540 37.660 83.140 40.720 ;
        RECT 86.460 37.660 88.060 40.720 ;
        RECT 81.540 37.650 83.270 37.660 ;
        RECT 69.530 37.530 83.270 37.650 ;
        RECT 86.330 37.650 88.060 37.660 ;
        RECT 90.800 37.650 92.400 40.730 ;
        RECT 95.140 40.720 100.070 40.730 ;
        RECT 95.140 37.660 96.740 40.720 ;
        RECT 98.470 37.660 100.070 40.720 ;
        RECT 95.140 37.650 100.070 37.660 ;
        RECT 86.330 37.530 100.070 37.650 ;
        RECT 69.530 36.060 100.070 37.530 ;
        RECT 69.530 34.925 71.130 36.060 ;
        RECT 66.330 33.325 71.130 34.925 ;
        RECT 66.330 33.190 67.930 33.325 ;
        RECT 5.060 32.850 67.930 33.190 ;
        RECT 1.860 31.250 6.660 32.850 ;
        RECT 10.190 31.590 67.930 32.850 ;
        RECT 0.560 29.650 3.460 31.250 ;
        RECT 5.060 29.650 7.960 31.250 ;
        RECT 1.860 28.050 6.660 29.650 ;
        RECT 10.190 28.720 11.790 31.590 ;
        RECT 13.400 28.850 23.920 31.590 ;
        RECT 27.000 28.850 37.520 31.590 ;
        RECT 40.600 28.850 51.120 31.590 ;
        RECT 54.200 28.850 64.720 31.590 ;
        RECT 13.400 28.720 64.720 28.850 ;
        RECT 66.330 30.465 67.930 31.590 ;
        RECT 69.530 33.190 71.130 33.325 ;
        RECT 72.740 35.930 96.860 36.060 ;
        RECT 72.740 33.190 83.260 35.930 ;
        RECT 86.340 33.190 96.860 35.930 ;
        RECT 98.470 33.190 100.070 36.060 ;
        RECT 69.530 31.590 100.070 33.190 ;
        RECT 69.530 30.465 71.130 31.590 ;
        RECT 66.330 28.865 71.130 30.465 ;
        RECT 66.330 28.720 67.930 28.865 ;
        RECT 10.190 28.050 67.930 28.720 ;
        RECT 0.560 26.450 3.460 28.050 ;
        RECT 5.060 27.250 67.930 28.050 ;
        RECT 5.060 27.130 23.930 27.250 ;
        RECT 5.060 27.120 15.120 27.130 ;
        RECT 5.060 26.450 11.790 27.120 ;
        RECT 1.860 24.850 6.660 26.450 ;
        RECT 0.560 23.250 3.460 24.850 ;
        RECT 5.060 23.250 7.960 24.850 ;
        RECT 10.190 24.060 11.790 26.450 ;
        RECT 13.520 24.060 15.120 27.120 ;
        RECT 10.190 24.050 15.120 24.060 ;
        RECT 17.860 24.050 19.460 27.130 ;
        RECT 22.200 27.120 23.930 27.130 ;
        RECT 26.990 27.130 37.530 27.250 ;
        RECT 26.990 27.120 28.720 27.130 ;
        RECT 22.200 24.060 23.800 27.120 ;
        RECT 27.120 24.060 28.720 27.120 ;
        RECT 22.200 24.050 23.930 24.060 ;
        RECT 10.190 23.930 23.930 24.050 ;
        RECT 26.990 24.050 28.720 24.060 ;
        RECT 31.460 24.050 33.060 27.130 ;
        RECT 35.800 27.120 37.530 27.130 ;
        RECT 40.590 27.130 51.130 27.250 ;
        RECT 40.590 27.120 42.320 27.130 ;
        RECT 35.800 24.060 37.400 27.120 ;
        RECT 40.720 24.060 42.320 27.120 ;
        RECT 35.800 24.050 37.530 24.060 ;
        RECT 26.990 23.930 37.530 24.050 ;
        RECT 40.590 24.050 42.320 24.060 ;
        RECT 45.060 24.050 46.660 27.130 ;
        RECT 49.400 27.120 51.130 27.130 ;
        RECT 54.190 27.130 67.930 27.250 ;
        RECT 54.190 27.120 55.920 27.130 ;
        RECT 49.400 24.060 51.000 27.120 ;
        RECT 54.320 24.060 55.920 27.120 ;
        RECT 49.400 24.050 51.130 24.060 ;
        RECT 40.590 23.930 51.130 24.050 ;
        RECT 54.190 24.050 55.920 24.060 ;
        RECT 58.660 24.050 60.260 27.130 ;
        RECT 63.000 27.120 67.930 27.130 ;
        RECT 63.000 24.060 64.600 27.120 ;
        RECT 66.330 24.060 67.930 27.120 ;
        RECT 63.000 24.050 67.930 24.060 ;
        RECT 54.190 23.930 67.930 24.050 ;
        RECT 1.860 21.650 6.660 23.250 ;
        RECT 10.190 22.460 67.930 23.930 ;
        RECT 10.190 21.650 11.790 22.460 ;
        RECT 0.560 20.050 3.460 21.650 ;
        RECT 5.060 20.050 11.790 21.650 ;
        RECT 1.860 18.450 6.660 20.050 ;
        RECT 10.190 19.800 11.790 20.050 ;
        RECT 13.400 22.330 64.720 22.460 ;
        RECT 13.400 19.800 23.920 22.330 ;
        RECT 10.190 19.590 23.920 19.800 ;
        RECT 27.000 19.590 37.520 22.330 ;
        RECT 40.600 19.590 51.120 22.330 ;
        RECT 54.200 19.595 64.720 22.330 ;
        RECT 66.330 21.985 67.930 22.460 ;
        RECT 69.530 28.720 71.130 28.865 ;
        RECT 72.740 28.850 83.260 31.590 ;
        RECT 86.340 28.850 96.860 31.590 ;
        RECT 72.740 28.720 96.860 28.850 ;
        RECT 98.470 28.720 100.070 31.590 ;
        RECT 69.530 27.250 100.070 28.720 ;
        RECT 69.530 27.130 83.270 27.250 ;
        RECT 69.530 27.120 74.460 27.130 ;
        RECT 69.530 24.060 71.130 27.120 ;
        RECT 72.860 24.060 74.460 27.120 ;
        RECT 69.530 24.050 74.460 24.060 ;
        RECT 77.200 24.050 78.800 27.130 ;
        RECT 81.540 27.120 83.270 27.130 ;
        RECT 86.330 27.130 100.070 27.250 ;
        RECT 86.330 27.120 88.060 27.130 ;
        RECT 81.540 24.060 83.140 27.120 ;
        RECT 86.460 24.060 88.060 27.120 ;
        RECT 81.540 24.050 83.270 24.060 ;
        RECT 69.530 23.930 83.270 24.050 ;
        RECT 86.330 24.050 88.060 24.060 ;
        RECT 90.800 24.050 92.400 27.130 ;
        RECT 95.140 27.120 100.070 27.130 ;
        RECT 95.140 24.060 96.740 27.120 ;
        RECT 98.470 24.060 100.070 27.120 ;
        RECT 95.140 24.050 100.070 24.060 ;
        RECT 86.330 23.930 100.070 24.050 ;
        RECT 69.530 22.460 100.070 23.930 ;
        RECT 69.530 21.985 71.130 22.460 ;
        RECT 66.330 20.385 71.130 21.985 ;
        RECT 66.330 19.595 67.930 20.385 ;
        RECT 54.200 19.590 67.930 19.595 ;
        RECT 0.560 16.850 3.460 18.450 ;
        RECT 5.060 16.850 7.960 18.450 ;
        RECT 10.190 18.195 67.930 19.590 ;
        RECT 1.860 15.250 6.660 16.850 ;
        RECT 10.190 15.530 11.790 18.195 ;
        RECT 13.400 17.995 67.930 18.195 ;
        RECT 13.400 17.990 64.720 17.995 ;
        RECT 13.400 15.530 23.920 17.990 ;
        RECT 10.190 15.250 23.920 15.530 ;
        RECT 27.000 15.250 37.520 17.990 ;
        RECT 40.600 15.250 51.120 17.990 ;
        RECT 54.200 15.250 64.720 17.990 ;
        RECT 0.560 13.650 3.460 15.250 ;
        RECT 1.860 6.100 3.460 13.650 ;
        RECT 5.060 15.130 64.720 15.250 ;
        RECT 66.330 17.515 67.930 17.995 ;
        RECT 69.530 19.800 71.130 20.385 ;
        RECT 72.740 22.330 96.860 22.460 ;
        RECT 72.740 19.800 83.260 22.330 ;
        RECT 69.530 19.590 83.260 19.800 ;
        RECT 86.340 19.595 96.860 22.330 ;
        RECT 98.470 19.595 100.070 22.460 ;
        RECT 86.340 19.590 100.070 19.595 ;
        RECT 69.530 18.195 100.070 19.590 ;
        RECT 69.530 17.515 71.130 18.195 ;
        RECT 66.330 15.915 71.130 17.515 ;
        RECT 66.330 15.130 67.930 15.915 ;
        RECT 5.060 13.930 67.930 15.130 ;
        RECT 5.060 13.650 11.790 13.930 ;
        RECT 5.060 6.100 6.660 13.650 ;
        RECT 10.190 11.920 11.790 13.650 ;
        RECT 13.400 13.650 67.930 13.930 ;
        RECT 13.400 13.530 23.930 13.650 ;
        RECT 13.400 11.920 15.000 13.530 ;
        RECT 17.865 11.920 19.465 13.530 ;
        RECT 22.330 11.920 23.930 13.530 ;
        RECT 26.990 13.530 37.530 13.650 ;
        RECT 26.990 11.920 28.590 13.530 ;
        RECT 31.460 11.920 33.060 13.530 ;
        RECT 35.930 11.920 37.530 13.530 ;
        RECT 40.590 13.530 51.130 13.650 ;
        RECT 40.590 11.920 42.190 13.530 ;
        RECT 45.060 11.920 46.660 13.530 ;
        RECT 49.530 11.920 51.130 13.530 ;
        RECT 54.190 13.530 67.930 13.650 ;
        RECT 54.190 11.920 55.790 13.530 ;
        RECT 58.450 11.920 60.055 13.530 ;
        RECT 62.720 11.920 64.320 13.530 ;
        RECT 66.330 13.045 67.930 13.530 ;
        RECT 69.530 15.530 71.130 15.915 ;
        RECT 72.740 17.995 100.070 18.195 ;
        RECT 72.740 17.990 96.860 17.995 ;
        RECT 72.740 15.530 83.260 17.990 ;
        RECT 69.530 15.250 83.260 15.530 ;
        RECT 86.340 15.250 96.860 17.990 ;
        RECT 69.530 15.130 96.860 15.250 ;
        RECT 98.470 15.130 100.070 17.995 ;
        RECT 69.530 13.930 100.070 15.130 ;
        RECT 69.530 13.045 71.130 13.930 ;
        RECT 66.330 11.920 71.130 13.045 ;
        RECT 72.740 13.650 100.070 13.930 ;
        RECT 72.740 13.530 83.270 13.650 ;
        RECT 72.740 11.920 74.340 13.530 ;
        RECT 77.205 11.920 78.805 13.530 ;
        RECT 81.670 11.920 83.270 13.530 ;
        RECT 86.330 13.530 100.070 13.650 ;
        RECT 86.330 11.920 87.930 13.530 ;
        RECT 90.590 11.920 92.195 13.530 ;
        RECT 94.860 11.920 96.460 13.530 ;
        RECT 98.470 11.920 100.070 13.530 ;
        RECT 10.190 11.445 100.070 11.920 ;
        RECT 10.190 10.320 67.930 11.445 ;
        RECT 69.530 10.320 100.070 11.445 ;
        RECT 140.310 121.790 170.850 122.460 ;
        RECT 172.450 121.790 230.190 122.460 ;
        RECT 232.420 122.450 235.320 124.050 ;
        RECT 236.920 122.450 239.820 124.050 ;
        RECT 140.310 120.860 230.190 121.790 ;
        RECT 140.310 118.850 141.910 120.860 ;
        RECT 143.520 119.250 145.120 120.860 ;
        RECT 147.985 119.250 149.585 120.860 ;
        RECT 152.450 119.250 154.050 120.860 ;
        RECT 143.520 119.130 154.050 119.250 ;
        RECT 157.110 119.250 158.710 120.860 ;
        RECT 161.370 119.250 162.975 120.860 ;
        RECT 165.640 119.250 167.240 120.860 ;
        RECT 169.250 120.190 174.050 120.860 ;
        RECT 169.250 119.250 170.850 120.190 ;
        RECT 157.110 119.130 170.850 119.250 ;
        RECT 143.520 118.850 170.850 119.130 ;
        RECT 140.310 117.650 170.850 118.850 ;
        RECT 140.310 117.530 167.640 117.650 ;
        RECT 140.310 117.250 154.040 117.530 ;
        RECT 140.310 114.585 141.910 117.250 ;
        RECT 143.520 114.790 154.040 117.250 ;
        RECT 157.120 114.790 167.640 117.530 ;
        RECT 143.520 114.785 167.640 114.790 ;
        RECT 169.250 114.785 170.850 117.650 ;
        RECT 143.520 114.635 170.850 114.785 ;
        RECT 172.450 118.850 174.050 120.190 ;
        RECT 175.660 119.250 177.260 120.860 ;
        RECT 180.125 119.250 181.725 120.860 ;
        RECT 184.590 119.250 186.190 120.860 ;
        RECT 175.660 119.130 186.190 119.250 ;
        RECT 189.250 119.250 190.850 120.860 ;
        RECT 193.720 119.250 195.320 120.860 ;
        RECT 198.190 119.250 199.790 120.860 ;
        RECT 189.250 119.130 199.790 119.250 ;
        RECT 202.850 119.250 204.450 120.860 ;
        RECT 207.320 119.250 208.920 120.860 ;
        RECT 211.790 119.250 213.390 120.860 ;
        RECT 202.850 119.130 213.390 119.250 ;
        RECT 216.450 119.250 218.050 120.860 ;
        RECT 220.710 119.250 222.315 120.860 ;
        RECT 224.980 119.250 226.580 120.860 ;
        RECT 228.590 119.250 230.190 120.860 ;
        RECT 233.720 120.850 238.520 122.450 ;
        RECT 232.420 119.250 235.320 120.850 ;
        RECT 236.920 119.250 239.820 120.850 ;
        RECT 216.450 119.130 230.190 119.250 ;
        RECT 175.660 118.850 230.190 119.130 ;
        RECT 172.450 117.650 230.190 118.850 ;
        RECT 233.720 117.650 238.520 119.250 ;
        RECT 172.450 117.530 226.980 117.650 ;
        RECT 172.450 117.250 186.180 117.530 ;
        RECT 172.450 114.635 174.050 117.250 ;
        RECT 143.520 114.585 174.050 114.635 ;
        RECT 175.660 114.790 186.180 117.250 ;
        RECT 189.260 114.790 199.780 117.530 ;
        RECT 202.860 114.790 213.380 117.530 ;
        RECT 216.460 114.790 226.980 117.530 ;
        RECT 175.660 114.785 226.980 114.790 ;
        RECT 228.590 116.050 235.320 117.650 ;
        RECT 236.920 116.050 239.820 117.650 ;
        RECT 228.590 114.785 230.190 116.050 ;
        RECT 175.660 114.585 230.190 114.785 ;
        RECT 140.310 113.190 230.190 114.585 ;
        RECT 233.720 114.450 238.520 116.050 ;
        RECT 140.310 112.980 154.040 113.190 ;
        RECT 140.310 110.320 141.910 112.980 ;
        RECT 143.520 110.450 154.040 112.980 ;
        RECT 157.120 113.185 186.180 113.190 ;
        RECT 157.120 110.450 167.640 113.185 ;
        RECT 143.520 110.320 167.640 110.450 ;
        RECT 169.250 113.035 186.180 113.185 ;
        RECT 169.250 110.320 170.850 113.035 ;
        RECT 140.310 109.025 170.850 110.320 ;
        RECT 172.450 112.980 186.180 113.035 ;
        RECT 172.450 110.320 174.050 112.980 ;
        RECT 175.660 110.450 186.180 112.980 ;
        RECT 189.260 110.450 199.780 113.190 ;
        RECT 202.860 110.450 213.380 113.190 ;
        RECT 216.460 113.185 230.190 113.190 ;
        RECT 216.460 110.450 226.980 113.185 ;
        RECT 175.660 110.320 226.980 110.450 ;
        RECT 228.590 111.250 230.190 113.185 ;
        RECT 232.420 112.850 235.320 114.450 ;
        RECT 236.920 112.850 239.820 114.450 ;
        RECT 233.720 111.250 238.520 112.850 ;
        RECT 228.590 110.320 235.320 111.250 ;
        RECT 172.450 109.650 235.320 110.320 ;
        RECT 236.920 109.650 239.820 111.250 ;
        RECT 172.450 109.025 230.190 109.650 ;
        RECT 140.310 108.850 230.190 109.025 ;
        RECT 140.310 108.730 154.050 108.850 ;
        RECT 140.310 108.720 145.240 108.730 ;
        RECT 140.310 105.660 141.910 108.720 ;
        RECT 143.640 105.660 145.240 108.720 ;
        RECT 140.310 105.650 145.240 105.660 ;
        RECT 147.980 105.650 149.580 108.730 ;
        RECT 152.320 108.720 154.050 108.730 ;
        RECT 157.110 108.730 186.190 108.850 ;
        RECT 157.110 108.720 158.840 108.730 ;
        RECT 152.320 105.660 153.920 108.720 ;
        RECT 157.240 105.660 158.840 108.720 ;
        RECT 152.320 105.650 154.050 105.660 ;
        RECT 140.310 105.530 154.050 105.650 ;
        RECT 157.110 105.650 158.840 105.660 ;
        RECT 161.580 105.650 163.180 108.730 ;
        RECT 165.920 108.720 177.380 108.730 ;
        RECT 165.920 105.660 167.520 108.720 ;
        RECT 169.250 107.425 174.050 108.720 ;
        RECT 169.250 105.660 170.850 107.425 ;
        RECT 165.920 105.650 170.850 105.660 ;
        RECT 157.110 105.530 170.850 105.650 ;
        RECT 140.310 104.550 170.850 105.530 ;
        RECT 172.450 105.660 174.050 107.425 ;
        RECT 175.780 105.660 177.380 108.720 ;
        RECT 172.450 105.650 177.380 105.660 ;
        RECT 180.120 105.650 181.720 108.730 ;
        RECT 184.460 108.720 186.190 108.730 ;
        RECT 189.250 108.730 199.790 108.850 ;
        RECT 189.250 108.720 190.980 108.730 ;
        RECT 184.460 105.660 186.060 108.720 ;
        RECT 189.380 105.660 190.980 108.720 ;
        RECT 184.460 105.650 186.190 105.660 ;
        RECT 172.450 105.530 186.190 105.650 ;
        RECT 189.250 105.650 190.980 105.660 ;
        RECT 193.720 105.650 195.320 108.730 ;
        RECT 198.060 108.720 199.790 108.730 ;
        RECT 202.850 108.730 213.390 108.850 ;
        RECT 202.850 108.720 204.580 108.730 ;
        RECT 198.060 105.660 199.660 108.720 ;
        RECT 202.980 105.660 204.580 108.720 ;
        RECT 198.060 105.650 199.790 105.660 ;
        RECT 189.250 105.530 199.790 105.650 ;
        RECT 202.850 105.650 204.580 105.660 ;
        RECT 207.320 105.650 208.920 108.730 ;
        RECT 211.660 108.720 213.390 108.730 ;
        RECT 216.450 108.730 230.190 108.850 ;
        RECT 216.450 108.720 218.180 108.730 ;
        RECT 211.660 105.660 213.260 108.720 ;
        RECT 216.580 105.660 218.180 108.720 ;
        RECT 211.660 105.650 213.390 105.660 ;
        RECT 202.850 105.530 213.390 105.650 ;
        RECT 216.450 105.650 218.180 105.660 ;
        RECT 220.920 105.650 222.520 108.730 ;
        RECT 225.260 108.720 230.190 108.730 ;
        RECT 225.260 105.660 226.860 108.720 ;
        RECT 228.590 105.660 230.190 108.720 ;
        RECT 233.720 108.050 238.520 109.650 ;
        RECT 232.420 106.450 235.320 108.050 ;
        RECT 236.920 106.450 239.820 108.050 ;
        RECT 225.260 105.650 230.190 105.660 ;
        RECT 216.450 105.530 230.190 105.650 ;
        RECT 172.450 104.850 230.190 105.530 ;
        RECT 233.720 104.850 238.520 106.450 ;
        RECT 172.450 104.550 235.320 104.850 ;
        RECT 140.310 104.060 235.320 104.550 ;
        RECT 140.310 101.190 141.910 104.060 ;
        RECT 143.520 103.930 167.640 104.060 ;
        RECT 143.520 101.190 154.040 103.930 ;
        RECT 157.120 101.190 167.640 103.930 ;
        RECT 169.250 102.950 174.050 104.060 ;
        RECT 169.250 101.190 170.850 102.950 ;
        RECT 140.310 100.135 170.850 101.190 ;
        RECT 172.450 101.190 174.050 102.950 ;
        RECT 175.660 103.930 226.980 104.060 ;
        RECT 175.660 101.190 186.180 103.930 ;
        RECT 189.260 101.190 199.780 103.930 ;
        RECT 202.860 101.190 213.380 103.930 ;
        RECT 216.460 101.190 226.980 103.930 ;
        RECT 228.590 103.250 235.320 104.060 ;
        RECT 236.920 103.250 239.820 104.850 ;
        RECT 228.590 101.190 230.190 103.250 ;
        RECT 233.720 101.650 238.520 103.250 ;
        RECT 172.450 100.135 230.190 101.190 ;
        RECT 140.310 99.590 230.190 100.135 ;
        RECT 232.420 100.050 235.320 101.650 ;
        RECT 236.920 100.050 239.820 101.650 ;
        RECT 140.310 96.720 141.910 99.590 ;
        RECT 143.520 96.850 154.040 99.590 ;
        RECT 157.120 96.850 167.640 99.590 ;
        RECT 143.520 96.720 167.640 96.850 ;
        RECT 169.250 98.535 174.050 99.590 ;
        RECT 169.250 96.720 170.850 98.535 ;
        RECT 140.310 95.250 170.850 96.720 ;
        RECT 140.310 95.130 154.050 95.250 ;
        RECT 140.310 95.120 145.240 95.130 ;
        RECT 140.310 92.060 141.910 95.120 ;
        RECT 143.640 92.060 145.240 95.120 ;
        RECT 140.310 92.050 145.240 92.060 ;
        RECT 147.980 92.050 149.580 95.130 ;
        RECT 152.320 95.120 154.050 95.130 ;
        RECT 157.110 95.130 170.850 95.250 ;
        RECT 157.110 95.120 158.840 95.130 ;
        RECT 152.320 92.060 153.920 95.120 ;
        RECT 157.240 92.060 158.840 95.120 ;
        RECT 152.320 92.050 154.050 92.060 ;
        RECT 140.310 91.930 154.050 92.050 ;
        RECT 157.110 92.050 158.840 92.060 ;
        RECT 161.580 92.050 163.180 95.130 ;
        RECT 165.920 95.120 170.850 95.130 ;
        RECT 165.920 92.060 167.520 95.120 ;
        RECT 169.250 92.060 170.850 95.120 ;
        RECT 165.920 92.050 170.850 92.060 ;
        RECT 157.110 91.930 170.850 92.050 ;
        RECT 140.310 91.615 170.850 91.930 ;
        RECT 172.450 96.720 174.050 98.535 ;
        RECT 175.660 96.850 186.180 99.590 ;
        RECT 189.260 96.850 199.780 99.590 ;
        RECT 202.860 96.850 213.380 99.590 ;
        RECT 216.460 96.850 226.980 99.590 ;
        RECT 175.660 96.720 226.980 96.850 ;
        RECT 228.590 98.450 230.190 99.590 ;
        RECT 233.720 98.450 238.520 100.050 ;
        RECT 228.590 96.850 235.320 98.450 ;
        RECT 236.920 96.850 239.820 98.450 ;
        RECT 228.590 96.720 230.190 96.850 ;
        RECT 172.450 95.250 230.190 96.720 ;
        RECT 233.720 95.250 238.520 96.850 ;
        RECT 172.450 95.130 186.190 95.250 ;
        RECT 172.450 95.120 177.380 95.130 ;
        RECT 172.450 92.060 174.050 95.120 ;
        RECT 175.780 92.060 177.380 95.120 ;
        RECT 172.450 92.050 177.380 92.060 ;
        RECT 180.120 92.050 181.720 95.130 ;
        RECT 184.460 95.120 186.190 95.130 ;
        RECT 189.250 95.130 199.790 95.250 ;
        RECT 189.250 95.120 190.980 95.130 ;
        RECT 184.460 92.060 186.060 95.120 ;
        RECT 189.380 92.060 190.980 95.120 ;
        RECT 184.460 92.050 186.190 92.060 ;
        RECT 172.450 91.930 186.190 92.050 ;
        RECT 189.250 92.050 190.980 92.060 ;
        RECT 193.720 92.050 195.320 95.130 ;
        RECT 198.060 95.120 199.790 95.130 ;
        RECT 202.850 95.130 213.390 95.250 ;
        RECT 202.850 95.120 204.580 95.130 ;
        RECT 198.060 92.060 199.660 95.120 ;
        RECT 202.980 92.060 204.580 95.120 ;
        RECT 198.060 92.050 199.790 92.060 ;
        RECT 189.250 91.930 199.790 92.050 ;
        RECT 202.850 92.050 204.580 92.060 ;
        RECT 207.320 92.050 208.920 95.130 ;
        RECT 211.660 95.120 213.390 95.130 ;
        RECT 216.450 95.130 230.190 95.250 ;
        RECT 216.450 95.120 218.180 95.130 ;
        RECT 211.660 92.060 213.260 95.120 ;
        RECT 216.580 92.060 218.180 95.120 ;
        RECT 211.660 92.050 213.390 92.060 ;
        RECT 202.850 91.930 213.390 92.050 ;
        RECT 216.450 92.050 218.180 92.060 ;
        RECT 220.920 92.050 222.520 95.130 ;
        RECT 225.260 95.120 230.190 95.130 ;
        RECT 225.260 92.060 226.860 95.120 ;
        RECT 228.590 92.060 230.190 95.120 ;
        RECT 232.420 93.650 235.320 95.250 ;
        RECT 236.920 93.650 239.820 95.250 ;
        RECT 225.260 92.050 230.190 92.060 ;
        RECT 233.720 92.050 238.520 93.650 ;
        RECT 216.450 91.930 235.320 92.050 ;
        RECT 172.450 91.615 235.320 91.930 ;
        RECT 140.310 90.460 235.320 91.615 ;
        RECT 140.310 87.590 141.910 90.460 ;
        RECT 143.520 90.330 167.640 90.460 ;
        RECT 143.520 87.590 154.040 90.330 ;
        RECT 157.120 87.590 167.640 90.330 ;
        RECT 169.250 90.015 174.050 90.460 ;
        RECT 169.250 87.590 170.850 90.015 ;
        RECT 140.310 87.205 170.850 87.590 ;
        RECT 172.450 87.590 174.050 90.015 ;
        RECT 175.660 90.330 226.980 90.460 ;
        RECT 175.660 87.590 186.180 90.330 ;
        RECT 189.260 87.590 199.780 90.330 ;
        RECT 202.860 87.590 213.380 90.330 ;
        RECT 216.460 87.590 226.980 90.330 ;
        RECT 228.590 90.450 235.320 90.460 ;
        RECT 236.920 90.450 239.820 92.050 ;
        RECT 228.590 87.590 230.190 90.450 ;
        RECT 233.720 88.850 238.520 90.450 ;
        RECT 172.450 87.205 230.190 87.590 ;
        RECT 232.420 87.250 235.320 88.850 ;
        RECT 236.920 87.250 239.820 88.850 ;
        RECT 140.310 85.990 230.190 87.205 ;
        RECT 140.310 83.120 141.910 85.990 ;
        RECT 143.520 83.250 154.040 85.990 ;
        RECT 157.120 83.250 167.640 85.990 ;
        RECT 143.520 83.120 167.640 83.250 ;
        RECT 169.250 85.605 174.050 85.990 ;
        RECT 169.250 83.120 170.850 85.605 ;
        RECT 140.310 82.720 170.850 83.120 ;
        RECT 172.450 83.120 174.050 85.605 ;
        RECT 175.660 83.250 186.180 85.990 ;
        RECT 189.260 83.250 199.780 85.990 ;
        RECT 202.860 83.250 213.380 85.990 ;
        RECT 216.460 83.250 226.980 85.990 ;
        RECT 175.660 83.120 226.980 83.250 ;
        RECT 228.590 85.650 230.190 85.990 ;
        RECT 233.720 85.650 238.520 87.250 ;
        RECT 228.590 84.050 235.320 85.650 ;
        RECT 236.920 84.050 239.820 85.650 ;
        RECT 228.590 83.120 230.190 84.050 ;
        RECT 172.450 82.720 230.190 83.120 ;
        RECT 140.310 81.650 230.190 82.720 ;
        RECT 233.720 82.450 238.520 84.050 ;
        RECT 140.310 81.530 154.050 81.650 ;
        RECT 140.310 81.520 145.240 81.530 ;
        RECT 140.310 78.460 141.910 81.520 ;
        RECT 143.640 78.460 145.240 81.520 ;
        RECT 140.310 78.450 145.240 78.460 ;
        RECT 147.980 78.450 149.580 81.530 ;
        RECT 152.320 81.520 154.050 81.530 ;
        RECT 157.110 81.530 186.190 81.650 ;
        RECT 157.110 81.520 158.840 81.530 ;
        RECT 152.320 78.460 153.920 81.520 ;
        RECT 157.240 78.460 158.840 81.520 ;
        RECT 152.320 78.450 154.050 78.460 ;
        RECT 140.310 78.330 154.050 78.450 ;
        RECT 157.110 78.450 158.840 78.460 ;
        RECT 161.580 78.450 163.180 81.530 ;
        RECT 165.920 81.520 177.380 81.530 ;
        RECT 165.920 78.460 167.520 81.520 ;
        RECT 169.250 81.120 174.050 81.520 ;
        RECT 169.250 78.460 170.850 81.120 ;
        RECT 165.920 78.450 170.850 78.460 ;
        RECT 157.110 78.330 170.850 78.450 ;
        RECT 140.310 76.860 170.850 78.330 ;
        RECT 140.310 73.990 141.910 76.860 ;
        RECT 143.520 76.730 167.640 76.860 ;
        RECT 143.520 73.990 154.040 76.730 ;
        RECT 157.120 73.990 167.640 76.730 ;
        RECT 169.250 74.255 170.850 76.860 ;
        RECT 172.450 78.460 174.050 81.120 ;
        RECT 175.780 78.460 177.380 81.520 ;
        RECT 172.450 78.450 177.380 78.460 ;
        RECT 180.120 78.450 181.720 81.530 ;
        RECT 184.460 81.520 186.190 81.530 ;
        RECT 189.250 81.530 199.790 81.650 ;
        RECT 189.250 81.520 190.980 81.530 ;
        RECT 184.460 78.460 186.060 81.520 ;
        RECT 189.380 78.460 190.980 81.520 ;
        RECT 184.460 78.450 186.190 78.460 ;
        RECT 172.450 78.330 186.190 78.450 ;
        RECT 189.250 78.450 190.980 78.460 ;
        RECT 193.720 78.450 195.320 81.530 ;
        RECT 198.060 81.520 199.790 81.530 ;
        RECT 202.850 81.530 213.390 81.650 ;
        RECT 202.850 81.520 204.580 81.530 ;
        RECT 198.060 78.460 199.660 81.520 ;
        RECT 202.980 78.460 204.580 81.520 ;
        RECT 198.060 78.450 199.790 78.460 ;
        RECT 189.250 78.330 199.790 78.450 ;
        RECT 202.850 78.450 204.580 78.460 ;
        RECT 207.320 78.450 208.920 81.530 ;
        RECT 211.660 81.520 213.390 81.530 ;
        RECT 216.450 81.530 230.190 81.650 ;
        RECT 216.450 81.520 218.180 81.530 ;
        RECT 211.660 78.460 213.260 81.520 ;
        RECT 216.580 78.460 218.180 81.520 ;
        RECT 211.660 78.450 213.390 78.460 ;
        RECT 202.850 78.330 213.390 78.450 ;
        RECT 216.450 78.450 218.180 78.460 ;
        RECT 220.920 78.450 222.520 81.530 ;
        RECT 225.260 81.520 230.190 81.530 ;
        RECT 225.260 78.460 226.860 81.520 ;
        RECT 228.590 79.250 230.190 81.520 ;
        RECT 232.420 80.850 235.320 82.450 ;
        RECT 236.920 80.850 239.820 82.450 ;
        RECT 233.720 79.250 238.520 80.850 ;
        RECT 228.590 78.460 235.320 79.250 ;
        RECT 225.260 78.450 235.320 78.460 ;
        RECT 216.450 78.330 235.320 78.450 ;
        RECT 172.450 77.650 235.320 78.330 ;
        RECT 236.920 77.650 239.820 79.250 ;
        RECT 172.450 76.860 230.190 77.650 ;
        RECT 172.450 74.255 174.050 76.860 ;
        RECT 169.250 73.990 174.050 74.255 ;
        RECT 175.660 76.730 226.980 76.860 ;
        RECT 175.660 73.990 186.180 76.730 ;
        RECT 189.260 73.990 199.780 76.730 ;
        RECT 202.860 73.990 213.380 76.730 ;
        RECT 216.460 73.990 226.980 76.730 ;
        RECT 228.590 73.990 230.190 76.860 ;
        RECT 233.720 76.050 238.520 77.650 ;
        RECT 232.420 74.450 235.320 76.050 ;
        RECT 236.920 74.450 239.820 76.050 ;
        RECT 140.310 72.850 230.190 73.990 ;
        RECT 233.720 72.850 238.520 74.450 ;
        RECT 140.310 72.655 235.320 72.850 ;
        RECT 140.310 72.390 170.850 72.655 ;
        RECT 140.310 69.520 141.910 72.390 ;
        RECT 143.520 69.650 154.040 72.390 ;
        RECT 157.120 69.650 167.640 72.390 ;
        RECT 143.520 69.520 167.640 69.650 ;
        RECT 169.250 69.765 170.850 72.390 ;
        RECT 172.450 72.390 235.320 72.655 ;
        RECT 172.450 69.765 174.050 72.390 ;
        RECT 169.250 69.520 174.050 69.765 ;
        RECT 175.660 69.650 186.180 72.390 ;
        RECT 189.260 69.650 199.780 72.390 ;
        RECT 202.860 69.650 213.380 72.390 ;
        RECT 216.460 69.650 226.980 72.390 ;
        RECT 175.660 69.520 226.980 69.650 ;
        RECT 228.590 71.250 235.320 72.390 ;
        RECT 236.920 71.250 239.820 72.850 ;
        RECT 228.590 69.520 230.190 71.250 ;
        RECT 233.720 69.650 238.520 71.250 ;
        RECT 140.310 68.165 230.190 69.520 ;
        RECT 140.310 68.050 170.850 68.165 ;
        RECT 140.310 67.930 154.050 68.050 ;
        RECT 140.310 67.920 145.240 67.930 ;
        RECT 140.310 64.860 141.910 67.920 ;
        RECT 143.640 64.860 145.240 67.920 ;
        RECT 140.310 64.850 145.240 64.860 ;
        RECT 147.980 64.850 149.580 67.930 ;
        RECT 152.320 67.920 154.050 67.930 ;
        RECT 157.110 67.930 170.850 68.050 ;
        RECT 157.110 67.920 158.840 67.930 ;
        RECT 152.320 64.860 153.920 67.920 ;
        RECT 157.240 64.860 158.840 67.920 ;
        RECT 152.320 64.850 154.050 64.860 ;
        RECT 140.310 64.730 154.050 64.850 ;
        RECT 157.110 64.850 158.840 64.860 ;
        RECT 161.580 64.850 163.180 67.930 ;
        RECT 165.920 67.920 170.850 67.930 ;
        RECT 165.920 64.860 167.520 67.920 ;
        RECT 169.250 65.300 170.850 67.920 ;
        RECT 172.450 68.050 230.190 68.165 ;
        RECT 232.420 68.050 235.320 69.650 ;
        RECT 236.920 68.050 239.820 69.650 ;
        RECT 172.450 67.930 186.190 68.050 ;
        RECT 172.450 67.920 177.380 67.930 ;
        RECT 172.450 65.300 174.050 67.920 ;
        RECT 169.250 64.860 174.050 65.300 ;
        RECT 175.780 64.860 177.380 67.920 ;
        RECT 165.920 64.850 177.380 64.860 ;
        RECT 180.120 64.850 181.720 67.930 ;
        RECT 184.460 67.920 186.190 67.930 ;
        RECT 189.250 67.930 199.790 68.050 ;
        RECT 189.250 67.920 190.980 67.930 ;
        RECT 184.460 64.860 186.060 67.920 ;
        RECT 189.380 64.860 190.980 67.920 ;
        RECT 184.460 64.850 186.190 64.860 ;
        RECT 157.110 64.730 186.190 64.850 ;
        RECT 189.250 64.850 190.980 64.860 ;
        RECT 193.720 64.850 195.320 67.930 ;
        RECT 198.060 67.920 199.790 67.930 ;
        RECT 202.850 67.930 213.390 68.050 ;
        RECT 202.850 67.920 204.580 67.930 ;
        RECT 198.060 64.860 199.660 67.920 ;
        RECT 202.980 64.860 204.580 67.920 ;
        RECT 198.060 64.850 199.790 64.860 ;
        RECT 189.250 64.730 199.790 64.850 ;
        RECT 202.850 64.850 204.580 64.860 ;
        RECT 207.320 64.850 208.920 67.930 ;
        RECT 211.660 67.920 213.390 67.930 ;
        RECT 216.450 67.930 230.190 68.050 ;
        RECT 216.450 67.920 218.180 67.930 ;
        RECT 211.660 64.860 213.260 67.920 ;
        RECT 216.580 64.860 218.180 67.920 ;
        RECT 211.660 64.850 213.390 64.860 ;
        RECT 202.850 64.730 213.390 64.850 ;
        RECT 216.450 64.850 218.180 64.860 ;
        RECT 220.920 64.850 222.520 67.930 ;
        RECT 225.260 67.920 230.190 67.930 ;
        RECT 225.260 64.860 226.860 67.920 ;
        RECT 228.590 66.450 230.190 67.920 ;
        RECT 233.720 66.450 238.520 68.050 ;
        RECT 228.590 64.860 235.320 66.450 ;
        RECT 225.260 64.850 235.320 64.860 ;
        RECT 236.920 64.850 239.820 66.450 ;
        RECT 216.450 64.730 230.190 64.850 ;
        RECT 140.310 63.700 230.190 64.730 ;
        RECT 140.310 63.260 170.850 63.700 ;
        RECT 140.310 60.390 141.910 63.260 ;
        RECT 143.520 63.130 167.640 63.260 ;
        RECT 143.520 60.390 154.040 63.130 ;
        RECT 157.120 60.390 167.640 63.130 ;
        RECT 169.250 60.390 170.850 63.260 ;
        RECT 140.310 58.790 170.850 60.390 ;
        RECT 140.310 55.920 141.910 58.790 ;
        RECT 143.520 56.050 154.040 58.790 ;
        RECT 157.120 56.050 167.640 58.790 ;
        RECT 143.520 55.920 167.640 56.050 ;
        RECT 169.250 56.820 170.850 58.790 ;
        RECT 172.450 63.260 230.190 63.700 ;
        RECT 172.450 60.390 174.050 63.260 ;
        RECT 175.660 63.130 226.980 63.260 ;
        RECT 175.660 60.390 186.180 63.130 ;
        RECT 189.260 60.390 199.780 63.130 ;
        RECT 202.860 60.390 213.380 63.130 ;
        RECT 216.460 60.390 226.980 63.130 ;
        RECT 228.590 60.390 230.190 63.260 ;
        RECT 233.720 63.250 238.520 64.850 ;
        RECT 232.420 61.650 235.320 63.250 ;
        RECT 236.920 61.650 239.820 63.250 ;
        RECT 172.450 60.050 230.190 60.390 ;
        RECT 233.720 60.050 238.520 61.650 ;
        RECT 172.450 58.790 235.320 60.050 ;
        RECT 172.450 56.820 174.050 58.790 ;
        RECT 169.250 55.920 174.050 56.820 ;
        RECT 175.660 56.050 186.180 58.790 ;
        RECT 189.260 56.050 199.780 58.790 ;
        RECT 202.860 56.050 213.380 58.790 ;
        RECT 216.460 56.050 226.980 58.790 ;
        RECT 175.660 55.920 226.980 56.050 ;
        RECT 228.590 58.450 235.320 58.790 ;
        RECT 236.920 58.450 239.820 60.050 ;
        RECT 228.590 55.920 230.190 58.450 ;
        RECT 233.720 56.850 238.520 58.450 ;
        RECT 140.310 55.220 230.190 55.920 ;
        RECT 232.420 55.250 235.320 56.850 ;
        RECT 236.920 55.250 239.820 56.850 ;
        RECT 140.310 54.450 170.850 55.220 ;
        RECT 140.310 54.330 154.050 54.450 ;
        RECT 140.310 54.320 145.240 54.330 ;
        RECT 140.310 51.260 141.910 54.320 ;
        RECT 143.640 51.260 145.240 54.320 ;
        RECT 140.310 51.250 145.240 51.260 ;
        RECT 147.980 51.250 149.580 54.330 ;
        RECT 152.320 54.320 154.050 54.330 ;
        RECT 157.110 54.330 170.850 54.450 ;
        RECT 157.110 54.320 158.840 54.330 ;
        RECT 152.320 51.260 153.920 54.320 ;
        RECT 157.240 51.260 158.840 54.320 ;
        RECT 152.320 51.250 154.050 51.260 ;
        RECT 140.310 51.130 154.050 51.250 ;
        RECT 157.110 51.250 158.840 51.260 ;
        RECT 161.580 51.250 163.180 54.330 ;
        RECT 165.920 54.320 170.850 54.330 ;
        RECT 165.920 51.260 167.520 54.320 ;
        RECT 169.250 52.355 170.850 54.320 ;
        RECT 172.450 54.450 230.190 55.220 ;
        RECT 172.450 54.330 186.190 54.450 ;
        RECT 172.450 54.320 177.380 54.330 ;
        RECT 172.450 52.355 174.050 54.320 ;
        RECT 169.250 51.260 174.050 52.355 ;
        RECT 175.780 51.260 177.380 54.320 ;
        RECT 165.920 51.250 177.380 51.260 ;
        RECT 180.120 51.250 181.720 54.330 ;
        RECT 184.460 54.320 186.190 54.330 ;
        RECT 189.250 54.330 199.790 54.450 ;
        RECT 189.250 54.320 190.980 54.330 ;
        RECT 184.460 51.260 186.060 54.320 ;
        RECT 189.380 51.260 190.980 54.320 ;
        RECT 184.460 51.250 186.190 51.260 ;
        RECT 157.110 51.130 186.190 51.250 ;
        RECT 189.250 51.250 190.980 51.260 ;
        RECT 193.720 51.250 195.320 54.330 ;
        RECT 198.060 54.320 199.790 54.330 ;
        RECT 202.850 54.330 213.390 54.450 ;
        RECT 202.850 54.320 204.580 54.330 ;
        RECT 198.060 51.260 199.660 54.320 ;
        RECT 202.980 51.260 204.580 54.320 ;
        RECT 198.060 51.250 199.790 51.260 ;
        RECT 189.250 51.130 199.790 51.250 ;
        RECT 202.850 51.250 204.580 51.260 ;
        RECT 207.320 51.250 208.920 54.330 ;
        RECT 211.660 54.320 213.390 54.330 ;
        RECT 216.450 54.330 230.190 54.450 ;
        RECT 216.450 54.320 218.180 54.330 ;
        RECT 211.660 51.260 213.260 54.320 ;
        RECT 216.580 51.260 218.180 54.320 ;
        RECT 211.660 51.250 213.390 51.260 ;
        RECT 202.850 51.130 213.390 51.250 ;
        RECT 216.450 51.250 218.180 51.260 ;
        RECT 220.920 51.250 222.520 54.330 ;
        RECT 225.260 54.320 230.190 54.330 ;
        RECT 225.260 51.260 226.860 54.320 ;
        RECT 228.590 53.650 230.190 54.320 ;
        RECT 233.720 53.650 238.520 55.250 ;
        RECT 228.590 52.050 235.320 53.650 ;
        RECT 236.920 52.050 239.820 53.650 ;
        RECT 228.590 51.260 230.190 52.050 ;
        RECT 225.260 51.250 230.190 51.260 ;
        RECT 216.450 51.130 230.190 51.250 ;
        RECT 140.310 50.755 230.190 51.130 ;
        RECT 140.310 49.660 170.850 50.755 ;
        RECT 140.310 46.790 141.910 49.660 ;
        RECT 143.520 49.530 167.640 49.660 ;
        RECT 143.520 46.790 154.040 49.530 ;
        RECT 157.120 46.790 167.640 49.530 ;
        RECT 169.250 47.880 170.850 49.660 ;
        RECT 172.450 49.660 230.190 50.755 ;
        RECT 233.720 50.450 238.520 52.050 ;
        RECT 172.450 47.880 174.050 49.660 ;
        RECT 169.250 46.790 174.050 47.880 ;
        RECT 175.660 49.530 226.980 49.660 ;
        RECT 175.660 46.790 186.180 49.530 ;
        RECT 189.260 46.790 199.780 49.530 ;
        RECT 202.860 46.790 213.380 49.530 ;
        RECT 216.460 46.790 226.980 49.530 ;
        RECT 228.590 47.250 230.190 49.660 ;
        RECT 232.420 48.850 235.320 50.450 ;
        RECT 236.920 48.850 239.820 50.450 ;
        RECT 233.720 47.250 238.520 48.850 ;
        RECT 228.590 46.790 235.320 47.250 ;
        RECT 140.310 46.280 235.320 46.790 ;
        RECT 140.310 45.190 170.850 46.280 ;
        RECT 140.310 42.320 141.910 45.190 ;
        RECT 143.520 42.450 154.040 45.190 ;
        RECT 157.120 42.450 167.640 45.190 ;
        RECT 143.520 42.320 167.640 42.450 ;
        RECT 169.250 42.320 170.850 45.190 ;
        RECT 140.310 40.850 170.850 42.320 ;
        RECT 140.310 40.730 154.050 40.850 ;
        RECT 140.310 40.720 145.240 40.730 ;
        RECT 140.310 37.660 141.910 40.720 ;
        RECT 143.640 37.660 145.240 40.720 ;
        RECT 140.310 37.650 145.240 37.660 ;
        RECT 147.980 37.650 149.580 40.730 ;
        RECT 152.320 40.720 154.050 40.730 ;
        RECT 157.110 40.730 170.850 40.850 ;
        RECT 157.110 40.720 158.840 40.730 ;
        RECT 152.320 37.660 153.920 40.720 ;
        RECT 157.240 37.660 158.840 40.720 ;
        RECT 152.320 37.650 154.050 37.660 ;
        RECT 140.310 37.530 154.050 37.650 ;
        RECT 157.110 37.650 158.840 37.660 ;
        RECT 161.580 37.650 163.180 40.730 ;
        RECT 165.920 40.720 170.850 40.730 ;
        RECT 165.920 37.660 167.520 40.720 ;
        RECT 169.250 39.390 170.850 40.720 ;
        RECT 172.450 45.650 235.320 46.280 ;
        RECT 236.920 45.650 239.820 47.250 ;
        RECT 172.450 45.190 230.190 45.650 ;
        RECT 172.450 42.320 174.050 45.190 ;
        RECT 175.660 42.450 186.180 45.190 ;
        RECT 189.260 42.450 199.780 45.190 ;
        RECT 202.860 42.450 213.380 45.190 ;
        RECT 216.460 42.450 226.980 45.190 ;
        RECT 175.660 42.320 226.980 42.450 ;
        RECT 228.590 42.320 230.190 45.190 ;
        RECT 233.720 44.050 238.520 45.650 ;
        RECT 232.420 42.450 235.320 44.050 ;
        RECT 236.920 42.450 239.820 44.050 ;
        RECT 172.450 40.850 230.190 42.320 ;
        RECT 233.720 40.850 238.520 42.450 ;
        RECT 172.450 40.730 186.190 40.850 ;
        RECT 172.450 40.720 177.380 40.730 ;
        RECT 172.450 39.390 174.050 40.720 ;
        RECT 169.250 37.790 174.050 39.390 ;
        RECT 169.250 37.660 170.850 37.790 ;
        RECT 165.920 37.650 170.850 37.660 ;
        RECT 157.110 37.530 170.850 37.650 ;
        RECT 140.310 36.060 170.850 37.530 ;
        RECT 140.310 33.190 141.910 36.060 ;
        RECT 143.520 35.930 167.640 36.060 ;
        RECT 143.520 33.190 154.040 35.930 ;
        RECT 157.120 33.190 167.640 35.930 ;
        RECT 169.250 34.925 170.850 36.060 ;
        RECT 172.450 37.660 174.050 37.790 ;
        RECT 175.780 37.660 177.380 40.720 ;
        RECT 172.450 37.650 177.380 37.660 ;
        RECT 180.120 37.650 181.720 40.730 ;
        RECT 184.460 40.720 186.190 40.730 ;
        RECT 189.250 40.730 199.790 40.850 ;
        RECT 189.250 40.720 190.980 40.730 ;
        RECT 184.460 37.660 186.060 40.720 ;
        RECT 189.380 37.660 190.980 40.720 ;
        RECT 184.460 37.650 186.190 37.660 ;
        RECT 172.450 37.530 186.190 37.650 ;
        RECT 189.250 37.650 190.980 37.660 ;
        RECT 193.720 37.650 195.320 40.730 ;
        RECT 198.060 40.720 199.790 40.730 ;
        RECT 202.850 40.730 213.390 40.850 ;
        RECT 202.850 40.720 204.580 40.730 ;
        RECT 198.060 37.660 199.660 40.720 ;
        RECT 202.980 37.660 204.580 40.720 ;
        RECT 198.060 37.650 199.790 37.660 ;
        RECT 189.250 37.530 199.790 37.650 ;
        RECT 202.850 37.650 204.580 37.660 ;
        RECT 207.320 37.650 208.920 40.730 ;
        RECT 211.660 40.720 213.390 40.730 ;
        RECT 216.450 40.730 235.320 40.850 ;
        RECT 216.450 40.720 218.180 40.730 ;
        RECT 211.660 37.660 213.260 40.720 ;
        RECT 216.580 37.660 218.180 40.720 ;
        RECT 211.660 37.650 213.390 37.660 ;
        RECT 202.850 37.530 213.390 37.650 ;
        RECT 216.450 37.650 218.180 37.660 ;
        RECT 220.920 37.650 222.520 40.730 ;
        RECT 225.260 40.720 235.320 40.730 ;
        RECT 225.260 37.660 226.860 40.720 ;
        RECT 228.590 39.250 235.320 40.720 ;
        RECT 236.920 39.250 239.820 40.850 ;
        RECT 228.590 37.660 230.190 39.250 ;
        RECT 225.260 37.650 230.190 37.660 ;
        RECT 233.720 37.650 238.520 39.250 ;
        RECT 216.450 37.530 230.190 37.650 ;
        RECT 172.450 36.060 230.190 37.530 ;
        RECT 172.450 34.925 174.050 36.060 ;
        RECT 169.250 33.325 174.050 34.925 ;
        RECT 169.250 33.190 170.850 33.325 ;
        RECT 140.310 31.590 170.850 33.190 ;
        RECT 140.310 28.720 141.910 31.590 ;
        RECT 143.520 28.850 154.040 31.590 ;
        RECT 157.120 28.850 167.640 31.590 ;
        RECT 143.520 28.720 167.640 28.850 ;
        RECT 169.250 30.465 170.850 31.590 ;
        RECT 172.450 33.190 174.050 33.325 ;
        RECT 175.660 35.930 226.980 36.060 ;
        RECT 175.660 33.190 186.180 35.930 ;
        RECT 189.260 33.190 199.780 35.930 ;
        RECT 202.860 33.190 213.380 35.930 ;
        RECT 216.460 33.190 226.980 35.930 ;
        RECT 228.590 34.450 230.190 36.060 ;
        RECT 232.420 36.050 235.320 37.650 ;
        RECT 236.920 36.050 239.820 37.650 ;
        RECT 233.720 34.450 238.520 36.050 ;
        RECT 228.590 33.190 235.320 34.450 ;
        RECT 172.450 32.850 235.320 33.190 ;
        RECT 236.920 32.850 239.820 34.450 ;
        RECT 172.450 31.590 230.190 32.850 ;
        RECT 172.450 30.465 174.050 31.590 ;
        RECT 169.250 28.865 174.050 30.465 ;
        RECT 169.250 28.720 170.850 28.865 ;
        RECT 140.310 27.250 170.850 28.720 ;
        RECT 140.310 27.130 154.050 27.250 ;
        RECT 140.310 27.120 145.240 27.130 ;
        RECT 140.310 24.060 141.910 27.120 ;
        RECT 143.640 24.060 145.240 27.120 ;
        RECT 140.310 24.050 145.240 24.060 ;
        RECT 147.980 24.050 149.580 27.130 ;
        RECT 152.320 27.120 154.050 27.130 ;
        RECT 157.110 27.130 170.850 27.250 ;
        RECT 157.110 27.120 158.840 27.130 ;
        RECT 152.320 24.060 153.920 27.120 ;
        RECT 157.240 24.060 158.840 27.120 ;
        RECT 152.320 24.050 154.050 24.060 ;
        RECT 140.310 23.930 154.050 24.050 ;
        RECT 157.110 24.050 158.840 24.060 ;
        RECT 161.580 24.050 163.180 27.130 ;
        RECT 165.920 27.120 170.850 27.130 ;
        RECT 165.920 24.060 167.520 27.120 ;
        RECT 169.250 24.060 170.850 27.120 ;
        RECT 165.920 24.050 170.850 24.060 ;
        RECT 157.110 23.930 170.850 24.050 ;
        RECT 140.310 22.460 170.850 23.930 ;
        RECT 140.310 19.595 141.910 22.460 ;
        RECT 143.520 22.330 167.640 22.460 ;
        RECT 143.520 19.595 154.040 22.330 ;
        RECT 140.310 19.590 154.040 19.595 ;
        RECT 157.120 19.800 167.640 22.330 ;
        RECT 169.250 21.985 170.850 22.460 ;
        RECT 172.450 28.720 174.050 28.865 ;
        RECT 175.660 28.850 186.180 31.590 ;
        RECT 189.260 28.850 199.780 31.590 ;
        RECT 202.860 28.850 213.380 31.590 ;
        RECT 216.460 28.850 226.980 31.590 ;
        RECT 175.660 28.720 226.980 28.850 ;
        RECT 228.590 28.720 230.190 31.590 ;
        RECT 233.720 31.250 238.520 32.850 ;
        RECT 232.420 29.650 235.320 31.250 ;
        RECT 236.920 29.650 239.820 31.250 ;
        RECT 172.450 28.050 230.190 28.720 ;
        RECT 233.720 28.050 238.520 29.650 ;
        RECT 172.450 27.250 235.320 28.050 ;
        RECT 172.450 27.130 186.190 27.250 ;
        RECT 172.450 27.120 177.380 27.130 ;
        RECT 172.450 24.060 174.050 27.120 ;
        RECT 175.780 24.060 177.380 27.120 ;
        RECT 172.450 24.050 177.380 24.060 ;
        RECT 180.120 24.050 181.720 27.130 ;
        RECT 184.460 27.120 186.190 27.130 ;
        RECT 189.250 27.130 199.790 27.250 ;
        RECT 189.250 27.120 190.980 27.130 ;
        RECT 184.460 24.060 186.060 27.120 ;
        RECT 189.380 24.060 190.980 27.120 ;
        RECT 184.460 24.050 186.190 24.060 ;
        RECT 172.450 23.930 186.190 24.050 ;
        RECT 189.250 24.050 190.980 24.060 ;
        RECT 193.720 24.050 195.320 27.130 ;
        RECT 198.060 27.120 199.790 27.130 ;
        RECT 202.850 27.130 213.390 27.250 ;
        RECT 202.850 27.120 204.580 27.130 ;
        RECT 198.060 24.060 199.660 27.120 ;
        RECT 202.980 24.060 204.580 27.120 ;
        RECT 198.060 24.050 199.790 24.060 ;
        RECT 189.250 23.930 199.790 24.050 ;
        RECT 202.850 24.050 204.580 24.060 ;
        RECT 207.320 24.050 208.920 27.130 ;
        RECT 211.660 27.120 213.390 27.130 ;
        RECT 216.450 27.130 235.320 27.250 ;
        RECT 216.450 27.120 218.180 27.130 ;
        RECT 211.660 24.060 213.260 27.120 ;
        RECT 216.580 24.060 218.180 27.120 ;
        RECT 211.660 24.050 213.390 24.060 ;
        RECT 202.850 23.930 213.390 24.050 ;
        RECT 216.450 24.050 218.180 24.060 ;
        RECT 220.920 24.050 222.520 27.130 ;
        RECT 225.260 27.120 235.320 27.130 ;
        RECT 225.260 24.060 226.860 27.120 ;
        RECT 228.590 26.450 235.320 27.120 ;
        RECT 236.920 26.450 239.820 28.050 ;
        RECT 228.590 24.060 230.190 26.450 ;
        RECT 233.720 24.850 238.520 26.450 ;
        RECT 225.260 24.050 230.190 24.060 ;
        RECT 216.450 23.930 230.190 24.050 ;
        RECT 172.450 22.460 230.190 23.930 ;
        RECT 232.420 23.250 235.320 24.850 ;
        RECT 236.920 23.250 239.820 24.850 ;
        RECT 172.450 21.985 174.050 22.460 ;
        RECT 169.250 20.385 174.050 21.985 ;
        RECT 169.250 19.800 170.850 20.385 ;
        RECT 157.120 19.590 170.850 19.800 ;
        RECT 140.310 18.195 170.850 19.590 ;
        RECT 140.310 17.995 167.640 18.195 ;
        RECT 140.310 15.130 141.910 17.995 ;
        RECT 143.520 17.990 167.640 17.995 ;
        RECT 143.520 15.250 154.040 17.990 ;
        RECT 157.120 15.530 167.640 17.990 ;
        RECT 169.250 17.515 170.850 18.195 ;
        RECT 172.450 19.595 174.050 20.385 ;
        RECT 175.660 22.330 226.980 22.460 ;
        RECT 175.660 19.595 186.180 22.330 ;
        RECT 172.450 19.590 186.180 19.595 ;
        RECT 189.260 19.590 199.780 22.330 ;
        RECT 202.860 19.590 213.380 22.330 ;
        RECT 216.460 19.800 226.980 22.330 ;
        RECT 228.590 21.650 230.190 22.460 ;
        RECT 233.720 21.650 238.520 23.250 ;
        RECT 228.590 20.050 235.320 21.650 ;
        RECT 236.920 20.050 239.820 21.650 ;
        RECT 228.590 19.800 230.190 20.050 ;
        RECT 216.460 19.590 230.190 19.800 ;
        RECT 172.450 18.195 230.190 19.590 ;
        RECT 233.720 18.450 238.520 20.050 ;
        RECT 172.450 17.995 226.980 18.195 ;
        RECT 172.450 17.515 174.050 17.995 ;
        RECT 169.250 15.915 174.050 17.515 ;
        RECT 169.250 15.530 170.850 15.915 ;
        RECT 157.120 15.250 170.850 15.530 ;
        RECT 143.520 15.130 170.850 15.250 ;
        RECT 140.310 13.930 170.850 15.130 ;
        RECT 140.310 13.650 167.640 13.930 ;
        RECT 140.310 13.530 154.050 13.650 ;
        RECT 140.310 11.920 141.910 13.530 ;
        RECT 143.920 11.920 145.520 13.530 ;
        RECT 148.185 11.920 149.790 13.530 ;
        RECT 152.450 11.920 154.050 13.530 ;
        RECT 157.110 13.530 167.640 13.650 ;
        RECT 157.110 11.920 158.710 13.530 ;
        RECT 161.575 11.920 163.175 13.530 ;
        RECT 166.040 11.920 167.640 13.530 ;
        RECT 169.250 13.045 170.850 13.930 ;
        RECT 172.450 15.130 174.050 15.915 ;
        RECT 175.660 17.990 226.980 17.995 ;
        RECT 175.660 15.250 186.180 17.990 ;
        RECT 189.260 15.250 199.780 17.990 ;
        RECT 202.860 15.250 213.380 17.990 ;
        RECT 216.460 15.530 226.980 17.990 ;
        RECT 228.590 15.530 230.190 18.195 ;
        RECT 232.420 16.850 235.320 18.450 ;
        RECT 236.920 16.850 239.820 18.450 ;
        RECT 216.460 15.250 230.190 15.530 ;
        RECT 233.720 15.250 238.520 16.850 ;
        RECT 175.660 15.130 235.320 15.250 ;
        RECT 172.450 13.930 235.320 15.130 ;
        RECT 172.450 13.650 226.980 13.930 ;
        RECT 172.450 13.530 186.190 13.650 ;
        RECT 172.450 13.045 174.050 13.530 ;
        RECT 169.250 11.920 174.050 13.045 ;
        RECT 176.060 11.920 177.660 13.530 ;
        RECT 180.325 11.920 181.930 13.530 ;
        RECT 184.590 11.920 186.190 13.530 ;
        RECT 189.250 13.530 199.790 13.650 ;
        RECT 189.250 11.920 190.850 13.530 ;
        RECT 193.720 11.920 195.320 13.530 ;
        RECT 198.190 11.920 199.790 13.530 ;
        RECT 202.850 13.530 213.390 13.650 ;
        RECT 202.850 11.920 204.450 13.530 ;
        RECT 207.320 11.920 208.920 13.530 ;
        RECT 211.790 11.920 213.390 13.530 ;
        RECT 216.450 13.530 226.980 13.650 ;
        RECT 216.450 11.920 218.050 13.530 ;
        RECT 220.915 11.920 222.515 13.530 ;
        RECT 225.380 11.920 226.980 13.530 ;
        RECT 228.590 13.650 235.320 13.930 ;
        RECT 228.590 11.920 230.190 13.650 ;
        RECT 140.310 11.445 230.190 11.920 ;
        RECT 140.310 10.320 170.850 11.445 ;
        RECT 172.450 10.320 230.190 11.445 ;
        RECT 9.570 6.100 11.170 7.400 ;
        RECT 12.770 6.100 14.370 10.320 ;
        RECT 15.970 6.100 17.570 7.400 ;
        RECT 19.170 6.100 20.770 10.320 ;
        RECT 22.370 6.100 23.970 7.400 ;
        RECT 25.570 6.100 27.170 10.320 ;
        RECT 28.770 6.100 30.370 7.400 ;
        RECT 31.970 6.100 33.570 10.320 ;
        RECT 35.170 6.100 36.770 7.400 ;
        RECT 38.370 6.100 39.970 10.320 ;
        RECT 41.570 6.100 43.170 7.400 ;
        RECT 44.770 6.100 46.370 10.320 ;
        RECT 47.970 6.100 49.570 7.400 ;
        RECT 51.170 6.100 52.770 10.320 ;
        RECT 54.370 6.100 55.970 7.400 ;
        RECT 57.570 6.100 59.170 10.320 ;
        RECT 60.770 6.100 62.370 7.400 ;
        RECT 63.970 6.100 65.570 10.320 ;
        RECT 67.170 6.100 68.770 7.400 ;
        RECT 70.370 6.100 71.970 10.320 ;
        RECT 73.570 6.100 75.170 7.400 ;
        RECT 76.770 6.100 78.370 7.400 ;
        RECT 79.970 6.100 81.570 7.400 ;
        RECT 83.170 6.100 84.770 10.320 ;
        RECT 86.370 6.100 87.970 7.400 ;
        RECT 89.570 6.100 91.170 10.320 ;
        RECT 92.770 6.100 94.370 7.400 ;
        RECT 95.970 6.100 97.570 10.320 ;
        RECT 99.170 6.100 100.770 7.400 ;
        RECT 102.370 6.100 103.970 7.400 ;
        RECT 105.570 6.100 107.170 7.400 ;
        RECT 108.770 6.100 110.370 7.400 ;
        RECT 111.970 6.100 113.570 7.400 ;
        RECT 115.170 6.100 116.770 7.400 ;
        RECT 123.610 6.100 125.210 7.400 ;
        RECT 126.810 6.100 128.410 7.400 ;
        RECT 130.010 6.100 131.610 7.400 ;
        RECT 133.210 6.100 134.810 7.400 ;
        RECT 136.410 6.100 138.010 7.400 ;
        RECT 139.610 6.100 141.210 7.400 ;
        RECT 142.810 6.100 144.410 10.320 ;
        RECT 146.010 6.100 147.610 7.400 ;
        RECT 149.210 6.100 150.810 10.320 ;
        RECT 152.410 6.100 154.010 7.400 ;
        RECT 155.610 6.100 157.210 10.320 ;
        RECT 158.810 6.100 160.410 7.400 ;
        RECT 162.010 6.100 163.610 7.400 ;
        RECT 165.210 6.100 166.810 7.400 ;
        RECT 168.410 6.100 170.010 10.320 ;
        RECT 171.610 6.100 173.210 7.400 ;
        RECT 174.810 6.100 176.410 10.320 ;
        RECT 178.010 6.100 179.610 7.400 ;
        RECT 181.210 6.100 182.810 10.320 ;
        RECT 184.410 6.100 186.010 7.400 ;
        RECT 187.610 6.100 189.210 10.320 ;
        RECT 190.810 6.100 192.410 7.400 ;
        RECT 194.010 6.100 195.610 10.320 ;
        RECT 197.210 6.100 198.810 7.400 ;
        RECT 200.410 6.100 202.010 10.320 ;
        RECT 203.610 6.100 205.210 7.400 ;
        RECT 206.810 6.100 208.410 10.320 ;
        RECT 210.010 6.100 211.610 7.400 ;
        RECT 213.210 6.100 214.810 10.320 ;
        RECT 216.410 6.100 218.010 7.400 ;
        RECT 219.610 6.100 221.210 10.320 ;
        RECT 222.810 6.100 224.410 7.400 ;
        RECT 226.010 6.100 227.610 10.320 ;
        RECT 229.210 6.100 230.810 7.400 ;
        RECT 233.720 6.100 235.320 13.650 ;
        RECT 236.920 13.650 239.820 15.250 ;
        RECT 236.920 6.100 238.520 13.650 ;
        RECT -0.130 4.500 253.790 6.100 ;
        RECT 1.860 2.900 3.460 4.500 ;
        RECT 7.970 2.900 9.570 4.500 ;
        RECT 11.170 2.900 12.770 4.500 ;
        RECT 14.370 2.900 15.970 4.500 ;
        RECT 17.570 2.900 19.170 4.500 ;
        RECT 20.770 2.900 22.370 4.500 ;
        RECT 23.970 2.900 25.570 4.500 ;
        RECT 27.170 2.900 28.770 4.500 ;
        RECT 30.370 2.900 31.970 4.500 ;
        RECT 33.570 2.900 35.170 4.500 ;
        RECT 36.770 2.900 38.370 4.500 ;
        RECT 39.970 2.900 41.570 4.500 ;
        RECT 43.170 2.900 44.770 4.500 ;
        RECT 46.370 2.900 47.970 4.500 ;
        RECT 49.570 2.900 51.170 4.500 ;
        RECT 52.770 2.900 54.370 4.500 ;
        RECT 55.970 2.900 57.570 4.500 ;
        RECT 59.170 2.900 60.770 4.500 ;
        RECT 62.370 2.900 63.970 4.500 ;
        RECT 65.570 2.900 67.170 4.500 ;
        RECT 68.770 2.900 70.370 4.500 ;
        RECT 71.970 2.900 73.570 4.500 ;
        RECT 75.170 2.900 76.770 4.500 ;
        RECT 78.370 2.900 79.970 4.500 ;
        RECT 81.570 2.900 83.170 4.500 ;
        RECT 84.770 2.900 86.370 4.500 ;
        RECT 87.970 2.900 89.570 4.500 ;
        RECT 91.170 2.900 92.770 4.500 ;
        RECT 94.370 2.900 95.970 4.500 ;
        RECT 97.570 2.900 99.170 4.500 ;
        RECT 100.770 2.900 102.370 4.500 ;
        RECT 103.970 2.900 105.570 4.500 ;
        RECT 107.170 2.900 108.770 4.500 ;
        RECT 110.370 2.900 111.970 4.500 ;
        RECT 113.570 2.900 115.170 4.500 ;
        RECT 116.770 2.900 118.370 4.500 ;
        RECT 122.010 2.900 123.610 4.500 ;
        RECT 125.210 2.900 126.810 4.500 ;
        RECT 128.410 2.900 130.010 4.500 ;
        RECT 131.610 2.900 133.210 4.500 ;
        RECT 134.810 2.900 136.410 4.500 ;
        RECT 138.010 2.900 139.610 4.500 ;
        RECT 141.210 2.900 142.810 4.500 ;
        RECT 144.410 2.900 146.010 4.500 ;
        RECT 147.610 2.900 149.210 4.500 ;
        RECT 150.810 2.900 152.410 4.500 ;
        RECT 154.010 2.900 155.610 4.500 ;
        RECT 157.210 2.900 158.810 4.500 ;
        RECT 160.410 2.900 162.010 4.500 ;
        RECT 163.610 2.900 165.210 4.500 ;
        RECT 166.810 2.900 168.410 4.500 ;
        RECT 170.010 2.900 171.610 4.500 ;
        RECT 173.210 2.900 174.810 4.500 ;
        RECT 176.410 2.900 178.010 4.500 ;
        RECT 179.610 2.900 181.210 4.500 ;
        RECT 182.810 2.900 184.410 4.500 ;
        RECT 186.010 2.900 187.610 4.500 ;
        RECT 189.210 2.900 190.810 4.500 ;
        RECT 192.410 2.900 194.010 4.500 ;
        RECT 195.610 2.900 197.210 4.500 ;
        RECT 198.810 2.900 200.410 4.500 ;
        RECT 202.010 2.900 203.610 4.500 ;
        RECT 205.210 2.900 206.810 4.500 ;
        RECT 208.410 2.900 210.010 4.500 ;
        RECT 211.610 2.900 213.210 4.500 ;
        RECT 214.810 2.900 216.410 4.500 ;
        RECT 218.010 2.900 219.610 4.500 ;
        RECT 221.210 2.900 222.810 4.500 ;
        RECT 224.410 2.900 226.010 4.500 ;
        RECT 227.610 2.900 229.210 4.500 ;
        RECT 230.810 2.900 232.410 4.500 ;
        RECT 236.920 2.900 238.520 4.500 ;
        RECT -0.130 1.300 253.790 2.900 ;
        RECT 9.570 0.000 11.170 1.300 ;
        RECT 12.770 0.000 14.370 1.300 ;
        RECT 15.970 0.000 17.570 1.300 ;
        RECT 19.170 0.000 20.770 1.300 ;
        RECT 22.370 0.000 23.970 1.300 ;
        RECT 25.570 0.000 27.170 1.300 ;
        RECT 28.770 0.000 30.370 1.300 ;
        RECT 31.970 0.000 33.570 1.300 ;
        RECT 35.170 0.000 36.770 1.300 ;
        RECT 38.370 0.000 39.970 1.300 ;
        RECT 41.570 0.000 43.170 1.300 ;
        RECT 44.770 0.000 46.370 1.300 ;
        RECT 47.970 0.000 49.570 1.300 ;
        RECT 51.170 0.000 52.770 1.300 ;
        RECT 54.370 0.000 55.970 1.300 ;
        RECT 57.570 0.000 59.170 1.300 ;
        RECT 60.770 0.000 62.370 1.300 ;
        RECT 63.970 0.000 65.570 1.300 ;
        RECT 67.170 0.000 68.770 1.300 ;
        RECT 70.370 0.000 71.970 1.300 ;
        RECT 73.570 0.000 75.170 1.300 ;
        RECT 76.770 0.000 78.370 1.300 ;
        RECT 79.970 0.000 81.570 1.300 ;
        RECT 83.170 0.000 84.770 1.300 ;
        RECT 86.370 0.000 87.970 1.300 ;
        RECT 89.570 0.000 91.170 1.300 ;
        RECT 92.770 0.000 94.370 1.300 ;
        RECT 95.970 0.000 97.570 1.300 ;
        RECT 99.170 0.000 100.770 1.300 ;
        RECT 102.370 0.000 103.970 1.300 ;
        RECT 105.570 0.000 107.170 1.300 ;
        RECT 108.770 0.000 110.370 1.300 ;
        RECT 111.970 0.000 113.570 1.300 ;
        RECT 115.170 0.000 116.770 1.300 ;
        RECT 123.610 0.000 125.210 1.300 ;
        RECT 126.810 0.000 128.410 1.300 ;
        RECT 130.010 0.000 131.610 1.300 ;
        RECT 133.210 0.000 134.810 1.300 ;
        RECT 136.410 0.000 138.010 1.300 ;
        RECT 139.610 0.000 141.210 1.300 ;
        RECT 142.810 0.000 144.410 1.300 ;
        RECT 146.010 0.000 147.610 1.300 ;
        RECT 149.210 0.000 150.810 1.300 ;
        RECT 152.410 0.000 154.010 1.300 ;
        RECT 155.610 0.000 157.210 1.300 ;
        RECT 158.810 0.000 160.410 1.300 ;
        RECT 162.010 0.000 163.610 1.300 ;
        RECT 165.210 0.000 166.810 1.300 ;
        RECT 168.410 0.000 170.010 1.300 ;
        RECT 171.610 0.000 173.210 1.300 ;
        RECT 174.810 0.000 176.410 1.300 ;
        RECT 178.010 0.000 179.610 1.300 ;
        RECT 181.210 0.000 182.810 1.300 ;
        RECT 184.410 0.000 186.010 1.300 ;
        RECT 187.610 0.000 189.210 1.300 ;
        RECT 190.810 0.000 192.410 1.300 ;
        RECT 194.010 0.000 195.610 1.300 ;
        RECT 197.210 0.000 198.810 1.300 ;
        RECT 200.410 0.000 202.010 1.300 ;
        RECT 203.610 0.000 205.210 1.300 ;
        RECT 206.810 0.000 208.410 1.300 ;
        RECT 210.010 0.000 211.610 1.300 ;
        RECT 213.210 0.000 214.810 1.300 ;
        RECT 216.410 0.000 218.010 1.300 ;
        RECT 219.610 0.000 221.210 1.300 ;
        RECT 222.810 0.000 224.410 1.300 ;
        RECT 226.010 0.000 227.610 1.300 ;
        RECT 229.210 0.000 230.810 1.300 ;
    END
  END vssd
  PIN vccd
    DIRECTION INOUT ;
    ANTENNAGATEAREA 0.302400 ;
    ANTENNADIFFAREA 10.175475 ;
    PORT
      LAYER nwell ;
        RECT 43.885 170.800 46.660 171.865 ;
        RECT 92.780 170.680 95.555 171.745 ;
        RECT 127.065 170.255 131.590 171.110 ;
        RECT 194.860 170.800 197.635 171.865 ;
        RECT 127.065 168.815 131.585 170.255 ;
        RECT 44.130 166.895 46.660 167.960 ;
        RECT 93.025 165.240 95.555 167.840 ;
        RECT 194.860 166.895 197.390 167.960 ;
        RECT 127.065 164.765 131.585 166.205 ;
        RECT 127.065 163.910 131.590 164.765 ;
        RECT 92.780 161.335 95.555 162.400 ;
        RECT 111.145 132.175 116.160 134.530 ;
        RECT 117.695 130.340 122.745 132.300 ;
        RECT 124.280 132.175 129.295 134.580 ;
      LAYER li1 ;
        RECT 43.770 172.015 46.990 172.185 ;
        RECT 44.155 171.600 44.325 172.015 ;
        RECT 92.665 171.895 95.885 172.065 ;
        RECT 194.530 172.015 197.750 172.185 ;
        RECT 44.060 170.980 44.435 171.600 ;
        RECT 93.050 171.480 93.220 171.895 ;
        RECT 197.195 171.600 197.365 172.015 ;
        RECT 92.955 170.860 93.330 171.480 ;
        RECT 197.085 170.980 197.460 171.600 ;
        RECT 45.930 170.310 46.100 170.640 ;
        RECT 94.825 170.190 94.995 170.520 ;
        RECT 128.830 170.315 129.080 170.685 ;
        RECT 127.255 170.145 131.395 170.315 ;
        RECT 195.420 170.310 195.590 170.640 ;
        RECT 127.510 169.345 127.765 170.145 ;
        RECT 128.435 169.345 128.605 170.145 ;
        RECT 129.275 169.345 129.445 170.145 ;
        RECT 130.115 169.345 130.285 170.145 ;
        RECT 130.955 169.345 131.255 170.145 ;
        RECT 44.775 167.755 45.065 167.765 ;
        RECT 45.940 167.760 46.230 167.770 ;
        RECT 195.290 167.760 195.580 167.770 ;
        RECT 44.390 167.150 45.100 167.755 ;
        RECT 44.410 167.110 45.100 167.150 ;
        RECT 45.895 167.155 46.265 167.760 ;
        RECT 93.670 167.635 93.960 167.645 ;
        RECT 94.835 167.640 95.125 167.650 ;
        RECT 45.895 167.115 46.260 167.155 ;
        RECT 44.410 166.745 44.960 167.110 ;
        RECT 45.970 166.745 46.150 167.115 ;
        RECT 93.285 167.030 93.995 167.635 ;
        RECT 93.305 166.990 93.995 167.030 ;
        RECT 94.790 167.035 95.160 167.640 ;
        RECT 195.255 167.155 195.625 167.760 ;
        RECT 196.455 167.755 196.745 167.765 ;
        RECT 195.260 167.115 195.625 167.155 ;
        RECT 196.420 167.150 197.130 167.755 ;
        RECT 94.790 166.995 95.155 167.035 ;
        RECT 43.770 166.575 46.990 166.745 ;
        RECT 93.305 166.625 93.855 166.990 ;
        RECT 94.865 166.625 95.045 166.995 ;
        RECT 195.370 166.745 195.550 167.115 ;
        RECT 196.420 167.110 197.110 167.150 ;
        RECT 196.560 166.745 197.110 167.110 ;
        RECT 92.665 166.455 95.885 166.625 ;
        RECT 194.530 166.575 197.750 166.745 ;
        RECT 93.305 166.090 93.855 166.455 ;
        RECT 93.305 166.050 93.995 166.090 ;
        RECT 94.865 166.085 95.045 166.455 ;
        RECT 93.285 165.445 93.995 166.050 ;
        RECT 94.790 166.045 95.155 166.085 ;
        RECT 93.670 165.435 93.960 165.445 ;
        RECT 94.790 165.440 95.160 166.045 ;
        RECT 94.835 165.430 95.125 165.440 ;
        RECT 127.510 164.875 127.765 165.675 ;
        RECT 128.435 164.875 128.605 165.675 ;
        RECT 129.275 164.875 129.445 165.675 ;
        RECT 130.115 164.875 130.285 165.675 ;
        RECT 130.955 164.875 131.255 165.675 ;
        RECT 127.255 164.705 131.395 164.875 ;
        RECT 128.830 164.335 129.080 164.705 ;
        RECT 94.825 162.560 94.995 162.890 ;
        RECT 92.955 161.600 93.330 162.220 ;
        RECT 93.050 161.185 93.220 161.600 ;
        RECT 92.665 161.015 95.885 161.185 ;
        RECT 114.285 133.295 114.515 134.130 ;
        RECT 125.295 133.815 125.615 134.250 ;
        RECT 119.220 133.530 121.220 133.700 ;
        RECT 111.910 132.915 112.260 133.295 ;
        RECT 113.070 132.915 113.420 133.295 ;
        RECT 114.230 132.915 114.580 133.295 ;
        RECT 115.390 132.915 115.740 133.295 ;
        RECT 118.105 131.430 118.330 131.810 ;
        RECT 120.135 131.790 120.305 133.530 ;
        RECT 124.700 132.915 125.050 133.295 ;
        RECT 125.860 132.915 126.210 133.295 ;
        RECT 127.020 132.915 127.370 133.295 ;
        RECT 128.180 132.915 128.530 133.295 ;
        RECT 120.080 131.510 120.360 131.790 ;
        RECT 120.135 130.615 120.305 131.510 ;
        RECT 122.110 131.430 122.335 131.810 ;
      LAYER mcon ;
        RECT 43.915 172.015 44.085 172.185 ;
        RECT 44.375 172.015 44.545 172.185 ;
        RECT 44.835 172.015 45.005 172.185 ;
        RECT 45.295 172.015 45.465 172.185 ;
        RECT 45.755 172.015 45.925 172.185 ;
        RECT 46.215 172.015 46.385 172.185 ;
        RECT 46.675 172.015 46.845 172.185 ;
        RECT 92.810 171.895 92.980 172.065 ;
        RECT 93.270 171.895 93.440 172.065 ;
        RECT 93.730 171.895 93.900 172.065 ;
        RECT 94.190 171.895 94.360 172.065 ;
        RECT 94.650 171.895 94.820 172.065 ;
        RECT 95.110 171.895 95.280 172.065 ;
        RECT 95.570 171.895 95.740 172.065 ;
        RECT 194.675 172.015 194.845 172.185 ;
        RECT 195.135 172.015 195.305 172.185 ;
        RECT 195.595 172.015 195.765 172.185 ;
        RECT 196.055 172.015 196.225 172.185 ;
        RECT 196.515 172.015 196.685 172.185 ;
        RECT 196.975 172.015 197.145 172.185 ;
        RECT 197.435 172.015 197.605 172.185 ;
        RECT 45.930 170.390 46.100 170.560 ;
        RECT 94.825 170.270 94.995 170.440 ;
        RECT 195.420 170.390 195.590 170.560 ;
        RECT 127.400 170.145 127.570 170.315 ;
        RECT 127.860 170.145 128.030 170.315 ;
        RECT 128.320 170.145 128.490 170.315 ;
        RECT 128.780 170.145 128.950 170.315 ;
        RECT 129.240 170.145 129.410 170.315 ;
        RECT 129.700 170.145 129.870 170.315 ;
        RECT 130.160 170.145 130.330 170.315 ;
        RECT 130.620 170.145 130.790 170.315 ;
        RECT 131.080 170.145 131.250 170.315 ;
        RECT 43.915 166.575 44.085 166.745 ;
        RECT 44.375 166.575 44.545 166.745 ;
        RECT 44.835 166.575 45.005 166.745 ;
        RECT 45.295 166.575 45.465 166.745 ;
        RECT 45.755 166.575 45.925 166.745 ;
        RECT 46.215 166.575 46.385 166.745 ;
        RECT 46.675 166.575 46.845 166.745 ;
        RECT 92.810 166.455 92.980 166.625 ;
        RECT 93.270 166.455 93.440 166.625 ;
        RECT 93.730 166.455 93.900 166.625 ;
        RECT 94.190 166.455 94.360 166.625 ;
        RECT 94.650 166.455 94.820 166.625 ;
        RECT 95.110 166.455 95.280 166.625 ;
        RECT 95.570 166.455 95.740 166.625 ;
        RECT 194.675 166.575 194.845 166.745 ;
        RECT 195.135 166.575 195.305 166.745 ;
        RECT 195.595 166.575 195.765 166.745 ;
        RECT 196.055 166.575 196.225 166.745 ;
        RECT 196.515 166.575 196.685 166.745 ;
        RECT 196.975 166.575 197.145 166.745 ;
        RECT 197.435 166.575 197.605 166.745 ;
        RECT 127.400 164.705 127.570 164.875 ;
        RECT 127.860 164.705 128.030 164.875 ;
        RECT 128.320 164.705 128.490 164.875 ;
        RECT 128.780 164.705 128.950 164.875 ;
        RECT 129.240 164.705 129.410 164.875 ;
        RECT 129.700 164.705 129.870 164.875 ;
        RECT 130.160 164.705 130.330 164.875 ;
        RECT 130.620 164.705 130.790 164.875 ;
        RECT 131.080 164.705 131.250 164.875 ;
        RECT 94.825 162.640 94.995 162.810 ;
        RECT 92.810 161.015 92.980 161.185 ;
        RECT 93.270 161.015 93.440 161.185 ;
        RECT 93.730 161.015 93.900 161.185 ;
        RECT 94.190 161.015 94.360 161.185 ;
        RECT 94.650 161.015 94.820 161.185 ;
        RECT 95.110 161.015 95.280 161.185 ;
        RECT 95.570 161.015 95.740 161.185 ;
        RECT 125.300 133.920 125.605 134.175 ;
        RECT 111.990 132.965 112.160 133.255 ;
        RECT 113.150 132.965 113.320 133.255 ;
        RECT 114.310 132.965 114.480 133.255 ;
        RECT 115.470 132.965 115.640 133.255 ;
        RECT 124.800 132.965 124.970 133.255 ;
        RECT 125.960 132.965 126.130 133.255 ;
        RECT 127.120 132.965 127.290 133.255 ;
        RECT 128.280 132.965 128.450 133.255 ;
        RECT 118.120 131.550 118.290 131.720 ;
        RECT 120.135 131.565 120.305 131.735 ;
        RECT 122.150 131.550 122.320 131.720 ;
        RECT 120.135 130.695 120.305 130.865 ;
      LAYER met1 ;
        RECT 46.685 172.340 46.905 172.345 ;
        RECT 194.615 172.340 194.835 172.345 ;
        RECT 42.450 171.860 46.990 172.340 ;
        RECT 92.665 172.220 95.800 172.225 ;
        RECT 42.450 166.900 42.950 171.860 ;
        RECT 45.880 170.575 46.150 170.645 ;
        RECT 46.685 170.575 46.905 171.860 ;
        RECT 92.665 171.740 95.885 172.220 ;
        RECT 194.530 171.860 199.070 172.340 ;
        RECT 45.880 170.375 46.905 170.575 ;
        RECT 94.775 170.455 95.045 170.525 ;
        RECT 95.580 170.455 95.800 171.740 ;
        RECT 194.615 170.575 194.835 171.860 ;
        RECT 195.370 170.575 195.640 170.645 ;
        RECT 45.880 170.305 46.150 170.375 ;
        RECT 94.775 170.255 95.800 170.455 ;
        RECT 94.775 170.185 95.045 170.255 ;
        RECT 127.255 169.990 131.395 170.470 ;
        RECT 194.615 170.375 195.640 170.575 ;
        RECT 195.370 170.305 195.640 170.375 ;
        RECT 198.570 166.900 199.070 171.860 ;
        RECT 42.450 166.420 46.990 166.900 ;
        RECT 92.665 166.300 95.885 166.780 ;
        RECT 194.530 166.420 199.070 166.900 ;
        RECT 127.255 164.550 131.395 165.030 ;
        RECT 94.775 162.825 95.045 162.895 ;
        RECT 94.775 162.625 95.800 162.825 ;
        RECT 94.775 162.555 95.045 162.625 ;
        RECT 95.580 161.340 95.800 162.625 ;
        RECT 92.665 160.860 95.885 161.340 ;
        RECT 95.580 160.855 95.800 160.860 ;
        RECT 125.270 133.920 125.660 134.240 ;
        RECT 111.910 133.720 128.530 133.920 ;
        RECT 111.910 133.485 112.260 133.720 ;
        RECT 113.070 133.485 113.420 133.720 ;
        RECT 114.230 133.485 114.580 133.720 ;
        RECT 115.390 133.485 115.740 133.720 ;
        RECT 111.990 133.295 112.160 133.485 ;
        RECT 113.150 133.295 113.320 133.485 ;
        RECT 114.310 133.295 114.480 133.485 ;
        RECT 115.470 133.295 115.640 133.485 ;
        RECT 116.400 133.440 124.040 133.720 ;
        RECT 124.700 133.485 125.050 133.720 ;
        RECT 125.860 133.485 126.210 133.720 ;
        RECT 127.020 133.485 127.370 133.720 ;
        RECT 128.180 133.485 128.530 133.720 ;
        RECT 124.800 133.295 124.970 133.485 ;
        RECT 125.960 133.295 126.130 133.485 ;
        RECT 127.120 133.295 127.290 133.485 ;
        RECT 128.280 133.295 128.450 133.485 ;
        RECT 111.930 132.915 112.220 133.295 ;
        RECT 113.090 132.915 113.380 133.295 ;
        RECT 114.250 132.915 114.540 133.295 ;
        RECT 115.410 132.915 115.700 133.295 ;
        RECT 124.740 132.915 125.030 133.295 ;
        RECT 125.900 132.915 126.190 133.295 ;
        RECT 127.060 132.915 127.350 133.295 ;
        RECT 128.220 132.915 128.510 133.295 ;
        RECT 118.090 131.720 118.325 131.750 ;
        RECT 120.105 131.735 120.335 131.770 ;
        RECT 118.060 131.705 118.350 131.720 ;
        RECT 120.075 131.705 120.365 131.735 ;
        RECT 122.120 131.720 122.355 131.765 ;
        RECT 122.085 131.705 122.380 131.720 ;
        RECT 118.060 131.565 122.380 131.705 ;
        RECT 118.060 131.550 118.350 131.565 ;
        RECT 118.090 131.520 118.325 131.550 ;
        RECT 120.105 131.535 120.335 131.565 ;
        RECT 122.085 131.550 122.380 131.565 ;
        RECT 122.120 131.520 122.355 131.550 ;
        RECT 120.085 130.615 120.355 130.945 ;
      LAYER via ;
        RECT 93.240 171.875 93.500 172.135 ;
        RECT 127.810 170.095 128.070 170.355 ;
        RECT 44.810 166.460 45.970 166.850 ;
        RECT 93.220 166.430 93.480 166.690 ;
        RECT 195.550 166.460 196.710 166.850 ;
        RECT 127.390 164.590 128.450 165.030 ;
        RECT 93.215 160.955 93.490 161.240 ;
        RECT 120.090 133.530 120.350 133.790 ;
      LAYER met2 ;
        RECT 93.230 171.820 93.510 172.190 ;
        RECT 127.800 170.040 128.090 170.420 ;
        RECT 44.810 154.990 45.970 166.900 ;
        RECT 93.210 166.375 93.490 166.745 ;
        RECT 93.200 160.890 93.500 161.300 ;
        RECT 44.760 154.380 46.020 154.990 ;
        RECT 120.045 133.500 120.400 154.850 ;
        RECT 127.340 154.380 128.500 165.070 ;
        RECT 195.550 154.990 196.710 166.900 ;
        RECT 195.500 154.380 196.760 154.990 ;
      LAYER via2 ;
        RECT 93.230 171.865 93.510 172.145 ;
        RECT 127.800 170.085 128.090 170.375 ;
        RECT 93.210 166.420 93.490 166.700 ;
        RECT 127.390 164.590 128.450 165.030 ;
        RECT 93.200 160.935 93.500 161.255 ;
        RECT 44.810 154.430 45.970 154.950 ;
        RECT 120.085 154.510 120.365 154.790 ;
        RECT 127.370 154.430 128.470 154.930 ;
        RECT 195.550 154.430 196.710 154.950 ;
      LAYER met3 ;
        RECT 93.125 171.750 93.615 172.240 ;
        RECT 127.700 169.980 128.200 170.475 ;
        RECT 93.105 166.305 93.595 166.795 ;
        RECT 127.340 164.550 128.500 165.070 ;
        RECT 93.055 160.785 93.680 161.410 ;
        RECT 44.760 154.930 46.020 154.990 ;
        RECT 127.340 154.930 128.500 154.980 ;
        RECT 195.500 154.930 196.760 154.990 ;
        RECT -0.130 154.430 253.790 154.930 ;
        RECT 44.760 154.380 46.020 154.430 ;
        RECT 127.340 154.380 128.500 154.430 ;
        RECT 195.500 154.380 196.760 154.430 ;
      LAYER via3 ;
        RECT 93.210 171.845 93.530 172.165 ;
        RECT 127.780 170.070 128.100 170.390 ;
        RECT 93.190 166.400 93.510 166.720 ;
        RECT 127.390 164.590 128.450 165.030 ;
        RECT 93.190 160.935 93.510 161.255 ;
        RECT 93.120 154.475 93.550 154.855 ;
      LAYER met4 ;
        RECT 93.105 161.305 93.575 172.245 ;
        RECT 127.750 165.070 128.125 170.395 ;
        RECT 127.340 164.550 128.500 165.070 ;
        RECT 93.090 154.430 93.580 161.305 ;
    END
  END vccd
  OBS
      LAYER pwell ;
        RECT 121.635 167.615 125.505 168.525 ;
        RECT 127.425 167.615 131.295 168.525 ;
        RECT 121.635 167.595 121.780 167.615 ;
        RECT 127.425 167.595 127.570 167.615 ;
        RECT 121.610 167.425 121.780 167.595 ;
        RECT 127.400 167.425 127.570 167.595 ;
        RECT 121.635 167.405 121.780 167.425 ;
        RECT 127.425 167.405 127.570 167.425 ;
        RECT 121.635 166.495 125.505 167.405 ;
        RECT 127.425 166.495 131.295 167.405 ;
      LAYER li1 ;
        RECT 113.330 175.275 113.695 175.315 ;
        RECT 116.090 175.275 116.455 175.315 ;
        RECT 106.890 173.700 107.260 174.890 ;
        RECT 110.840 173.960 111.185 175.205 ;
        RECT 113.330 174.670 113.700 175.275 ;
        RECT 116.090 174.670 116.460 175.275 ;
        RECT 113.375 174.660 113.665 174.670 ;
        RECT 116.135 174.660 116.425 174.670 ;
        RECT 112.385 174.170 112.715 174.340 ;
        RECT 113.410 173.865 113.580 174.660 ;
        RECT 115.145 174.170 115.475 174.340 ;
        RECT 116.170 173.865 116.340 174.660 ;
        RECT 106.935 173.690 107.225 173.700 ;
        RECT 113.330 173.445 113.630 173.865 ;
        RECT 116.090 173.445 116.390 173.865 ;
        RECT 113.395 172.640 113.665 172.665 ;
        RECT 105.980 172.395 106.310 172.565 ;
        RECT 110.000 171.980 110.170 172.310 ;
        RECT 113.395 172.285 113.945 172.640 ;
        RECT 114.160 172.285 114.460 172.645 ;
        RECT 44.730 171.005 45.100 171.650 ;
        RECT 44.775 170.995 45.065 171.005 ;
        RECT 45.895 171.000 46.440 171.645 ;
        RECT 50.815 171.460 52.610 171.630 ;
        RECT 45.940 170.990 46.440 171.000 ;
        RECT 46.270 170.195 46.440 170.990 ;
        RECT 50.675 170.570 50.845 171.185 ;
        RECT 51.635 170.855 51.805 171.460 ;
        RECT 50.675 170.400 51.650 170.570 ;
        RECT 46.270 170.140 48.110 170.195 ;
        RECT 46.140 170.025 48.110 170.140 ;
        RECT 46.140 169.780 46.440 170.025 ;
        RECT 48.115 169.210 48.285 169.540 ;
        RECT 48.980 169.210 49.150 169.540 ;
        RECT 49.845 169.210 50.015 169.540 ;
        RECT 50.710 169.210 50.880 170.400 ;
        RECT 51.575 169.210 51.745 169.540 ;
        RECT 52.440 169.210 52.610 171.460 ;
        RECT 93.625 170.885 93.995 171.530 ;
        RECT 93.670 170.875 93.960 170.885 ;
        RECT 94.790 170.880 95.335 171.525 ;
        RECT 99.710 171.340 101.505 171.510 ;
        RECT 107.790 171.390 108.000 171.425 ;
        RECT 110.015 171.400 110.295 171.525 ;
        RECT 110.820 171.400 111.140 171.445 ;
        RECT 113.550 171.430 113.720 172.285 ;
        RECT 114.290 171.920 114.460 172.285 ;
        RECT 116.090 172.225 116.390 172.645 ;
        RECT 114.290 171.750 115.475 171.920 ;
        RECT 114.290 171.435 114.460 171.750 ;
        RECT 112.795 171.420 113.085 171.430 ;
        RECT 113.375 171.420 113.720 171.430 ;
        RECT 113.960 171.425 114.460 171.435 ;
        RECT 116.170 171.430 116.340 172.225 ;
        RECT 188.910 171.460 190.705 171.630 ;
        RECT 94.835 170.870 95.335 170.880 ;
        RECT 95.165 170.075 95.335 170.870 ;
        RECT 99.570 170.450 99.740 171.065 ;
        RECT 100.530 170.735 100.700 171.340 ;
        RECT 99.570 170.280 100.545 170.450 ;
        RECT 95.165 170.020 97.005 170.075 ;
        RECT 95.035 169.905 97.005 170.020 ;
        RECT 95.035 169.660 95.335 169.905 ;
        RECT 53.305 169.210 53.475 169.540 ;
        RECT 54.170 169.210 54.340 169.540 ;
        RECT 97.010 169.090 97.180 169.420 ;
        RECT 97.875 169.090 98.045 169.420 ;
        RECT 98.740 169.090 98.910 169.420 ;
        RECT 99.605 169.090 99.775 170.280 ;
        RECT 100.470 169.090 100.640 169.420 ;
        RECT 101.335 169.090 101.505 171.340 ;
        RECT 107.740 170.980 108.045 171.390 ;
        RECT 110.015 171.230 111.140 171.400 ;
        RECT 110.015 171.105 110.295 171.230 ;
        RECT 110.820 171.185 111.140 171.230 ;
        RECT 107.790 170.965 108.000 170.980 ;
        RECT 112.750 170.775 113.120 171.420 ;
        RECT 113.330 171.260 113.720 171.420 ;
        RECT 113.330 170.815 113.700 171.260 ;
        RECT 113.330 170.775 113.695 170.815 ;
        RECT 113.915 170.780 114.460 171.425 ;
        RECT 116.135 171.420 116.425 171.430 ;
        RECT 116.090 170.815 116.460 171.420 ;
        RECT 116.090 170.775 116.455 170.815 ;
        RECT 113.330 169.835 113.695 169.875 ;
        RECT 116.090 169.835 116.455 169.875 ;
        RECT 102.200 169.090 102.370 169.420 ;
        RECT 103.065 169.090 103.235 169.420 ;
        RECT 45.310 168.560 45.610 168.980 ;
        RECT 50.620 168.780 50.955 168.950 ;
        RECT 45.390 168.360 45.560 168.560 ;
        RECT 45.390 168.185 48.160 168.360 ;
        RECT 45.390 167.765 45.560 168.185 ;
        RECT 47.985 167.780 48.160 168.185 ;
        RECT 50.700 168.080 50.875 168.780 ;
        RECT 94.205 168.440 94.505 168.860 ;
        RECT 99.515 168.660 99.850 168.830 ;
        RECT 94.285 168.240 94.455 168.440 ;
        RECT 50.700 167.910 51.950 168.080 ;
        RECT 94.285 168.065 97.055 168.240 ;
        RECT 45.355 167.755 45.645 167.765 ;
        RECT 45.310 167.150 45.680 167.755 ;
        RECT 94.285 167.645 94.455 168.065 ;
        RECT 96.880 167.660 97.055 168.065 ;
        RECT 99.595 167.960 99.770 168.660 ;
        RECT 106.890 168.260 107.260 169.450 ;
        RECT 110.840 168.520 111.185 169.765 ;
        RECT 113.330 169.230 113.700 169.835 ;
        RECT 116.090 169.230 116.460 169.835 ;
        RECT 113.375 169.220 113.665 169.230 ;
        RECT 116.135 169.220 116.425 169.230 ;
        RECT 112.385 168.730 112.715 168.900 ;
        RECT 113.410 168.425 113.580 169.220 ;
        RECT 115.145 168.730 115.475 168.900 ;
        RECT 116.170 168.425 116.340 169.220 ;
        RECT 122.145 169.175 122.475 169.975 ;
        RECT 122.985 169.175 123.315 169.975 ;
        RECT 123.825 169.175 124.155 169.975 ;
        RECT 124.665 169.175 124.995 169.975 ;
        RECT 127.935 169.175 128.265 169.975 ;
        RECT 128.775 169.175 129.105 169.975 ;
        RECT 129.615 169.175 129.945 169.975 ;
        RECT 130.455 169.175 130.785 169.975 ;
        RECT 187.180 169.210 187.350 169.540 ;
        RECT 188.045 169.210 188.215 169.540 ;
        RECT 188.910 169.210 189.080 171.460 ;
        RECT 189.715 170.855 189.885 171.460 ;
        RECT 190.675 170.570 190.845 171.185 ;
        RECT 189.870 170.400 190.845 170.570 ;
        RECT 195.080 171.000 195.625 171.645 ;
        RECT 196.420 171.005 196.790 171.650 ;
        RECT 195.080 170.990 195.580 171.000 ;
        RECT 196.455 170.995 196.745 171.005 ;
        RECT 189.775 169.210 189.945 169.540 ;
        RECT 190.640 169.210 190.810 170.400 ;
        RECT 195.080 170.195 195.250 170.990 ;
        RECT 193.410 170.140 195.250 170.195 ;
        RECT 193.410 170.025 195.380 170.140 ;
        RECT 195.080 169.780 195.380 170.025 ;
        RECT 191.505 169.210 191.675 169.540 ;
        RECT 192.370 169.210 192.540 169.540 ;
        RECT 193.235 169.210 193.405 169.540 ;
        RECT 121.550 169.005 125.520 169.175 ;
        RECT 106.935 168.250 107.225 168.260 ;
        RECT 113.330 168.005 113.630 168.425 ;
        RECT 116.090 168.005 116.390 168.425 ;
        RECT 121.550 168.415 121.895 169.005 ;
        RECT 122.145 168.585 125.000 168.835 ;
        RECT 125.200 168.415 125.520 169.005 ;
        RECT 121.550 168.225 125.520 168.415 ;
        RECT 127.340 169.005 131.310 169.175 ;
        RECT 127.340 168.415 127.685 169.005 ;
        RECT 127.935 168.585 130.790 168.835 ;
        RECT 130.990 168.415 131.310 169.005 ;
        RECT 190.565 168.780 190.900 168.950 ;
        RECT 127.340 168.225 131.310 168.415 ;
        RECT 99.595 167.790 100.845 167.960 ;
        RECT 122.145 167.765 122.475 168.225 ;
        RECT 122.985 167.765 123.315 168.225 ;
        RECT 123.825 167.765 124.155 168.225 ;
        RECT 124.665 167.765 124.995 168.225 ;
        RECT 127.935 167.765 128.265 168.225 ;
        RECT 128.775 167.765 129.105 168.225 ;
        RECT 129.615 167.765 129.945 168.225 ;
        RECT 130.455 167.765 130.785 168.225 ;
        RECT 190.645 168.080 190.820 168.780 ;
        RECT 195.910 168.560 196.210 168.980 ;
        RECT 195.960 168.360 196.130 168.560 ;
        RECT 189.570 167.910 190.820 168.080 ;
        RECT 193.360 168.185 196.130 168.360 ;
        RECT 193.360 167.780 193.535 168.185 ;
        RECT 195.960 167.765 196.130 168.185 ;
        RECT 195.875 167.755 196.165 167.765 ;
        RECT 94.250 167.635 94.540 167.645 ;
        RECT 45.310 167.110 45.675 167.150 ;
        RECT 48.115 167.010 48.285 167.340 ;
        RECT 48.980 167.010 49.150 167.340 ;
        RECT 49.845 167.010 50.015 167.345 ;
        RECT 50.710 167.010 50.880 167.340 ;
        RECT 51.575 167.010 51.745 167.340 ;
        RECT 52.440 167.010 52.610 167.340 ;
        RECT 53.305 167.010 53.475 167.340 ;
        RECT 54.170 167.010 54.340 167.340 ;
        RECT 94.205 167.030 94.575 167.635 ;
        RECT 94.205 166.990 94.570 167.030 ;
        RECT 97.010 166.890 97.180 167.220 ;
        RECT 97.875 166.890 98.045 167.220 ;
        RECT 98.740 166.890 98.910 167.225 ;
        RECT 99.605 166.890 99.775 167.220 ;
        RECT 100.470 166.890 100.640 167.220 ;
        RECT 101.335 166.890 101.505 167.220 ;
        RECT 102.200 166.890 102.370 167.220 ;
        RECT 103.065 166.890 103.235 167.220 ;
        RECT 113.395 167.200 113.665 167.225 ;
        RECT 105.980 166.955 106.310 167.125 ;
        RECT 110.000 166.540 110.170 166.870 ;
        RECT 113.395 166.845 113.945 167.200 ;
        RECT 114.160 166.845 114.460 167.205 ;
        RECT 94.205 166.050 94.570 166.090 ;
        RECT 94.205 165.445 94.575 166.050 ;
        RECT 97.010 165.860 97.180 166.190 ;
        RECT 97.875 165.860 98.045 166.190 ;
        RECT 98.740 165.855 98.910 166.190 ;
        RECT 99.605 165.860 99.775 166.190 ;
        RECT 100.470 165.860 100.640 166.190 ;
        RECT 101.335 165.860 101.505 166.190 ;
        RECT 102.200 165.860 102.370 166.190 ;
        RECT 103.065 165.860 103.235 166.190 ;
        RECT 107.790 165.950 108.000 165.985 ;
        RECT 110.015 165.960 110.295 166.085 ;
        RECT 110.820 165.960 111.140 166.005 ;
        RECT 113.550 165.990 113.720 166.845 ;
        RECT 114.290 166.480 114.460 166.845 ;
        RECT 116.090 166.785 116.390 167.205 ;
        RECT 122.145 166.795 122.475 167.255 ;
        RECT 122.985 166.795 123.315 167.255 ;
        RECT 123.825 166.795 124.155 167.255 ;
        RECT 124.665 166.795 124.995 167.255 ;
        RECT 187.180 167.010 187.350 167.340 ;
        RECT 188.045 167.010 188.215 167.340 ;
        RECT 188.910 167.010 189.080 167.340 ;
        RECT 189.775 167.010 189.945 167.340 ;
        RECT 190.640 167.010 190.810 167.340 ;
        RECT 191.505 167.010 191.675 167.345 ;
        RECT 192.370 167.010 192.540 167.340 ;
        RECT 193.235 167.010 193.405 167.340 ;
        RECT 195.840 167.150 196.210 167.755 ;
        RECT 195.845 167.110 196.210 167.150 ;
        RECT 114.290 166.310 115.475 166.480 ;
        RECT 114.290 165.995 114.460 166.310 ;
        RECT 112.795 165.980 113.085 165.990 ;
        RECT 113.375 165.980 113.720 165.990 ;
        RECT 113.960 165.985 114.460 165.995 ;
        RECT 116.170 165.990 116.340 166.785 ;
        RECT 121.550 166.605 125.520 166.795 ;
        RECT 121.550 166.015 121.895 166.605 ;
        RECT 122.145 166.185 125.000 166.435 ;
        RECT 125.200 166.015 125.520 166.605 ;
        RECT 127.935 166.185 130.790 166.435 ;
        RECT 107.740 165.540 108.045 165.950 ;
        RECT 110.015 165.790 111.140 165.960 ;
        RECT 110.015 165.665 110.295 165.790 ;
        RECT 110.820 165.745 111.140 165.790 ;
        RECT 107.790 165.525 108.000 165.540 ;
        RECT 94.250 165.435 94.540 165.445 ;
        RECT 94.285 165.015 94.455 165.435 ;
        RECT 96.880 165.015 97.055 165.420 ;
        RECT 112.750 165.335 113.120 165.980 ;
        RECT 113.330 165.820 113.720 165.980 ;
        RECT 113.330 165.375 113.700 165.820 ;
        RECT 113.330 165.335 113.695 165.375 ;
        RECT 113.915 165.340 114.460 165.985 ;
        RECT 116.135 165.980 116.425 165.990 ;
        RECT 116.090 165.375 116.460 165.980 ;
        RECT 121.550 165.845 125.520 166.015 ;
        RECT 116.090 165.335 116.455 165.375 ;
        RECT 94.285 164.840 97.055 165.015 ;
        RECT 99.595 165.120 100.845 165.290 ;
        RECT 94.285 164.640 94.455 164.840 ;
        RECT 94.205 164.220 94.505 164.640 ;
        RECT 99.595 164.420 99.770 165.120 ;
        RECT 122.145 165.045 122.475 165.845 ;
        RECT 122.985 165.045 123.315 165.845 ;
        RECT 123.825 165.045 124.155 165.845 ;
        RECT 124.665 165.045 124.995 165.845 ;
        RECT 99.515 164.250 99.850 164.420 ;
        RECT 113.330 164.395 113.695 164.435 ;
        RECT 116.090 164.395 116.455 164.435 ;
        RECT 97.010 163.660 97.180 163.990 ;
        RECT 97.875 163.660 98.045 163.990 ;
        RECT 98.740 163.660 98.910 163.990 ;
        RECT 95.035 163.175 95.335 163.420 ;
        RECT 95.035 163.060 97.005 163.175 ;
        RECT 95.165 163.005 97.005 163.060 ;
        RECT 95.165 162.210 95.335 163.005 ;
        RECT 99.605 162.800 99.775 163.990 ;
        RECT 100.470 163.660 100.640 163.990 ;
        RECT 93.670 162.195 93.960 162.205 ;
        RECT 94.835 162.200 95.335 162.210 ;
        RECT 93.625 161.550 93.995 162.195 ;
        RECT 94.790 161.555 95.335 162.200 ;
        RECT 99.570 162.630 100.545 162.800 ;
        RECT 99.570 162.015 99.740 162.630 ;
        RECT 100.530 161.740 100.700 162.345 ;
        RECT 101.335 161.740 101.505 163.990 ;
        RECT 102.200 163.660 102.370 163.990 ;
        RECT 103.065 163.660 103.235 163.990 ;
        RECT 106.890 162.820 107.260 164.010 ;
        RECT 110.110 162.820 110.480 164.010 ;
        RECT 113.330 163.790 113.700 164.395 ;
        RECT 116.090 163.790 116.460 164.395 ;
        RECT 113.375 163.780 113.665 163.790 ;
        RECT 116.135 163.780 116.425 163.790 ;
        RECT 112.385 163.290 112.715 163.460 ;
        RECT 113.410 162.985 113.580 163.780 ;
        RECT 115.145 163.290 115.475 163.460 ;
        RECT 116.170 162.985 116.340 163.780 ;
        RECT 106.935 162.810 107.225 162.820 ;
        RECT 110.155 162.810 110.445 162.820 ;
        RECT 113.330 162.565 113.630 162.985 ;
        RECT 116.090 162.565 116.390 162.985 ;
        RECT 99.710 161.570 101.505 161.740 ;
        RECT 113.395 161.760 113.665 161.785 ;
        RECT 105.980 161.515 106.310 161.685 ;
        RECT 109.200 161.515 109.530 161.685 ;
        RECT 113.395 161.405 113.945 161.760 ;
        RECT 114.160 161.405 114.460 161.765 ;
        RECT 113.550 160.550 113.720 161.405 ;
        RECT 114.290 161.040 114.460 161.405 ;
        RECT 116.090 161.345 116.390 161.765 ;
        RECT 114.290 160.870 115.475 161.040 ;
        RECT 114.290 160.555 114.460 160.870 ;
        RECT 107.790 160.510 108.000 160.545 ;
        RECT 111.010 160.510 111.220 160.545 ;
        RECT 112.795 160.540 113.085 160.550 ;
        RECT 113.375 160.540 113.720 160.550 ;
        RECT 113.960 160.545 114.460 160.555 ;
        RECT 116.170 160.550 116.340 161.345 ;
        RECT 107.740 160.100 108.045 160.510 ;
        RECT 110.960 160.100 111.265 160.510 ;
        RECT 107.790 160.085 108.000 160.100 ;
        RECT 111.010 160.085 111.220 160.100 ;
        RECT 112.750 159.895 113.120 160.540 ;
        RECT 113.330 160.380 113.720 160.540 ;
        RECT 113.330 159.935 113.700 160.380 ;
        RECT 113.330 159.895 113.695 159.935 ;
        RECT 113.915 159.900 114.460 160.545 ;
        RECT 116.135 160.540 116.425 160.550 ;
        RECT 116.090 159.935 116.460 160.540 ;
        RECT 116.090 159.895 116.455 159.935 ;
        RECT 109.925 143.815 110.155 144.195 ;
        RECT 130.225 143.815 130.455 144.195 ;
        RECT 109.575 143.370 109.905 143.540 ;
        RECT 110.175 143.370 111.235 143.540 ;
        RECT 129.145 143.370 130.205 143.540 ;
        RECT 130.475 143.370 130.805 143.540 ;
        RECT 110.195 143.120 110.365 143.370 ;
        RECT 109.655 142.950 110.365 143.120 ;
        RECT 130.015 143.120 130.185 143.370 ;
        RECT 130.015 142.950 130.725 143.120 ;
        RECT 109.655 142.680 109.825 142.950 ;
        RECT 130.555 142.680 130.725 142.950 ;
        RECT 109.575 142.510 109.905 142.680 ;
        RECT 110.175 142.510 111.900 142.680 ;
        RECT 128.480 142.510 130.205 142.680 ;
        RECT 130.475 142.510 130.805 142.680 ;
        RECT 109.925 141.900 110.155 142.280 ;
        RECT 111.045 141.950 111.215 142.280 ;
        RECT 129.165 141.950 129.335 142.280 ;
        RECT 130.225 141.900 130.455 142.280 ;
        RECT 3.755 131.945 3.925 133.010 ;
        RECT 4.655 131.945 4.825 133.010 ;
        RECT 112.550 132.915 112.880 133.295 ;
        RECT 113.710 132.915 114.040 133.295 ;
        RECT 114.870 132.915 115.200 133.295 ;
        RECT 125.240 132.915 125.570 133.295 ;
        RECT 126.400 132.915 126.730 133.295 ;
        RECT 127.560 132.915 127.890 133.295 ;
        RECT 128.720 132.915 129.050 133.295 ;
        RECT 111.660 132.265 111.990 132.565 ;
        RECT 112.820 132.265 113.150 132.565 ;
        RECT 113.980 132.265 114.310 132.565 ;
        RECT 115.140 132.265 115.470 132.565 ;
        RECT 124.970 132.265 125.300 132.565 ;
        RECT 126.130 132.265 126.460 132.565 ;
        RECT 127.290 132.265 127.620 132.565 ;
        RECT 128.450 132.265 128.780 132.565 ;
        RECT 3.675 131.775 4.005 131.945 ;
        RECT 4.205 131.775 4.905 131.945 ;
        RECT 111.740 131.915 111.910 132.265 ;
        RECT 112.900 131.915 113.070 132.265 ;
        RECT 114.060 131.915 114.230 132.265 ;
        RECT 115.220 131.915 115.390 132.265 ;
        RECT 116.830 132.230 117.330 132.245 ;
        RECT 123.110 132.230 123.610 132.245 ;
        RECT 116.315 132.060 119.265 132.230 ;
        RECT 116.315 132.055 117.330 132.060 ;
        RECT 116.830 131.960 117.330 132.055 ;
        RECT 111.660 131.865 111.990 131.915 ;
        RECT 112.820 131.865 113.150 131.915 ;
        RECT 113.980 131.865 114.310 131.915 ;
        RECT 115.140 131.865 115.470 131.915 ;
        RECT 3.100 131.340 3.470 131.600 ;
        RECT 4.205 131.165 4.375 131.775 ;
        RECT 111.660 131.685 112.435 131.865 ;
        RECT 112.820 131.685 113.595 131.865 ;
        RECT 113.980 131.685 114.755 131.865 ;
        RECT 115.140 131.685 115.915 131.865 ;
        RECT 111.660 131.625 111.990 131.685 ;
        RECT 112.820 131.625 113.150 131.685 ;
        RECT 113.980 131.625 114.310 131.685 ;
        RECT 115.140 131.625 115.470 131.685 ;
        RECT 5.075 131.340 5.445 131.600 ;
        RECT 3.675 130.995 4.375 131.165 ;
        RECT 4.575 130.995 4.905 131.165 ;
        RECT 4.205 130.610 4.375 130.995 ;
        RECT 9.135 130.955 9.305 131.285 ;
        RECT 19.285 130.955 19.455 131.285 ;
        RECT 30.435 130.955 30.605 131.285 ;
        RECT 37.135 130.955 37.305 131.285 ;
        RECT 67.885 130.955 68.055 131.285 ;
        RECT 75.825 130.955 75.995 131.285 ;
        RECT 98.935 130.955 99.105 131.285 ;
        RECT 106.585 130.955 106.755 131.285 ;
        RECT 112.560 131.065 112.890 131.445 ;
        RECT 113.720 131.065 114.050 131.445 ;
        RECT 114.880 131.065 115.210 131.445 ;
        RECT 117.480 130.890 117.650 131.525 ;
        RECT 118.995 131.130 119.265 132.060 ;
        RECT 121.175 132.060 124.125 132.230 ;
        RECT 121.175 131.130 121.445 132.060 ;
        RECT 123.110 132.055 124.125 132.060 ;
        RECT 123.110 131.960 123.610 132.055 ;
        RECT 125.050 131.915 125.220 132.265 ;
        RECT 126.210 131.915 126.380 132.265 ;
        RECT 127.370 131.915 127.540 132.265 ;
        RECT 128.530 131.915 128.700 132.265 ;
        RECT 235.555 131.945 235.725 133.010 ;
        RECT 236.455 131.945 236.625 133.010 ;
        RECT 124.970 131.865 125.300 131.915 ;
        RECT 126.130 131.865 126.460 131.915 ;
        RECT 127.290 131.865 127.620 131.915 ;
        RECT 128.450 131.865 128.780 131.915 ;
        RECT 124.525 131.685 125.300 131.865 ;
        RECT 125.685 131.685 126.460 131.865 ;
        RECT 126.845 131.685 127.620 131.865 ;
        RECT 128.005 131.685 128.780 131.865 ;
        RECT 235.475 131.775 236.175 131.945 ;
        RECT 236.375 131.775 236.705 131.945 ;
        RECT 124.970 131.625 125.300 131.685 ;
        RECT 126.130 131.625 126.460 131.685 ;
        RECT 127.290 131.625 127.620 131.685 ;
        RECT 128.450 131.625 128.780 131.685 ;
        RECT 119.030 131.120 119.260 131.130 ;
        RECT 119.060 131.100 119.230 131.120 ;
        RECT 121.210 131.100 121.380 131.130 ;
        RECT 119.690 130.885 119.860 130.945 ;
        RECT 3.675 130.440 4.005 130.610 ;
        RECT 4.205 130.440 4.905 130.610 ;
        RECT 3.100 130.005 3.470 130.265 ;
        RECT 4.205 129.830 4.375 130.440 ;
        RECT 5.075 130.005 5.445 130.265 ;
        RECT 3.675 129.660 4.375 129.830 ;
        RECT 4.575 129.660 4.905 129.830 ;
        RECT 8.425 129.480 9.065 130.745 ;
        RECT 9.375 130.230 9.545 130.745 ;
        RECT 19.045 130.230 19.215 130.745 ;
        RECT 9.375 130.060 10.315 130.230 ;
        RECT 18.275 130.060 19.215 130.230 ;
        RECT 9.375 129.480 9.545 130.060 ;
        RECT 19.045 129.480 19.215 130.060 ;
        RECT 19.525 129.480 20.165 130.745 ;
        RECT 29.725 129.480 30.365 130.745 ;
        RECT 30.675 130.230 30.845 130.745 ;
        RECT 36.895 130.230 37.065 130.745 ;
        RECT 30.675 130.060 31.615 130.230 ;
        RECT 36.125 130.060 37.065 130.230 ;
        RECT 30.675 129.480 30.845 130.060 ;
        RECT 36.895 129.480 37.065 130.060 ;
        RECT 37.375 129.480 38.015 130.745 ;
        RECT 67.175 129.480 67.815 130.745 ;
        RECT 68.125 130.230 68.295 130.745 ;
        RECT 75.585 130.230 75.755 130.745 ;
        RECT 68.125 130.060 69.065 130.230 ;
        RECT 74.815 130.060 75.755 130.230 ;
        RECT 68.125 129.480 68.295 130.060 ;
        RECT 75.585 129.480 75.755 130.060 ;
        RECT 76.065 129.480 76.705 130.745 ;
        RECT 98.225 129.480 98.865 130.745 ;
        RECT 99.175 130.230 99.345 130.745 ;
        RECT 106.345 130.230 106.515 130.745 ;
        RECT 99.175 130.060 100.115 130.230 ;
        RECT 105.575 130.060 106.515 130.230 ;
        RECT 99.175 129.480 99.345 130.060 ;
        RECT 106.345 129.480 106.515 130.060 ;
        RECT 106.825 129.480 107.465 130.745 ;
        RECT 118.735 130.715 119.860 130.885 ;
        RECT 118.815 129.490 118.985 130.715 ;
        RECT 119.690 130.615 119.860 130.715 ;
        RECT 120.580 130.885 120.750 130.945 ;
        RECT 122.790 130.890 122.960 131.525 ;
        RECT 125.230 131.065 125.560 131.445 ;
        RECT 126.390 131.065 126.720 131.445 ;
        RECT 127.550 131.065 127.880 131.445 ;
        RECT 128.710 131.065 129.040 131.445 ;
        RECT 234.935 131.340 235.305 131.600 ;
        RECT 133.625 130.955 133.795 131.285 ;
        RECT 141.275 130.955 141.445 131.285 ;
        RECT 164.385 130.955 164.555 131.285 ;
        RECT 172.325 130.955 172.495 131.285 ;
        RECT 203.075 130.955 203.245 131.285 ;
        RECT 209.775 130.955 209.945 131.285 ;
        RECT 220.925 130.955 221.095 131.285 ;
        RECT 231.075 130.955 231.245 131.285 ;
        RECT 236.005 131.165 236.175 131.775 ;
        RECT 236.910 131.340 237.280 131.600 ;
        RECT 235.475 130.995 235.805 131.165 ;
        RECT 236.005 130.995 236.705 131.165 ;
        RECT 120.580 130.715 121.705 130.885 ;
        RECT 120.580 130.615 120.750 130.715 ;
        RECT 120.050 130.160 120.385 130.340 ;
        RECT 121.455 129.490 121.625 130.715 ;
        RECT 9.135 128.990 9.305 129.320 ;
        RECT 19.285 128.990 19.455 129.320 ;
        RECT 30.435 128.990 30.605 129.320 ;
        RECT 37.135 128.990 37.305 129.320 ;
        RECT 67.885 128.990 68.055 129.320 ;
        RECT 75.825 128.990 75.995 129.320 ;
        RECT 98.935 128.990 99.105 129.320 ;
        RECT 106.585 128.990 106.755 129.320 ;
        RECT 118.430 129.220 119.400 129.490 ;
        RECT 121.040 129.220 122.010 129.490 ;
        RECT 132.915 129.480 133.555 130.745 ;
        RECT 133.865 130.230 134.035 130.745 ;
        RECT 141.035 130.230 141.205 130.745 ;
        RECT 133.865 130.060 134.805 130.230 ;
        RECT 140.265 130.060 141.205 130.230 ;
        RECT 133.865 129.480 134.035 130.060 ;
        RECT 141.035 129.480 141.205 130.060 ;
        RECT 141.515 129.480 142.155 130.745 ;
        RECT 163.675 129.480 164.315 130.745 ;
        RECT 164.625 130.230 164.795 130.745 ;
        RECT 172.085 130.230 172.255 130.745 ;
        RECT 164.625 130.060 165.565 130.230 ;
        RECT 171.315 130.060 172.255 130.230 ;
        RECT 164.625 129.480 164.795 130.060 ;
        RECT 172.085 129.480 172.255 130.060 ;
        RECT 172.565 129.480 173.205 130.745 ;
        RECT 202.365 129.480 203.005 130.745 ;
        RECT 203.315 130.230 203.485 130.745 ;
        RECT 209.535 130.230 209.705 130.745 ;
        RECT 203.315 130.060 204.255 130.230 ;
        RECT 208.765 130.060 209.705 130.230 ;
        RECT 203.315 129.480 203.485 130.060 ;
        RECT 209.535 129.480 209.705 130.060 ;
        RECT 210.015 129.480 210.655 130.745 ;
        RECT 220.215 129.480 220.855 130.745 ;
        RECT 221.165 130.230 221.335 130.745 ;
        RECT 230.835 130.230 231.005 130.745 ;
        RECT 221.165 130.060 222.105 130.230 ;
        RECT 230.065 130.060 231.005 130.230 ;
        RECT 221.165 129.480 221.335 130.060 ;
        RECT 230.835 129.480 231.005 130.060 ;
        RECT 231.315 129.480 231.955 130.745 ;
        RECT 236.005 130.610 236.175 130.995 ;
        RECT 235.475 130.440 236.175 130.610 ;
        RECT 236.375 130.440 236.705 130.610 ;
        RECT 234.935 130.005 235.305 130.265 ;
        RECT 236.005 129.830 236.175 130.440 ;
        RECT 236.910 130.005 237.280 130.265 ;
        RECT 235.475 129.660 235.805 129.830 ;
        RECT 236.005 129.660 236.705 129.830 ;
        RECT 117.100 128.710 118.260 129.210 ;
        RECT 122.180 128.710 123.340 129.210 ;
        RECT 133.625 128.990 133.795 129.320 ;
        RECT 141.275 128.990 141.445 129.320 ;
        RECT 164.385 128.990 164.555 129.320 ;
        RECT 172.325 128.990 172.495 129.320 ;
        RECT 203.075 128.990 203.245 129.320 ;
        RECT 209.775 128.990 209.945 129.320 ;
        RECT 220.925 128.990 221.095 129.320 ;
        RECT 231.075 128.990 231.245 129.320 ;
        RECT 119.380 128.705 121.065 128.710 ;
        RECT 118.485 128.435 121.980 128.705 ;
        RECT 120.050 128.025 120.390 128.435 ;
        RECT 119.970 127.760 120.470 128.025 ;
        RECT 119.650 126.195 119.820 126.830 ;
        RECT 120.620 126.195 120.790 126.830 ;
      LAYER mcon ;
        RECT 106.935 173.770 107.225 174.805 ;
        RECT 110.895 174.060 111.135 175.125 ;
        RECT 112.465 174.170 112.635 174.340 ;
        RECT 115.225 174.170 115.395 174.340 ;
        RECT 106.060 172.395 106.230 172.565 ;
        RECT 113.445 172.375 113.865 172.545 ;
        RECT 110.000 172.060 110.170 172.230 ;
        RECT 44.775 171.075 45.065 171.550 ;
        RECT 45.940 171.070 46.230 171.545 ;
        RECT 48.115 169.290 48.285 169.460 ;
        RECT 48.980 169.290 49.150 169.460 ;
        RECT 49.845 169.290 50.015 169.460 ;
        RECT 50.710 169.290 50.880 169.460 ;
        RECT 51.575 169.290 51.745 169.460 ;
        RECT 93.670 170.955 93.960 171.430 ;
        RECT 94.835 170.950 95.125 171.425 ;
        RECT 101.335 171.340 101.505 171.510 ;
        RECT 115.225 171.750 115.395 171.920 ;
        RECT 52.440 169.290 52.610 169.460 ;
        RECT 53.305 169.290 53.475 169.460 ;
        RECT 54.170 169.290 54.340 169.460 ;
        RECT 97.010 169.170 97.180 169.340 ;
        RECT 97.875 169.170 98.045 169.340 ;
        RECT 98.740 169.170 98.910 169.340 ;
        RECT 99.605 169.170 99.775 169.340 ;
        RECT 100.470 169.170 100.640 169.340 ;
        RECT 107.790 171.045 108.000 171.335 ;
        RECT 110.895 171.230 111.065 171.400 ;
        RECT 112.795 170.875 113.085 171.350 ;
        RECT 113.960 170.880 114.250 171.355 ;
        RECT 101.335 169.170 101.505 169.340 ;
        RECT 102.200 169.170 102.370 169.340 ;
        RECT 103.065 169.170 103.235 169.340 ;
        RECT 106.935 168.330 107.225 169.365 ;
        RECT 110.895 168.620 111.135 169.685 ;
        RECT 112.465 168.730 112.635 168.900 ;
        RECT 115.225 168.730 115.395 168.900 ;
        RECT 187.180 169.290 187.350 169.460 ;
        RECT 188.045 169.290 188.215 169.460 ;
        RECT 195.290 171.070 195.580 171.545 ;
        RECT 196.455 171.075 196.745 171.550 ;
        RECT 188.910 169.290 189.080 169.460 ;
        RECT 189.775 169.290 189.945 169.460 ;
        RECT 190.640 169.290 190.810 169.460 ;
        RECT 191.505 169.290 191.675 169.460 ;
        RECT 192.370 169.290 192.540 169.460 ;
        RECT 193.235 169.290 193.405 169.460 ;
        RECT 122.225 168.635 122.395 168.805 ;
        RECT 122.645 168.640 122.815 168.810 ;
        RECT 123.060 168.635 123.230 168.805 ;
        RECT 125.290 168.615 125.460 168.785 ;
        RECT 128.320 168.615 128.490 168.785 ;
        RECT 131.085 168.615 131.255 168.785 ;
        RECT 48.115 167.090 48.285 167.260 ;
        RECT 48.980 167.090 49.150 167.260 ;
        RECT 49.845 167.095 50.015 167.265 ;
        RECT 50.710 167.090 50.880 167.260 ;
        RECT 51.575 167.090 51.745 167.260 ;
        RECT 52.440 167.090 52.610 167.260 ;
        RECT 53.305 167.090 53.475 167.260 ;
        RECT 54.170 167.090 54.340 167.260 ;
        RECT 97.010 166.970 97.180 167.140 ;
        RECT 97.875 166.970 98.045 167.140 ;
        RECT 98.740 166.975 98.910 167.145 ;
        RECT 99.605 166.970 99.775 167.140 ;
        RECT 100.470 166.970 100.640 167.140 ;
        RECT 101.335 166.970 101.505 167.140 ;
        RECT 102.200 166.970 102.370 167.140 ;
        RECT 103.065 166.970 103.235 167.140 ;
        RECT 106.060 166.955 106.230 167.125 ;
        RECT 113.445 166.935 113.865 167.105 ;
        RECT 110.000 166.620 110.170 166.790 ;
        RECT 97.010 165.940 97.180 166.110 ;
        RECT 97.875 165.940 98.045 166.110 ;
        RECT 98.740 165.935 98.910 166.105 ;
        RECT 99.605 165.940 99.775 166.110 ;
        RECT 100.470 165.940 100.640 166.110 ;
        RECT 101.335 165.940 101.505 166.110 ;
        RECT 102.200 165.940 102.370 166.110 ;
        RECT 103.065 165.940 103.235 166.110 ;
        RECT 187.180 167.090 187.350 167.260 ;
        RECT 188.045 167.090 188.215 167.260 ;
        RECT 188.910 167.090 189.080 167.260 ;
        RECT 189.775 167.090 189.945 167.260 ;
        RECT 190.640 167.090 190.810 167.260 ;
        RECT 191.505 167.095 191.675 167.265 ;
        RECT 192.370 167.090 192.540 167.260 ;
        RECT 193.235 167.090 193.405 167.260 ;
        RECT 115.225 166.310 115.395 166.480 ;
        RECT 122.225 166.215 122.395 166.385 ;
        RECT 122.645 166.210 122.815 166.380 ;
        RECT 123.060 166.215 123.230 166.385 ;
        RECT 125.290 166.235 125.460 166.405 ;
        RECT 128.320 166.235 128.490 166.405 ;
        RECT 107.790 165.605 108.000 165.895 ;
        RECT 110.895 165.790 111.065 165.960 ;
        RECT 112.795 165.435 113.085 165.910 ;
        RECT 113.960 165.440 114.250 165.915 ;
        RECT 97.010 163.740 97.180 163.910 ;
        RECT 97.875 163.740 98.045 163.910 ;
        RECT 98.740 163.740 98.910 163.910 ;
        RECT 99.605 163.740 99.775 163.910 ;
        RECT 100.470 163.740 100.640 163.910 ;
        RECT 101.335 163.740 101.505 163.910 ;
        RECT 93.670 161.650 93.960 162.125 ;
        RECT 94.835 161.655 95.125 162.130 ;
        RECT 102.200 163.740 102.370 163.910 ;
        RECT 103.065 163.740 103.235 163.910 ;
        RECT 106.935 162.890 107.225 163.925 ;
        RECT 110.155 162.890 110.445 163.925 ;
        RECT 112.465 163.290 112.635 163.460 ;
        RECT 115.225 163.290 115.395 163.460 ;
        RECT 101.330 161.570 101.500 161.740 ;
        RECT 106.060 161.515 106.230 161.685 ;
        RECT 109.280 161.515 109.450 161.685 ;
        RECT 113.445 161.495 113.865 161.665 ;
        RECT 115.225 160.870 115.395 161.040 ;
        RECT 107.790 160.165 108.000 160.455 ;
        RECT 111.010 160.165 111.220 160.455 ;
        RECT 112.795 159.995 113.085 160.470 ;
        RECT 113.960 160.000 114.250 160.475 ;
        RECT 109.970 143.900 110.140 144.070 ;
        RECT 130.240 143.900 130.410 144.070 ;
        RECT 111.050 143.370 111.220 143.540 ;
        RECT 129.160 143.370 129.330 143.540 ;
        RECT 111.700 142.510 111.870 142.680 ;
        RECT 128.510 142.510 128.680 142.680 ;
        RECT 109.970 142.025 110.140 142.195 ;
        RECT 130.240 142.025 130.410 142.195 ;
        RECT 3.755 132.840 3.925 133.010 ;
        RECT 4.655 132.840 4.825 133.010 ;
        RECT 112.630 132.965 112.800 133.255 ;
        RECT 113.790 132.965 113.960 133.255 ;
        RECT 114.950 132.965 115.120 133.255 ;
        RECT 125.320 132.965 125.490 133.255 ;
        RECT 126.480 132.965 126.650 133.255 ;
        RECT 127.640 132.965 127.810 133.255 ;
        RECT 128.800 132.965 128.970 133.255 ;
        RECT 235.555 132.840 235.725 133.010 ;
        RECT 3.220 131.380 3.390 131.560 ;
        RECT 112.225 131.685 112.415 131.865 ;
        RECT 113.385 131.685 113.575 131.865 ;
        RECT 114.545 131.685 114.735 131.865 ;
        RECT 115.705 131.685 115.895 131.865 ;
        RECT 5.155 131.380 5.325 131.560 ;
        RECT 9.135 131.030 9.305 131.200 ;
        RECT 19.285 131.030 19.455 131.200 ;
        RECT 30.435 131.030 30.605 131.200 ;
        RECT 37.135 131.030 37.305 131.200 ;
        RECT 67.885 131.030 68.055 131.200 ;
        RECT 75.825 131.030 75.995 131.200 ;
        RECT 98.935 131.030 99.105 131.200 ;
        RECT 106.585 131.030 106.755 131.200 ;
        RECT 112.640 131.115 112.810 131.405 ;
        RECT 113.800 131.115 113.970 131.405 ;
        RECT 114.960 131.115 115.130 131.405 ;
        RECT 117.480 130.970 117.650 131.445 ;
        RECT 119.060 131.110 119.230 131.280 ;
        RECT 121.205 132.035 121.380 132.205 ;
        RECT 123.955 132.055 124.125 132.225 ;
        RECT 236.455 132.840 236.625 133.010 ;
        RECT 124.545 131.685 124.735 131.865 ;
        RECT 125.705 131.685 125.895 131.865 ;
        RECT 126.865 131.685 127.055 131.865 ;
        RECT 128.025 131.685 128.215 131.865 ;
        RECT 122.790 130.970 122.960 131.445 ;
        RECT 125.310 131.115 125.480 131.405 ;
        RECT 126.470 131.115 126.640 131.405 ;
        RECT 127.630 131.115 127.800 131.405 ;
        RECT 128.790 131.115 128.960 131.405 ;
        RECT 235.055 131.380 235.225 131.560 ;
        RECT 3.220 130.045 3.390 130.225 ;
        RECT 5.155 130.045 5.325 130.225 ;
        RECT 8.675 129.665 8.845 130.600 ;
        RECT 9.595 130.060 10.285 130.230 ;
        RECT 18.305 130.060 18.995 130.230 ;
        RECT 19.745 129.665 19.915 130.600 ;
        RECT 29.975 129.665 30.145 130.600 ;
        RECT 30.895 130.060 31.585 130.230 ;
        RECT 36.155 130.060 36.845 130.230 ;
        RECT 37.595 129.665 37.765 130.600 ;
        RECT 67.425 129.665 67.595 130.600 ;
        RECT 68.345 130.060 69.035 130.230 ;
        RECT 74.845 130.060 75.535 130.230 ;
        RECT 76.285 129.665 76.455 130.600 ;
        RECT 98.475 129.665 98.645 130.600 ;
        RECT 99.395 130.060 100.085 130.230 ;
        RECT 105.605 130.060 106.295 130.230 ;
        RECT 107.045 129.665 107.215 130.600 ;
        RECT 133.625 131.030 133.795 131.200 ;
        RECT 141.275 131.030 141.445 131.200 ;
        RECT 164.385 131.030 164.555 131.200 ;
        RECT 172.325 131.030 172.495 131.200 ;
        RECT 203.075 131.030 203.245 131.200 ;
        RECT 209.775 131.030 209.945 131.200 ;
        RECT 220.925 131.030 221.095 131.200 ;
        RECT 231.075 131.030 231.245 131.200 ;
        RECT 236.990 131.380 237.160 131.560 ;
        RECT 120.130 130.170 120.305 130.340 ;
        RECT 133.165 129.665 133.335 130.600 ;
        RECT 9.135 129.070 9.305 129.240 ;
        RECT 19.285 129.070 19.455 129.240 ;
        RECT 30.435 129.070 30.605 129.240 ;
        RECT 37.135 129.070 37.305 129.240 ;
        RECT 67.885 129.070 68.055 129.240 ;
        RECT 75.825 129.070 75.995 129.240 ;
        RECT 98.935 129.070 99.105 129.240 ;
        RECT 106.585 129.070 106.755 129.240 ;
        RECT 134.085 130.060 134.775 130.230 ;
        RECT 140.295 130.060 140.985 130.230 ;
        RECT 141.735 129.665 141.905 130.600 ;
        RECT 163.925 129.665 164.095 130.600 ;
        RECT 164.845 130.060 165.535 130.230 ;
        RECT 171.345 130.060 172.035 130.230 ;
        RECT 172.785 129.665 172.955 130.600 ;
        RECT 202.615 129.665 202.785 130.600 ;
        RECT 203.535 130.060 204.225 130.230 ;
        RECT 208.795 130.060 209.485 130.230 ;
        RECT 210.235 129.665 210.405 130.600 ;
        RECT 220.465 129.665 220.635 130.600 ;
        RECT 221.385 130.060 222.075 130.230 ;
        RECT 230.095 130.060 230.785 130.230 ;
        RECT 231.535 129.665 231.705 130.600 ;
        RECT 235.055 130.045 235.225 130.225 ;
        RECT 236.990 130.045 237.160 130.225 ;
        RECT 117.180 128.760 118.180 129.150 ;
        RECT 122.260 128.770 123.260 129.160 ;
        RECT 133.625 129.070 133.795 129.240 ;
        RECT 141.275 129.070 141.445 129.240 ;
        RECT 164.385 129.070 164.555 129.240 ;
        RECT 172.325 129.070 172.495 129.240 ;
        RECT 203.075 129.070 203.245 129.240 ;
        RECT 209.775 129.070 209.945 129.240 ;
        RECT 220.925 129.070 221.095 129.240 ;
        RECT 231.075 129.070 231.245 129.240 ;
        RECT 119.650 126.275 119.820 126.750 ;
        RECT 120.620 126.275 120.790 126.750 ;
      LAYER met1 ;
        RECT 106.905 174.035 107.255 174.865 ;
        RECT 110.865 174.370 111.165 175.185 ;
        RECT 112.400 174.385 112.715 174.390 ;
        RECT 112.390 174.370 112.715 174.385 ;
        RECT 110.865 174.130 112.715 174.370 ;
        RECT 107.810 174.035 108.070 174.095 ;
        RECT 106.905 173.865 108.070 174.035 ;
        RECT 110.865 174.000 111.165 174.130 ;
        RECT 112.390 174.125 112.715 174.130 ;
        RECT 112.400 174.120 112.715 174.125 ;
        RECT 113.365 174.360 113.620 174.725 ;
        RECT 115.160 174.385 115.475 174.390 ;
        RECT 115.150 174.360 115.475 174.385 ;
        RECT 113.365 174.145 115.475 174.360 ;
        RECT 106.905 173.740 107.255 173.865 ;
        RECT 107.810 173.775 108.070 173.865 ;
        RECT 113.365 173.805 113.620 174.145 ;
        RECT 115.150 174.125 115.475 174.145 ;
        RECT 115.160 174.120 115.475 174.125 ;
        RECT 116.125 174.360 116.380 174.725 ;
        RECT 123.230 174.360 123.490 174.420 ;
        RECT 116.125 174.140 123.490 174.360 ;
        RECT 116.125 173.805 116.380 174.140 ;
        RECT 123.230 174.100 123.490 174.140 ;
        RECT 106.935 173.710 107.225 173.740 ;
        RECT 105.995 172.610 106.310 172.615 ;
        RECT 105.985 172.350 106.310 172.610 ;
        RECT 105.995 172.345 106.310 172.350 ;
        RECT 113.385 172.330 113.925 172.590 ;
        RECT 109.950 171.980 110.220 172.310 ;
        RECT 44.740 171.415 45.120 171.615 ;
        RECT 45.900 171.415 46.280 171.605 ;
        RECT 44.740 171.165 46.280 171.415 ;
        RECT 44.740 171.015 45.120 171.165 ;
        RECT 45.900 171.010 46.280 171.165 ;
        RECT 93.635 171.295 94.015 171.495 ;
        RECT 94.795 171.295 95.175 171.485 ;
        RECT 93.635 171.045 95.175 171.295 ;
        RECT 101.265 171.275 101.590 171.570 ;
        RECT 107.790 171.365 108.000 171.395 ;
        RECT 107.760 171.345 108.030 171.365 ;
        RECT 109.990 171.345 110.160 171.980 ;
        RECT 115.160 171.965 115.475 171.970 ;
        RECT 115.150 171.705 115.475 171.965 ;
        RECT 115.160 171.700 115.475 171.705 ;
        RECT 116.125 171.925 116.380 172.285 ;
        RECT 122.015 171.925 122.275 171.980 ;
        RECT 116.125 171.705 122.275 171.925 ;
        RECT 110.835 171.445 111.125 171.460 ;
        RECT 93.635 170.895 94.015 171.045 ;
        RECT 94.795 170.890 95.175 171.045 ;
        RECT 107.760 171.175 110.160 171.345 ;
        RECT 110.820 171.185 111.140 171.445 ;
        RECT 112.760 171.260 113.140 171.410 ;
        RECT 113.920 171.260 114.300 171.415 ;
        RECT 116.125 171.365 116.380 171.705 ;
        RECT 122.015 171.660 122.275 171.705 ;
        RECT 195.240 171.415 195.620 171.605 ;
        RECT 196.400 171.415 196.780 171.615 ;
        RECT 107.760 171.015 108.030 171.175 ;
        RECT 110.835 171.170 111.125 171.185 ;
        RECT 107.790 170.985 108.000 171.015 ;
        RECT 112.760 171.010 114.300 171.260 ;
        RECT 195.240 171.165 196.780 171.415 ;
        RECT 195.240 171.010 195.620 171.165 ;
        RECT 196.400 171.015 196.780 171.165 ;
        RECT 112.760 170.810 113.140 171.010 ;
        RECT 113.920 170.820 114.300 171.010 ;
        RECT 48.055 169.415 48.360 169.500 ;
        RECT 48.920 169.415 49.225 169.500 ;
        RECT 49.775 169.415 50.095 169.500 ;
        RECT 50.650 169.415 50.955 169.500 ;
        RECT 51.515 169.415 51.820 169.500 ;
        RECT 52.365 169.415 52.685 169.500 ;
        RECT 53.245 169.415 53.550 169.500 ;
        RECT 54.110 169.415 54.415 169.500 ;
        RECT 48.055 169.260 50.955 169.415 ;
        RECT 51.510 169.260 54.830 169.415 ;
        RECT 96.950 169.295 97.255 169.380 ;
        RECT 97.815 169.295 98.120 169.380 ;
        RECT 98.670 169.295 98.990 169.380 ;
        RECT 99.545 169.295 99.850 169.380 ;
        RECT 100.410 169.295 100.715 169.380 ;
        RECT 101.260 169.295 101.580 169.380 ;
        RECT 102.140 169.295 102.445 169.380 ;
        RECT 103.005 169.295 103.310 169.380 ;
        RECT 49.775 169.235 50.095 169.260 ;
        RECT 52.365 169.240 52.685 169.260 ;
        RECT 96.950 169.140 99.850 169.295 ;
        RECT 100.405 169.140 103.725 169.295 ;
        RECT 98.670 169.115 98.990 169.140 ;
        RECT 101.260 169.120 101.580 169.140 ;
        RECT 45.345 167.700 45.600 168.620 ;
        RECT 106.905 168.595 107.255 169.425 ;
        RECT 110.865 168.930 111.165 169.745 ;
        RECT 187.105 169.415 187.410 169.500 ;
        RECT 187.970 169.415 188.275 169.500 ;
        RECT 188.835 169.415 189.155 169.500 ;
        RECT 189.700 169.415 190.005 169.500 ;
        RECT 190.565 169.415 190.870 169.500 ;
        RECT 191.425 169.415 191.745 169.500 ;
        RECT 192.295 169.415 192.600 169.500 ;
        RECT 193.160 169.415 193.465 169.500 ;
        RECT 112.400 168.945 112.715 168.950 ;
        RECT 112.390 168.930 112.715 168.945 ;
        RECT 110.865 168.690 112.715 168.930 ;
        RECT 107.810 168.595 108.070 168.655 ;
        RECT 94.240 167.580 94.495 168.500 ;
        RECT 106.905 168.425 108.070 168.595 ;
        RECT 110.865 168.560 111.165 168.690 ;
        RECT 112.390 168.685 112.715 168.690 ;
        RECT 112.400 168.680 112.715 168.685 ;
        RECT 113.365 168.920 113.620 169.285 ;
        RECT 115.160 168.945 115.475 168.950 ;
        RECT 115.150 168.920 115.475 168.945 ;
        RECT 113.365 168.705 115.475 168.920 ;
        RECT 106.905 168.300 107.255 168.425 ;
        RECT 107.810 168.335 108.070 168.425 ;
        RECT 113.365 168.365 113.620 168.705 ;
        RECT 115.150 168.685 115.475 168.705 ;
        RECT 115.160 168.680 115.475 168.685 ;
        RECT 116.125 168.825 116.380 169.285 ;
        RECT 186.690 169.260 190.010 169.415 ;
        RECT 190.565 169.260 193.465 169.415 ;
        RECT 188.835 169.240 189.155 169.260 ;
        RECT 191.425 169.235 191.745 169.260 ;
        RECT 121.050 168.860 121.310 168.875 ;
        RECT 121.050 168.825 123.555 168.860 ;
        RECT 116.125 168.605 123.555 168.825 ;
        RECT 116.125 168.365 116.380 168.605 ;
        RECT 121.050 168.570 123.555 168.605 ;
        RECT 121.050 168.555 121.310 168.570 ;
        RECT 125.210 168.560 128.660 168.835 ;
        RECT 130.920 168.535 132.250 168.855 ;
        RECT 106.935 168.270 107.225 168.300 ;
        RECT 195.920 167.700 196.175 168.620 ;
        RECT 48.055 167.215 48.360 167.300 ;
        RECT 48.920 167.215 49.225 167.300 ;
        RECT 49.775 167.215 50.095 167.305 ;
        RECT 50.650 167.215 50.955 167.300 ;
        RECT 51.515 167.215 51.820 167.300 ;
        RECT 52.375 167.215 52.695 167.300 ;
        RECT 53.245 167.215 53.550 167.300 ;
        RECT 54.110 167.215 54.415 167.300 ;
        RECT 48.055 167.060 50.955 167.215 ;
        RECT 51.510 167.060 54.415 167.215 ;
        RECT 187.105 167.215 187.410 167.300 ;
        RECT 187.970 167.215 188.275 167.300 ;
        RECT 188.825 167.215 189.145 167.300 ;
        RECT 189.700 167.215 190.005 167.300 ;
        RECT 190.565 167.215 190.870 167.300 ;
        RECT 191.425 167.215 191.745 167.305 ;
        RECT 192.295 167.215 192.600 167.300 ;
        RECT 193.160 167.215 193.465 167.300 ;
        RECT 96.950 167.095 97.255 167.180 ;
        RECT 97.815 167.095 98.120 167.180 ;
        RECT 98.670 167.095 98.990 167.185 ;
        RECT 99.545 167.095 99.850 167.180 ;
        RECT 100.410 167.095 100.715 167.180 ;
        RECT 101.270 167.095 101.590 167.180 ;
        RECT 102.140 167.095 102.445 167.180 ;
        RECT 103.005 167.095 103.310 167.180 ;
        RECT 105.995 167.170 106.310 167.175 ;
        RECT 49.775 167.040 50.095 167.060 ;
        RECT 52.375 167.040 52.695 167.060 ;
        RECT 96.950 166.940 99.850 167.095 ;
        RECT 100.405 166.940 103.310 167.095 ;
        RECT 98.670 166.920 98.990 166.940 ;
        RECT 101.270 166.920 101.590 166.940 ;
        RECT 105.985 166.910 106.310 167.170 ;
        RECT 105.995 166.905 106.310 166.910 ;
        RECT 113.385 166.890 113.925 167.150 ;
        RECT 187.105 167.060 190.010 167.215 ;
        RECT 190.565 167.060 193.465 167.215 ;
        RECT 188.825 167.040 189.145 167.060 ;
        RECT 191.425 167.040 191.745 167.060 ;
        RECT 109.950 166.540 110.220 166.870 ;
        RECT 98.670 166.140 98.990 166.160 ;
        RECT 101.270 166.140 101.590 166.160 ;
        RECT 96.950 165.985 99.850 166.140 ;
        RECT 100.405 165.985 103.310 166.140 ;
        RECT 96.950 165.900 97.255 165.985 ;
        RECT 97.815 165.900 98.120 165.985 ;
        RECT 98.670 165.895 98.990 165.985 ;
        RECT 99.545 165.900 99.850 165.985 ;
        RECT 100.410 165.900 100.715 165.985 ;
        RECT 101.270 165.900 101.590 165.985 ;
        RECT 102.140 165.900 102.445 165.985 ;
        RECT 103.005 165.900 103.310 165.985 ;
        RECT 107.790 165.925 108.000 165.955 ;
        RECT 107.760 165.905 108.030 165.925 ;
        RECT 109.990 165.905 110.160 166.540 ;
        RECT 115.160 166.525 115.475 166.530 ;
        RECT 115.150 166.265 115.475 166.525 ;
        RECT 115.160 166.260 115.475 166.265 ;
        RECT 116.125 166.485 116.380 166.845 ;
        RECT 118.785 166.485 119.050 166.515 ;
        RECT 116.125 166.455 119.050 166.485 ;
        RECT 116.125 166.450 121.500 166.455 ;
        RECT 116.125 166.265 123.555 166.450 ;
        RECT 110.835 166.005 111.125 166.020 ;
        RECT 107.760 165.735 110.160 165.905 ;
        RECT 110.820 165.745 111.140 166.005 ;
        RECT 112.760 165.820 113.140 165.970 ;
        RECT 113.920 165.820 114.300 165.975 ;
        RECT 116.125 165.925 116.380 166.265 ;
        RECT 118.785 166.195 123.555 166.265 ;
        RECT 118.945 166.185 123.555 166.195 ;
        RECT 125.210 166.185 128.660 166.460 ;
        RECT 121.200 166.160 123.555 166.185 ;
        RECT 107.760 165.575 108.030 165.735 ;
        RECT 110.835 165.730 111.125 165.745 ;
        RECT 107.790 165.545 108.000 165.575 ;
        RECT 112.760 165.570 114.300 165.820 ;
        RECT 94.240 164.580 94.495 165.500 ;
        RECT 112.760 165.370 113.140 165.570 ;
        RECT 113.920 165.380 114.300 165.570 ;
        RECT 98.670 163.940 98.990 163.965 ;
        RECT 101.260 163.940 101.580 163.960 ;
        RECT 96.950 163.785 99.850 163.940 ;
        RECT 100.405 163.785 103.725 163.940 ;
        RECT 96.950 163.700 97.255 163.785 ;
        RECT 97.815 163.700 98.120 163.785 ;
        RECT 98.670 163.700 98.990 163.785 ;
        RECT 99.545 163.700 99.850 163.785 ;
        RECT 100.410 163.700 100.715 163.785 ;
        RECT 101.260 163.700 101.580 163.785 ;
        RECT 102.140 163.700 102.445 163.785 ;
        RECT 103.005 163.700 103.310 163.785 ;
        RECT 106.905 163.155 107.255 163.985 ;
        RECT 110.125 163.815 112.635 163.985 ;
        RECT 107.810 163.155 108.070 163.215 ;
        RECT 106.905 162.985 108.070 163.155 ;
        RECT 106.905 162.860 107.255 162.985 ;
        RECT 107.810 162.895 108.070 162.985 ;
        RECT 110.125 163.155 110.475 163.815 ;
        RECT 112.465 163.510 112.635 163.815 ;
        RECT 112.400 163.505 112.715 163.510 ;
        RECT 112.390 163.245 112.715 163.505 ;
        RECT 112.400 163.240 112.715 163.245 ;
        RECT 113.365 163.480 113.620 163.845 ;
        RECT 115.160 163.505 115.475 163.510 ;
        RECT 115.150 163.480 115.475 163.505 ;
        RECT 113.365 163.265 115.475 163.480 ;
        RECT 111.030 163.155 111.290 163.215 ;
        RECT 110.125 162.985 111.290 163.155 ;
        RECT 110.125 162.860 110.475 162.985 ;
        RECT 111.030 162.895 111.290 162.985 ;
        RECT 113.365 162.925 113.620 163.265 ;
        RECT 115.150 163.245 115.475 163.265 ;
        RECT 115.160 163.240 115.475 163.245 ;
        RECT 116.125 163.360 116.380 163.845 ;
        RECT 117.965 163.360 118.230 163.390 ;
        RECT 116.125 163.075 118.230 163.360 ;
        RECT 116.125 162.925 116.380 163.075 ;
        RECT 117.965 163.045 118.230 163.075 ;
        RECT 106.935 162.830 107.225 162.860 ;
        RECT 110.155 162.830 110.445 162.860 ;
        RECT 93.635 162.035 94.015 162.185 ;
        RECT 94.795 162.035 95.175 162.190 ;
        RECT 93.635 161.785 95.175 162.035 ;
        RECT 93.635 161.585 94.015 161.785 ;
        RECT 94.795 161.595 95.175 161.785 ;
        RECT 101.265 161.780 101.580 161.790 ;
        RECT 101.255 161.520 101.580 161.780 ;
        RECT 105.995 161.730 106.310 161.735 ;
        RECT 109.215 161.730 109.530 161.735 ;
        RECT 101.265 161.515 101.580 161.520 ;
        RECT 105.985 161.470 106.310 161.730 ;
        RECT 109.205 161.470 109.530 161.730 ;
        RECT 105.995 161.465 106.310 161.470 ;
        RECT 109.215 161.465 109.530 161.470 ;
        RECT 113.385 161.450 113.925 161.710 ;
        RECT 116.125 161.380 116.380 161.405 ;
        RECT 115.160 161.085 115.475 161.090 ;
        RECT 115.150 160.825 115.475 161.085 ;
        RECT 115.160 160.820 115.475 160.825 ;
        RECT 107.790 160.485 108.000 160.515 ;
        RECT 111.010 160.485 111.220 160.515 ;
        RECT 107.760 160.135 108.030 160.485 ;
        RECT 110.980 160.135 111.250 160.485 ;
        RECT 112.760 160.380 113.140 160.530 ;
        RECT 113.920 160.380 114.300 160.535 ;
        RECT 116.125 160.515 116.385 161.380 ;
        RECT 116.125 160.485 116.380 160.515 ;
        RECT 107.790 160.105 108.000 160.135 ;
        RECT 111.010 160.105 111.220 160.135 ;
        RECT 112.760 160.130 114.300 160.380 ;
        RECT 112.760 159.930 113.140 160.130 ;
        RECT 113.920 159.940 114.300 160.130 ;
        RECT 4.620 151.750 4.880 151.825 ;
        RECT 191.430 151.750 191.750 151.780 ;
        RECT 235.500 151.750 235.760 151.825 ;
        RECT 4.615 151.550 235.765 151.750 ;
        RECT 4.620 151.505 4.880 151.550 ;
        RECT 191.430 151.520 191.750 151.550 ;
        RECT 235.500 151.505 235.760 151.550 ;
        RECT 3.710 151.150 3.970 151.200 ;
        RECT 188.865 151.150 189.125 151.210 ;
        RECT 236.410 151.150 236.670 151.200 ;
        RECT 3.705 150.950 236.675 151.150 ;
        RECT 3.710 150.880 3.970 150.950 ;
        RECT 188.865 150.890 189.125 150.950 ;
        RECT 236.410 150.880 236.670 150.950 ;
        RECT 19.235 150.550 19.495 150.595 ;
        RECT 37.115 150.550 37.375 150.580 ;
        RECT 75.780 150.550 76.040 150.605 ;
        RECT 106.525 150.550 106.785 150.620 ;
        RECT 122.010 150.550 122.280 150.630 ;
        RECT 133.595 150.550 133.855 150.620 ;
        RECT 164.340 150.550 164.600 150.605 ;
        RECT 203.005 150.550 203.265 150.580 ;
        RECT 220.885 150.550 221.145 150.595 ;
        RECT 19.225 150.350 221.155 150.550 ;
        RECT 19.235 150.275 19.495 150.350 ;
        RECT 37.115 150.260 37.375 150.350 ;
        RECT 75.780 150.285 76.040 150.350 ;
        RECT 106.525 150.300 106.785 150.350 ;
        RECT 122.010 150.310 122.280 150.350 ;
        RECT 133.595 150.300 133.855 150.350 ;
        RECT 164.340 150.285 164.600 150.350 ;
        RECT 203.005 150.260 203.265 150.350 ;
        RECT 220.885 150.275 221.145 150.350 ;
        RECT 18.800 149.950 19.060 149.995 ;
        RECT 36.725 149.950 36.985 150.000 ;
        RECT 75.390 149.950 75.650 150.035 ;
        RECT 106.195 149.950 106.455 149.970 ;
        RECT 123.225 149.950 123.485 150.015 ;
        RECT 133.925 149.950 134.185 149.970 ;
        RECT 164.730 149.950 164.990 150.035 ;
        RECT 203.395 149.950 203.655 150.000 ;
        RECT 221.320 149.950 221.580 149.995 ;
        RECT 18.795 149.750 221.585 149.950 ;
        RECT 18.800 149.675 19.060 149.750 ;
        RECT 36.725 149.680 36.985 149.750 ;
        RECT 75.390 149.715 75.650 149.750 ;
        RECT 106.195 149.650 106.455 149.750 ;
        RECT 123.225 149.695 123.485 149.750 ;
        RECT 133.925 149.650 134.185 149.750 ;
        RECT 164.730 149.715 164.990 149.750 ;
        RECT 203.395 149.680 203.655 149.750 ;
        RECT 221.320 149.675 221.580 149.750 ;
        RECT 9.090 149.350 9.350 149.415 ;
        RECT 30.395 149.350 30.655 149.415 ;
        RECT 67.855 149.350 68.115 149.390 ;
        RECT 98.900 149.350 99.160 149.380 ;
        RECT 118.790 149.350 119.050 149.430 ;
        RECT 141.220 149.350 141.480 149.380 ;
        RECT 172.265 149.350 172.525 149.390 ;
        RECT 209.725 149.350 209.985 149.415 ;
        RECT 231.030 149.350 231.290 149.415 ;
        RECT 9.085 149.150 231.295 149.350 ;
        RECT 9.090 149.095 9.350 149.150 ;
        RECT 30.395 149.095 30.655 149.150 ;
        RECT 67.855 149.070 68.115 149.150 ;
        RECT 98.900 149.060 99.160 149.150 ;
        RECT 118.790 149.110 119.050 149.150 ;
        RECT 141.220 149.060 141.480 149.150 ;
        RECT 172.265 149.070 172.525 149.150 ;
        RECT 209.725 149.095 209.985 149.150 ;
        RECT 231.030 149.095 231.290 149.150 ;
        RECT 9.520 148.750 9.780 148.835 ;
        RECT 30.815 148.750 31.075 148.800 ;
        RECT 68.285 148.750 68.545 148.830 ;
        RECT 99.335 148.750 99.595 148.825 ;
        RECT 121.045 148.750 121.305 148.810 ;
        RECT 140.785 148.750 141.045 148.825 ;
        RECT 171.835 148.750 172.095 148.830 ;
        RECT 209.305 148.750 209.565 148.800 ;
        RECT 230.600 148.750 230.860 148.835 ;
        RECT 9.515 148.550 230.865 148.750 ;
        RECT 9.520 148.515 9.780 148.550 ;
        RECT 30.815 148.480 31.075 148.550 ;
        RECT 68.285 148.510 68.545 148.550 ;
        RECT 99.335 148.505 99.595 148.550 ;
        RECT 121.045 148.490 121.305 148.550 ;
        RECT 140.785 148.505 141.045 148.550 ;
        RECT 171.835 148.510 172.095 148.550 ;
        RECT 209.305 148.480 209.565 148.550 ;
        RECT 230.600 148.515 230.860 148.550 ;
        RECT 109.900 143.840 110.195 144.150 ;
        RECT 130.185 143.840 130.480 144.150 ;
        RECT 109.970 142.255 110.140 143.840 ;
        RECT 110.995 143.585 111.295 143.605 ;
        RECT 110.985 143.555 111.305 143.585 ;
        RECT 117.965 143.555 118.225 143.595 ;
        RECT 129.085 143.585 129.385 143.605 ;
        RECT 129.075 143.555 129.395 143.585 ;
        RECT 110.985 143.330 129.395 143.555 ;
        RECT 110.985 143.325 111.305 143.330 ;
        RECT 110.995 143.300 111.295 143.325 ;
        RECT 117.965 143.270 118.225 143.330 ;
        RECT 129.075 143.325 129.395 143.330 ;
        RECT 129.085 143.300 129.385 143.325 ;
        RECT 111.645 142.725 111.945 142.740 ;
        RECT 111.635 142.705 111.955 142.725 ;
        RECT 116.120 142.705 116.380 142.750 ;
        RECT 128.435 142.725 128.735 142.740 ;
        RECT 128.425 142.705 128.745 142.725 ;
        RECT 111.395 142.480 128.965 142.705 ;
        RECT 111.635 142.465 111.955 142.480 ;
        RECT 111.645 142.440 111.945 142.465 ;
        RECT 116.120 142.430 116.380 142.480 ;
        RECT 128.425 142.465 128.745 142.480 ;
        RECT 128.435 142.440 128.735 142.465 ;
        RECT 130.240 142.255 130.410 143.840 ;
        RECT 109.910 141.965 110.200 142.255 ;
        RECT 130.180 141.965 130.470 142.255 ;
        RECT 109.940 140.315 110.150 141.965 ;
        RECT 130.230 140.315 130.440 141.965 ;
        RECT 109.530 138.755 111.125 140.315 ;
        RECT 129.255 138.755 130.850 140.315 ;
        RECT 3.680 132.760 4.000 133.100 ;
        RECT 4.580 132.760 4.900 133.100 ;
        RECT 112.570 132.915 112.860 133.295 ;
        RECT 113.730 132.915 114.020 133.295 ;
        RECT 114.890 132.915 115.180 133.295 ;
        RECT 125.260 132.915 125.550 133.295 ;
        RECT 126.420 132.915 126.710 133.295 ;
        RECT 127.580 132.915 127.870 133.295 ;
        RECT 128.740 132.915 129.030 133.295 ;
        RECT 112.580 131.935 112.750 132.915 ;
        RECT 113.740 131.935 113.910 132.915 ;
        RECT 114.900 131.935 115.070 132.915 ;
        RECT 3.145 131.560 3.465 131.600 ;
        RECT 3.145 131.380 3.470 131.560 ;
        RECT 3.145 131.340 3.465 131.380 ;
        RECT 4.545 131.310 4.805 131.630 ;
        RECT 112.155 131.615 112.750 131.935 ;
        RECT 113.315 131.615 113.910 131.935 ;
        RECT 114.475 131.615 115.070 131.935 ;
        RECT 115.635 132.015 116.545 132.285 ;
        RECT 121.175 132.205 121.410 132.235 ;
        RECT 121.145 132.195 121.440 132.205 ;
        RECT 117.480 132.045 121.440 132.195 ;
        RECT 115.635 131.615 115.965 132.015 ;
        RECT 5.080 131.340 5.400 131.600 ;
        RECT 112.580 131.445 112.750 131.615 ;
        RECT 113.740 131.445 113.910 131.615 ;
        RECT 114.900 131.445 115.070 131.615 ;
        RECT 117.480 131.475 117.650 132.045 ;
        RECT 121.145 132.035 121.440 132.045 ;
        RECT 121.175 132.005 121.410 132.035 ;
        RECT 123.895 132.005 124.805 132.275 ;
        RECT 124.475 131.615 124.805 132.005 ;
        RECT 125.370 131.935 125.540 132.915 ;
        RECT 126.530 131.935 126.700 132.915 ;
        RECT 127.690 131.935 127.860 132.915 ;
        RECT 125.370 131.615 125.965 131.935 ;
        RECT 126.530 131.615 127.125 131.935 ;
        RECT 127.690 131.615 128.285 131.935 ;
        RECT 122.790 131.475 122.960 131.505 ;
        RECT 9.090 131.270 9.350 131.275 ;
        RECT 19.240 131.270 19.500 131.275 ;
        RECT 30.390 131.270 30.650 131.275 ;
        RECT 37.090 131.270 37.350 131.275 ;
        RECT 67.840 131.270 68.100 131.275 ;
        RECT 75.780 131.270 76.040 131.275 ;
        RECT 98.890 131.270 99.150 131.275 ;
        RECT 106.540 131.270 106.800 131.275 ;
        RECT 9.065 130.950 9.375 131.270 ;
        RECT 19.215 130.950 19.525 131.270 ;
        RECT 30.365 130.950 30.675 131.270 ;
        RECT 37.065 130.950 37.375 131.270 ;
        RECT 67.815 130.950 68.125 131.270 ;
        RECT 75.755 130.950 76.065 131.270 ;
        RECT 98.865 130.950 99.175 131.270 ;
        RECT 106.515 130.950 106.825 131.270 ;
        RECT 112.580 131.065 112.870 131.445 ;
        RECT 113.740 131.065 114.030 131.445 ;
        RECT 114.900 131.065 115.190 131.445 ;
        RECT 117.450 130.940 117.680 131.475 ;
        RECT 119.030 131.280 119.290 131.310 ;
        RECT 119.000 131.235 119.290 131.280 ;
        RECT 122.760 131.235 122.990 131.475 ;
        RECT 125.370 131.445 125.540 131.615 ;
        RECT 126.530 131.445 126.700 131.615 ;
        RECT 127.690 131.445 127.860 131.615 ;
        RECT 128.850 131.445 129.020 132.915 ;
        RECT 235.480 132.760 235.800 133.100 ;
        RECT 236.380 132.760 236.700 133.100 ;
        RECT 118.770 131.085 122.990 131.235 ;
        RECT 119.030 131.080 119.290 131.085 ;
        RECT 122.760 130.940 122.990 131.085 ;
        RECT 125.250 131.065 125.540 131.445 ;
        RECT 126.410 131.065 126.700 131.445 ;
        RECT 127.570 131.065 127.860 131.445 ;
        RECT 128.730 131.065 129.020 131.445 ;
        RECT 234.980 131.340 235.300 131.600 ;
        RECT 235.575 131.310 235.835 131.630 ;
        RECT 236.915 131.560 237.235 131.600 ;
        RECT 236.910 131.380 237.235 131.560 ;
        RECT 236.915 131.340 237.235 131.380 ;
        RECT 133.580 131.270 133.840 131.275 ;
        RECT 141.230 131.270 141.490 131.275 ;
        RECT 164.340 131.270 164.600 131.275 ;
        RECT 172.280 131.270 172.540 131.275 ;
        RECT 203.030 131.270 203.290 131.275 ;
        RECT 209.730 131.270 209.990 131.275 ;
        RECT 220.880 131.270 221.140 131.275 ;
        RECT 231.030 131.270 231.290 131.275 ;
        RECT 133.555 130.950 133.865 131.270 ;
        RECT 141.205 130.950 141.515 131.270 ;
        RECT 164.315 130.950 164.625 131.270 ;
        RECT 172.255 130.950 172.565 131.270 ;
        RECT 203.005 130.950 203.315 131.270 ;
        RECT 209.705 130.950 210.015 131.270 ;
        RECT 220.855 130.950 221.165 131.270 ;
        RECT 231.005 130.950 231.315 131.270 ;
        RECT 117.480 130.910 117.650 130.940 ;
        RECT 122.790 130.910 122.960 130.940 ;
        RECT 3.145 130.225 3.465 130.265 ;
        RECT 3.145 130.045 3.470 130.225 ;
        RECT 3.145 130.005 3.465 130.045 ;
        RECT 3.915 130.005 4.235 130.265 ;
        RECT 5.080 130.005 5.400 130.265 ;
        RECT 8.600 129.590 8.920 130.680 ;
        RECT 9.520 129.990 10.315 130.300 ;
        RECT 18.275 129.990 19.070 130.300 ;
        RECT 19.670 129.590 19.990 130.680 ;
        RECT 29.900 129.590 30.220 130.680 ;
        RECT 30.820 129.990 31.615 130.300 ;
        RECT 36.125 129.990 36.920 130.300 ;
        RECT 37.520 129.590 37.840 130.680 ;
        RECT 67.350 129.590 67.670 130.680 ;
        RECT 68.270 129.990 69.065 130.300 ;
        RECT 74.815 129.990 75.610 130.300 ;
        RECT 76.210 129.590 76.530 130.680 ;
        RECT 98.400 129.590 98.720 130.680 ;
        RECT 99.320 129.990 100.115 130.300 ;
        RECT 105.575 129.990 106.370 130.300 ;
        RECT 106.970 129.590 107.290 130.680 ;
        RECT 120.085 130.400 120.345 130.415 ;
        RECT 120.075 130.070 120.360 130.400 ;
        RECT 133.090 129.590 133.410 130.680 ;
        RECT 134.010 129.990 134.805 130.300 ;
        RECT 140.265 129.990 141.060 130.300 ;
        RECT 141.660 129.590 141.980 130.680 ;
        RECT 163.850 129.590 164.170 130.680 ;
        RECT 164.770 129.990 165.565 130.300 ;
        RECT 171.315 129.990 172.110 130.300 ;
        RECT 172.710 129.590 173.030 130.680 ;
        RECT 202.540 129.590 202.860 130.680 ;
        RECT 203.460 129.990 204.255 130.300 ;
        RECT 208.765 129.990 209.560 130.300 ;
        RECT 210.160 129.590 210.480 130.680 ;
        RECT 220.390 129.590 220.710 130.680 ;
        RECT 221.310 129.990 222.105 130.300 ;
        RECT 230.065 129.990 230.860 130.300 ;
        RECT 231.460 129.590 231.780 130.680 ;
        RECT 234.980 130.005 235.300 130.265 ;
        RECT 236.145 130.005 236.465 130.265 ;
        RECT 236.915 130.225 237.235 130.265 ;
        RECT 236.910 130.045 237.235 130.225 ;
        RECT 236.915 130.005 237.235 130.045 ;
        RECT 9.065 129.000 9.375 129.320 ;
        RECT 19.215 129.000 19.525 129.320 ;
        RECT 30.365 129.000 30.675 129.320 ;
        RECT 37.065 129.000 37.375 129.320 ;
        RECT 67.815 129.000 68.125 129.320 ;
        RECT 75.755 129.000 76.065 129.320 ;
        RECT 98.865 129.000 99.175 129.320 ;
        RECT 106.515 129.000 106.825 129.320 ;
        RECT 117.120 128.730 118.240 129.180 ;
        RECT 122.200 128.740 123.320 129.190 ;
        RECT 133.555 129.000 133.865 129.320 ;
        RECT 141.205 129.000 141.515 129.320 ;
        RECT 164.315 129.000 164.625 129.320 ;
        RECT 172.255 129.000 172.565 129.320 ;
        RECT 203.005 129.000 203.315 129.320 ;
        RECT 209.705 129.000 210.015 129.320 ;
        RECT 220.855 129.000 221.165 129.320 ;
        RECT 231.005 129.000 231.315 129.320 ;
        RECT 119.620 126.750 119.850 126.810 ;
        RECT 120.590 126.750 120.820 126.810 ;
        RECT 119.620 126.275 120.820 126.750 ;
        RECT 119.620 126.215 119.850 126.275 ;
        RECT 120.590 126.215 120.820 126.275 ;
      LAYER via ;
        RECT 106.935 173.770 107.225 174.805 ;
        RECT 107.810 173.805 108.070 174.065 ;
        RECT 110.885 174.060 111.145 175.125 ;
        RECT 112.420 174.125 112.680 174.385 ;
        RECT 115.180 174.125 115.440 174.385 ;
        RECT 123.230 174.130 123.490 174.390 ;
        RECT 106.015 172.350 106.275 172.610 ;
        RECT 113.445 172.330 113.865 172.590 ;
        RECT 109.955 172.020 110.215 172.280 ;
        RECT 101.300 171.295 101.560 171.555 ;
        RECT 115.180 171.705 115.440 171.965 ;
        RECT 107.765 171.060 108.025 171.320 ;
        RECT 110.850 171.185 111.110 171.445 ;
        RECT 122.015 171.690 122.275 171.950 ;
        RECT 49.805 169.240 50.065 169.500 ;
        RECT 52.395 169.240 52.655 169.500 ;
        RECT 98.700 169.120 98.960 169.380 ;
        RECT 101.290 169.120 101.550 169.380 ;
        RECT 106.935 168.330 107.225 169.365 ;
        RECT 107.810 168.365 108.070 168.625 ;
        RECT 110.885 168.620 111.145 169.685 ;
        RECT 112.420 168.685 112.680 168.945 ;
        RECT 115.180 168.685 115.440 168.945 ;
        RECT 188.865 169.240 189.125 169.500 ;
        RECT 191.455 169.240 191.715 169.500 ;
        RECT 121.050 168.585 121.310 168.845 ;
        RECT 131.035 168.570 131.295 168.830 ;
        RECT 49.805 167.045 50.065 167.305 ;
        RECT 52.405 167.040 52.665 167.300 ;
        RECT 98.700 166.925 98.960 167.185 ;
        RECT 101.300 166.920 101.560 167.180 ;
        RECT 106.015 166.910 106.275 167.170 ;
        RECT 113.445 166.890 113.865 167.150 ;
        RECT 188.855 167.040 189.115 167.300 ;
        RECT 191.455 167.045 191.715 167.305 ;
        RECT 109.955 166.580 110.215 166.840 ;
        RECT 98.700 165.895 98.960 166.155 ;
        RECT 101.300 165.900 101.560 166.160 ;
        RECT 115.180 166.265 115.440 166.525 ;
        RECT 107.765 165.620 108.025 165.880 ;
        RECT 110.850 165.745 111.110 166.005 ;
        RECT 118.785 166.225 119.050 166.485 ;
        RECT 98.700 163.700 98.960 163.960 ;
        RECT 101.290 163.700 101.550 163.960 ;
        RECT 106.935 162.890 107.225 163.925 ;
        RECT 107.810 162.925 108.070 163.185 ;
        RECT 110.155 162.890 110.445 163.925 ;
        RECT 112.420 163.245 112.680 163.505 ;
        RECT 111.030 162.925 111.290 163.185 ;
        RECT 115.180 163.245 115.440 163.505 ;
        RECT 117.965 163.075 118.225 163.360 ;
        RECT 101.285 161.520 101.545 161.780 ;
        RECT 106.015 161.470 106.275 161.730 ;
        RECT 109.235 161.470 109.495 161.730 ;
        RECT 113.445 161.450 113.865 161.710 ;
        RECT 115.180 160.825 115.440 161.085 ;
        RECT 116.125 160.545 116.385 161.350 ;
        RECT 107.765 160.180 108.025 160.440 ;
        RECT 110.985 160.180 111.245 160.440 ;
        RECT 4.620 151.535 4.880 151.795 ;
        RECT 191.460 151.520 191.720 151.780 ;
        RECT 235.500 151.535 235.760 151.795 ;
        RECT 3.710 150.910 3.970 151.170 ;
        RECT 188.865 150.920 189.125 151.180 ;
        RECT 236.410 150.910 236.670 151.170 ;
        RECT 19.235 150.305 19.495 150.565 ;
        RECT 37.115 150.290 37.375 150.550 ;
        RECT 75.780 150.315 76.040 150.575 ;
        RECT 106.525 150.330 106.785 150.590 ;
        RECT 122.015 150.340 122.275 150.600 ;
        RECT 133.595 150.330 133.855 150.590 ;
        RECT 164.340 150.315 164.600 150.575 ;
        RECT 203.005 150.290 203.265 150.550 ;
        RECT 220.885 150.305 221.145 150.565 ;
        RECT 18.800 149.705 19.060 149.965 ;
        RECT 36.725 149.710 36.985 149.970 ;
        RECT 75.390 149.745 75.650 150.005 ;
        RECT 106.195 149.680 106.455 149.940 ;
        RECT 123.225 149.725 123.485 149.985 ;
        RECT 133.925 149.680 134.185 149.940 ;
        RECT 164.730 149.745 164.990 150.005 ;
        RECT 203.395 149.710 203.655 149.970 ;
        RECT 221.320 149.705 221.580 149.965 ;
        RECT 9.090 149.125 9.350 149.385 ;
        RECT 30.395 149.125 30.655 149.385 ;
        RECT 67.855 149.100 68.115 149.360 ;
        RECT 98.900 149.090 99.160 149.350 ;
        RECT 118.790 149.140 119.050 149.400 ;
        RECT 141.220 149.090 141.480 149.350 ;
        RECT 172.265 149.100 172.525 149.360 ;
        RECT 209.725 149.125 209.985 149.385 ;
        RECT 231.030 149.125 231.290 149.385 ;
        RECT 9.520 148.545 9.780 148.805 ;
        RECT 30.815 148.510 31.075 148.770 ;
        RECT 68.285 148.540 68.545 148.800 ;
        RECT 99.335 148.535 99.595 148.795 ;
        RECT 121.045 148.520 121.305 148.780 ;
        RECT 140.785 148.535 141.045 148.795 ;
        RECT 171.835 148.540 172.095 148.800 ;
        RECT 209.305 148.510 209.565 148.770 ;
        RECT 230.600 148.545 230.860 148.805 ;
        RECT 111.015 143.325 111.275 143.585 ;
        RECT 117.965 143.305 118.225 143.565 ;
        RECT 129.105 143.325 129.365 143.585 ;
        RECT 111.665 142.465 111.925 142.725 ;
        RECT 116.120 142.460 116.380 142.720 ;
        RECT 128.455 142.465 128.715 142.725 ;
        RECT 109.595 138.840 111.045 140.190 ;
        RECT 129.335 138.840 130.785 140.190 ;
        RECT 3.710 132.810 3.970 133.070 ;
        RECT 4.610 132.800 4.870 133.060 ;
        RECT 3.175 131.340 3.435 131.600 ;
        RECT 4.545 131.340 4.805 131.600 ;
        RECT 5.110 131.340 5.370 131.600 ;
        RECT 9.090 130.985 9.350 131.245 ;
        RECT 19.240 130.985 19.500 131.245 ;
        RECT 30.390 130.985 30.650 131.245 ;
        RECT 37.090 130.985 37.350 131.245 ;
        RECT 67.840 130.985 68.100 131.245 ;
        RECT 75.780 130.985 76.040 131.245 ;
        RECT 98.890 130.985 99.150 131.245 ;
        RECT 106.540 130.985 106.800 131.245 ;
        RECT 235.510 132.800 235.770 133.060 ;
        RECT 236.410 132.810 236.670 133.070 ;
        RECT 235.010 131.340 235.270 131.600 ;
        RECT 235.575 131.340 235.835 131.600 ;
        RECT 236.945 131.340 237.205 131.600 ;
        RECT 133.580 130.985 133.840 131.245 ;
        RECT 141.230 130.985 141.490 131.245 ;
        RECT 164.340 130.985 164.600 131.245 ;
        RECT 172.280 130.985 172.540 131.245 ;
        RECT 203.030 130.985 203.290 131.245 ;
        RECT 209.730 130.985 209.990 131.245 ;
        RECT 220.880 130.985 221.140 131.245 ;
        RECT 231.030 130.985 231.290 131.245 ;
        RECT 3.175 130.005 3.435 130.265 ;
        RECT 3.945 130.005 4.205 130.265 ;
        RECT 5.110 130.005 5.370 130.265 ;
        RECT 8.630 129.620 8.890 130.650 ;
        RECT 9.550 130.015 10.285 130.275 ;
        RECT 18.305 130.015 19.040 130.275 ;
        RECT 19.700 129.620 19.960 130.650 ;
        RECT 29.930 129.620 30.190 130.650 ;
        RECT 30.850 130.015 31.585 130.275 ;
        RECT 36.155 130.015 36.890 130.275 ;
        RECT 37.550 129.620 37.810 130.650 ;
        RECT 67.380 129.620 67.640 130.650 ;
        RECT 68.300 130.015 69.035 130.275 ;
        RECT 74.845 130.015 75.580 130.275 ;
        RECT 76.240 129.620 76.500 130.650 ;
        RECT 98.430 129.620 98.690 130.650 ;
        RECT 99.350 130.015 100.085 130.275 ;
        RECT 105.605 130.015 106.340 130.275 ;
        RECT 107.000 129.620 107.260 130.650 ;
        RECT 120.085 130.125 120.345 130.385 ;
        RECT 133.120 129.620 133.380 130.650 ;
        RECT 134.040 130.015 134.775 130.275 ;
        RECT 140.295 130.015 141.030 130.275 ;
        RECT 141.690 129.620 141.950 130.650 ;
        RECT 163.880 129.620 164.140 130.650 ;
        RECT 164.800 130.015 165.535 130.275 ;
        RECT 171.345 130.015 172.080 130.275 ;
        RECT 172.740 129.620 173.000 130.650 ;
        RECT 202.570 129.620 202.830 130.650 ;
        RECT 203.490 130.015 204.225 130.275 ;
        RECT 208.795 130.015 209.530 130.275 ;
        RECT 210.190 129.620 210.450 130.650 ;
        RECT 220.420 129.620 220.680 130.650 ;
        RECT 221.340 130.015 222.075 130.275 ;
        RECT 230.095 130.015 230.830 130.275 ;
        RECT 231.490 129.620 231.750 130.650 ;
        RECT 235.010 130.005 235.270 130.265 ;
        RECT 236.175 130.005 236.435 130.265 ;
        RECT 236.945 130.005 237.205 130.265 ;
        RECT 9.090 129.030 9.350 129.290 ;
        RECT 19.240 129.030 19.500 129.290 ;
        RECT 30.390 129.030 30.650 129.290 ;
        RECT 37.090 129.030 37.350 129.290 ;
        RECT 67.840 129.030 68.100 129.290 ;
        RECT 75.780 129.030 76.040 129.290 ;
        RECT 98.890 129.030 99.150 129.290 ;
        RECT 106.540 129.030 106.800 129.290 ;
        RECT 117.180 128.760 118.180 129.150 ;
        RECT 122.260 128.770 123.260 129.160 ;
        RECT 133.580 129.030 133.840 129.290 ;
        RECT 141.230 129.030 141.490 129.290 ;
        RECT 164.340 129.030 164.600 129.290 ;
        RECT 172.280 129.030 172.540 129.290 ;
        RECT 203.030 129.030 203.290 129.290 ;
        RECT 209.730 129.030 209.990 129.290 ;
        RECT 220.880 129.030 221.140 129.290 ;
        RECT 231.030 129.030 231.290 129.290 ;
        RECT 120.090 126.380 120.350 126.640 ;
      LAYER met2 ;
        RECT 106.935 173.740 107.225 174.835 ;
        RECT 107.810 173.775 108.070 174.095 ;
        RECT 110.885 174.030 111.145 175.155 ;
        RECT 112.390 174.330 112.710 174.385 ;
        RECT 112.390 174.170 113.790 174.330 ;
        RECT 112.390 174.125 112.710 174.170 ;
        RECT 105.960 172.340 106.330 172.620 ;
        RECT 101.245 171.285 101.615 171.565 ;
        RECT 107.810 171.350 107.980 173.775 ;
        RECT 109.955 171.990 110.215 172.310 ;
        RECT 110.905 171.445 111.065 174.030 ;
        RECT 113.625 172.590 113.790 174.170 ;
        RECT 115.150 174.125 115.470 174.385 ;
        RECT 123.230 174.100 123.490 174.420 ;
        RECT 113.415 172.330 113.895 172.590 ;
        RECT 115.150 171.705 115.470 171.965 ;
        RECT 122.015 171.660 122.275 171.980 ;
        RECT 107.765 171.030 108.025 171.350 ;
        RECT 110.820 171.185 111.140 171.445 ;
        RECT 49.775 169.240 50.095 169.500 ;
        RECT 52.365 169.240 52.685 169.500 ;
        RECT 49.845 167.305 50.015 169.240 ;
        RECT 49.775 167.040 50.095 167.305 ;
        RECT 52.440 167.300 52.610 169.240 ;
        RECT 98.670 169.120 98.990 169.380 ;
        RECT 101.260 169.120 101.580 169.380 ;
        RECT 49.845 155.800 50.015 167.040 ;
        RECT 52.375 167.030 52.695 167.300 ;
        RECT 98.740 167.195 98.910 169.120 ;
        RECT 52.440 156.680 52.610 167.030 ;
        RECT 98.645 166.915 99.015 167.195 ;
        RECT 101.335 167.180 101.505 169.120 ;
        RECT 106.935 168.300 107.225 169.395 ;
        RECT 107.810 168.335 108.070 168.655 ;
        RECT 110.885 168.590 111.145 169.715 ;
        RECT 112.390 168.890 112.710 168.945 ;
        RECT 112.390 168.730 113.790 168.890 ;
        RECT 112.390 168.685 112.710 168.730 ;
        RECT 101.270 166.910 101.590 167.180 ;
        RECT 105.960 166.900 106.330 167.180 ;
        RECT 98.670 165.895 98.990 166.160 ;
        RECT 101.270 165.900 101.590 166.170 ;
        RECT 107.810 165.910 107.980 168.335 ;
        RECT 109.955 166.550 110.215 166.870 ;
        RECT 110.905 166.005 111.065 168.590 ;
        RECT 113.625 167.150 113.790 168.730 ;
        RECT 115.150 168.685 115.470 168.945 ;
        RECT 121.050 168.555 121.310 168.875 ;
        RECT 113.415 166.890 113.895 167.150 ;
        RECT 115.150 166.265 115.470 166.525 ;
        RECT 118.785 166.195 119.050 166.515 ;
        RECT 98.740 163.960 98.910 165.895 ;
        RECT 101.335 163.960 101.505 165.900 ;
        RECT 107.765 165.590 108.025 165.910 ;
        RECT 110.820 165.745 111.140 166.005 ;
        RECT 98.670 163.700 98.990 163.960 ;
        RECT 101.260 163.700 101.580 163.960 ;
        RECT 106.935 162.860 107.225 163.955 ;
        RECT 107.810 162.895 108.070 163.215 ;
        RECT 101.230 161.510 101.600 161.790 ;
        RECT 105.960 161.460 106.330 161.745 ;
        RECT 107.810 161.685 107.980 162.895 ;
        RECT 110.155 162.860 110.445 163.955 ;
        RECT 112.390 163.450 112.710 163.505 ;
        RECT 112.390 163.290 113.790 163.450 ;
        RECT 112.390 163.245 112.710 163.290 ;
        RECT 111.030 162.895 111.290 163.215 ;
        RECT 109.205 161.685 109.525 161.730 ;
        RECT 107.810 161.495 109.525 161.685 ;
        RECT 107.810 160.470 107.980 161.495 ;
        RECT 109.205 161.470 109.525 161.495 ;
        RECT 111.030 160.470 111.200 162.895 ;
        RECT 113.625 161.710 113.790 163.290 ;
        RECT 115.150 163.245 115.470 163.505 ;
        RECT 117.965 163.045 118.230 163.390 ;
        RECT 113.415 161.450 113.895 161.710 ;
        RECT 115.150 160.825 115.470 161.085 ;
        RECT 116.125 160.515 116.385 161.380 ;
        RECT 107.765 160.150 108.025 160.470 ;
        RECT 110.985 160.150 111.245 160.470 ;
        RECT 52.300 156.250 52.750 156.680 ;
        RECT 49.700 155.370 50.150 155.800 ;
        RECT 4.620 151.505 4.880 151.825 ;
        RECT 3.710 150.880 3.970 151.200 ;
        RECT 3.770 133.100 3.920 150.880 ;
        RECT 3.710 132.780 3.970 133.100 ;
        RECT 4.665 133.090 4.815 151.505 ;
        RECT 19.235 150.275 19.495 150.595 ;
        RECT 18.800 149.675 19.060 149.995 ;
        RECT 9.090 149.095 9.350 149.415 ;
        RECT 4.610 132.770 4.870 133.090 ;
        RECT 3.145 131.555 3.465 131.600 ;
        RECT 4.545 131.555 4.805 131.630 ;
        RECT 5.080 131.555 5.400 131.600 ;
        RECT 3.145 131.385 5.400 131.555 ;
        RECT 3.145 131.340 3.465 131.385 ;
        RECT 4.545 131.310 4.805 131.385 ;
        RECT 5.080 131.340 5.400 131.385 ;
        RECT 9.145 131.275 9.295 149.095 ;
        RECT 9.520 148.515 9.780 148.835 ;
        RECT 9.090 130.955 9.350 131.275 ;
        RECT 9.145 130.950 9.295 130.955 ;
        RECT 3.145 130.220 3.465 130.265 ;
        RECT 3.915 130.220 4.235 130.265 ;
        RECT 5.080 130.255 5.400 130.265 ;
        RECT 8.620 130.255 8.900 130.680 ;
        RECT 9.540 130.640 9.690 148.515 ;
        RECT 5.080 130.220 8.900 130.255 ;
        RECT 3.145 130.050 8.900 130.220 ;
        RECT 3.145 130.005 3.465 130.050 ;
        RECT 3.915 130.005 4.235 130.050 ;
        RECT 5.080 130.035 8.900 130.050 ;
        RECT 5.080 130.005 5.400 130.035 ;
        RECT 8.620 129.565 8.900 130.035 ;
        RECT 9.145 130.490 9.690 130.640 ;
        RECT 18.900 130.640 19.050 149.675 ;
        RECT 19.295 131.275 19.445 150.275 ;
        RECT 37.115 150.260 37.375 150.580 ;
        RECT 75.780 150.285 76.040 150.605 ;
        RECT 106.525 150.300 106.785 150.620 ;
        RECT 36.725 149.680 36.985 150.000 ;
        RECT 30.395 149.095 30.655 149.415 ;
        RECT 30.445 131.275 30.595 149.095 ;
        RECT 30.815 148.480 31.075 148.800 ;
        RECT 19.240 130.955 19.500 131.275 ;
        RECT 30.390 130.955 30.650 131.275 ;
        RECT 19.295 130.950 19.445 130.955 ;
        RECT 30.445 130.950 30.595 130.955 ;
        RECT 18.900 130.490 19.445 130.640 ;
        RECT 9.145 129.320 9.295 130.490 ;
        RECT 9.540 129.960 10.315 130.330 ;
        RECT 18.275 129.960 19.050 130.330 ;
        RECT 19.295 129.320 19.445 130.490 ;
        RECT 19.690 129.565 19.970 130.680 ;
        RECT 29.920 129.565 30.200 130.680 ;
        RECT 30.840 130.640 30.990 148.480 ;
        RECT 30.445 130.490 30.990 130.640 ;
        RECT 36.750 130.640 36.900 149.680 ;
        RECT 37.145 131.275 37.295 150.260 ;
        RECT 75.390 149.715 75.650 150.035 ;
        RECT 67.855 149.070 68.115 149.390 ;
        RECT 67.895 131.275 68.045 149.070 ;
        RECT 68.285 148.510 68.545 148.830 ;
        RECT 37.090 130.955 37.350 131.275 ;
        RECT 67.840 130.955 68.100 131.275 ;
        RECT 37.145 130.950 37.295 130.955 ;
        RECT 67.895 130.950 68.045 130.955 ;
        RECT 36.750 130.490 37.295 130.640 ;
        RECT 30.445 129.320 30.595 130.490 ;
        RECT 30.840 129.960 31.615 130.330 ;
        RECT 36.125 129.960 36.900 130.330 ;
        RECT 37.145 129.320 37.295 130.490 ;
        RECT 37.540 129.565 37.820 130.680 ;
        RECT 67.370 129.565 67.650 130.680 ;
        RECT 68.290 130.640 68.440 148.510 ;
        RECT 67.895 130.490 68.440 130.640 ;
        RECT 75.440 130.640 75.590 149.715 ;
        RECT 75.835 131.275 75.985 150.285 ;
        RECT 106.195 149.650 106.455 149.970 ;
        RECT 98.900 149.060 99.160 149.380 ;
        RECT 98.945 131.275 99.095 149.060 ;
        RECT 99.335 148.505 99.595 148.825 ;
        RECT 75.780 130.955 76.040 131.275 ;
        RECT 98.890 130.955 99.150 131.275 ;
        RECT 75.835 130.950 75.985 130.955 ;
        RECT 98.945 130.950 99.095 130.955 ;
        RECT 75.440 130.490 75.985 130.640 ;
        RECT 67.895 129.320 68.045 130.490 ;
        RECT 68.290 129.960 69.065 130.330 ;
        RECT 74.815 129.960 75.590 130.330 ;
        RECT 75.835 129.320 75.985 130.490 ;
        RECT 76.230 129.565 76.510 130.680 ;
        RECT 98.420 129.565 98.700 130.680 ;
        RECT 99.340 130.640 99.490 148.505 ;
        RECT 98.945 130.490 99.490 130.640 ;
        RECT 106.200 130.640 106.350 149.650 ;
        RECT 106.595 131.275 106.745 150.300 ;
        RECT 110.985 143.325 111.305 143.585 ;
        RECT 116.135 142.755 116.375 160.515 ;
        RECT 117.970 143.595 118.220 163.045 ;
        RECT 118.790 149.045 119.050 166.195 ;
        RECT 121.055 148.810 121.300 168.555 ;
        RECT 122.020 150.630 122.270 171.660 ;
        RECT 122.010 150.310 122.280 150.630 ;
        RECT 122.020 150.300 122.270 150.310 ;
        RECT 123.235 150.015 123.480 174.100 ;
        RECT 188.835 169.240 189.155 169.500 ;
        RECT 191.425 169.240 191.745 169.500 ;
        RECT 130.975 168.510 131.375 168.915 ;
        RECT 188.910 167.300 189.080 169.240 ;
        RECT 191.505 167.305 191.675 169.240 ;
        RECT 188.825 167.030 189.145 167.300 ;
        RECT 191.425 167.040 191.745 167.305 ;
        RECT 188.910 151.180 189.080 167.030 ;
        RECT 191.505 151.810 191.675 167.040 ;
        RECT 191.460 151.490 191.720 151.810 ;
        RECT 235.500 151.505 235.760 151.825 ;
        RECT 188.835 150.920 189.155 151.180 ;
        RECT 133.595 150.300 133.855 150.620 ;
        RECT 123.225 149.695 123.485 150.015 ;
        RECT 123.235 149.625 123.480 149.695 ;
        RECT 121.045 148.490 121.305 148.810 ;
        RECT 117.965 143.270 118.225 143.595 ;
        RECT 129.075 143.325 129.395 143.585 ;
        RECT 111.635 142.465 111.955 142.725 ;
        RECT 116.120 142.430 116.380 142.755 ;
        RECT 128.425 142.465 128.745 142.725 ;
        RECT 109.530 138.755 111.125 140.315 ;
        RECT 129.255 138.755 130.850 140.315 ;
        RECT 133.635 131.275 133.785 150.300 ;
        RECT 164.340 150.285 164.600 150.605 ;
        RECT 133.925 149.650 134.185 149.970 ;
        RECT 106.540 130.955 106.800 131.275 ;
        RECT 133.580 130.955 133.840 131.275 ;
        RECT 106.595 130.950 106.745 130.955 ;
        RECT 133.635 130.950 133.785 130.955 ;
        RECT 106.200 130.490 106.745 130.640 ;
        RECT 98.945 129.320 99.095 130.490 ;
        RECT 99.340 129.960 100.115 130.330 ;
        RECT 105.575 129.960 106.350 130.330 ;
        RECT 106.595 129.320 106.745 130.490 ;
        RECT 106.990 129.565 107.270 130.680 ;
        RECT 120.075 130.070 120.355 130.440 ;
        RECT 133.110 129.565 133.390 130.680 ;
        RECT 134.030 130.640 134.180 149.650 ;
        RECT 141.220 149.060 141.480 149.380 ;
        RECT 140.785 148.505 141.045 148.825 ;
        RECT 133.635 130.490 134.180 130.640 ;
        RECT 140.890 130.640 141.040 148.505 ;
        RECT 141.285 131.275 141.435 149.060 ;
        RECT 164.395 131.275 164.545 150.285 ;
        RECT 203.005 150.260 203.265 150.580 ;
        RECT 220.885 150.275 221.145 150.595 ;
        RECT 164.730 149.715 164.990 150.035 ;
        RECT 141.230 130.955 141.490 131.275 ;
        RECT 164.340 130.955 164.600 131.275 ;
        RECT 141.285 130.950 141.435 130.955 ;
        RECT 164.395 130.950 164.545 130.955 ;
        RECT 140.890 130.490 141.435 130.640 ;
        RECT 133.635 129.320 133.785 130.490 ;
        RECT 134.030 129.960 134.805 130.330 ;
        RECT 140.265 129.960 141.040 130.330 ;
        RECT 141.285 129.320 141.435 130.490 ;
        RECT 141.680 129.565 141.960 130.680 ;
        RECT 163.870 129.565 164.150 130.680 ;
        RECT 164.790 130.640 164.940 149.715 ;
        RECT 172.265 149.070 172.525 149.390 ;
        RECT 171.835 148.510 172.095 148.830 ;
        RECT 164.395 130.490 164.940 130.640 ;
        RECT 171.940 130.640 172.090 148.510 ;
        RECT 172.335 131.275 172.485 149.070 ;
        RECT 203.085 131.275 203.235 150.260 ;
        RECT 203.395 149.680 203.655 150.000 ;
        RECT 172.280 130.955 172.540 131.275 ;
        RECT 203.030 130.955 203.290 131.275 ;
        RECT 172.335 130.950 172.485 130.955 ;
        RECT 203.085 130.950 203.235 130.955 ;
        RECT 171.940 130.490 172.485 130.640 ;
        RECT 164.395 129.320 164.545 130.490 ;
        RECT 164.790 129.960 165.565 130.330 ;
        RECT 171.315 129.960 172.090 130.330 ;
        RECT 172.335 129.320 172.485 130.490 ;
        RECT 172.730 129.565 173.010 130.680 ;
        RECT 202.560 129.565 202.840 130.680 ;
        RECT 203.480 130.640 203.630 149.680 ;
        RECT 209.725 149.095 209.985 149.415 ;
        RECT 209.305 148.480 209.565 148.800 ;
        RECT 203.085 130.490 203.630 130.640 ;
        RECT 209.390 130.640 209.540 148.480 ;
        RECT 209.785 131.275 209.935 149.095 ;
        RECT 220.935 131.275 221.085 150.275 ;
        RECT 221.320 149.675 221.580 149.995 ;
        RECT 209.730 130.955 209.990 131.275 ;
        RECT 220.880 130.955 221.140 131.275 ;
        RECT 209.785 130.950 209.935 130.955 ;
        RECT 220.935 130.950 221.085 130.955 ;
        RECT 209.390 130.490 209.935 130.640 ;
        RECT 203.085 129.320 203.235 130.490 ;
        RECT 203.480 129.960 204.255 130.330 ;
        RECT 208.765 129.960 209.540 130.330 ;
        RECT 209.785 129.320 209.935 130.490 ;
        RECT 210.180 129.565 210.460 130.680 ;
        RECT 220.410 129.565 220.690 130.680 ;
        RECT 221.330 130.640 221.480 149.675 ;
        RECT 231.030 149.095 231.290 149.415 ;
        RECT 230.600 148.515 230.860 148.835 ;
        RECT 220.935 130.490 221.480 130.640 ;
        RECT 230.690 130.640 230.840 148.515 ;
        RECT 231.085 131.275 231.235 149.095 ;
        RECT 235.565 133.090 235.715 151.505 ;
        RECT 236.410 150.880 236.670 151.200 ;
        RECT 236.460 133.100 236.610 150.880 ;
        RECT 235.510 132.770 235.770 133.090 ;
        RECT 236.410 132.780 236.670 133.100 ;
        RECT 234.980 131.570 235.300 131.600 ;
        RECT 231.550 131.555 235.300 131.570 ;
        RECT 235.575 131.555 235.835 131.630 ;
        RECT 236.915 131.555 237.235 131.600 ;
        RECT 231.550 131.385 237.235 131.555 ;
        RECT 231.550 131.350 235.300 131.385 ;
        RECT 231.030 130.955 231.290 131.275 ;
        RECT 231.085 130.950 231.235 130.955 ;
        RECT 231.550 130.680 231.775 131.350 ;
        RECT 234.980 131.340 235.300 131.350 ;
        RECT 235.575 131.310 235.835 131.385 ;
        RECT 236.915 131.340 237.235 131.385 ;
        RECT 230.690 130.490 231.235 130.640 ;
        RECT 220.935 129.320 221.085 130.490 ;
        RECT 221.330 129.960 222.105 130.330 ;
        RECT 230.065 129.960 230.840 130.330 ;
        RECT 231.085 129.320 231.235 130.490 ;
        RECT 231.480 130.320 231.775 130.680 ;
        RECT 231.480 129.565 231.760 130.320 ;
        RECT 234.980 130.220 235.300 130.265 ;
        RECT 236.145 130.220 236.465 130.265 ;
        RECT 236.915 130.220 237.235 130.265 ;
        RECT 234.980 130.050 237.235 130.220 ;
        RECT 234.980 130.005 235.300 130.050 ;
        RECT 236.145 130.005 236.465 130.050 ;
        RECT 236.915 130.005 237.235 130.050 ;
        RECT 9.090 129.000 9.350 129.320 ;
        RECT 19.240 129.000 19.500 129.320 ;
        RECT 30.390 129.000 30.650 129.320 ;
        RECT 37.090 129.000 37.350 129.320 ;
        RECT 67.840 129.000 68.100 129.320 ;
        RECT 75.780 129.000 76.040 129.320 ;
        RECT 98.890 129.000 99.150 129.320 ;
        RECT 106.540 129.000 106.800 129.320 ;
        RECT 117.120 128.730 118.240 129.180 ;
        RECT 122.200 128.740 123.320 129.190 ;
        RECT 133.580 129.000 133.840 129.320 ;
        RECT 141.230 129.000 141.490 129.320 ;
        RECT 164.340 129.000 164.600 129.320 ;
        RECT 172.280 129.000 172.540 129.320 ;
        RECT 203.030 129.000 203.290 129.320 ;
        RECT 209.730 129.000 209.990 129.320 ;
        RECT 220.880 129.000 221.140 129.320 ;
        RECT 231.030 129.000 231.290 129.320 ;
        RECT 120.080 126.325 120.360 126.695 ;
      LAYER via2 ;
        RECT 106.005 172.340 106.285 172.620 ;
        RECT 101.290 171.285 101.570 171.565 ;
        RECT 98.690 166.915 98.970 167.195 ;
        RECT 106.005 166.900 106.285 167.180 ;
        RECT 101.275 161.510 101.555 161.790 ;
        RECT 106.005 161.460 106.285 161.745 ;
        RECT 52.350 156.290 52.700 156.640 ;
        RECT 49.750 155.410 50.100 155.760 ;
        RECT 8.620 129.610 8.900 130.625 ;
        RECT 9.540 130.005 10.285 130.285 ;
        RECT 18.305 130.005 19.050 130.285 ;
        RECT 19.690 129.610 19.970 130.625 ;
        RECT 29.920 129.610 30.200 130.625 ;
        RECT 30.840 130.005 31.585 130.285 ;
        RECT 36.155 130.005 36.900 130.285 ;
        RECT 37.540 129.610 37.820 130.625 ;
        RECT 67.370 129.610 67.650 130.625 ;
        RECT 68.290 130.005 69.035 130.285 ;
        RECT 74.845 130.005 75.590 130.285 ;
        RECT 76.230 129.610 76.510 130.625 ;
        RECT 98.420 129.610 98.700 130.625 ;
        RECT 131.020 168.555 131.330 168.870 ;
        RECT 109.595 138.840 111.045 140.190 ;
        RECT 129.335 138.840 130.785 140.190 ;
        RECT 99.340 130.005 100.085 130.285 ;
        RECT 105.605 130.005 106.350 130.285 ;
        RECT 106.990 129.610 107.270 130.625 ;
        RECT 120.075 130.115 120.355 130.395 ;
        RECT 133.110 129.610 133.390 130.625 ;
        RECT 134.030 130.005 134.775 130.285 ;
        RECT 140.295 130.005 141.040 130.285 ;
        RECT 141.680 129.610 141.960 130.625 ;
        RECT 163.870 129.610 164.150 130.625 ;
        RECT 164.790 130.005 165.535 130.285 ;
        RECT 171.345 130.005 172.090 130.285 ;
        RECT 172.730 129.610 173.010 130.625 ;
        RECT 202.560 129.610 202.840 130.625 ;
        RECT 203.480 130.005 204.225 130.285 ;
        RECT 208.795 130.005 209.540 130.285 ;
        RECT 210.180 129.610 210.460 130.625 ;
        RECT 220.410 129.610 220.690 130.625 ;
        RECT 221.330 130.005 222.075 130.285 ;
        RECT 230.095 130.005 230.840 130.285 ;
        RECT 231.480 129.610 231.760 130.625 ;
        RECT 117.180 128.760 118.180 129.150 ;
        RECT 122.260 128.770 123.260 129.160 ;
        RECT 120.080 126.370 120.360 126.650 ;
      LAYER met3 ;
        RECT 101.245 171.585 101.725 171.590 ;
        RECT 105.965 171.585 106.320 172.725 ;
        RECT 101.245 171.260 106.320 171.585 ;
        RECT 130.895 168.460 131.440 169.000 ;
        RECT 98.615 167.210 99.015 167.220 ;
        RECT 105.960 167.210 106.330 167.215 ;
        RECT 98.615 166.890 106.330 167.210 ;
        RECT 105.960 166.875 106.330 166.890 ;
        RECT 101.230 161.805 101.600 161.815 ;
        RECT 101.230 161.485 106.335 161.805 ;
        RECT 105.955 161.415 106.335 161.485 ;
        RECT 29.170 156.610 29.600 156.630 ;
        RECT 52.300 156.610 52.750 156.680 ;
        RECT 29.170 156.310 52.750 156.610 ;
        RECT 29.170 156.290 29.600 156.310 ;
        RECT 52.300 156.250 52.750 156.310 ;
        RECT 49.700 155.730 50.150 155.800 ;
        RECT 210.780 155.730 211.210 155.750 ;
        RECT 49.700 155.430 211.210 155.730 ;
        RECT 49.700 155.370 50.150 155.430 ;
        RECT 210.780 155.410 211.210 155.430 ;
        RECT 8.560 130.395 8.955 130.705 ;
        RECT 8.445 129.895 8.955 130.395 ;
        RECT 19.635 130.395 20.030 130.705 ;
        RECT 29.860 130.395 30.255 130.705 ;
        RECT 8.560 129.555 8.955 129.895 ;
        RECT 9.495 129.890 10.315 130.390 ;
        RECT 18.275 129.890 19.095 130.390 ;
        RECT 19.635 129.895 20.145 130.395 ;
        RECT 29.745 129.895 30.255 130.395 ;
        RECT 37.485 130.395 37.880 130.705 ;
        RECT 67.310 130.395 67.705 130.705 ;
        RECT 19.635 129.555 20.030 129.895 ;
        RECT 29.860 129.555 30.255 129.895 ;
        RECT 30.795 129.890 31.615 130.390 ;
        RECT 36.125 129.890 36.945 130.390 ;
        RECT 37.485 129.895 37.995 130.395 ;
        RECT 67.195 129.895 67.705 130.395 ;
        RECT 76.175 130.395 76.570 130.705 ;
        RECT 98.360 130.395 98.755 130.705 ;
        RECT 37.485 129.555 37.880 129.895 ;
        RECT 67.310 129.555 67.705 129.895 ;
        RECT 68.245 129.890 69.065 130.390 ;
        RECT 74.815 129.890 75.635 130.390 ;
        RECT 76.175 129.895 76.685 130.395 ;
        RECT 98.245 129.895 98.755 130.395 ;
        RECT 106.935 130.395 107.330 130.705 ;
        RECT 76.175 129.555 76.570 129.895 ;
        RECT 98.360 129.555 98.755 129.895 ;
        RECT 99.295 129.890 100.115 130.390 ;
        RECT 105.575 129.890 106.395 130.390 ;
        RECT 106.935 129.895 107.445 130.395 ;
        RECT 106.935 129.555 107.330 129.895 ;
        RECT 109.530 122.450 111.130 140.315 ;
        RECT 120.070 130.460 120.370 130.570 ;
        RECT 120.020 130.065 120.405 130.460 ;
        RECT 117.150 128.730 118.210 129.180 ;
        RECT 120.070 126.675 120.370 130.065 ;
        RECT 122.230 128.740 123.290 129.190 ;
        RECT 120.055 126.345 120.385 126.675 ;
        RECT 120.070 126.325 120.370 126.345 ;
        RECT 129.250 122.450 130.850 140.315 ;
        RECT 133.050 130.395 133.445 130.705 ;
        RECT 132.935 129.895 133.445 130.395 ;
        RECT 141.625 130.395 142.020 130.705 ;
        RECT 163.810 130.395 164.205 130.705 ;
        RECT 133.050 129.555 133.445 129.895 ;
        RECT 133.985 129.890 134.805 130.390 ;
        RECT 140.265 129.890 141.085 130.390 ;
        RECT 141.625 129.895 142.135 130.395 ;
        RECT 163.695 129.895 164.205 130.395 ;
        RECT 172.675 130.395 173.070 130.705 ;
        RECT 202.500 130.395 202.895 130.705 ;
        RECT 141.625 129.555 142.020 129.895 ;
        RECT 163.810 129.555 164.205 129.895 ;
        RECT 164.745 129.890 165.565 130.390 ;
        RECT 171.315 129.890 172.135 130.390 ;
        RECT 172.675 129.895 173.185 130.395 ;
        RECT 202.385 129.895 202.895 130.395 ;
        RECT 210.125 130.395 210.520 130.705 ;
        RECT 220.350 130.395 220.745 130.705 ;
        RECT 172.675 129.555 173.070 129.895 ;
        RECT 202.500 129.555 202.895 129.895 ;
        RECT 203.435 129.890 204.255 130.390 ;
        RECT 208.765 129.890 209.585 130.390 ;
        RECT 210.125 129.895 210.635 130.395 ;
        RECT 220.235 129.895 220.745 130.395 ;
        RECT 231.425 130.395 231.820 130.705 ;
        RECT 210.125 129.555 210.520 129.895 ;
        RECT 220.350 129.555 220.745 129.895 ;
        RECT 221.285 129.890 222.105 130.390 ;
        RECT 230.065 129.890 230.885 130.390 ;
        RECT 231.425 129.895 231.935 130.395 ;
        RECT 231.425 129.555 231.820 129.895 ;
        RECT 101.665 120.840 118.605 122.450 ;
        RECT 101.665 116.715 103.275 120.840 ;
        RECT 104.875 116.715 115.395 119.240 ;
        RECT 116.995 116.715 118.605 120.840 ;
        RECT 101.665 115.115 118.605 116.715 ;
        RECT 101.665 110.890 103.275 115.115 ;
        RECT 104.875 110.890 115.395 115.115 ;
        RECT 116.995 110.890 118.605 115.115 ;
        RECT 101.665 109.290 118.605 110.890 ;
        RECT 101.665 104.660 103.275 109.290 ;
        RECT 104.875 108.720 115.395 109.290 ;
        RECT 104.875 108.710 106.595 108.720 ;
        RECT 104.995 105.650 106.595 108.710 ;
        RECT 104.875 105.640 106.595 105.650 ;
        RECT 109.335 105.640 110.935 108.720 ;
        RECT 113.675 108.710 115.395 108.720 ;
        RECT 113.675 105.650 115.275 108.710 ;
        RECT 113.675 105.640 115.395 105.650 ;
        RECT 104.875 104.660 115.395 105.640 ;
        RECT 116.995 104.660 118.605 109.290 ;
        RECT 101.665 103.045 118.605 104.660 ;
        RECT 101.665 97.925 103.275 103.045 ;
        RECT 104.875 97.925 115.395 103.045 ;
        RECT 116.995 97.925 118.605 103.045 ;
        RECT 101.665 96.310 118.605 97.925 ;
        RECT 101.665 91.060 103.275 96.310 ;
        RECT 104.875 95.120 115.395 96.310 ;
        RECT 104.875 95.110 106.595 95.120 ;
        RECT 104.995 92.050 106.595 95.110 ;
        RECT 104.875 92.040 106.595 92.050 ;
        RECT 109.335 92.040 110.935 95.120 ;
        RECT 113.675 95.110 115.395 95.120 ;
        RECT 113.675 92.050 115.275 95.110 ;
        RECT 113.675 92.040 115.395 92.050 ;
        RECT 104.875 91.060 115.395 92.040 ;
        RECT 116.995 91.060 118.605 96.310 ;
        RECT 101.665 89.445 118.605 91.060 ;
        RECT 101.665 84.325 103.275 89.445 ;
        RECT 104.875 84.325 115.395 89.445 ;
        RECT 116.995 84.325 118.605 89.445 ;
        RECT 101.665 82.710 118.605 84.325 ;
        RECT 101.665 77.460 103.275 82.710 ;
        RECT 104.875 81.520 115.395 82.710 ;
        RECT 104.875 81.510 106.595 81.520 ;
        RECT 104.995 78.450 106.595 81.510 ;
        RECT 104.875 78.440 106.595 78.450 ;
        RECT 109.335 78.440 110.935 81.520 ;
        RECT 113.675 81.510 115.395 81.520 ;
        RECT 113.675 78.450 115.275 81.510 ;
        RECT 113.675 78.440 115.395 78.450 ;
        RECT 104.875 77.460 115.395 78.440 ;
        RECT 116.995 77.460 118.605 82.710 ;
        RECT 101.665 75.845 118.605 77.460 ;
        RECT 101.665 70.725 103.275 75.845 ;
        RECT 104.875 70.725 115.395 75.845 ;
        RECT 116.995 70.725 118.605 75.845 ;
        RECT 101.665 69.110 118.605 70.725 ;
        RECT 101.665 63.860 103.275 69.110 ;
        RECT 104.875 67.920 115.395 69.110 ;
        RECT 104.875 67.910 106.595 67.920 ;
        RECT 104.995 64.850 106.595 67.910 ;
        RECT 104.875 64.840 106.595 64.850 ;
        RECT 109.335 64.840 110.935 67.920 ;
        RECT 113.675 67.910 115.395 67.920 ;
        RECT 113.675 64.850 115.275 67.910 ;
        RECT 113.675 64.840 115.395 64.850 ;
        RECT 104.875 63.860 115.395 64.840 ;
        RECT 116.995 63.860 118.605 69.110 ;
        RECT 101.665 62.245 118.605 63.860 ;
        RECT 101.665 57.125 103.275 62.245 ;
        RECT 104.875 57.125 115.395 62.245 ;
        RECT 116.995 57.125 118.605 62.245 ;
        RECT 101.665 55.510 118.605 57.125 ;
        RECT 101.665 50.260 103.275 55.510 ;
        RECT 104.875 54.320 115.395 55.510 ;
        RECT 104.875 54.310 106.595 54.320 ;
        RECT 104.995 51.250 106.595 54.310 ;
        RECT 104.875 51.240 106.595 51.250 ;
        RECT 109.335 51.240 110.935 54.320 ;
        RECT 113.675 54.310 115.395 54.320 ;
        RECT 113.675 51.250 115.275 54.310 ;
        RECT 113.675 51.240 115.395 51.250 ;
        RECT 104.875 50.260 115.395 51.240 ;
        RECT 116.995 50.260 118.605 55.510 ;
        RECT 101.665 48.645 118.605 50.260 ;
        RECT 101.665 43.525 103.275 48.645 ;
        RECT 104.875 43.525 115.395 48.645 ;
        RECT 116.995 43.525 118.605 48.645 ;
        RECT 101.665 41.910 118.605 43.525 ;
        RECT 101.665 36.660 103.275 41.910 ;
        RECT 104.875 40.720 115.395 41.910 ;
        RECT 104.875 40.710 106.595 40.720 ;
        RECT 104.995 37.650 106.595 40.710 ;
        RECT 104.875 37.640 106.595 37.650 ;
        RECT 109.335 37.640 110.935 40.720 ;
        RECT 113.675 40.710 115.395 40.720 ;
        RECT 113.675 37.650 115.275 40.710 ;
        RECT 113.675 37.640 115.395 37.650 ;
        RECT 104.875 36.660 115.395 37.640 ;
        RECT 116.995 36.660 118.605 41.910 ;
        RECT 101.665 35.045 118.605 36.660 ;
        RECT 101.665 29.925 103.275 35.045 ;
        RECT 104.875 29.925 115.395 35.045 ;
        RECT 116.995 29.925 118.605 35.045 ;
        RECT 101.665 28.310 118.605 29.925 ;
        RECT 101.665 23.470 103.275 28.310 ;
        RECT 104.875 27.120 115.395 28.310 ;
        RECT 104.875 27.110 106.595 27.120 ;
        RECT 104.995 24.050 106.595 27.110 ;
        RECT 104.875 24.040 106.595 24.050 ;
        RECT 109.335 24.040 110.935 27.120 ;
        RECT 113.675 27.110 115.395 27.120 ;
        RECT 113.675 24.050 115.275 27.110 ;
        RECT 113.675 24.040 115.395 24.050 ;
        RECT 104.875 23.470 115.395 24.040 ;
        RECT 116.995 23.470 118.605 28.310 ;
        RECT 101.665 21.870 118.605 23.470 ;
        RECT 101.665 17.645 103.275 21.870 ;
        RECT 104.875 17.645 115.395 21.870 ;
        RECT 116.995 17.645 118.605 21.870 ;
        RECT 101.665 16.045 118.605 17.645 ;
        RECT 101.665 11.920 103.275 16.045 ;
        RECT 104.875 13.520 115.395 16.045 ;
        RECT 116.995 11.920 118.605 16.045 ;
        RECT 101.665 10.310 118.605 11.920 ;
        RECT 121.775 120.840 138.715 122.450 ;
        RECT 121.775 116.715 123.385 120.840 ;
        RECT 124.985 116.715 135.505 119.240 ;
        RECT 137.105 116.715 138.715 120.840 ;
        RECT 121.775 115.115 138.715 116.715 ;
        RECT 121.775 110.890 123.385 115.115 ;
        RECT 124.985 110.890 135.505 115.115 ;
        RECT 137.105 110.890 138.715 115.115 ;
        RECT 121.775 109.290 138.715 110.890 ;
        RECT 121.775 104.660 123.385 109.290 ;
        RECT 124.985 108.720 135.505 109.290 ;
        RECT 124.985 108.710 126.705 108.720 ;
        RECT 125.105 105.650 126.705 108.710 ;
        RECT 124.985 105.640 126.705 105.650 ;
        RECT 129.445 105.640 131.045 108.720 ;
        RECT 133.785 108.710 135.505 108.720 ;
        RECT 133.785 105.650 135.385 108.710 ;
        RECT 133.785 105.640 135.505 105.650 ;
        RECT 124.985 104.660 135.505 105.640 ;
        RECT 137.105 104.660 138.715 109.290 ;
        RECT 121.775 103.045 138.715 104.660 ;
        RECT 121.775 97.925 123.385 103.045 ;
        RECT 124.985 97.925 135.505 103.045 ;
        RECT 137.105 97.925 138.715 103.045 ;
        RECT 121.775 96.310 138.715 97.925 ;
        RECT 121.775 91.060 123.385 96.310 ;
        RECT 124.985 95.120 135.505 96.310 ;
        RECT 124.985 95.110 126.705 95.120 ;
        RECT 125.105 92.050 126.705 95.110 ;
        RECT 124.985 92.040 126.705 92.050 ;
        RECT 129.445 92.040 131.045 95.120 ;
        RECT 133.785 95.110 135.505 95.120 ;
        RECT 133.785 92.050 135.385 95.110 ;
        RECT 133.785 92.040 135.505 92.050 ;
        RECT 124.985 91.060 135.505 92.040 ;
        RECT 137.105 91.060 138.715 96.310 ;
        RECT 121.775 89.445 138.715 91.060 ;
        RECT 121.775 84.325 123.385 89.445 ;
        RECT 124.985 84.325 135.505 89.445 ;
        RECT 137.105 84.325 138.715 89.445 ;
        RECT 121.775 82.710 138.715 84.325 ;
        RECT 121.775 77.460 123.385 82.710 ;
        RECT 124.985 81.520 135.505 82.710 ;
        RECT 124.985 81.510 126.705 81.520 ;
        RECT 125.105 78.450 126.705 81.510 ;
        RECT 124.985 78.440 126.705 78.450 ;
        RECT 129.445 78.440 131.045 81.520 ;
        RECT 133.785 81.510 135.505 81.520 ;
        RECT 133.785 78.450 135.385 81.510 ;
        RECT 133.785 78.440 135.505 78.450 ;
        RECT 124.985 77.460 135.505 78.440 ;
        RECT 137.105 77.460 138.715 82.710 ;
        RECT 121.775 75.845 138.715 77.460 ;
        RECT 121.775 70.725 123.385 75.845 ;
        RECT 124.985 70.725 135.505 75.845 ;
        RECT 137.105 70.725 138.715 75.845 ;
        RECT 121.775 69.110 138.715 70.725 ;
        RECT 121.775 63.860 123.385 69.110 ;
        RECT 124.985 67.920 135.505 69.110 ;
        RECT 124.985 67.910 126.705 67.920 ;
        RECT 125.105 64.850 126.705 67.910 ;
        RECT 124.985 64.840 126.705 64.850 ;
        RECT 129.445 64.840 131.045 67.920 ;
        RECT 133.785 67.910 135.505 67.920 ;
        RECT 133.785 64.850 135.385 67.910 ;
        RECT 133.785 64.840 135.505 64.850 ;
        RECT 124.985 63.860 135.505 64.840 ;
        RECT 137.105 63.860 138.715 69.110 ;
        RECT 121.775 62.245 138.715 63.860 ;
        RECT 121.775 57.125 123.385 62.245 ;
        RECT 124.985 57.125 135.505 62.245 ;
        RECT 137.105 57.125 138.715 62.245 ;
        RECT 121.775 55.510 138.715 57.125 ;
        RECT 121.775 50.260 123.385 55.510 ;
        RECT 124.985 54.320 135.505 55.510 ;
        RECT 124.985 54.310 126.705 54.320 ;
        RECT 125.105 51.250 126.705 54.310 ;
        RECT 124.985 51.240 126.705 51.250 ;
        RECT 129.445 51.240 131.045 54.320 ;
        RECT 133.785 54.310 135.505 54.320 ;
        RECT 133.785 51.250 135.385 54.310 ;
        RECT 133.785 51.240 135.505 51.250 ;
        RECT 124.985 50.260 135.505 51.240 ;
        RECT 137.105 50.260 138.715 55.510 ;
        RECT 121.775 48.645 138.715 50.260 ;
        RECT 121.775 43.525 123.385 48.645 ;
        RECT 124.985 43.525 135.505 48.645 ;
        RECT 137.105 43.525 138.715 48.645 ;
        RECT 121.775 41.910 138.715 43.525 ;
        RECT 121.775 36.660 123.385 41.910 ;
        RECT 124.985 40.720 135.505 41.910 ;
        RECT 124.985 40.710 126.705 40.720 ;
        RECT 125.105 37.650 126.705 40.710 ;
        RECT 124.985 37.640 126.705 37.650 ;
        RECT 129.445 37.640 131.045 40.720 ;
        RECT 133.785 40.710 135.505 40.720 ;
        RECT 133.785 37.650 135.385 40.710 ;
        RECT 133.785 37.640 135.505 37.650 ;
        RECT 124.985 36.660 135.505 37.640 ;
        RECT 137.105 36.660 138.715 41.910 ;
        RECT 121.775 35.045 138.715 36.660 ;
        RECT 121.775 29.925 123.385 35.045 ;
        RECT 124.985 29.925 135.505 35.045 ;
        RECT 137.105 29.925 138.715 35.045 ;
        RECT 121.775 28.310 138.715 29.925 ;
        RECT 121.775 23.470 123.385 28.310 ;
        RECT 124.985 27.120 135.505 28.310 ;
        RECT 124.985 27.110 126.705 27.120 ;
        RECT 125.105 24.050 126.705 27.110 ;
        RECT 124.985 24.040 126.705 24.050 ;
        RECT 129.445 24.040 131.045 27.120 ;
        RECT 133.785 27.110 135.505 27.120 ;
        RECT 133.785 24.050 135.385 27.110 ;
        RECT 133.785 24.040 135.505 24.050 ;
        RECT 124.985 23.470 135.505 24.040 ;
        RECT 137.105 23.470 138.715 28.310 ;
        RECT 121.775 21.870 138.715 23.470 ;
        RECT 121.775 17.645 123.385 21.870 ;
        RECT 124.985 17.645 135.505 21.870 ;
        RECT 137.105 17.645 138.715 21.870 ;
        RECT 121.775 16.045 138.715 17.645 ;
        RECT 121.775 11.920 123.385 16.045 ;
        RECT 124.985 13.520 135.505 16.045 ;
        RECT 137.105 11.920 138.715 16.045 ;
        RECT 121.775 10.310 138.715 11.920 ;
      LAYER via3 ;
        RECT 130.975 168.510 131.375 168.915 ;
        RECT 29.200 156.300 29.570 156.620 ;
        RECT 210.810 155.420 211.180 155.740 ;
        RECT 109.595 138.840 111.045 140.190 ;
        RECT 8.600 129.590 8.920 130.690 ;
        RECT 9.520 129.985 10.315 130.305 ;
        RECT 18.275 129.985 19.070 130.305 ;
        RECT 19.670 129.590 19.990 130.690 ;
        RECT 29.900 129.590 30.220 130.690 ;
        RECT 30.820 129.985 31.615 130.305 ;
        RECT 36.125 129.985 36.920 130.305 ;
        RECT 37.520 129.590 37.840 130.690 ;
        RECT 67.350 129.590 67.670 130.690 ;
        RECT 68.270 129.985 69.065 130.305 ;
        RECT 74.815 129.985 75.610 130.305 ;
        RECT 76.210 129.590 76.530 130.690 ;
        RECT 98.400 129.590 98.720 130.690 ;
        RECT 99.320 129.985 100.115 130.305 ;
        RECT 105.575 129.985 106.370 130.305 ;
        RECT 106.970 129.590 107.290 130.690 ;
        RECT 129.335 138.840 130.785 140.190 ;
        RECT 120.050 130.095 120.370 130.415 ;
        RECT 117.180 128.760 118.180 129.150 ;
        RECT 122.260 128.770 123.260 129.160 ;
        RECT 133.090 129.590 133.410 130.690 ;
        RECT 134.010 129.985 134.805 130.305 ;
        RECT 140.265 129.985 141.060 130.305 ;
        RECT 141.660 129.590 141.980 130.690 ;
        RECT 163.850 129.590 164.170 130.690 ;
        RECT 164.770 129.985 165.565 130.305 ;
        RECT 171.315 129.985 172.110 130.305 ;
        RECT 172.710 129.590 173.030 130.690 ;
        RECT 202.540 129.590 202.860 130.690 ;
        RECT 203.460 129.985 204.255 130.305 ;
        RECT 208.765 129.985 209.560 130.305 ;
        RECT 210.160 129.590 210.480 130.690 ;
        RECT 220.390 129.590 220.710 130.690 ;
        RECT 221.310 129.985 222.105 130.305 ;
        RECT 230.065 129.985 230.860 130.305 ;
        RECT 231.460 129.590 231.780 130.690 ;
        RECT 101.830 120.995 106.620 122.285 ;
        RECT 115.200 120.995 118.440 122.285 ;
        RECT 101.830 107.925 103.120 120.995 ;
        RECT 101.830 94.230 103.120 106.250 ;
        RECT 117.150 107.925 118.440 120.995 ;
        RECT 101.830 80.630 103.120 92.650 ;
        RECT 117.150 94.230 118.440 106.250 ;
        RECT 101.830 67.030 103.120 79.050 ;
        RECT 117.150 80.630 118.440 92.650 ;
        RECT 101.830 53.430 103.120 65.450 ;
        RECT 117.150 67.030 118.440 79.050 ;
        RECT 101.830 39.830 103.120 51.850 ;
        RECT 117.150 53.430 118.440 65.450 ;
        RECT 101.830 26.230 103.120 38.250 ;
        RECT 117.150 39.830 118.440 51.850 ;
        RECT 101.830 11.765 103.120 24.835 ;
        RECT 117.150 26.230 118.440 38.250 ;
        RECT 117.150 11.765 118.440 24.835 ;
        RECT 101.830 10.475 105.070 11.765 ;
        RECT 113.650 10.475 118.440 11.765 ;
        RECT 121.940 120.995 125.180 122.285 ;
        RECT 133.760 120.995 138.550 122.285 ;
        RECT 121.940 107.925 123.230 120.995 ;
        RECT 121.940 94.230 123.230 106.250 ;
        RECT 137.260 107.925 138.550 120.995 ;
        RECT 121.940 80.630 123.230 92.650 ;
        RECT 137.260 94.230 138.550 106.250 ;
        RECT 121.940 67.030 123.230 79.050 ;
        RECT 137.260 80.630 138.550 92.650 ;
        RECT 121.940 53.430 123.230 65.450 ;
        RECT 137.260 67.030 138.550 79.050 ;
        RECT 121.940 39.830 123.230 51.850 ;
        RECT 137.260 53.430 138.550 65.450 ;
        RECT 121.940 26.230 123.230 38.250 ;
        RECT 137.260 39.830 138.550 51.850 ;
        RECT 121.940 11.765 123.230 24.835 ;
        RECT 137.260 26.230 138.550 38.250 ;
        RECT 137.260 11.765 138.550 24.835 ;
        RECT 121.940 10.475 126.730 11.765 ;
        RECT 135.310 10.475 138.550 11.765 ;
      LAYER met4 ;
        RECT 130.895 168.885 131.440 169.000 ;
        RECT 130.215 168.520 131.440 168.885 ;
        RECT 130.220 162.520 130.555 168.520 ;
        RECT 130.895 168.460 131.440 168.520 ;
        RECT 121.205 162.160 130.555 162.520 ;
        RECT 29.170 156.290 29.600 156.630 ;
        RECT 10.935 135.820 11.455 136.340 ;
        RECT 11.935 135.820 12.455 136.340 ;
        RECT 12.935 135.820 13.455 136.340 ;
        RECT 13.935 135.820 14.455 136.340 ;
        RECT 14.935 135.820 15.455 136.340 ;
        RECT 15.935 135.820 16.455 136.340 ;
        RECT 16.935 135.820 17.455 136.340 ;
        RECT 10.935 134.820 11.455 135.340 ;
        RECT 16.935 134.820 17.455 135.340 ;
        RECT 10.935 133.820 11.455 134.340 ;
        RECT 16.935 133.820 17.455 134.340 ;
        RECT 10.935 132.820 11.455 133.340 ;
        RECT 16.935 132.820 17.455 133.340 ;
        RECT 10.935 131.820 11.455 132.340 ;
        RECT 16.935 131.820 17.455 132.340 ;
        RECT 10.935 131.335 11.455 131.340 ;
        RECT 11.935 131.335 12.455 131.340 ;
        RECT 10.295 130.820 12.455 131.335 ;
        RECT 12.935 130.820 13.455 131.340 ;
        RECT 13.935 130.820 14.455 131.340 ;
        RECT 14.935 130.820 15.455 131.340 ;
        RECT 15.935 130.820 16.455 131.340 ;
        RECT 16.935 131.090 17.455 131.340 ;
        RECT 16.935 130.820 17.705 131.090 ;
        RECT 8.595 130.325 8.940 130.695 ;
        RECT 10.295 130.325 12.185 130.820 ;
        RECT 8.270 129.965 8.940 130.325 ;
        RECT 9.500 129.965 12.185 130.325 ;
        RECT 16.970 130.325 17.705 130.820 ;
        RECT 19.650 130.325 19.995 130.695 ;
        RECT 29.200 130.325 29.570 156.290 ;
        RECT 109.530 138.755 111.125 140.315 ;
        RECT 121.205 136.050 121.580 162.160 ;
        RECT 210.780 155.410 211.210 155.750 ;
        RECT 129.255 138.755 130.850 140.315 ;
        RECT 32.040 130.790 35.720 133.840 ;
        RECT 69.895 131.045 74.175 135.855 ;
        RECT 119.120 135.620 121.580 136.050 ;
        RECT 69.895 130.940 74.645 131.045 ;
        RECT 32.030 130.780 35.720 130.790 ;
        RECT 29.895 130.325 30.240 130.695 ;
        RECT 32.030 130.560 35.890 130.780 ;
        RECT 32.030 130.325 32.585 130.560 ;
        RECT 16.970 129.965 19.090 130.325 ;
        RECT 8.595 129.570 8.940 129.965 ;
        RECT 10.295 129.880 12.185 129.965 ;
        RECT 19.650 129.570 21.095 130.325 ;
        RECT 29.200 129.965 30.240 130.325 ;
        RECT 30.800 129.965 32.585 130.325 ;
        RECT 35.350 130.325 35.890 130.560 ;
        RECT 37.500 130.325 37.845 130.695 ;
        RECT 67.345 130.325 67.690 130.695 ;
        RECT 69.815 130.575 74.645 130.940 ;
        RECT 69.815 130.325 70.485 130.575 ;
        RECT 35.350 129.965 36.940 130.325 ;
        RECT 29.895 129.570 30.240 129.965 ;
        RECT 35.350 129.955 35.890 129.965 ;
        RECT 37.500 129.570 39.240 130.325 ;
        RECT 20.555 119.130 21.095 129.570 ;
        RECT 13.520 118.730 23.800 119.130 ;
        RECT 27.120 118.730 37.400 119.130 ;
        RECT 38.640 118.730 39.240 129.570 ;
        RECT 61.240 129.965 67.690 130.325 ;
        RECT 68.250 129.965 70.485 130.325 ;
        RECT 74.335 130.325 74.645 130.575 ;
        RECT 76.190 130.325 76.535 130.695 ;
        RECT 98.395 130.325 98.740 130.695 ;
        RECT 100.905 130.470 104.585 133.750 ;
        RECT 100.905 130.325 101.635 130.470 ;
        RECT 74.335 129.965 75.630 130.325 ;
        RECT 76.190 129.965 80.460 130.325 ;
        RECT 61.240 119.130 62.175 129.965 ;
        RECT 67.345 129.570 67.690 129.965 ;
        RECT 69.815 129.960 70.485 129.965 ;
        RECT 76.190 129.570 76.535 129.965 ;
        RECT 79.790 119.130 80.460 129.965 ;
        RECT 93.825 129.965 98.740 130.325 ;
        RECT 99.300 129.965 101.635 130.325 ;
        RECT 93.825 119.130 94.710 129.965 ;
        RECT 98.395 129.570 98.740 129.965 ;
        RECT 100.905 129.940 101.635 129.965 ;
        RECT 104.030 130.325 104.585 130.470 ;
        RECT 106.950 130.325 107.295 130.695 ;
        RECT 120.050 130.445 120.380 135.620 ;
        RECT 104.030 129.965 106.390 130.325 ;
        RECT 106.950 129.995 108.250 130.325 ;
        RECT 120.020 130.065 120.405 130.445 ;
        RECT 133.085 130.325 133.430 130.695 ;
        RECT 135.795 130.470 139.475 133.750 ;
        RECT 166.205 131.045 170.485 135.855 ;
        RECT 165.735 130.940 170.485 131.045 ;
        RECT 135.795 130.325 136.350 130.470 ;
        RECT 104.030 129.950 104.585 129.965 ;
        RECT 106.945 129.570 108.250 129.995 ;
        RECT 101.790 122.320 103.155 122.440 ;
        RECT 101.675 120.960 106.625 122.320 ;
        RECT 101.675 120.955 103.155 120.960 ;
        RECT 40.720 118.730 51.000 119.130 ;
        RECT 54.320 118.730 64.600 119.130 ;
        RECT 13.520 117.930 64.600 118.730 ;
        RECT 13.520 114.390 23.800 117.930 ;
        RECT 27.120 114.390 37.400 117.930 ;
        RECT 40.720 114.390 51.000 117.930 ;
        RECT 54.320 114.390 64.600 117.930 ;
        RECT 13.520 113.590 64.600 114.390 ;
        RECT 13.520 110.050 23.800 113.590 ;
        RECT 27.120 110.050 37.400 113.590 ;
        RECT 40.720 110.050 51.000 113.590 ;
        RECT 54.320 110.050 64.600 113.590 ;
        RECT 13.520 109.250 64.600 110.050 ;
        RECT 13.520 108.850 23.800 109.250 ;
        RECT 27.120 108.850 37.400 109.250 ;
        RECT 40.720 108.850 51.000 109.250 ;
        RECT 54.320 108.850 64.600 109.250 ;
        RECT 72.860 118.730 83.140 119.130 ;
        RECT 86.460 118.730 96.740 119.130 ;
        RECT 72.860 117.930 96.740 118.730 ;
        RECT 72.860 114.390 83.140 117.930 ;
        RECT 86.460 114.390 96.740 117.930 ;
        RECT 72.860 113.590 96.740 114.390 ;
        RECT 72.860 110.050 83.140 113.590 ;
        RECT 86.460 110.050 96.740 113.590 ;
        RECT 72.860 109.250 96.740 110.050 ;
        RECT 72.860 108.850 83.140 109.250 ;
        RECT 86.460 108.850 96.740 109.250 ;
        RECT 13.920 105.530 14.720 108.850 ;
        RECT 18.260 105.530 19.060 108.850 ;
        RECT 22.600 105.530 23.400 108.850 ;
        RECT 27.520 105.530 28.320 108.850 ;
        RECT 31.860 105.530 32.660 108.850 ;
        RECT 36.200 105.530 37.000 108.850 ;
        RECT 41.120 105.530 41.920 108.850 ;
        RECT 45.460 105.530 46.260 108.850 ;
        RECT 49.800 105.530 50.600 108.850 ;
        RECT 54.720 105.530 55.520 108.850 ;
        RECT 59.060 105.530 59.860 108.850 ;
        RECT 63.400 105.530 64.200 108.850 ;
        RECT 73.260 105.530 74.060 108.850 ;
        RECT 77.600 105.530 78.400 108.850 ;
        RECT 81.940 105.530 82.740 108.850 ;
        RECT 86.860 105.530 87.660 108.850 ;
        RECT 91.200 105.530 92.000 108.850 ;
        RECT 95.540 105.530 96.340 108.850 ;
        RECT 101.795 107.180 103.155 120.955 ;
        RECT 107.625 119.120 108.250 129.570 ;
        RECT 132.130 129.995 133.430 130.325 ;
        RECT 132.130 129.570 133.435 129.995 ;
        RECT 133.990 129.965 136.350 130.325 ;
        RECT 135.795 129.950 136.350 129.965 ;
        RECT 138.745 130.325 139.475 130.470 ;
        RECT 141.640 130.325 141.985 130.695 ;
        RECT 163.845 130.325 164.190 130.695 ;
        RECT 165.735 130.575 170.565 130.940 ;
        RECT 204.660 130.790 208.340 133.840 ;
        RECT 204.660 130.780 208.350 130.790 ;
        RECT 165.735 130.325 166.045 130.575 ;
        RECT 138.745 129.965 141.080 130.325 ;
        RECT 141.640 129.965 146.555 130.325 ;
        RECT 138.745 129.940 139.475 129.965 ;
        RECT 141.640 129.570 141.985 129.965 ;
        RECT 113.310 128.710 118.260 129.210 ;
        RECT 122.180 128.710 127.070 129.210 ;
        RECT 113.310 119.120 113.910 128.710 ;
        RECT 115.195 120.960 118.475 122.320 ;
        RECT 104.995 118.720 115.275 119.120 ;
        RECT 104.990 117.920 115.275 118.720 ;
        RECT 104.995 114.380 115.275 117.920 ;
        RECT 104.990 113.580 115.275 114.380 ;
        RECT 104.995 110.040 115.275 113.580 ;
        RECT 104.990 109.240 115.275 110.040 ;
        RECT 104.995 108.840 115.275 109.240 ;
        RECT 101.790 106.250 103.155 107.180 ;
        RECT 13.520 105.130 23.800 105.530 ;
        RECT 27.120 105.130 37.400 105.530 ;
        RECT 40.720 105.130 51.000 105.530 ;
        RECT 54.320 105.130 64.600 105.530 ;
        RECT 13.520 104.330 64.600 105.130 ;
        RECT 13.520 100.790 23.800 104.330 ;
        RECT 27.120 100.790 37.400 104.330 ;
        RECT 40.720 100.790 51.000 104.330 ;
        RECT 54.320 100.790 64.600 104.330 ;
        RECT 13.520 99.990 64.600 100.790 ;
        RECT 13.520 96.450 23.800 99.990 ;
        RECT 27.120 96.450 37.400 99.990 ;
        RECT 40.720 96.450 51.000 99.990 ;
        RECT 54.320 96.450 64.600 99.990 ;
        RECT 13.520 95.650 64.600 96.450 ;
        RECT 13.520 95.250 23.800 95.650 ;
        RECT 27.120 95.250 37.400 95.650 ;
        RECT 40.720 95.250 51.000 95.650 ;
        RECT 54.320 95.250 64.600 95.650 ;
        RECT 72.860 105.130 83.140 105.530 ;
        RECT 86.460 105.130 96.740 105.530 ;
        RECT 72.860 104.330 96.740 105.130 ;
        RECT 72.860 100.790 83.140 104.330 ;
        RECT 86.460 100.790 96.740 104.330 ;
        RECT 72.860 99.990 96.740 100.790 ;
        RECT 72.860 96.450 83.140 99.990 ;
        RECT 86.460 96.450 96.740 99.990 ;
        RECT 72.860 95.650 96.740 96.450 ;
        RECT 72.860 95.250 83.140 95.650 ;
        RECT 86.460 95.250 96.740 95.650 ;
        RECT 13.920 91.930 14.720 95.250 ;
        RECT 18.260 91.930 19.060 95.250 ;
        RECT 22.600 91.930 23.400 95.250 ;
        RECT 27.520 91.930 28.320 95.250 ;
        RECT 31.860 91.930 32.660 95.250 ;
        RECT 36.200 91.930 37.000 95.250 ;
        RECT 41.120 91.930 41.920 95.250 ;
        RECT 45.460 91.930 46.260 95.250 ;
        RECT 49.800 91.930 50.600 95.250 ;
        RECT 54.720 91.930 55.520 95.250 ;
        RECT 59.060 91.930 59.860 95.250 ;
        RECT 63.400 91.930 64.200 95.250 ;
        RECT 73.260 91.930 74.060 95.250 ;
        RECT 77.600 91.930 78.400 95.250 ;
        RECT 81.940 91.930 82.740 95.250 ;
        RECT 86.860 91.930 87.660 95.250 ;
        RECT 91.200 91.930 92.000 95.250 ;
        RECT 95.540 91.930 96.340 95.250 ;
        RECT 101.795 94.510 103.155 106.250 ;
        RECT 105.395 105.520 106.195 108.840 ;
        RECT 109.735 105.520 110.535 108.840 ;
        RECT 114.075 105.520 114.875 108.840 ;
        RECT 117.115 107.180 118.475 120.960 ;
        RECT 117.110 106.250 118.475 107.180 ;
        RECT 104.995 95.240 115.275 105.520 ;
        RECT 101.795 93.580 103.160 94.510 ;
        RECT 101.790 92.650 103.155 93.580 ;
        RECT 13.520 91.530 23.800 91.930 ;
        RECT 27.120 91.530 37.400 91.930 ;
        RECT 40.720 91.530 51.000 91.930 ;
        RECT 54.320 91.530 64.600 91.930 ;
        RECT 13.520 90.730 64.600 91.530 ;
        RECT 13.520 87.190 23.800 90.730 ;
        RECT 27.120 87.190 37.400 90.730 ;
        RECT 40.720 87.190 51.000 90.730 ;
        RECT 54.320 87.190 64.600 90.730 ;
        RECT 13.520 86.390 64.600 87.190 ;
        RECT 13.520 82.850 23.800 86.390 ;
        RECT 27.120 82.850 37.400 86.390 ;
        RECT 40.720 82.850 51.000 86.390 ;
        RECT 54.320 82.850 64.600 86.390 ;
        RECT 13.520 82.050 64.600 82.850 ;
        RECT 13.520 81.650 23.800 82.050 ;
        RECT 27.120 81.650 37.400 82.050 ;
        RECT 40.720 81.650 51.000 82.050 ;
        RECT 54.320 81.650 64.600 82.050 ;
        RECT 72.860 91.530 83.140 91.930 ;
        RECT 86.460 91.530 96.740 91.930 ;
        RECT 72.860 90.730 96.740 91.530 ;
        RECT 72.860 87.190 83.140 90.730 ;
        RECT 86.460 87.190 96.740 90.730 ;
        RECT 72.860 86.390 96.740 87.190 ;
        RECT 72.860 82.850 83.140 86.390 ;
        RECT 86.460 82.850 96.740 86.390 ;
        RECT 72.860 82.050 96.740 82.850 ;
        RECT 72.860 81.650 83.140 82.050 ;
        RECT 86.460 81.650 96.740 82.050 ;
        RECT 13.920 78.330 14.720 81.650 ;
        RECT 18.260 78.330 19.060 81.650 ;
        RECT 22.600 78.330 23.400 81.650 ;
        RECT 27.520 78.330 28.320 81.650 ;
        RECT 31.860 78.330 32.660 81.650 ;
        RECT 36.200 78.330 37.000 81.650 ;
        RECT 41.120 78.330 41.920 81.650 ;
        RECT 45.460 78.330 46.260 81.650 ;
        RECT 49.800 78.330 50.600 81.650 ;
        RECT 54.720 78.330 55.520 81.650 ;
        RECT 59.060 78.330 59.860 81.650 ;
        RECT 63.400 78.330 64.200 81.650 ;
        RECT 73.260 78.330 74.060 81.650 ;
        RECT 77.600 78.330 78.400 81.650 ;
        RECT 81.940 78.330 82.740 81.650 ;
        RECT 86.860 78.330 87.660 81.650 ;
        RECT 91.200 78.330 92.000 81.650 ;
        RECT 95.540 78.330 96.340 81.650 ;
        RECT 101.795 80.910 103.155 92.650 ;
        RECT 105.395 91.920 106.195 95.240 ;
        RECT 109.735 91.920 110.535 95.240 ;
        RECT 114.075 91.920 114.875 95.240 ;
        RECT 117.115 94.510 118.475 106.250 ;
        RECT 121.905 120.960 125.185 122.320 ;
        RECT 121.905 107.180 123.265 120.960 ;
        RECT 126.470 119.120 127.070 128.710 ;
        RECT 132.130 119.120 132.755 129.570 ;
        RECT 137.225 122.320 138.590 122.440 ;
        RECT 133.755 120.960 138.705 122.320 ;
        RECT 137.225 120.955 138.705 120.960 ;
        RECT 125.105 118.720 135.385 119.120 ;
        RECT 125.105 117.920 135.390 118.720 ;
        RECT 125.105 114.380 135.385 117.920 ;
        RECT 125.105 113.580 135.390 114.380 ;
        RECT 125.105 110.040 135.385 113.580 ;
        RECT 125.105 109.240 135.390 110.040 ;
        RECT 125.105 108.840 135.385 109.240 ;
        RECT 121.905 106.250 123.270 107.180 ;
        RECT 121.905 94.510 123.265 106.250 ;
        RECT 125.505 105.520 126.305 108.840 ;
        RECT 129.845 105.520 130.645 108.840 ;
        RECT 134.185 105.520 134.985 108.840 ;
        RECT 137.225 107.180 138.585 120.955 ;
        RECT 145.670 119.130 146.555 129.965 ;
        RECT 159.920 129.965 164.190 130.325 ;
        RECT 164.750 129.965 166.045 130.325 ;
        RECT 169.895 130.325 170.565 130.575 ;
        RECT 172.690 130.325 173.035 130.695 ;
        RECT 202.535 130.325 202.880 130.695 ;
        RECT 204.490 130.560 208.350 130.780 ;
        RECT 204.490 130.325 205.030 130.560 ;
        RECT 169.895 129.965 172.130 130.325 ;
        RECT 172.690 129.965 179.140 130.325 ;
        RECT 159.920 119.130 160.590 129.965 ;
        RECT 163.845 129.570 164.190 129.965 ;
        RECT 169.895 129.960 170.565 129.965 ;
        RECT 172.690 129.570 173.035 129.965 ;
        RECT 178.205 119.130 179.140 129.965 ;
        RECT 201.140 129.570 202.880 130.325 ;
        RECT 203.440 129.965 205.030 130.325 ;
        RECT 207.795 130.325 208.350 130.560 ;
        RECT 210.140 130.325 210.485 130.695 ;
        RECT 210.810 130.325 211.180 155.410 ;
        RECT 222.925 135.820 223.445 136.340 ;
        RECT 223.925 135.820 224.445 136.340 ;
        RECT 224.925 135.820 225.445 136.340 ;
        RECT 225.925 135.820 226.445 136.340 ;
        RECT 226.925 135.820 227.445 136.340 ;
        RECT 227.925 135.820 228.445 136.340 ;
        RECT 228.925 135.820 229.445 136.340 ;
        RECT 222.925 134.820 223.445 135.340 ;
        RECT 228.925 134.820 229.445 135.340 ;
        RECT 222.925 133.820 223.445 134.340 ;
        RECT 228.925 133.820 229.445 134.340 ;
        RECT 222.925 132.820 223.445 133.340 ;
        RECT 228.925 132.820 229.445 133.340 ;
        RECT 222.925 131.820 223.445 132.340 ;
        RECT 228.925 131.820 229.445 132.340 ;
        RECT 222.925 131.090 223.445 131.340 ;
        RECT 222.675 130.820 223.445 131.090 ;
        RECT 223.925 130.820 224.445 131.340 ;
        RECT 224.925 130.820 225.445 131.340 ;
        RECT 225.925 130.820 226.445 131.340 ;
        RECT 226.925 130.820 227.445 131.340 ;
        RECT 227.925 131.335 228.445 131.340 ;
        RECT 228.925 131.335 229.445 131.340 ;
        RECT 227.925 130.820 230.085 131.335 ;
        RECT 220.385 130.325 220.730 130.695 ;
        RECT 222.675 130.325 223.410 130.820 ;
        RECT 207.795 129.965 209.580 130.325 ;
        RECT 210.140 129.965 211.180 130.325 ;
        RECT 204.490 129.955 205.030 129.965 ;
        RECT 210.140 129.570 210.485 129.965 ;
        RECT 219.285 129.570 220.730 130.325 ;
        RECT 221.290 129.965 223.410 130.325 ;
        RECT 228.195 130.325 230.085 130.820 ;
        RECT 231.440 130.325 231.785 130.695 ;
        RECT 228.195 129.965 230.880 130.325 ;
        RECT 231.440 129.965 232.110 130.325 ;
        RECT 228.195 129.880 230.085 129.965 ;
        RECT 231.440 129.570 231.785 129.965 ;
        RECT 143.640 118.730 153.920 119.130 ;
        RECT 157.240 118.730 167.520 119.130 ;
        RECT 143.640 117.930 167.520 118.730 ;
        RECT 143.640 114.390 153.920 117.930 ;
        RECT 157.240 114.390 167.520 117.930 ;
        RECT 143.640 113.590 167.520 114.390 ;
        RECT 143.640 110.050 153.920 113.590 ;
        RECT 157.240 110.050 167.520 113.590 ;
        RECT 143.640 109.250 167.520 110.050 ;
        RECT 143.640 108.850 153.920 109.250 ;
        RECT 157.240 108.850 167.520 109.250 ;
        RECT 175.780 118.730 186.060 119.130 ;
        RECT 189.380 118.730 199.660 119.130 ;
        RECT 201.140 118.730 201.740 129.570 ;
        RECT 219.285 119.130 219.825 129.570 ;
        RECT 202.980 118.730 213.260 119.130 ;
        RECT 216.580 118.730 226.860 119.130 ;
        RECT 175.780 117.930 226.860 118.730 ;
        RECT 175.780 114.390 186.060 117.930 ;
        RECT 189.380 114.390 199.660 117.930 ;
        RECT 202.980 114.390 213.260 117.930 ;
        RECT 216.580 114.390 226.860 117.930 ;
        RECT 175.780 113.590 226.860 114.390 ;
        RECT 175.780 110.050 186.060 113.590 ;
        RECT 189.380 110.050 199.660 113.590 ;
        RECT 202.980 110.050 213.260 113.590 ;
        RECT 216.580 110.050 226.860 113.590 ;
        RECT 175.780 109.250 226.860 110.050 ;
        RECT 175.780 108.850 186.060 109.250 ;
        RECT 189.380 108.850 199.660 109.250 ;
        RECT 202.980 108.850 213.260 109.250 ;
        RECT 216.580 108.850 226.860 109.250 ;
        RECT 137.225 106.250 138.590 107.180 ;
        RECT 125.105 95.240 135.385 105.520 ;
        RECT 117.115 93.580 118.480 94.510 ;
        RECT 121.900 93.580 123.265 94.510 ;
        RECT 117.110 92.650 118.475 93.580 ;
        RECT 104.995 81.640 115.275 91.920 ;
        RECT 101.795 79.980 103.160 80.910 ;
        RECT 101.790 79.050 103.155 79.980 ;
        RECT 13.520 77.930 23.800 78.330 ;
        RECT 27.120 77.930 37.400 78.330 ;
        RECT 40.720 77.930 51.000 78.330 ;
        RECT 54.320 77.930 64.600 78.330 ;
        RECT 13.520 77.130 64.600 77.930 ;
        RECT 13.520 73.590 23.800 77.130 ;
        RECT 27.120 73.590 37.400 77.130 ;
        RECT 40.720 73.590 51.000 77.130 ;
        RECT 54.320 73.590 64.600 77.130 ;
        RECT 13.520 72.790 64.600 73.590 ;
        RECT 13.520 69.250 23.800 72.790 ;
        RECT 27.120 69.250 37.400 72.790 ;
        RECT 40.720 69.250 51.000 72.790 ;
        RECT 54.320 69.250 64.600 72.790 ;
        RECT 13.520 68.450 64.600 69.250 ;
        RECT 13.520 68.050 23.800 68.450 ;
        RECT 27.120 68.050 37.400 68.450 ;
        RECT 40.720 68.050 51.000 68.450 ;
        RECT 54.320 68.050 64.600 68.450 ;
        RECT 72.860 77.930 83.140 78.330 ;
        RECT 86.460 77.930 96.740 78.330 ;
        RECT 72.860 77.130 96.740 77.930 ;
        RECT 72.860 73.590 83.140 77.130 ;
        RECT 86.460 73.590 96.740 77.130 ;
        RECT 72.860 72.790 96.740 73.590 ;
        RECT 72.860 69.250 83.140 72.790 ;
        RECT 86.460 69.250 96.740 72.790 ;
        RECT 72.860 68.450 96.740 69.250 ;
        RECT 72.860 68.050 83.140 68.450 ;
        RECT 86.460 68.050 96.740 68.450 ;
        RECT 13.920 64.730 14.720 68.050 ;
        RECT 18.260 64.730 19.060 68.050 ;
        RECT 22.600 64.730 23.400 68.050 ;
        RECT 27.520 64.730 28.320 68.050 ;
        RECT 31.860 64.730 32.660 68.050 ;
        RECT 36.200 64.730 37.000 68.050 ;
        RECT 41.120 64.730 41.920 68.050 ;
        RECT 45.460 64.730 46.260 68.050 ;
        RECT 49.800 64.730 50.600 68.050 ;
        RECT 54.720 64.730 55.520 68.050 ;
        RECT 59.060 64.730 59.860 68.050 ;
        RECT 63.400 64.730 64.200 68.050 ;
        RECT 73.260 64.730 74.060 68.050 ;
        RECT 77.600 64.730 78.400 68.050 ;
        RECT 81.940 64.730 82.740 68.050 ;
        RECT 86.860 64.730 87.660 68.050 ;
        RECT 91.200 64.730 92.000 68.050 ;
        RECT 95.540 64.730 96.340 68.050 ;
        RECT 101.795 67.310 103.155 79.050 ;
        RECT 105.395 78.320 106.195 81.640 ;
        RECT 109.735 78.320 110.535 81.640 ;
        RECT 114.075 78.320 114.875 81.640 ;
        RECT 117.115 80.910 118.475 92.650 ;
        RECT 121.905 92.650 123.270 93.580 ;
        RECT 121.905 80.910 123.265 92.650 ;
        RECT 125.505 91.920 126.305 95.240 ;
        RECT 129.845 91.920 130.645 95.240 ;
        RECT 134.185 91.920 134.985 95.240 ;
        RECT 137.225 94.510 138.585 106.250 ;
        RECT 144.040 105.530 144.840 108.850 ;
        RECT 148.380 105.530 149.180 108.850 ;
        RECT 152.720 105.530 153.520 108.850 ;
        RECT 157.640 105.530 158.440 108.850 ;
        RECT 161.980 105.530 162.780 108.850 ;
        RECT 166.320 105.530 167.120 108.850 ;
        RECT 176.180 105.530 176.980 108.850 ;
        RECT 180.520 105.530 181.320 108.850 ;
        RECT 184.860 105.530 185.660 108.850 ;
        RECT 189.780 105.530 190.580 108.850 ;
        RECT 194.120 105.530 194.920 108.850 ;
        RECT 198.460 105.530 199.260 108.850 ;
        RECT 203.380 105.530 204.180 108.850 ;
        RECT 207.720 105.530 208.520 108.850 ;
        RECT 212.060 105.530 212.860 108.850 ;
        RECT 216.980 105.530 217.780 108.850 ;
        RECT 221.320 105.530 222.120 108.850 ;
        RECT 225.660 105.530 226.460 108.850 ;
        RECT 143.640 105.130 153.920 105.530 ;
        RECT 157.240 105.130 167.520 105.530 ;
        RECT 143.640 104.330 167.520 105.130 ;
        RECT 143.640 100.790 153.920 104.330 ;
        RECT 157.240 100.790 167.520 104.330 ;
        RECT 143.640 99.990 167.520 100.790 ;
        RECT 143.640 96.450 153.920 99.990 ;
        RECT 157.240 96.450 167.520 99.990 ;
        RECT 143.640 95.650 167.520 96.450 ;
        RECT 143.640 95.250 153.920 95.650 ;
        RECT 157.240 95.250 167.520 95.650 ;
        RECT 175.780 105.130 186.060 105.530 ;
        RECT 189.380 105.130 199.660 105.530 ;
        RECT 202.980 105.130 213.260 105.530 ;
        RECT 216.580 105.130 226.860 105.530 ;
        RECT 175.780 104.330 226.860 105.130 ;
        RECT 175.780 100.790 186.060 104.330 ;
        RECT 189.380 100.790 199.660 104.330 ;
        RECT 202.980 100.790 213.260 104.330 ;
        RECT 216.580 100.790 226.860 104.330 ;
        RECT 175.780 99.990 226.860 100.790 ;
        RECT 175.780 96.450 186.060 99.990 ;
        RECT 189.380 96.450 199.660 99.990 ;
        RECT 202.980 96.450 213.260 99.990 ;
        RECT 216.580 96.450 226.860 99.990 ;
        RECT 175.780 95.650 226.860 96.450 ;
        RECT 175.780 95.250 186.060 95.650 ;
        RECT 189.380 95.250 199.660 95.650 ;
        RECT 202.980 95.250 213.260 95.650 ;
        RECT 216.580 95.250 226.860 95.650 ;
        RECT 137.220 93.580 138.585 94.510 ;
        RECT 137.225 92.650 138.590 93.580 ;
        RECT 125.105 81.640 135.385 91.920 ;
        RECT 117.115 79.980 118.480 80.910 ;
        RECT 121.900 79.980 123.265 80.910 ;
        RECT 117.110 79.050 118.475 79.980 ;
        RECT 104.995 68.040 115.275 78.320 ;
        RECT 101.795 66.380 103.160 67.310 ;
        RECT 101.790 65.450 103.155 66.380 ;
        RECT 13.520 64.330 23.800 64.730 ;
        RECT 27.120 64.330 37.400 64.730 ;
        RECT 40.720 64.330 51.000 64.730 ;
        RECT 54.320 64.330 64.600 64.730 ;
        RECT 13.520 63.530 64.600 64.330 ;
        RECT 13.520 59.990 23.800 63.530 ;
        RECT 27.120 59.990 37.400 63.530 ;
        RECT 40.720 59.990 51.000 63.530 ;
        RECT 54.320 59.990 64.600 63.530 ;
        RECT 13.520 59.190 64.600 59.990 ;
        RECT 13.520 55.650 23.800 59.190 ;
        RECT 27.120 55.650 37.400 59.190 ;
        RECT 40.720 55.650 51.000 59.190 ;
        RECT 54.320 55.650 64.600 59.190 ;
        RECT 13.520 54.850 64.600 55.650 ;
        RECT 13.520 54.450 23.800 54.850 ;
        RECT 27.120 54.450 37.400 54.850 ;
        RECT 40.720 54.450 51.000 54.850 ;
        RECT 54.320 54.450 64.600 54.850 ;
        RECT 72.860 64.330 83.140 64.730 ;
        RECT 86.460 64.330 96.740 64.730 ;
        RECT 72.860 63.530 96.740 64.330 ;
        RECT 72.860 59.990 83.140 63.530 ;
        RECT 86.460 59.990 96.740 63.530 ;
        RECT 72.860 59.190 96.740 59.990 ;
        RECT 72.860 55.650 83.140 59.190 ;
        RECT 86.460 55.650 96.740 59.190 ;
        RECT 72.860 54.850 96.740 55.650 ;
        RECT 72.860 54.450 83.140 54.850 ;
        RECT 86.460 54.450 96.740 54.850 ;
        RECT 13.920 51.130 14.720 54.450 ;
        RECT 18.260 51.130 19.060 54.450 ;
        RECT 22.600 51.130 23.400 54.450 ;
        RECT 27.520 51.130 28.320 54.450 ;
        RECT 31.860 51.130 32.660 54.450 ;
        RECT 36.200 51.130 37.000 54.450 ;
        RECT 41.120 51.130 41.920 54.450 ;
        RECT 45.460 51.130 46.260 54.450 ;
        RECT 49.800 51.130 50.600 54.450 ;
        RECT 54.720 51.130 55.520 54.450 ;
        RECT 59.060 51.130 59.860 54.450 ;
        RECT 63.400 51.130 64.200 54.450 ;
        RECT 73.260 51.130 74.060 54.450 ;
        RECT 77.600 51.130 78.400 54.450 ;
        RECT 81.940 51.130 82.740 54.450 ;
        RECT 86.860 51.130 87.660 54.450 ;
        RECT 91.200 51.130 92.000 54.450 ;
        RECT 95.540 51.130 96.340 54.450 ;
        RECT 101.795 53.710 103.155 65.450 ;
        RECT 105.395 64.720 106.195 68.040 ;
        RECT 109.735 64.720 110.535 68.040 ;
        RECT 114.075 64.720 114.875 68.040 ;
        RECT 117.115 67.310 118.475 79.050 ;
        RECT 121.905 79.050 123.270 79.980 ;
        RECT 121.905 67.310 123.265 79.050 ;
        RECT 125.505 78.320 126.305 81.640 ;
        RECT 129.845 78.320 130.645 81.640 ;
        RECT 134.185 78.320 134.985 81.640 ;
        RECT 137.225 80.910 138.585 92.650 ;
        RECT 144.040 91.930 144.840 95.250 ;
        RECT 148.380 91.930 149.180 95.250 ;
        RECT 152.720 91.930 153.520 95.250 ;
        RECT 157.640 91.930 158.440 95.250 ;
        RECT 161.980 91.930 162.780 95.250 ;
        RECT 166.320 91.930 167.120 95.250 ;
        RECT 176.180 91.930 176.980 95.250 ;
        RECT 180.520 91.930 181.320 95.250 ;
        RECT 184.860 91.930 185.660 95.250 ;
        RECT 189.780 91.930 190.580 95.250 ;
        RECT 194.120 91.930 194.920 95.250 ;
        RECT 198.460 91.930 199.260 95.250 ;
        RECT 203.380 91.930 204.180 95.250 ;
        RECT 207.720 91.930 208.520 95.250 ;
        RECT 212.060 91.930 212.860 95.250 ;
        RECT 216.980 91.930 217.780 95.250 ;
        RECT 221.320 91.930 222.120 95.250 ;
        RECT 225.660 91.930 226.460 95.250 ;
        RECT 143.640 91.530 153.920 91.930 ;
        RECT 157.240 91.530 167.520 91.930 ;
        RECT 143.640 90.730 167.520 91.530 ;
        RECT 143.640 87.190 153.920 90.730 ;
        RECT 157.240 87.190 167.520 90.730 ;
        RECT 143.640 86.390 167.520 87.190 ;
        RECT 143.640 82.850 153.920 86.390 ;
        RECT 157.240 82.850 167.520 86.390 ;
        RECT 143.640 82.050 167.520 82.850 ;
        RECT 143.640 81.650 153.920 82.050 ;
        RECT 157.240 81.650 167.520 82.050 ;
        RECT 175.780 91.530 186.060 91.930 ;
        RECT 189.380 91.530 199.660 91.930 ;
        RECT 202.980 91.530 213.260 91.930 ;
        RECT 216.580 91.530 226.860 91.930 ;
        RECT 175.780 90.730 226.860 91.530 ;
        RECT 175.780 87.190 186.060 90.730 ;
        RECT 189.380 87.190 199.660 90.730 ;
        RECT 202.980 87.190 213.260 90.730 ;
        RECT 216.580 87.190 226.860 90.730 ;
        RECT 175.780 86.390 226.860 87.190 ;
        RECT 175.780 82.850 186.060 86.390 ;
        RECT 189.380 82.850 199.660 86.390 ;
        RECT 202.980 82.850 213.260 86.390 ;
        RECT 216.580 82.850 226.860 86.390 ;
        RECT 175.780 82.050 226.860 82.850 ;
        RECT 175.780 81.650 186.060 82.050 ;
        RECT 189.380 81.650 199.660 82.050 ;
        RECT 202.980 81.650 213.260 82.050 ;
        RECT 216.580 81.650 226.860 82.050 ;
        RECT 137.220 79.980 138.585 80.910 ;
        RECT 137.225 79.050 138.590 79.980 ;
        RECT 125.105 68.040 135.385 78.320 ;
        RECT 117.115 66.380 118.480 67.310 ;
        RECT 121.900 66.380 123.265 67.310 ;
        RECT 117.110 65.450 118.475 66.380 ;
        RECT 104.995 54.440 115.275 64.720 ;
        RECT 101.795 52.780 103.160 53.710 ;
        RECT 101.790 51.850 103.155 52.780 ;
        RECT 13.520 50.730 23.800 51.130 ;
        RECT 27.120 50.730 37.400 51.130 ;
        RECT 40.720 50.730 51.000 51.130 ;
        RECT 54.320 50.730 64.600 51.130 ;
        RECT 13.520 49.930 64.600 50.730 ;
        RECT 13.520 46.390 23.800 49.930 ;
        RECT 27.120 46.390 37.400 49.930 ;
        RECT 40.720 46.390 51.000 49.930 ;
        RECT 54.320 46.390 64.600 49.930 ;
        RECT 13.520 45.590 64.600 46.390 ;
        RECT 13.520 42.050 23.800 45.590 ;
        RECT 27.120 42.050 37.400 45.590 ;
        RECT 40.720 42.050 51.000 45.590 ;
        RECT 54.320 42.050 64.600 45.590 ;
        RECT 13.520 41.250 64.600 42.050 ;
        RECT 13.520 40.850 23.800 41.250 ;
        RECT 27.120 40.850 37.400 41.250 ;
        RECT 40.720 40.850 51.000 41.250 ;
        RECT 54.320 40.850 64.600 41.250 ;
        RECT 72.860 50.730 83.140 51.130 ;
        RECT 86.460 50.730 96.740 51.130 ;
        RECT 72.860 49.930 96.740 50.730 ;
        RECT 72.860 46.390 83.140 49.930 ;
        RECT 86.460 46.390 96.740 49.930 ;
        RECT 72.860 45.590 96.740 46.390 ;
        RECT 72.860 42.050 83.140 45.590 ;
        RECT 86.460 42.050 96.740 45.590 ;
        RECT 72.860 41.250 96.740 42.050 ;
        RECT 72.860 40.850 83.140 41.250 ;
        RECT 86.460 40.850 96.740 41.250 ;
        RECT 13.920 37.530 14.720 40.850 ;
        RECT 18.260 37.530 19.060 40.850 ;
        RECT 22.600 37.530 23.400 40.850 ;
        RECT 27.520 37.530 28.320 40.850 ;
        RECT 31.860 37.530 32.660 40.850 ;
        RECT 36.200 37.530 37.000 40.850 ;
        RECT 41.120 37.530 41.920 40.850 ;
        RECT 45.460 37.530 46.260 40.850 ;
        RECT 49.800 37.530 50.600 40.850 ;
        RECT 54.720 37.530 55.520 40.850 ;
        RECT 59.060 37.530 59.860 40.850 ;
        RECT 63.400 37.530 64.200 40.850 ;
        RECT 73.260 37.530 74.060 40.850 ;
        RECT 77.600 37.530 78.400 40.850 ;
        RECT 81.940 37.530 82.740 40.850 ;
        RECT 86.860 37.530 87.660 40.850 ;
        RECT 91.200 37.530 92.000 40.850 ;
        RECT 95.540 37.530 96.340 40.850 ;
        RECT 101.795 40.110 103.155 51.850 ;
        RECT 105.395 51.120 106.195 54.440 ;
        RECT 109.735 51.120 110.535 54.440 ;
        RECT 114.075 51.120 114.875 54.440 ;
        RECT 117.115 53.710 118.475 65.450 ;
        RECT 121.905 65.450 123.270 66.380 ;
        RECT 121.905 53.710 123.265 65.450 ;
        RECT 125.505 64.720 126.305 68.040 ;
        RECT 129.845 64.720 130.645 68.040 ;
        RECT 134.185 64.720 134.985 68.040 ;
        RECT 137.225 67.310 138.585 79.050 ;
        RECT 144.040 78.330 144.840 81.650 ;
        RECT 148.380 78.330 149.180 81.650 ;
        RECT 152.720 78.330 153.520 81.650 ;
        RECT 157.640 78.330 158.440 81.650 ;
        RECT 161.980 78.330 162.780 81.650 ;
        RECT 166.320 78.330 167.120 81.650 ;
        RECT 176.180 78.330 176.980 81.650 ;
        RECT 180.520 78.330 181.320 81.650 ;
        RECT 184.860 78.330 185.660 81.650 ;
        RECT 189.780 78.330 190.580 81.650 ;
        RECT 194.120 78.330 194.920 81.650 ;
        RECT 198.460 78.330 199.260 81.650 ;
        RECT 203.380 78.330 204.180 81.650 ;
        RECT 207.720 78.330 208.520 81.650 ;
        RECT 212.060 78.330 212.860 81.650 ;
        RECT 216.980 78.330 217.780 81.650 ;
        RECT 221.320 78.330 222.120 81.650 ;
        RECT 225.660 78.330 226.460 81.650 ;
        RECT 143.640 77.930 153.920 78.330 ;
        RECT 157.240 77.930 167.520 78.330 ;
        RECT 143.640 77.130 167.520 77.930 ;
        RECT 143.640 73.590 153.920 77.130 ;
        RECT 157.240 73.590 167.520 77.130 ;
        RECT 143.640 72.790 167.520 73.590 ;
        RECT 143.640 69.250 153.920 72.790 ;
        RECT 157.240 69.250 167.520 72.790 ;
        RECT 143.640 68.450 167.520 69.250 ;
        RECT 143.640 68.050 153.920 68.450 ;
        RECT 157.240 68.050 167.520 68.450 ;
        RECT 175.780 77.930 186.060 78.330 ;
        RECT 189.380 77.930 199.660 78.330 ;
        RECT 202.980 77.930 213.260 78.330 ;
        RECT 216.580 77.930 226.860 78.330 ;
        RECT 175.780 77.130 226.860 77.930 ;
        RECT 175.780 73.590 186.060 77.130 ;
        RECT 189.380 73.590 199.660 77.130 ;
        RECT 202.980 73.590 213.260 77.130 ;
        RECT 216.580 73.590 226.860 77.130 ;
        RECT 175.780 72.790 226.860 73.590 ;
        RECT 175.780 69.250 186.060 72.790 ;
        RECT 189.380 69.250 199.660 72.790 ;
        RECT 202.980 69.250 213.260 72.790 ;
        RECT 216.580 69.250 226.860 72.790 ;
        RECT 175.780 68.450 226.860 69.250 ;
        RECT 175.780 68.050 186.060 68.450 ;
        RECT 189.380 68.050 199.660 68.450 ;
        RECT 202.980 68.050 213.260 68.450 ;
        RECT 216.580 68.050 226.860 68.450 ;
        RECT 137.220 66.380 138.585 67.310 ;
        RECT 137.225 65.450 138.590 66.380 ;
        RECT 125.105 54.440 135.385 64.720 ;
        RECT 117.115 52.780 118.480 53.710 ;
        RECT 121.900 52.780 123.265 53.710 ;
        RECT 117.110 51.850 118.475 52.780 ;
        RECT 104.995 40.840 115.275 51.120 ;
        RECT 101.795 39.180 103.160 40.110 ;
        RECT 101.790 38.250 103.155 39.180 ;
        RECT 13.520 37.130 23.800 37.530 ;
        RECT 27.120 37.130 37.400 37.530 ;
        RECT 40.720 37.130 51.000 37.530 ;
        RECT 54.320 37.130 64.600 37.530 ;
        RECT 13.520 36.330 64.600 37.130 ;
        RECT 13.520 32.790 23.800 36.330 ;
        RECT 27.120 32.790 37.400 36.330 ;
        RECT 40.720 32.790 51.000 36.330 ;
        RECT 54.320 32.790 64.600 36.330 ;
        RECT 13.520 31.990 64.600 32.790 ;
        RECT 13.520 28.450 23.800 31.990 ;
        RECT 27.120 28.450 37.400 31.990 ;
        RECT 40.720 28.450 51.000 31.990 ;
        RECT 54.320 28.450 64.600 31.990 ;
        RECT 13.520 27.650 64.600 28.450 ;
        RECT 13.520 27.250 23.800 27.650 ;
        RECT 27.120 27.250 37.400 27.650 ;
        RECT 40.720 27.250 51.000 27.650 ;
        RECT 54.320 27.250 64.600 27.650 ;
        RECT 72.860 37.130 83.140 37.530 ;
        RECT 86.460 37.130 96.740 37.530 ;
        RECT 72.860 36.330 96.740 37.130 ;
        RECT 72.860 32.790 83.140 36.330 ;
        RECT 86.460 32.790 96.740 36.330 ;
        RECT 72.860 31.990 96.740 32.790 ;
        RECT 72.860 28.450 83.140 31.990 ;
        RECT 86.460 28.450 96.740 31.990 ;
        RECT 72.860 27.650 96.740 28.450 ;
        RECT 72.860 27.250 83.140 27.650 ;
        RECT 86.460 27.250 96.740 27.650 ;
        RECT 13.920 23.930 14.720 27.250 ;
        RECT 18.260 23.930 19.060 27.250 ;
        RECT 22.600 23.930 23.400 27.250 ;
        RECT 27.520 23.930 28.320 27.250 ;
        RECT 31.860 23.930 32.660 27.250 ;
        RECT 36.200 23.930 37.000 27.250 ;
        RECT 41.120 23.930 41.920 27.250 ;
        RECT 45.460 23.930 46.260 27.250 ;
        RECT 49.800 23.930 50.600 27.250 ;
        RECT 54.720 23.930 55.520 27.250 ;
        RECT 59.060 23.930 59.860 27.250 ;
        RECT 63.400 23.930 64.200 27.250 ;
        RECT 73.260 23.930 74.060 27.250 ;
        RECT 77.600 23.930 78.400 27.250 ;
        RECT 81.940 23.930 82.740 27.250 ;
        RECT 86.860 23.930 87.660 27.250 ;
        RECT 91.200 23.930 92.000 27.250 ;
        RECT 95.540 23.930 96.340 27.250 ;
        RECT 101.795 26.510 103.155 38.250 ;
        RECT 105.395 37.520 106.195 40.840 ;
        RECT 109.735 37.520 110.535 40.840 ;
        RECT 114.075 37.520 114.875 40.840 ;
        RECT 117.115 40.110 118.475 51.850 ;
        RECT 121.905 51.850 123.270 52.780 ;
        RECT 121.905 40.110 123.265 51.850 ;
        RECT 125.505 51.120 126.305 54.440 ;
        RECT 129.845 51.120 130.645 54.440 ;
        RECT 134.185 51.120 134.985 54.440 ;
        RECT 137.225 53.710 138.585 65.450 ;
        RECT 144.040 64.730 144.840 68.050 ;
        RECT 148.380 64.730 149.180 68.050 ;
        RECT 152.720 64.730 153.520 68.050 ;
        RECT 157.640 64.730 158.440 68.050 ;
        RECT 161.980 64.730 162.780 68.050 ;
        RECT 166.320 64.730 167.120 68.050 ;
        RECT 176.180 64.730 176.980 68.050 ;
        RECT 180.520 64.730 181.320 68.050 ;
        RECT 184.860 64.730 185.660 68.050 ;
        RECT 189.780 64.730 190.580 68.050 ;
        RECT 194.120 64.730 194.920 68.050 ;
        RECT 198.460 64.730 199.260 68.050 ;
        RECT 203.380 64.730 204.180 68.050 ;
        RECT 207.720 64.730 208.520 68.050 ;
        RECT 212.060 64.730 212.860 68.050 ;
        RECT 216.980 64.730 217.780 68.050 ;
        RECT 221.320 64.730 222.120 68.050 ;
        RECT 225.660 64.730 226.460 68.050 ;
        RECT 143.640 64.330 153.920 64.730 ;
        RECT 157.240 64.330 167.520 64.730 ;
        RECT 143.640 63.530 167.520 64.330 ;
        RECT 143.640 59.990 153.920 63.530 ;
        RECT 157.240 59.990 167.520 63.530 ;
        RECT 143.640 59.190 167.520 59.990 ;
        RECT 143.640 55.650 153.920 59.190 ;
        RECT 157.240 55.650 167.520 59.190 ;
        RECT 143.640 54.850 167.520 55.650 ;
        RECT 143.640 54.450 153.920 54.850 ;
        RECT 157.240 54.450 167.520 54.850 ;
        RECT 175.780 64.330 186.060 64.730 ;
        RECT 189.380 64.330 199.660 64.730 ;
        RECT 202.980 64.330 213.260 64.730 ;
        RECT 216.580 64.330 226.860 64.730 ;
        RECT 175.780 63.530 226.860 64.330 ;
        RECT 175.780 59.990 186.060 63.530 ;
        RECT 189.380 59.990 199.660 63.530 ;
        RECT 202.980 59.990 213.260 63.530 ;
        RECT 216.580 59.990 226.860 63.530 ;
        RECT 175.780 59.190 226.860 59.990 ;
        RECT 175.780 55.650 186.060 59.190 ;
        RECT 189.380 55.650 199.660 59.190 ;
        RECT 202.980 55.650 213.260 59.190 ;
        RECT 216.580 55.650 226.860 59.190 ;
        RECT 175.780 54.850 226.860 55.650 ;
        RECT 175.780 54.450 186.060 54.850 ;
        RECT 189.380 54.450 199.660 54.850 ;
        RECT 202.980 54.450 213.260 54.850 ;
        RECT 216.580 54.450 226.860 54.850 ;
        RECT 137.220 52.780 138.585 53.710 ;
        RECT 137.225 51.850 138.590 52.780 ;
        RECT 125.105 40.840 135.385 51.120 ;
        RECT 117.115 39.180 118.480 40.110 ;
        RECT 121.900 39.180 123.265 40.110 ;
        RECT 117.110 38.250 118.475 39.180 ;
        RECT 104.995 27.240 115.275 37.520 ;
        RECT 101.795 25.580 103.160 26.510 ;
        RECT 13.520 23.530 23.800 23.930 ;
        RECT 27.120 23.530 37.400 23.930 ;
        RECT 40.720 23.530 51.000 23.930 ;
        RECT 54.320 23.530 64.600 23.930 ;
        RECT 13.520 22.730 64.600 23.530 ;
        RECT 13.520 19.190 23.800 22.730 ;
        RECT 27.120 19.190 37.400 22.730 ;
        RECT 40.720 19.190 51.000 22.730 ;
        RECT 54.320 19.190 64.600 22.730 ;
        RECT 13.520 18.390 64.600 19.190 ;
        RECT 13.520 14.850 23.800 18.390 ;
        RECT 27.120 14.850 37.400 18.390 ;
        RECT 40.720 14.850 51.000 18.390 ;
        RECT 54.320 14.850 64.600 18.390 ;
        RECT 13.520 14.050 64.600 14.850 ;
        RECT 13.520 13.650 23.800 14.050 ;
        RECT 27.120 13.650 37.400 14.050 ;
        RECT 40.720 13.650 51.000 14.050 ;
        RECT 54.320 13.650 64.600 14.050 ;
        RECT 72.860 23.530 83.140 23.930 ;
        RECT 86.460 23.530 96.740 23.930 ;
        RECT 72.860 22.730 96.740 23.530 ;
        RECT 72.860 19.190 83.140 22.730 ;
        RECT 86.460 19.190 96.740 22.730 ;
        RECT 72.860 18.390 96.740 19.190 ;
        RECT 72.860 14.850 83.140 18.390 ;
        RECT 86.460 14.850 96.740 18.390 ;
        RECT 72.860 14.050 96.740 14.850 ;
        RECT 72.860 13.650 83.140 14.050 ;
        RECT 86.460 13.650 96.740 14.050 ;
        RECT 101.795 11.800 103.155 25.580 ;
        RECT 105.395 23.920 106.195 27.240 ;
        RECT 109.735 23.920 110.535 27.240 ;
        RECT 114.075 23.920 114.875 27.240 ;
        RECT 117.115 26.510 118.475 38.250 ;
        RECT 121.905 38.250 123.270 39.180 ;
        RECT 121.905 26.510 123.265 38.250 ;
        RECT 125.505 37.520 126.305 40.840 ;
        RECT 129.845 37.520 130.645 40.840 ;
        RECT 134.185 37.520 134.985 40.840 ;
        RECT 137.225 40.110 138.585 51.850 ;
        RECT 144.040 51.130 144.840 54.450 ;
        RECT 148.380 51.130 149.180 54.450 ;
        RECT 152.720 51.130 153.520 54.450 ;
        RECT 157.640 51.130 158.440 54.450 ;
        RECT 161.980 51.130 162.780 54.450 ;
        RECT 166.320 51.130 167.120 54.450 ;
        RECT 176.180 51.130 176.980 54.450 ;
        RECT 180.520 51.130 181.320 54.450 ;
        RECT 184.860 51.130 185.660 54.450 ;
        RECT 189.780 51.130 190.580 54.450 ;
        RECT 194.120 51.130 194.920 54.450 ;
        RECT 198.460 51.130 199.260 54.450 ;
        RECT 203.380 51.130 204.180 54.450 ;
        RECT 207.720 51.130 208.520 54.450 ;
        RECT 212.060 51.130 212.860 54.450 ;
        RECT 216.980 51.130 217.780 54.450 ;
        RECT 221.320 51.130 222.120 54.450 ;
        RECT 225.660 51.130 226.460 54.450 ;
        RECT 143.640 50.730 153.920 51.130 ;
        RECT 157.240 50.730 167.520 51.130 ;
        RECT 143.640 49.930 167.520 50.730 ;
        RECT 143.640 46.390 153.920 49.930 ;
        RECT 157.240 46.390 167.520 49.930 ;
        RECT 143.640 45.590 167.520 46.390 ;
        RECT 143.640 42.050 153.920 45.590 ;
        RECT 157.240 42.050 167.520 45.590 ;
        RECT 143.640 41.250 167.520 42.050 ;
        RECT 143.640 40.850 153.920 41.250 ;
        RECT 157.240 40.850 167.520 41.250 ;
        RECT 175.780 50.730 186.060 51.130 ;
        RECT 189.380 50.730 199.660 51.130 ;
        RECT 202.980 50.730 213.260 51.130 ;
        RECT 216.580 50.730 226.860 51.130 ;
        RECT 175.780 49.930 226.860 50.730 ;
        RECT 175.780 46.390 186.060 49.930 ;
        RECT 189.380 46.390 199.660 49.930 ;
        RECT 202.980 46.390 213.260 49.930 ;
        RECT 216.580 46.390 226.860 49.930 ;
        RECT 175.780 45.590 226.860 46.390 ;
        RECT 175.780 42.050 186.060 45.590 ;
        RECT 189.380 42.050 199.660 45.590 ;
        RECT 202.980 42.050 213.260 45.590 ;
        RECT 216.580 42.050 226.860 45.590 ;
        RECT 175.780 41.250 226.860 42.050 ;
        RECT 175.780 40.850 186.060 41.250 ;
        RECT 189.380 40.850 199.660 41.250 ;
        RECT 202.980 40.850 213.260 41.250 ;
        RECT 216.580 40.850 226.860 41.250 ;
        RECT 137.220 39.180 138.585 40.110 ;
        RECT 137.225 38.250 138.590 39.180 ;
        RECT 125.105 27.240 135.385 37.520 ;
        RECT 117.115 25.580 118.480 26.510 ;
        RECT 121.900 25.580 123.265 26.510 ;
        RECT 104.995 23.520 115.275 23.920 ;
        RECT 104.995 22.720 115.280 23.520 ;
        RECT 104.995 19.180 115.275 22.720 ;
        RECT 104.995 18.380 115.280 19.180 ;
        RECT 104.995 14.840 115.275 18.380 ;
        RECT 104.995 14.040 115.280 14.840 ;
        RECT 104.995 13.640 115.275 14.040 ;
        RECT 117.115 11.805 118.475 25.580 ;
        RECT 121.905 11.805 123.265 25.580 ;
        RECT 125.505 23.920 126.305 27.240 ;
        RECT 129.845 23.920 130.645 27.240 ;
        RECT 134.185 23.920 134.985 27.240 ;
        RECT 137.225 26.510 138.585 38.250 ;
        RECT 144.040 37.530 144.840 40.850 ;
        RECT 148.380 37.530 149.180 40.850 ;
        RECT 152.720 37.530 153.520 40.850 ;
        RECT 157.640 37.530 158.440 40.850 ;
        RECT 161.980 37.530 162.780 40.850 ;
        RECT 166.320 37.530 167.120 40.850 ;
        RECT 176.180 37.530 176.980 40.850 ;
        RECT 180.520 37.530 181.320 40.850 ;
        RECT 184.860 37.530 185.660 40.850 ;
        RECT 189.780 37.530 190.580 40.850 ;
        RECT 194.120 37.530 194.920 40.850 ;
        RECT 198.460 37.530 199.260 40.850 ;
        RECT 203.380 37.530 204.180 40.850 ;
        RECT 207.720 37.530 208.520 40.850 ;
        RECT 212.060 37.530 212.860 40.850 ;
        RECT 216.980 37.530 217.780 40.850 ;
        RECT 221.320 37.530 222.120 40.850 ;
        RECT 225.660 37.530 226.460 40.850 ;
        RECT 143.640 37.130 153.920 37.530 ;
        RECT 157.240 37.130 167.520 37.530 ;
        RECT 143.640 36.330 167.520 37.130 ;
        RECT 143.640 32.790 153.920 36.330 ;
        RECT 157.240 32.790 167.520 36.330 ;
        RECT 143.640 31.990 167.520 32.790 ;
        RECT 143.640 28.450 153.920 31.990 ;
        RECT 157.240 28.450 167.520 31.990 ;
        RECT 143.640 27.650 167.520 28.450 ;
        RECT 143.640 27.250 153.920 27.650 ;
        RECT 157.240 27.250 167.520 27.650 ;
        RECT 175.780 37.130 186.060 37.530 ;
        RECT 189.380 37.130 199.660 37.530 ;
        RECT 202.980 37.130 213.260 37.530 ;
        RECT 216.580 37.130 226.860 37.530 ;
        RECT 175.780 36.330 226.860 37.130 ;
        RECT 175.780 32.790 186.060 36.330 ;
        RECT 189.380 32.790 199.660 36.330 ;
        RECT 202.980 32.790 213.260 36.330 ;
        RECT 216.580 32.790 226.860 36.330 ;
        RECT 175.780 31.990 226.860 32.790 ;
        RECT 175.780 28.450 186.060 31.990 ;
        RECT 189.380 28.450 199.660 31.990 ;
        RECT 202.980 28.450 213.260 31.990 ;
        RECT 216.580 28.450 226.860 31.990 ;
        RECT 175.780 27.650 226.860 28.450 ;
        RECT 175.780 27.250 186.060 27.650 ;
        RECT 189.380 27.250 199.660 27.650 ;
        RECT 202.980 27.250 213.260 27.650 ;
        RECT 216.580 27.250 226.860 27.650 ;
        RECT 137.220 25.580 138.585 26.510 ;
        RECT 125.105 23.520 135.385 23.920 ;
        RECT 125.100 22.720 135.385 23.520 ;
        RECT 125.105 19.180 135.385 22.720 ;
        RECT 125.100 18.380 135.385 19.180 ;
        RECT 125.105 14.840 135.385 18.380 ;
        RECT 125.100 14.040 135.385 14.840 ;
        RECT 125.105 13.640 135.385 14.040 ;
        RECT 117.115 11.800 118.595 11.805 ;
        RECT 101.795 10.440 105.075 11.800 ;
        RECT 113.645 10.440 118.595 11.800 ;
        RECT 121.785 11.800 123.265 11.805 ;
        RECT 137.225 11.800 138.585 25.580 ;
        RECT 144.040 23.930 144.840 27.250 ;
        RECT 148.380 23.930 149.180 27.250 ;
        RECT 152.720 23.930 153.520 27.250 ;
        RECT 157.640 23.930 158.440 27.250 ;
        RECT 161.980 23.930 162.780 27.250 ;
        RECT 166.320 23.930 167.120 27.250 ;
        RECT 176.180 23.930 176.980 27.250 ;
        RECT 180.520 23.930 181.320 27.250 ;
        RECT 184.860 23.930 185.660 27.250 ;
        RECT 189.780 23.930 190.580 27.250 ;
        RECT 194.120 23.930 194.920 27.250 ;
        RECT 198.460 23.930 199.260 27.250 ;
        RECT 203.380 23.930 204.180 27.250 ;
        RECT 207.720 23.930 208.520 27.250 ;
        RECT 212.060 23.930 212.860 27.250 ;
        RECT 216.980 23.930 217.780 27.250 ;
        RECT 221.320 23.930 222.120 27.250 ;
        RECT 225.660 23.930 226.460 27.250 ;
        RECT 143.640 23.530 153.920 23.930 ;
        RECT 157.240 23.530 167.520 23.930 ;
        RECT 143.640 22.730 167.520 23.530 ;
        RECT 143.640 19.190 153.920 22.730 ;
        RECT 157.240 19.190 167.520 22.730 ;
        RECT 143.640 18.390 167.520 19.190 ;
        RECT 143.640 14.850 153.920 18.390 ;
        RECT 157.240 14.850 167.520 18.390 ;
        RECT 143.640 14.050 167.520 14.850 ;
        RECT 143.640 13.650 153.920 14.050 ;
        RECT 157.240 13.650 167.520 14.050 ;
        RECT 175.780 23.530 186.060 23.930 ;
        RECT 189.380 23.530 199.660 23.930 ;
        RECT 202.980 23.530 213.260 23.930 ;
        RECT 216.580 23.530 226.860 23.930 ;
        RECT 175.780 22.730 226.860 23.530 ;
        RECT 175.780 19.190 186.060 22.730 ;
        RECT 189.380 19.190 199.660 22.730 ;
        RECT 202.980 19.190 213.260 22.730 ;
        RECT 216.580 19.190 226.860 22.730 ;
        RECT 175.780 18.390 226.860 19.190 ;
        RECT 175.780 14.850 186.060 18.390 ;
        RECT 189.380 14.850 199.660 18.390 ;
        RECT 202.980 14.850 213.260 18.390 ;
        RECT 216.580 14.850 226.860 18.390 ;
        RECT 175.780 14.050 226.860 14.850 ;
        RECT 175.780 13.650 186.060 14.050 ;
        RECT 189.380 13.650 199.660 14.050 ;
        RECT 202.980 13.650 213.260 14.050 ;
        RECT 216.580 13.650 226.860 14.050 ;
        RECT 121.785 10.440 126.735 11.800 ;
        RECT 135.305 10.440 138.585 11.800 ;
        RECT 117.115 10.320 118.480 10.440 ;
        RECT 121.900 10.320 123.265 10.440 ;
      LAYER met4 ;
        RECT -0.130 -1.640 253.790 -1.600 ;
      LAYER via4 ;
        RECT 109.655 138.890 110.835 140.075 ;
        RECT 129.545 138.890 130.725 140.075 ;
        RECT 101.795 120.960 106.620 122.320 ;
        RECT 101.795 107.925 103.155 120.960 ;
        RECT 115.200 120.960 118.475 122.320 ;
        RECT 101.795 94.230 103.155 106.250 ;
        RECT 117.115 107.925 118.475 120.960 ;
        RECT 101.795 80.630 103.155 92.650 ;
        RECT 117.115 94.230 118.475 106.250 ;
        RECT 121.905 120.960 125.180 122.320 ;
        RECT 121.905 107.925 123.265 120.960 ;
        RECT 133.760 120.960 138.585 122.320 ;
        RECT 121.905 94.230 123.265 106.250 ;
        RECT 137.225 107.925 138.585 120.960 ;
        RECT 101.795 67.030 103.155 79.050 ;
        RECT 117.115 80.630 118.475 92.650 ;
        RECT 121.905 80.630 123.265 92.650 ;
        RECT 137.225 94.230 138.585 106.250 ;
        RECT 101.795 53.430 103.155 65.450 ;
        RECT 117.115 67.030 118.475 79.050 ;
        RECT 121.905 67.030 123.265 79.050 ;
        RECT 137.225 80.630 138.585 92.650 ;
        RECT 101.795 39.830 103.155 51.850 ;
        RECT 117.115 53.430 118.475 65.450 ;
        RECT 121.905 53.430 123.265 65.450 ;
        RECT 137.225 67.030 138.585 79.050 ;
        RECT 101.795 26.230 103.155 38.250 ;
        RECT 117.115 39.830 118.475 51.850 ;
        RECT 121.905 39.830 123.265 51.850 ;
        RECT 137.225 53.430 138.585 65.450 ;
        RECT 101.795 11.800 103.155 24.835 ;
        RECT 117.115 26.230 118.475 38.250 ;
        RECT 121.905 26.230 123.265 38.250 ;
        RECT 137.225 39.830 138.585 51.850 ;
        RECT 117.115 11.800 118.475 24.835 ;
        RECT 113.650 10.440 118.475 11.800 ;
        RECT 121.905 11.800 123.265 24.835 ;
        RECT 137.225 26.230 138.585 38.250 ;
        RECT 137.225 11.800 138.585 24.835 ;
        RECT 121.905 10.440 126.730 11.800 ;
        RECT 135.310 10.440 138.585 11.800 ;
      LAYER met5 ;
        RECT 109.530 122.440 111.130 140.315 ;
        RECT 129.250 122.440 130.850 140.315 ;
        RECT 101.675 120.840 118.595 122.440 ;
        RECT 101.675 116.715 103.275 120.840 ;
        RECT 104.875 116.715 115.395 119.240 ;
        RECT 116.995 116.715 118.595 120.840 ;
        RECT 101.675 115.115 118.595 116.715 ;
        RECT 101.675 110.890 103.275 115.115 ;
        RECT 104.875 110.890 115.395 115.115 ;
        RECT 116.995 110.890 118.595 115.115 ;
        RECT 101.675 109.290 118.595 110.890 ;
        RECT 101.675 104.660 103.275 109.290 ;
        RECT 104.875 108.720 115.395 109.290 ;
        RECT 104.875 108.710 106.595 108.720 ;
        RECT 104.995 105.650 106.595 108.710 ;
        RECT 104.875 105.640 106.595 105.650 ;
        RECT 109.335 105.640 110.935 108.720 ;
        RECT 113.675 108.710 115.395 108.720 ;
        RECT 113.675 105.650 115.275 108.710 ;
        RECT 113.675 105.640 115.395 105.650 ;
        RECT 104.875 104.660 115.395 105.640 ;
        RECT 116.995 104.660 118.595 109.290 ;
        RECT 101.675 103.045 118.595 104.660 ;
        RECT 101.675 97.925 103.275 103.045 ;
        RECT 104.875 97.925 115.395 103.045 ;
        RECT 116.995 97.925 118.595 103.045 ;
        RECT 101.675 96.310 118.595 97.925 ;
        RECT 101.675 91.060 103.275 96.310 ;
        RECT 104.875 95.120 115.395 96.310 ;
        RECT 104.875 95.110 106.595 95.120 ;
        RECT 104.995 92.050 106.595 95.110 ;
        RECT 104.875 92.040 106.595 92.050 ;
        RECT 109.335 92.040 110.935 95.120 ;
        RECT 113.675 95.110 115.395 95.120 ;
        RECT 113.675 92.050 115.275 95.110 ;
        RECT 113.675 92.040 115.395 92.050 ;
        RECT 104.875 91.060 115.395 92.040 ;
        RECT 116.995 91.060 118.595 96.310 ;
        RECT 101.675 89.445 118.595 91.060 ;
        RECT 101.675 84.325 103.275 89.445 ;
        RECT 104.875 84.325 115.395 89.445 ;
        RECT 116.995 84.325 118.595 89.445 ;
        RECT 101.675 82.710 118.595 84.325 ;
        RECT 101.675 77.460 103.275 82.710 ;
        RECT 104.875 81.520 115.395 82.710 ;
        RECT 104.875 81.510 106.595 81.520 ;
        RECT 104.995 78.450 106.595 81.510 ;
        RECT 104.875 78.440 106.595 78.450 ;
        RECT 109.335 78.440 110.935 81.520 ;
        RECT 113.675 81.510 115.395 81.520 ;
        RECT 113.675 78.450 115.275 81.510 ;
        RECT 113.675 78.440 115.395 78.450 ;
        RECT 104.875 77.460 115.395 78.440 ;
        RECT 116.995 77.460 118.595 82.710 ;
        RECT 101.675 75.845 118.595 77.460 ;
        RECT 101.675 70.725 103.275 75.845 ;
        RECT 104.875 70.725 115.395 75.845 ;
        RECT 116.995 70.725 118.595 75.845 ;
        RECT 101.675 69.110 118.595 70.725 ;
        RECT 101.675 63.860 103.275 69.110 ;
        RECT 104.875 67.920 115.395 69.110 ;
        RECT 104.875 67.910 106.595 67.920 ;
        RECT 104.995 64.850 106.595 67.910 ;
        RECT 104.875 64.840 106.595 64.850 ;
        RECT 109.335 64.840 110.935 67.920 ;
        RECT 113.675 67.910 115.395 67.920 ;
        RECT 113.675 64.850 115.275 67.910 ;
        RECT 113.675 64.840 115.395 64.850 ;
        RECT 104.875 63.860 115.395 64.840 ;
        RECT 116.995 63.860 118.595 69.110 ;
        RECT 101.675 62.245 118.595 63.860 ;
        RECT 101.675 57.125 103.275 62.245 ;
        RECT 104.875 57.125 115.395 62.245 ;
        RECT 116.995 57.125 118.595 62.245 ;
        RECT 101.675 55.510 118.595 57.125 ;
        RECT 101.675 50.260 103.275 55.510 ;
        RECT 104.875 54.320 115.395 55.510 ;
        RECT 104.875 54.310 106.595 54.320 ;
        RECT 104.995 51.250 106.595 54.310 ;
        RECT 104.875 51.240 106.595 51.250 ;
        RECT 109.335 51.240 110.935 54.320 ;
        RECT 113.675 54.310 115.395 54.320 ;
        RECT 113.675 51.250 115.275 54.310 ;
        RECT 113.675 51.240 115.395 51.250 ;
        RECT 104.875 50.260 115.395 51.240 ;
        RECT 116.995 50.260 118.595 55.510 ;
        RECT 101.675 48.645 118.595 50.260 ;
        RECT 101.675 43.525 103.275 48.645 ;
        RECT 104.875 43.525 115.395 48.645 ;
        RECT 116.995 43.525 118.595 48.645 ;
        RECT 101.675 41.910 118.595 43.525 ;
        RECT 101.675 36.660 103.275 41.910 ;
        RECT 104.875 40.720 115.395 41.910 ;
        RECT 104.875 40.710 106.595 40.720 ;
        RECT 104.995 37.650 106.595 40.710 ;
        RECT 104.875 37.640 106.595 37.650 ;
        RECT 109.335 37.640 110.935 40.720 ;
        RECT 113.675 40.710 115.395 40.720 ;
        RECT 113.675 37.650 115.275 40.710 ;
        RECT 113.675 37.640 115.395 37.650 ;
        RECT 104.875 36.660 115.395 37.640 ;
        RECT 116.995 36.660 118.595 41.910 ;
        RECT 101.675 35.045 118.595 36.660 ;
        RECT 101.675 29.925 103.275 35.045 ;
        RECT 104.875 29.925 115.395 35.045 ;
        RECT 116.995 29.925 118.595 35.045 ;
        RECT 101.675 28.310 118.595 29.925 ;
        RECT 101.675 23.470 103.275 28.310 ;
        RECT 104.875 27.120 115.395 28.310 ;
        RECT 104.875 27.110 106.595 27.120 ;
        RECT 104.995 24.050 106.595 27.110 ;
        RECT 104.875 24.040 106.595 24.050 ;
        RECT 109.335 24.040 110.935 27.120 ;
        RECT 113.675 27.110 115.395 27.120 ;
        RECT 113.675 24.050 115.275 27.110 ;
        RECT 113.675 24.040 115.395 24.050 ;
        RECT 104.875 23.470 115.395 24.040 ;
        RECT 116.995 23.470 118.595 28.310 ;
        RECT 101.675 21.870 118.595 23.470 ;
        RECT 101.675 17.645 103.275 21.870 ;
        RECT 104.875 17.645 115.395 21.870 ;
        RECT 116.995 17.645 118.595 21.870 ;
        RECT 101.675 16.045 118.595 17.645 ;
        RECT 101.675 11.920 103.275 16.045 ;
        RECT 104.875 13.520 115.395 16.045 ;
        RECT 116.995 11.920 118.595 16.045 ;
        RECT 101.675 10.320 118.595 11.920 ;
        RECT 121.785 120.840 138.705 122.440 ;
        RECT 121.785 116.715 123.385 120.840 ;
        RECT 124.985 116.715 135.505 119.240 ;
        RECT 137.105 116.715 138.705 120.840 ;
        RECT 121.785 115.115 138.705 116.715 ;
        RECT 121.785 110.890 123.385 115.115 ;
        RECT 124.985 110.890 135.505 115.115 ;
        RECT 137.105 110.890 138.705 115.115 ;
        RECT 121.785 109.290 138.705 110.890 ;
        RECT 121.785 104.660 123.385 109.290 ;
        RECT 124.985 108.720 135.505 109.290 ;
        RECT 124.985 108.710 126.705 108.720 ;
        RECT 125.105 105.650 126.705 108.710 ;
        RECT 124.985 105.640 126.705 105.650 ;
        RECT 129.445 105.640 131.045 108.720 ;
        RECT 133.785 108.710 135.505 108.720 ;
        RECT 133.785 105.650 135.385 108.710 ;
        RECT 133.785 105.640 135.505 105.650 ;
        RECT 124.985 104.660 135.505 105.640 ;
        RECT 137.105 104.660 138.705 109.290 ;
        RECT 121.785 103.045 138.705 104.660 ;
        RECT 121.785 97.925 123.385 103.045 ;
        RECT 124.985 97.925 135.505 103.045 ;
        RECT 137.105 97.925 138.705 103.045 ;
        RECT 121.785 96.310 138.705 97.925 ;
        RECT 121.785 91.060 123.385 96.310 ;
        RECT 124.985 95.120 135.505 96.310 ;
        RECT 124.985 95.110 126.705 95.120 ;
        RECT 125.105 92.050 126.705 95.110 ;
        RECT 124.985 92.040 126.705 92.050 ;
        RECT 129.445 92.040 131.045 95.120 ;
        RECT 133.785 95.110 135.505 95.120 ;
        RECT 133.785 92.050 135.385 95.110 ;
        RECT 133.785 92.040 135.505 92.050 ;
        RECT 124.985 91.060 135.505 92.040 ;
        RECT 137.105 91.060 138.705 96.310 ;
        RECT 121.785 89.445 138.705 91.060 ;
        RECT 121.785 84.325 123.385 89.445 ;
        RECT 124.985 84.325 135.505 89.445 ;
        RECT 137.105 84.325 138.705 89.445 ;
        RECT 121.785 82.710 138.705 84.325 ;
        RECT 121.785 77.460 123.385 82.710 ;
        RECT 124.985 81.520 135.505 82.710 ;
        RECT 124.985 81.510 126.705 81.520 ;
        RECT 125.105 78.450 126.705 81.510 ;
        RECT 124.985 78.440 126.705 78.450 ;
        RECT 129.445 78.440 131.045 81.520 ;
        RECT 133.785 81.510 135.505 81.520 ;
        RECT 133.785 78.450 135.385 81.510 ;
        RECT 133.785 78.440 135.505 78.450 ;
        RECT 124.985 77.460 135.505 78.440 ;
        RECT 137.105 77.460 138.705 82.710 ;
        RECT 121.785 75.845 138.705 77.460 ;
        RECT 121.785 70.725 123.385 75.845 ;
        RECT 124.985 70.725 135.505 75.845 ;
        RECT 137.105 70.725 138.705 75.845 ;
        RECT 121.785 69.110 138.705 70.725 ;
        RECT 121.785 63.860 123.385 69.110 ;
        RECT 124.985 67.920 135.505 69.110 ;
        RECT 124.985 67.910 126.705 67.920 ;
        RECT 125.105 64.850 126.705 67.910 ;
        RECT 124.985 64.840 126.705 64.850 ;
        RECT 129.445 64.840 131.045 67.920 ;
        RECT 133.785 67.910 135.505 67.920 ;
        RECT 133.785 64.850 135.385 67.910 ;
        RECT 133.785 64.840 135.505 64.850 ;
        RECT 124.985 63.860 135.505 64.840 ;
        RECT 137.105 63.860 138.705 69.110 ;
        RECT 121.785 62.245 138.705 63.860 ;
        RECT 121.785 57.125 123.385 62.245 ;
        RECT 124.985 57.125 135.505 62.245 ;
        RECT 137.105 57.125 138.705 62.245 ;
        RECT 121.785 55.510 138.705 57.125 ;
        RECT 121.785 50.260 123.385 55.510 ;
        RECT 124.985 54.320 135.505 55.510 ;
        RECT 124.985 54.310 126.705 54.320 ;
        RECT 125.105 51.250 126.705 54.310 ;
        RECT 124.985 51.240 126.705 51.250 ;
        RECT 129.445 51.240 131.045 54.320 ;
        RECT 133.785 54.310 135.505 54.320 ;
        RECT 133.785 51.250 135.385 54.310 ;
        RECT 133.785 51.240 135.505 51.250 ;
        RECT 124.985 50.260 135.505 51.240 ;
        RECT 137.105 50.260 138.705 55.510 ;
        RECT 121.785 48.645 138.705 50.260 ;
        RECT 121.785 43.525 123.385 48.645 ;
        RECT 124.985 43.525 135.505 48.645 ;
        RECT 137.105 43.525 138.705 48.645 ;
        RECT 121.785 41.910 138.705 43.525 ;
        RECT 121.785 36.660 123.385 41.910 ;
        RECT 124.985 40.720 135.505 41.910 ;
        RECT 124.985 40.710 126.705 40.720 ;
        RECT 125.105 37.650 126.705 40.710 ;
        RECT 124.985 37.640 126.705 37.650 ;
        RECT 129.445 37.640 131.045 40.720 ;
        RECT 133.785 40.710 135.505 40.720 ;
        RECT 133.785 37.650 135.385 40.710 ;
        RECT 133.785 37.640 135.505 37.650 ;
        RECT 124.985 36.660 135.505 37.640 ;
        RECT 137.105 36.660 138.705 41.910 ;
        RECT 121.785 35.045 138.705 36.660 ;
        RECT 121.785 29.925 123.385 35.045 ;
        RECT 124.985 29.925 135.505 35.045 ;
        RECT 137.105 29.925 138.705 35.045 ;
        RECT 121.785 28.310 138.705 29.925 ;
        RECT 121.785 23.470 123.385 28.310 ;
        RECT 124.985 27.120 135.505 28.310 ;
        RECT 124.985 27.110 126.705 27.120 ;
        RECT 125.105 24.050 126.705 27.110 ;
        RECT 124.985 24.040 126.705 24.050 ;
        RECT 129.445 24.040 131.045 27.120 ;
        RECT 133.785 27.110 135.505 27.120 ;
        RECT 133.785 24.050 135.385 27.110 ;
        RECT 133.785 24.040 135.505 24.050 ;
        RECT 124.985 23.470 135.505 24.040 ;
        RECT 137.105 23.470 138.705 28.310 ;
        RECT 121.785 21.870 138.705 23.470 ;
        RECT 121.785 17.645 123.385 21.870 ;
        RECT 124.985 17.645 135.505 21.870 ;
        RECT 137.105 17.645 138.705 21.870 ;
        RECT 121.785 16.045 138.705 17.645 ;
        RECT 121.785 11.920 123.385 16.045 ;
        RECT 124.985 13.520 135.505 16.045 ;
        RECT 137.105 11.920 138.705 16.045 ;
        RECT 121.785 10.320 138.705 11.920 ;
      LAYER met5 ;
        RECT -0.130 -1.640 253.790 -1.600 ;
  END
END /local_disk/fossi_cochlea/mag/final_designs/filter_p_m
END LIBRARY

