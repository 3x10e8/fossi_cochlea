magic
tech sky130A
timestamp 1654307754
<< metal3 >>
rect -14 -14 684 614
<< mimcap >>
rect 0 549 670 600
rect 0 517 17 549
rect 49 517 117 549
rect 149 517 217 549
rect 249 517 317 549
rect 349 517 417 549
rect 449 517 517 549
rect 549 517 617 549
rect 649 517 670 549
rect 0 449 670 517
rect 0 417 17 449
rect 49 417 617 449
rect 649 417 670 449
rect 0 349 670 417
rect 0 317 17 349
rect 49 317 617 349
rect 649 317 670 349
rect 0 249 670 317
rect 0 217 17 249
rect 49 217 617 249
rect 649 217 670 249
rect 0 149 670 217
rect 0 117 17 149
rect 49 117 617 149
rect 649 117 670 149
rect 0 49 670 117
rect 0 17 17 49
rect 49 17 117 49
rect 149 17 217 49
rect 249 17 317 49
rect 349 17 417 49
rect 449 17 517 49
rect 549 17 617 49
rect 649 17 670 49
rect 0 0 670 17
<< mimcapcontact >>
rect 17 517 49 549
rect 117 517 149 549
rect 217 517 249 549
rect 317 517 349 549
rect 417 517 449 549
rect 517 517 549 549
rect 617 517 649 549
rect 17 417 49 449
rect 617 417 649 449
rect 17 317 49 349
rect 617 317 649 349
rect 17 217 49 249
rect 617 217 649 249
rect 17 117 49 149
rect 617 117 649 149
rect 17 17 49 49
rect 117 17 149 49
rect 217 17 249 49
rect 317 17 349 49
rect 417 17 449 49
rect 517 17 549 49
rect 617 17 649 49
<< metal4 >>
rect 7 549 59 559
rect 7 517 17 549
rect 49 517 59 549
rect 7 507 59 517
rect 107 549 159 559
rect 107 517 117 549
rect 149 517 159 549
rect 107 507 159 517
rect 207 549 259 559
rect 207 517 217 549
rect 249 517 259 549
rect 207 507 259 517
rect 307 549 359 559
rect 307 517 317 549
rect 349 517 359 549
rect 307 507 359 517
rect 407 549 459 559
rect 407 517 417 549
rect 449 517 459 549
rect 407 507 459 517
rect 507 549 559 559
rect 507 517 517 549
rect 549 517 559 549
rect 507 507 559 517
rect 607 549 659 559
rect 607 517 617 549
rect 649 517 659 549
rect 607 507 659 517
rect 7 449 59 459
rect 7 417 17 449
rect 49 417 59 449
rect 7 407 59 417
rect 607 449 659 459
rect 607 417 617 449
rect 649 417 659 449
rect 607 407 659 417
rect 7 349 59 359
rect 7 317 17 349
rect 49 317 59 349
rect 7 307 59 317
rect 607 349 659 359
rect 607 317 617 349
rect 649 317 659 349
rect 607 307 659 317
rect 7 249 59 259
rect 7 217 17 249
rect 49 217 59 249
rect 7 207 59 217
rect 607 249 659 259
rect 607 217 617 249
rect 649 217 659 249
rect 607 207 659 217
rect 7 149 59 159
rect 7 117 17 149
rect 49 117 59 149
rect 7 107 59 117
rect 607 149 659 159
rect 607 117 617 149
rect 649 117 659 149
rect 607 107 659 117
rect 7 49 59 59
rect 7 17 17 49
rect 49 17 59 49
rect 7 7 59 17
rect 107 49 159 59
rect 107 17 117 49
rect 149 17 159 49
rect 107 7 159 17
rect 207 49 259 59
rect 207 17 217 49
rect 249 17 259 49
rect 207 7 259 17
rect 307 49 359 59
rect 307 17 317 49
rect 349 17 359 49
rect 307 7 359 17
rect 407 49 459 59
rect 407 17 417 49
rect 449 17 459 49
rect 407 7 459 17
rect 507 49 559 59
rect 507 17 517 49
rect 549 17 559 49
rect 507 7 559 17
rect 607 49 659 59
rect 607 17 617 49
rect 649 17 659 49
rect 607 7 659 17
<< end >>
