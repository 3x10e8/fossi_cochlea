magic
tech sky130B
magscale 1 2
timestamp 1654741520
<< nwell >>
rect -94 162 185 330
<< nmos >>
rect 0 10 30 94
<< pmos >>
rect 0 199 30 283
<< ndiff >>
rect -58 70 0 94
rect -58 36 -50 70
rect -16 36 0 70
rect -58 10 0 36
rect 30 70 92 94
rect 30 36 46 70
rect 80 36 92 70
rect 30 10 92 36
<< pdiff >>
rect -58 257 0 283
rect -58 223 -50 257
rect -16 223 0 257
rect -58 199 0 223
rect 30 257 91 283
rect 30 223 46 257
rect 80 223 91 257
rect 30 199 91 223
<< ndiffc >>
rect -50 36 -16 70
rect 46 36 80 70
<< pdiffc >>
rect -50 223 -16 257
rect 46 223 80 257
<< psubdiff >>
rect 92 70 150 94
rect 92 36 116 70
rect 92 10 150 36
<< nsubdiff >>
rect 91 257 149 283
rect 91 223 114 257
rect 148 223 149 257
rect 91 199 149 223
<< psubdiffcont >>
rect 116 36 150 70
<< nsubdiffcont >>
rect 114 223 148 257
<< poly >>
rect -2 375 32 381
rect -12 365 42 375
rect -12 331 -2 365
rect 32 331 42 365
rect -12 319 42 331
rect -2 315 32 319
rect 0 283 30 315
rect 0 173 30 199
rect 0 94 30 120
rect 0 -12 30 10
rect -2 -16 32 -12
rect -12 -28 42 -16
rect -12 -62 -2 -28
rect 32 -62 42 -28
rect -12 -72 42 -62
rect -2 -78 32 -72
<< polycont >>
rect -2 331 32 365
rect -2 -62 32 -28
<< locali >>
rect -2 365 32 381
rect -2 315 32 330
rect 114 344 176 378
rect -144 257 -16 273
rect -144 244 -50 257
rect -144 57 -94 244
rect -60 223 -50 244
rect -60 70 -16 223
rect -60 57 -50 70
rect -144 36 -50 57
rect -144 20 -16 36
rect 46 257 80 273
rect 46 170 80 223
rect 114 257 148 344
rect 114 207 148 223
rect 46 136 90 170
rect 228 136 234 170
rect 46 70 80 136
rect 46 20 80 36
rect 116 70 150 86
rect -2 -28 32 -12
rect -2 -78 32 -62
rect 116 -45 150 36
<< viali >>
rect -2 331 32 364
rect -2 330 32 331
rect 176 344 210 378
rect -94 57 -60 244
rect 90 136 228 170
rect -2 -62 32 -28
rect 116 -79 150 -45
<< metal1 >>
rect 167 3564 219 3570
rect 167 3506 219 3512
rect 167 388 219 394
rect -11 378 41 379
rect -16 373 46 378
rect -16 321 -11 373
rect 41 321 46 373
rect 167 330 219 336
rect -16 314 46 321
rect -109 254 -45 260
rect -109 48 -103 254
rect -51 48 -45 254
rect 75 179 234 184
rect 75 127 81 179
rect 228 127 234 179
rect 75 122 234 127
rect -109 42 -45 48
rect -16 -18 46 -12
rect -16 -70 -11 -18
rect 41 -70 46 -18
rect -16 -76 46 -70
rect 100 -37 164 -33
rect 100 -89 106 -37
rect 158 -89 164 -37
rect 100 -91 164 -89
<< via1 >>
rect 167 3512 219 3564
rect 167 378 219 388
rect -11 364 41 373
rect -11 330 -2 364
rect -2 330 32 364
rect 32 330 41 364
rect -11 321 41 330
rect 167 344 176 378
rect 176 344 210 378
rect 210 344 219 378
rect 167 336 219 344
rect -103 244 -51 254
rect -103 57 -94 244
rect -94 57 -60 244
rect -60 57 -51 244
rect -103 48 -51 57
rect 81 170 228 179
rect 81 136 90 170
rect 90 136 228 170
rect 81 127 228 136
rect -11 -28 41 -18
rect -11 -62 -2 -28
rect -2 -62 32 -28
rect 32 -62 41 -28
rect -11 -70 41 -62
rect 106 -45 158 -37
rect 106 -79 116 -45
rect 116 -79 150 -45
rect 150 -79 158 -45
rect 106 -89 158 -79
<< metal2 >>
rect 167 3564 219 3570
rect 167 3506 219 3512
rect 176 394 210 3506
rect 0 379 30 393
rect -11 373 41 379
rect -11 315 41 321
rect 0 314 30 315
rect -105 254 -49 260
rect -105 249 -103 254
rect -51 249 -49 254
rect 79 252 109 393
rect 167 388 219 394
rect 167 330 219 336
rect -105 37 -49 46
rect 0 222 109 252
rect 0 -12 30 222
rect 79 181 234 190
rect 228 125 234 181
rect 79 116 234 125
rect -11 -18 41 -12
rect -11 -76 41 -70
rect 106 -37 158 -31
rect 106 -95 158 -89
<< via2 >>
rect -105 48 -103 249
rect -103 48 -51 249
rect -51 48 -49 249
rect -105 46 -49 48
rect 79 179 228 181
rect 79 127 81 179
rect 81 127 228 179
rect 79 125 228 127
<< metal3 >>
rect -117 262 -38 265
rect -117 203 -109 262
rect -140 103 -109 203
rect -117 42 -109 103
rect -45 42 -38 262
rect 70 185 234 202
rect 70 121 75 185
rect 70 102 234 121
rect -117 35 -38 42
<< via3 >>
rect -109 249 -45 262
rect -109 46 -105 249
rect -105 46 -49 249
rect -49 46 -45 249
rect -109 42 -45 46
rect 75 181 234 185
rect 75 125 79 181
rect 79 125 228 181
rect 228 125 234 181
rect 75 121 234 125
<< metal4 >>
rect -110 262 -41 263
rect -110 189 -109 262
rect -175 117 -109 189
rect -110 42 -109 117
rect -45 42 -41 262
rect 71 185 235 189
rect 71 121 75 185
rect 234 121 235 185
rect 71 117 235 121
rect -110 38 -41 42
<< labels >>
flabel via1 -2 330 32 364 0 FreeSans 80 0 0 0 phib
flabel viali -94 136 -60 170 0 FreeSans 80 0 0 0 in
flabel via1 -2 -62 32 -28 0 FreeSans 80 0 0 0 phi
flabel viali 90 136 124 170 0 FreeSans 80 0 0 0 out
flabel viali -94 57 -60 91 0 FreeSans 80 0 0 0 in
<< end >>
