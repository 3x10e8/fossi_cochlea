`timescale 1ns/10ps
`include "edge_ff_n.v"
`include "tbuf.v"
`include "u_d_bin_counter.v"
//To be included with testbenches
`include "gray_count.v"
`include "./../cclk/cclk_gen.v"


module dlrtn(//this is negative reset and active low enable latch.
	input d,
	input gate,
	input rstb,
	output reg q);
	always@(rstb,d,gate)begin
		if(!rstb) q<=0;
		else if(!gate) q<=d;
	end
endmodule

module gray_selector_fb( //clk_ext is the core's clock
input d,clk_ext,rstb_ext, //d has to be connected to vdd in our case
input [9:0]in,clk, //ext gray clocks are to be connected to the clk
output wire out_muxed); //rstb pin of eff has to be ext clk signal
wire [9:0]eff_out,eff_outb; //rstb_ext to be connected to rstb(global)
wire out_muxed_raw;
assign eff_outb[9:0]=~eff_out[9:0];
genvar i;
generate for(i=0;i<=9;i=i+1) begin: fb_gray_selector_loop
edge_ff_n eff(.d(d),.rstb(clk_ext),.clk(clk[i]),.out(eff_out[i]));
tbuf t_buf(.in(in[i]),.ctrlb(eff_outb[i]),.out(out_muxed_raw));
dlrtn dl(.d(out_muxed_raw),.gate(clk_ext),.rstb(rstb_ext),.q(out_muxed));
end
endgenerate
endmodule

module fb(
	input vpwr,clkdiv2,comp_out,cclk,rstb,ud_en, //clkdiv2 is the max clk frequency of the core
	input [9:0]gray_clk, //ud_en is the en port of the ud counter. extra control to the feedback.
	output wire fb_out);
	wire [15:0]c_count; //c_count is the bin counter's output

	u_d_bin_counter ud_c(.u_d(comp_out),.clk(cclk),.rstb(rstb),.en(ud_en),.q(c_count[15:0]));
	gray_selector_fb gs_f(.d(vpwr),.clk_ext(clkdiv2),.rstb_ext(rstb),.in({c_count[6],c_count[7],c_count[8],c_count[9],c_count[10],c_count[11],c_count[12],c_count[13],c_count[14],c_count[15]}),.clk(gray_clk[9:0]),.out_muxed(fb_out));

endmodule

/*
//Testbench parameterized for all the cores
//gc: Gray Counter
//gs: Gray Selector
//c: Counter
//clk_ext: external clock of the core
module tb_fb;
	reg vpwr,clkdiv2,comp_out,rstb,ud_en;
	wire fb_out,cclk;
	reg clk_master; //clk_master is the master clk of the whole chip 
	wire [18:0]gc_clk;
	parameter PERIOD_MASTER=400;
	real clk_master_half_pd=PERIOD_MASTER/2;
	parameter n=1;
	parameter PERIOD_CORE=400*(2**(n-1));
	real clk_core_half_pd=(PERIOD_CORE)/2;
	real comp_out_half_pd=PERIOD_CORE;//factor of 2 is multiplied here because the period of comput is double that of the core clock
	//module instantiation	
	gray_count gc_clock(
		.clk(clk_master), 
		.reset(rstb), 
		.gray_count(gc_clk[18:0]));

	fb fb_block(
		.vpwr(vpwr),
		.clkdiv2(clkdiv2),
		.comp_out(comp_out),
		.cclk(cclk),
		.rstb(rstb),
		.ud_en(ud_en),
		.gray_clk(gc_clk[n+9:n]),
		.fb_out(fb_out));// gray_clk is indexed from 10:1 here because 																		//	the feedback requires gray bit frequency
																		// to be 1/4 times that of the max freqency.
	cclk_gen cc(
		.clk(clkdiv2),
		.rstb(rstb),
		.cclk(cclk)); //cclk is used to model the cclk generated by the analog clcok generator.
	initial begin
	$dumpfile("fb.vcd");
	$dumpvars;
	end 	
	//signal generation
	initial begin
		clk_master=0;
		forever
			#(clk_master_half_pd)clk_master = ~clk_master; //ext_clk generation freq=2.56 MHz
	end

	initial begin
		clkdiv2=0;
		//#(clk_master_half_pd) clkdiv2=1;
		forever
			#(clk_core_half_pd)clkdiv2 = ~clkdiv2; //ext_clk generation freq=2.56 MHz
	end

		
	always @(posedge rstb or negedge rstb or negedge clkdiv2) begin
		//comp_out=0;
			if(rstb&~clkdiv2) begin
				#2 comp_out<=1;
				#(comp_out_half_pd) comp_out=~comp_out;
				end
			else comp_out<=comp_out;
	end 

	initial begin
		//comp_out=1;
		rstb=0;
		ud_en=1;
		vpwr=1;
		#5 rstb=1;
		#6476802 ud_en=0;
		repeat(2048) @(posedge clkdiv2);
		#2 ud_en=1;
		repeat(34000) @(negedge clkdiv2);
		rstb=0;
		repeat(10) @(negedge clkdiv2);
		#5 rstb=1;
        #100;
		$finish; 
	end
endmodule
*/

	
