VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital_unison
  CLASS BLOCK ;
  FOREIGN digital_unison ;
  ORIGIN 0.000 0.000 ;
  SIZE 480.000 BY 100.000 ;
  PIN cclk_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 96.000 141.130 100.000 ;
    END
  END cclk_I[0]
  PIN cclk_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 96.000 378.490 100.000 ;
    END
  END cclk_I[1]
  PIN cclk_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END cclk_Q[0]
  PIN cclk_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END cclk_Q[1]
  PIN clk_master
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END clk_master
  PIN clkdiv2_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 96.000 101.570 100.000 ;
    END
  END clkdiv2_I[0]
  PIN clkdiv2_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 96.000 338.930 100.000 ;
    END
  END clkdiv2_I[1]
  PIN clkdiv2_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END clkdiv2_Q[0]
  PIN clkdiv2_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END clkdiv2_Q[1]
  PIN comp_high_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 96.000 220.250 100.000 ;
    END
  END comp_high_I[0]
  PIN comp_high_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 96.000 457.610 100.000 ;
    END
  END comp_high_I[1]
  PIN comp_high_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END comp_high_Q[0]
  PIN comp_high_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END comp_high_Q[1]
  PIN cos_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 96.000 22.450 100.000 ;
    END
  END cos_out[0]
  PIN cos_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 96.000 259.810 100.000 ;
    END
  END cos_out[1]
  PIN fb1_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 96.000 62.010 100.000 ;
    END
  END fb1_I[0]
  PIN fb1_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 96.000 299.370 100.000 ;
    END
  END fb1_I[1]
  PIN fb1_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END fb1_Q[0]
  PIN fb1_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END fb1_Q[1]
  PIN phi1b_dig_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 96.000 180.690 100.000 ;
    END
  END phi1b_dig_I[0]
  PIN phi1b_dig_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 96.000 418.050 100.000 ;
    END
  END phi1b_dig_I[1]
  PIN phi1b_dig_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END phi1b_dig_Q[0]
  PIN phi1b_dig_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END phi1b_dig_Q[1]
  PIN read_out_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 86.400 480.000 87.000 ;
    END
  END read_out_I[0]
  PIN read_out_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 61.920 480.000 62.520 ;
    END
  END read_out_I[1]
  PIN read_out_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 37.440 480.000 38.040 ;
    END
  END read_out_Q[0]
  PIN read_out_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 12.960 480.000 13.560 ;
    END
  END read_out_Q[1]
  PIN rstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END rstb
  PIN sin_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END sin_out[0]
  PIN sin_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END sin_out[1]
  PIN ud_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END ud_en
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 63.310 10.640 64.910 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 180.495 10.640 182.095 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.680 10.640 299.280 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.865 10.640 416.465 87.280 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 121.900 10.640 123.500 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 239.085 10.640 240.685 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 356.270 10.640 357.870 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 473.455 10.640 475.055 87.280 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 474.260 87.125 ;
      LAYER met1 ;
        RECT 5.520 10.640 476.030 87.680 ;
      LAYER met2 ;
        RECT 7.910 95.720 21.890 96.000 ;
        RECT 22.730 95.720 61.450 96.000 ;
        RECT 62.290 95.720 101.010 96.000 ;
        RECT 101.850 95.720 140.570 96.000 ;
        RECT 141.410 95.720 180.130 96.000 ;
        RECT 180.970 95.720 219.690 96.000 ;
        RECT 220.530 95.720 259.250 96.000 ;
        RECT 260.090 95.720 298.810 96.000 ;
        RECT 299.650 95.720 338.370 96.000 ;
        RECT 339.210 95.720 377.930 96.000 ;
        RECT 378.770 95.720 417.490 96.000 ;
        RECT 418.330 95.720 457.050 96.000 ;
        RECT 457.890 95.720 476.010 96.000 ;
        RECT 7.910 4.280 476.010 95.720 ;
        RECT 7.910 4.000 21.890 4.280 ;
        RECT 22.730 4.000 61.450 4.280 ;
        RECT 62.290 4.000 101.010 4.280 ;
        RECT 101.850 4.000 140.570 4.280 ;
        RECT 141.410 4.000 180.130 4.280 ;
        RECT 180.970 4.000 219.690 4.280 ;
        RECT 220.530 4.000 259.250 4.280 ;
        RECT 260.090 4.000 298.810 4.280 ;
        RECT 299.650 4.000 338.370 4.280 ;
        RECT 339.210 4.000 377.930 4.280 ;
        RECT 378.770 4.000 417.490 4.280 ;
        RECT 418.330 4.000 457.050 4.280 ;
        RECT 457.890 4.000 476.010 4.280 ;
      LAYER met3 ;
        RECT 4.000 86.000 475.600 87.205 ;
        RECT 4.000 84.000 477.170 86.000 ;
        RECT 4.400 82.600 477.170 84.000 ;
        RECT 4.000 62.920 477.170 82.600 ;
        RECT 4.000 61.520 475.600 62.920 ;
        RECT 4.000 50.680 477.170 61.520 ;
        RECT 4.400 49.280 477.170 50.680 ;
        RECT 4.000 38.440 477.170 49.280 ;
        RECT 4.000 37.040 475.600 38.440 ;
        RECT 4.000 17.360 477.170 37.040 ;
        RECT 4.400 15.960 477.170 17.360 ;
        RECT 4.000 13.960 477.170 15.960 ;
        RECT 4.000 12.560 475.600 13.960 ;
        RECT 4.000 10.715 477.170 12.560 ;
      LAYER met4 ;
        RECT 296.535 23.975 297.280 65.785 ;
        RECT 299.680 23.975 318.025 65.785 ;
  END
END digital_unison
END LIBRARY

