magic
tech sky130A
magscale 1 2
timestamp 1647892206
<< metal1 >>
rect 11566 -2518 11618 -2512
rect 11192 -2570 11566 -2546
rect 11618 -2570 11724 -2546
rect 11192 -2574 11724 -2570
rect 11566 -2576 11618 -2574
rect 11494 -2608 11546 -2604
rect 11194 -2610 11744 -2608
rect 11194 -2636 11494 -2610
rect 11546 -2636 11744 -2610
rect 11494 -2668 11546 -2662
rect 11200 -2694 11252 -2688
rect 10316 -2734 11200 -2700
rect 11252 -2734 11744 -2700
rect 11200 -2752 11252 -2746
rect 11426 -3162 11478 -3156
rect 11194 -3198 11426 -3170
rect 11426 -3220 11478 -3214
rect 11634 -3162 11686 -3156
rect 11686 -3198 11722 -3170
rect 11634 -3220 11686 -3214
rect 11285 -3436 11337 -3430
rect 11192 -3488 11285 -3468
rect 11337 -3488 11718 -3468
rect 11192 -3496 11718 -3488
rect 11366 -3530 11418 -3524
rect 11194 -3560 11366 -3532
rect 11418 -3560 11722 -3532
rect 11366 -3588 11418 -3582
rect 11208 -9719 11308 -9704
rect 11208 -9773 11214 -9719
rect 11268 -9773 11308 -9719
rect 11208 -9802 11308 -9773
<< via1 >>
rect 11566 -2570 11618 -2518
rect 11494 -2662 11546 -2610
rect 11200 -2746 11252 -2694
rect 11426 -3214 11478 -3162
rect 11634 -3214 11686 -3162
rect 11285 -3488 11337 -3436
rect 11366 -3582 11418 -3530
rect 11214 -9773 11268 -9719
rect 19471 -10439 19525 -10387
<< metal2 >>
rect 11226 -2688 11256 6398
rect 11200 -2694 11256 -2688
rect 11252 -2746 11256 -2694
rect 11200 -2752 11256 -2746
rect 11226 -9704 11256 -2752
rect 11296 -3430 11326 6398
rect 11285 -3436 11337 -3430
rect 11285 -3494 11337 -3488
rect 11295 -3496 11337 -3494
rect 11296 -3497 11337 -3496
rect 11296 -9682 11326 -3497
rect 11366 -3524 11396 6398
rect 11436 -3156 11466 6398
rect 11506 -2604 11536 6398
rect 11576 -2512 11606 6398
rect 11566 -2518 11618 -2512
rect 11566 -2576 11618 -2570
rect 11494 -2610 11546 -2604
rect 11494 -2668 11546 -2662
rect 11426 -3162 11478 -3156
rect 11426 -3220 11478 -3214
rect 11366 -3530 11418 -3524
rect 11366 -3588 11418 -3582
rect 11506 -9680 11536 -2668
rect 11646 -3156 11676 6398
rect 11634 -3162 11686 -3156
rect 11634 -3220 11686 -3214
rect 11208 -9719 11268 -9704
rect 11208 -9773 11214 -9719
rect 11208 -9802 11268 -9773
rect 19459 -10387 19536 -10378
rect 19459 -10443 19469 -10387
rect 19525 -10443 19536 -10387
rect 19459 -10453 19536 -10443
<< via2 >>
rect 19469 -10439 19471 -10387
rect 19471 -10439 19525 -10387
rect 19469 -10443 19525 -10439
<< metal3 >>
rect 11120 5512 11761 5675
rect 11139 4857 11780 5020
rect 10991 3273 11899 3546
rect 11015 2017 11923 2290
rect 10976 820 11884 1093
rect 11049 -308 11957 -35
rect 10991 -1407 11899 -1134
rect 19415 -10387 19583 -9532
rect 19415 -10443 19469 -10387
rect 19525 -10443 19583 -10387
rect 19415 -10468 19583 -10443
<< metal4 >>
rect 11126 -9630 11184 -9628
rect 11126 -10112 11186 -9630
rect 11614 -9650 11720 -9552
rect 11614 -10048 11674 -9650
rect 11596 -10088 11674 -10048
rect 11126 -10172 11357 -10112
use comparator_final  comparator_final_0
timestamp 1647892206
transform 1 0 11870 0 1 -10038
box -574 -430 9938 401
use fitler_cell  fitler_cell_0
timestamp 1647840975
transform 1 0 4 0 1 0
box -5288 -9650 11208 6206
use fitler_cell  fitler_cell_1
timestamp 1647840975
transform -1 0 22898 0 1 0
box -5288 -9650 11208 6206
<< end >>
