magic
tech sky130A
magscale 1 2
timestamp 1654685496
<< nwell >>
rect -1347 690 -720 815
rect -1093 673 -1033 690
rect 1001 671 1625 823
rect -359 -11 651 381
<< pmos >>
rect -228 203 -198 287
rect -133 145 -103 345
rect 395 145 425 345
rect 490 203 520 287
rect 87 36 117 120
rect 176 36 206 120
<< nnmos >>
rect -217 -337 -17 -237
rect 309 -337 509 -237
<< nmoslvt >>
rect -524 370 -440 770
rect 732 370 816 770
rect -524 -87 -440 313
rect 732 -87 816 313
rect 104 -927 188 -527
<< ndiff >>
rect -524 815 -440 839
rect -524 781 -516 815
rect -448 781 -440 815
rect -524 770 -440 781
rect 732 815 816 839
rect 732 781 740 815
rect 808 781 816 815
rect 732 770 816 781
rect -524 359 -440 370
rect -524 324 -516 359
rect -448 324 -440 359
rect 732 359 816 370
rect -524 313 -440 324
rect 732 324 740 359
rect 808 324 816 359
rect 732 313 816 324
rect -524 -98 -440 -87
rect -524 -132 -516 -98
rect -448 -132 -440 -98
rect -524 -144 -440 -132
rect 732 -98 816 -87
rect 732 -132 740 -98
rect 808 -132 816 -98
rect 732 -144 816 -132
rect 104 -482 188 -470
rect 104 -516 112 -482
rect 180 -516 188 -482
rect 104 -527 188 -516
rect 104 -938 188 -927
rect 104 -972 112 -938
rect 180 -972 188 -938
rect 104 -994 188 -972
<< pdiff >>
rect -183 287 -133 345
rect -283 265 -228 287
rect -283 231 -274 265
rect -240 231 -228 265
rect -283 203 -228 231
rect -198 203 -133 287
rect -183 145 -133 203
rect -103 333 -44 345
rect -103 157 -86 333
rect -52 157 -44 333
rect 336 333 395 345
rect -103 145 -44 157
rect 336 157 344 333
rect 378 157 395 333
rect 336 145 395 157
rect 425 287 475 345
rect 425 203 490 287
rect 520 265 575 287
rect 520 231 532 265
rect 566 231 575 265
rect 520 203 575 231
rect 425 145 475 203
rect 32 94 87 120
rect 32 60 40 94
rect 74 60 87 94
rect 32 36 87 60
rect 117 94 176 120
rect 117 60 129 94
rect 163 60 176 94
rect 117 36 176 60
rect 206 94 261 120
rect 206 60 218 94
rect 252 60 261 94
rect 206 36 261 60
<< mvndiff >>
rect -217 -192 -17 -180
rect -217 -226 -196 -192
rect -34 -226 -17 -192
rect -217 -237 -17 -226
rect 309 -192 509 -180
rect 309 -226 326 -192
rect 488 -226 509 -192
rect 309 -237 509 -226
rect -217 -349 -17 -337
rect -217 -383 -185 -349
rect -34 -383 -17 -349
rect -217 -394 -17 -383
rect 309 -349 509 -337
rect 309 -383 326 -349
rect 482 -383 509 -349
rect 309 -394 509 -383
<< ndiffc >>
rect -516 781 -448 815
rect 740 781 808 815
rect -516 324 -448 359
rect 740 324 808 359
rect -516 -132 -448 -98
rect 740 -132 808 -98
rect 112 -516 180 -482
rect 112 -972 180 -938
<< pdiffc >>
rect -274 231 -240 265
rect -86 157 -52 333
rect 344 157 378 333
rect 532 231 566 265
rect 40 60 74 94
rect 129 60 163 94
rect 218 60 252 94
<< mvndiffc >>
rect -196 -226 -34 -192
rect 326 -226 488 -192
rect -185 -383 -34 -349
rect 326 -383 482 -349
<< psubdiff >>
rect -524 894 -440 897
rect -524 860 -498 894
rect -464 860 -440 894
rect -524 839 -440 860
rect 732 894 816 897
rect 732 860 758 894
rect 792 860 816 894
rect 732 839 816 860
rect -1086 78 -984 96
rect -1086 43 -1062 78
rect -1015 43 -984 78
rect -1086 28 -984 43
rect 1244 83 1386 96
rect 1244 27 1270 83
rect 1354 27 1386 83
rect 1244 11 1386 27
rect 104 -1017 188 -994
rect 104 -1051 130 -1017
rect 164 -1051 188 -1017
rect 104 -1057 188 -1051
<< nsubdiff >>
rect -1170 762 -948 779
rect -1170 722 -1093 762
rect -1034 722 -948 762
rect -1170 704 -948 722
rect 1209 755 1401 781
rect 1209 708 1263 755
rect 1353 708 1401 755
rect 1209 695 1401 708
rect 105 268 187 292
rect 105 234 129 268
rect 163 234 187 268
rect 105 210 187 234
<< psubdiffcont >>
rect -498 860 -464 894
rect 758 860 792 894
rect -1062 43 -1015 78
rect 1270 27 1354 83
rect 130 -1051 164 -1017
<< nsubdiffcont >>
rect -1093 722 -1034 762
rect 1263 708 1353 755
rect 129 234 163 268
<< poly >>
rect -550 578 -524 770
rect -606 568 -524 578
rect -618 473 -596 568
rect -562 473 -524 568
rect -606 463 -524 473
rect -550 370 -524 463
rect -440 370 -414 770
rect -133 345 -103 371
rect 395 345 425 371
rect 706 370 732 770
rect 816 578 842 770
rect 816 568 898 578
rect 816 473 854 568
rect 888 473 910 568
rect 816 463 898 473
rect 816 370 842 463
rect -550 -87 -524 313
rect -440 220 -414 313
rect -228 287 -198 313
rect -440 210 -358 220
rect -440 115 -402 210
rect -368 171 -346 210
rect -228 171 -198 203
rect -368 141 -198 171
rect -368 115 -346 141
rect -440 105 -358 115
rect -133 114 -103 145
rect 87 120 117 146
rect 176 120 206 146
rect 490 287 520 313
rect 706 220 732 313
rect 650 210 732 220
rect 490 171 520 203
rect 638 171 660 210
rect -135 108 -101 114
rect -440 -87 -414 105
rect -145 98 -91 108
rect -145 64 -135 98
rect -101 64 -91 98
rect -145 54 -91 64
rect -135 48 -101 54
rect 395 114 425 145
rect 490 141 660 171
rect 638 115 660 141
rect 694 115 732 210
rect 393 108 427 114
rect 383 98 437 108
rect 650 105 732 115
rect 383 64 393 98
rect 427 64 437 98
rect 383 54 437 64
rect 393 48 427 54
rect 87 21 117 36
rect 176 21 206 36
rect 87 -9 206 21
rect 112 -11 179 -9
rect 112 -45 128 -11
rect 163 -45 179 -11
rect 118 -55 173 -45
rect 128 -58 163 -55
rect 706 -87 732 105
rect 816 -87 842 313
rect -478 -249 -217 -237
rect -478 -327 -462 -249
rect -262 -327 -217 -249
rect -478 -337 -217 -327
rect -17 -337 12 -237
rect 280 -337 309 -237
rect 509 -247 770 -237
rect 509 -325 554 -247
rect 754 -325 770 -247
rect 509 -337 770 -325
rect 78 -719 104 -527
rect 22 -729 104 -719
rect 10 -824 32 -729
rect 66 -824 104 -729
rect 22 -834 104 -824
rect 78 -927 104 -834
rect 188 -719 214 -527
rect 188 -729 270 -719
rect 188 -824 226 -729
rect 260 -824 282 -729
rect 188 -834 270 -824
rect 188 -927 214 -834
<< polycont >>
rect -596 473 -562 568
rect 854 473 888 568
rect -402 115 -368 210
rect -135 64 -101 98
rect 660 115 694 210
rect 393 64 427 98
rect 128 -45 163 -11
rect -462 -327 -262 -249
rect 554 -325 754 -247
rect 32 -824 66 -729
rect 226 -824 260 -729
<< locali >>
rect -514 860 -498 894
rect -464 860 -448 894
rect 742 860 758 894
rect 792 860 808 894
rect -498 823 -464 860
rect 758 823 792 860
rect -532 815 -432 823
rect -532 781 -516 815
rect -448 781 -432 815
rect -1093 762 -1034 778
rect -532 770 -432 781
rect 724 815 824 823
rect 724 781 740 815
rect 808 781 824 815
rect 724 770 824 781
rect -1034 722 -1033 762
rect -1093 673 -1033 722
rect 1263 755 1353 772
rect 1263 672 1353 708
rect -596 568 -562 584
rect -596 457 -562 473
rect -1062 312 -1016 378
rect -532 367 -432 370
rect -532 366 -45 367
rect -779 359 -45 366
rect -779 332 -516 359
rect -532 324 -516 332
rect -448 333 -45 359
rect -448 324 -432 333
rect -532 313 -432 324
rect -277 265 -232 283
rect -277 231 -274 265
rect -240 231 -232 265
rect -402 210 -368 226
rect -1062 78 -1015 106
rect -759 96 -670 130
rect -277 207 -232 231
rect -99 147 -86 333
rect -92 145 -86 147
rect -52 147 -45 333
rect 129 279 163 627
rect 854 568 888 584
rect 854 457 888 473
rect 724 367 824 370
rect 337 362 1058 367
rect 337 328 343 362
rect 378 359 1058 362
rect 378 333 740 359
rect 118 268 174 279
rect 118 234 129 268
rect 163 234 174 268
rect 118 223 174 234
rect -52 145 -46 147
rect -86 141 -52 143
rect -402 99 -368 115
rect 40 98 74 110
rect -1062 27 -1015 43
rect -704 -87 -670 96
rect -151 64 -135 98
rect -101 94 74 98
rect -101 64 40 94
rect -704 -96 -432 -87
rect -670 -98 -432 -96
rect -670 -130 -516 -98
rect -704 -132 -516 -130
rect -448 -132 -432 -98
rect -704 -140 -432 -132
rect -135 -181 -101 64
rect 40 44 74 60
rect 129 94 163 223
rect 337 157 344 328
rect 378 157 391 333
rect 724 324 740 333
rect 808 332 1058 359
rect 808 324 824 332
rect 724 313 824 324
rect 1289 312 1362 378
rect 524 265 569 283
rect 524 231 532 265
rect 566 231 569 265
rect 524 207 569 231
rect 660 210 694 226
rect 337 147 391 157
rect 344 141 378 147
rect 129 44 163 60
rect 218 98 252 110
rect 660 99 694 115
rect 218 94 393 98
rect 252 64 393 94
rect 427 64 443 98
rect 962 96 1037 130
rect 218 44 252 60
rect 112 -45 128 -11
rect 163 -45 179 -11
rect 112 -47 179 -45
rect 393 -181 427 64
rect 962 -87 996 96
rect 1270 83 1354 102
rect 1270 11 1354 27
rect 724 -97 996 -87
rect 724 -98 962 -97
rect 724 -132 740 -98
rect 808 -131 962 -98
rect 808 -132 996 -131
rect 724 -140 996 -132
rect -212 -192 -18 -181
rect -212 -226 -196 -192
rect -34 -226 -18 -192
rect -212 -235 -18 -226
rect 310 -192 504 -181
rect 310 -226 326 -192
rect 488 -226 504 -192
rect 310 -235 504 -226
rect -478 -249 -246 -237
rect -478 -327 -462 -249
rect -262 -327 -246 -249
rect -478 -337 -246 -327
rect 538 -247 770 -237
rect 538 -325 554 -247
rect 754 -325 770 -247
rect 538 -337 770 -325
rect -22 -338 315 -337
rect -201 -349 498 -338
rect -201 -383 -185 -349
rect -34 -383 326 -349
rect 482 -383 498 -349
rect -201 -392 498 -383
rect 112 -474 180 -392
rect 96 -482 196 -474
rect 96 -516 112 -482
rect 180 -516 196 -482
rect 96 -527 196 -516
rect 32 -729 66 -713
rect 32 -840 66 -824
rect 226 -729 260 -713
rect 226 -840 260 -824
rect 96 -938 196 -927
rect 96 -972 112 -938
rect 180 -972 196 -938
rect 96 -980 196 -972
rect 130 -1017 164 -980
rect 114 -1051 130 -1017
rect 164 -1051 180 -1017
<< viali >>
rect -516 781 -448 815
rect 740 781 808 815
rect -54 627 346 661
rect -596 473 -562 568
rect -274 231 -240 265
rect -402 115 -368 210
rect -86 157 -52 177
rect -86 143 -52 157
rect 854 473 888 568
rect 343 333 378 362
rect 343 328 344 333
rect 344 328 378 333
rect 129 234 163 268
rect -704 -130 -670 -96
rect -516 -132 -448 -98
rect 532 231 566 265
rect 660 115 694 210
rect 129 60 163 94
rect 128 -45 163 -11
rect 740 -132 808 -98
rect 962 -131 996 -97
rect -462 -327 -262 -249
rect 554 -325 754 -247
rect 32 -824 66 -729
rect 226 -824 260 -729
rect 112 -972 180 -938
<< metal1 >>
rect -522 815 -516 824
rect -448 815 -442 824
rect 734 815 740 824
rect 808 815 814 824
rect -528 781 -516 815
rect -448 781 -436 815
rect 728 781 740 815
rect 808 781 820 815
rect -522 772 -516 781
rect -448 772 -442 781
rect 734 772 740 781
rect 808 772 814 781
rect -1093 673 -1033 762
rect -979 691 -972 700
rect -763 661 1346 705
rect -763 627 -54 661
rect 346 627 1346 661
rect -763 609 1346 627
rect -596 574 -562 580
rect 854 574 888 580
rect -602 568 -556 574
rect -602 556 -596 568
rect -605 550 -596 556
rect -562 556 -556 568
rect 848 568 894 574
rect 848 556 854 568
rect -562 550 -553 556
rect -690 510 -605 538
rect 845 550 854 556
rect 888 556 894 568
rect 888 550 897 556
rect -553 510 -551 538
rect 843 510 845 538
rect -605 492 -596 498
rect -602 473 -596 492
rect -562 492 -553 498
rect 897 510 969 538
rect 845 492 854 498
rect -562 473 -556 492
rect -602 467 -556 473
rect 848 473 854 492
rect 888 492 897 498
rect 888 473 894 492
rect 848 467 894 473
rect -596 461 -562 467
rect 854 461 888 467
rect 337 362 384 368
rect 331 360 343 362
rect -402 330 343 360
rect -402 216 -368 330
rect 331 328 343 330
rect 378 328 390 362
rect 337 322 384 328
rect -280 265 -233 271
rect 123 268 169 275
rect -286 231 -274 265
rect -240 262 -228 265
rect 117 262 129 268
rect -240 234 129 262
rect 163 262 175 268
rect 526 265 573 274
rect 519 262 532 265
rect 163 234 532 262
rect -240 231 -228 234
rect -280 225 -233 231
rect 123 228 169 234
rect 519 231 532 234
rect 566 231 578 265
rect 526 225 573 231
rect 660 216 694 222
rect -408 210 -362 216
rect -408 115 -402 210
rect -368 115 -362 210
rect 654 210 700 216
rect -92 177 -40 183
rect -98 168 -86 177
rect -144 143 -86 168
rect -52 168 -40 177
rect 654 168 660 210
rect -52 143 660 168
rect -144 138 660 143
rect -92 137 -40 138
rect -408 109 -362 115
rect 654 115 660 138
rect 694 115 700 210
rect -402 103 -368 109
rect 119 94 173 110
rect 654 109 700 115
rect 660 103 694 109
rect 119 60 129 94
rect 163 60 173 94
rect 119 44 173 60
rect 119 1 171 4
rect 117 -2 174 1
rect 117 -54 119 -2
rect 171 -54 174 -2
rect 117 -65 174 -54
rect -716 -96 -658 -87
rect -716 -130 -704 -96
rect -670 -130 -658 -96
rect -716 -140 -658 -130
rect -704 -935 -670 -140
rect -528 -141 -516 -89
rect -448 -141 -436 -89
rect 728 -141 740 -89
rect 808 -141 820 -89
rect 950 -97 1008 -87
rect 950 -131 962 -97
rect 996 -131 1008 -97
rect 950 -140 1008 -131
rect -474 -249 -250 -243
rect -474 -327 -462 -249
rect -262 -327 -250 -249
rect -474 -333 -250 -327
rect 542 -247 766 -241
rect 542 -325 554 -247
rect 754 -325 766 -247
rect 542 -331 766 -325
rect 26 -729 72 -717
rect 220 -729 266 -717
rect 26 -824 32 -729
rect 66 -751 226 -729
rect 66 -803 120 -751
rect 172 -803 226 -751
rect 66 -824 226 -803
rect 260 -824 266 -729
rect 26 -836 72 -824
rect 220 -836 266 -824
rect 106 -935 186 -932
rect 962 -935 996 -140
rect -704 -938 996 -935
rect -704 -972 112 -938
rect 180 -972 996 -938
rect -704 -973 996 -972
rect 106 -978 186 -973
<< via1 >>
rect -516 815 -448 824
rect 740 815 808 824
rect -516 781 -448 815
rect 740 781 808 815
rect -516 772 -448 781
rect 740 772 808 781
rect -605 498 -596 550
rect -596 498 -562 550
rect -562 498 -553 550
rect 845 498 854 550
rect 854 498 888 550
rect 888 498 897 550
rect 119 -11 171 -2
rect 119 -45 128 -11
rect 128 -45 163 -11
rect 163 -45 171 -11
rect 119 -54 171 -45
rect -516 -98 -448 -89
rect -516 -132 -448 -98
rect -516 -141 -448 -132
rect 740 -98 808 -89
rect 740 -132 808 -98
rect 740 -141 808 -132
rect -462 -327 -262 -249
rect 554 -325 754 -247
rect 120 -803 172 -751
<< metal2 >>
rect -522 772 -516 824
rect -448 772 -442 824
rect 734 772 740 824
rect 808 772 814 824
rect -607 553 -551 562
rect -607 488 -551 497
rect -498 -83 -466 772
rect 117 0 173 9
rect 117 -65 173 -56
rect 758 -83 790 772
rect 843 552 899 561
rect 843 487 899 496
rect -516 -89 -448 -83
rect -516 -147 -448 -141
rect 740 -89 808 -83
rect 740 -147 808 -141
rect -474 -249 -250 -243
rect -474 -327 -462 -249
rect -262 -327 -250 -249
rect -474 -333 -250 -327
rect 542 -247 766 -241
rect 542 -325 554 -247
rect 754 -325 766 -247
rect 542 -331 766 -325
rect 118 -749 174 -740
rect 118 -814 174 -805
<< via2 >>
rect -607 550 -551 553
rect -607 498 -605 550
rect -605 498 -553 550
rect -553 498 -551 550
rect -607 497 -551 498
rect 117 -2 173 0
rect 117 -54 119 -2
rect 119 -54 171 -2
rect 171 -54 173 -2
rect 117 -56 173 -54
rect 843 550 899 552
rect 843 498 845 550
rect 845 498 897 550
rect 897 498 899 550
rect 843 496 899 498
rect -462 -327 -262 -249
rect 554 -325 754 -247
rect 118 -751 174 -749
rect 118 -803 120 -751
rect 120 -803 172 -751
rect 172 -803 174 -751
rect 118 -805 174 -803
<< metal3 >>
rect -607 559 -547 562
rect -613 554 -545 559
rect 843 557 904 561
rect 838 554 904 557
rect -613 553 904 554
rect -613 497 -607 553
rect -551 552 904 553
rect -551 497 843 552
rect -613 496 843 497
rect 899 496 904 552
rect -613 494 904 496
rect -613 489 -545 494
rect 838 491 904 494
rect -607 488 -547 489
rect 843 487 904 491
rect 116 5 176 35
rect 112 0 178 5
rect 112 -56 117 0
rect 173 -56 178 0
rect 112 -62 178 -56
rect -468 -249 -256 -243
rect -468 -327 -462 -249
rect -262 -327 -256 -249
rect -468 -333 -256 -327
rect 116 -744 176 -62
rect 548 -247 760 -241
rect 548 -325 554 -247
rect 754 -325 760 -247
rect 548 -331 760 -325
rect 113 -749 179 -744
rect 113 -805 118 -749
rect 174 -805 179 -749
rect 113 -810 179 -805
rect 116 -814 176 -810
<< via3 >>
rect -462 -327 -262 -249
rect 554 -325 754 -247
<< metal4 >>
rect 553 -247 969 -246
rect -690 -249 -261 -248
rect -690 -327 -462 -249
rect -262 -327 -261 -249
rect 553 -325 554 -247
rect 754 -325 969 -247
rect 553 -326 969 -325
rect -690 -328 -261 -327
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1037 0 1 113
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_1
timestamp 1644511149
transform 1 0 1313 0 1 113
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_2
timestamp 1644511149
transform -1 0 -758 0 1 113
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_3
timestamp 1644511149
transform -1 0 -1034 0 1 113
box -38 -48 314 592
<< labels >>
rlabel metal1 -690 524 -690 524 7 phi1b
rlabel metal4 -690 -287 -690 -287 7 inp
rlabel locali -135 -111 -135 -111 7 FP
rlabel locali 427 -109 427 -109 3 FN
rlabel locali 144 -337 144 -337 1 tail
rlabel locali 824 342 824 342 3 low
rlabel locali -532 341 -532 341 7 high
rlabel pdiff -183 201 -183 201 7 pfetw
rlabel pdiff 475 195 475 195 3 pfete
<< end >>
