magic
tech sky130B
timestamp 1654741520
use cap_10_10__side_x2  cap_10_10__side_x2_0
array 0 0 1528 0 5 -1360
timestamp 1654741520
transform 0 1 7174 -1 0 4083
box -356 -183 1172 1177
use cap_10_10__side_x2  cap_10_10__side_x2_1
array 0 0 1528 0 5 -1360
timestamp 1654741520
transform 0 -1 1368 1 0 -981
box -356 -183 1172 1177
use cap_10_10__side_x2  cap_10_10__side_x2_2
timestamp 1654741520
transform 1 0 -981 0 1 374
box -356 -183 1172 1177
use cap_10_10__side_x2  cap_10_10__side_x2_3
timestamp 1654741520
transform -1 0 9523 0 -1 2728
box -356 -183 1172 1177
use cap_10_10__side_x2  cap_10_10__side_x2_4
timestamp 1654741520
transform -1 0 9523 0 -1 1368
box -356 -183 1172 1177
use cap_10_10__side_x2  cap_10_10__side_x2_5
timestamp 1654741520
transform 1 0 -981 0 1 1734
box -356 -183 1172 1177
use cap_10_10_edge_x2  cap_10_10_edge_x2_0
timestamp 1654741520
transform 1 0 -981 0 1 -986
box -356 -351 1172 1177
use cap_10_10_edge_x2  cap_10_10_edge_x2_1
timestamp 1654741520
transform 0 -1 9528 1 0 -981
box -356 -351 1172 1177
use cap_10_10_edge_x2  cap_10_10_edge_x2_2
timestamp 1654741520
transform -1 0 9523 0 -1 4088
box -356 -351 1172 1177
use cap_10_10_edge_x2  cap_10_10_edge_x2_3
timestamp 1654741520
transform 0 1 -986 -1 0 4083
box -356 -351 1172 1177
use cap_10_10_x2  cap_10_10_x2_0
array 0 5 1360 0 1 1360
timestamp 1654741520
transform 1 0 379 0 1 374
box -188 -183 1172 1177
<< end >>
