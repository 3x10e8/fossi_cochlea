magic
tech sky130A
magscale 1 2
timestamp 1654658877
<< error_s >>
rect 6859 27015 6986 27050
rect 6799 26955 7046 26990
rect 13789 26725 14198 27045
rect 13798 25875 14207 26195
rect 13790 25023 14199 25343
rect 13785 23322 14194 23642
rect 13795 22427 14204 22747
rect 13786 21544 14195 21864
rect 13805 19840 14214 20160
rect 13800 18958 14209 19278
rect 13811 18061 14220 18381
rect 13800 16368 14209 16688
rect 13806 15470 14215 15790
rect 13809 14577 14218 14897
rect 13814 12881 14223 13201
rect 13809 11988 14218 12308
rect 13815 11093 14224 11413
rect 13813 9395 14222 9715
rect 13810 8502 14219 8822
rect 13806 7610 14208 7930
rect 13808 5914 14210 6234
rect 13812 5020 14214 5340
rect 13804 4126 14206 4446
rect 13812 2430 14214 2750
rect 13803 1541 14212 1861
rect 13794 676 14203 996
<< metal2 >>
rect -1289 28654 -1280 28710
rect -1224 28654 -1215 28710
rect -901 28387 -892 28443
rect -836 28387 -827 28443
rect -87 28308 -78 28364
rect -22 28308 -13 28364
rect 1707 28304 1716 28365
rect 1776 28304 1785 28365
rect 13920 28363 13977 28372
rect 13920 28296 13977 28305
rect 15274 28364 15331 28373
rect 15274 28298 15331 28307
rect 20816 28365 20877 28374
rect 20816 28297 20877 28306
rect 22117 28363 22174 28372
rect 22117 28298 22174 28307
<< via2 >>
rect -1280 28654 -1224 28710
rect -892 28387 -836 28443
rect -78 28308 -22 28364
rect 1716 28304 1776 28365
rect 13920 28305 13977 28363
rect 15274 28307 15331 28364
rect 20816 28306 20877 28365
rect 22117 28307 22174 28363
<< metal3 >>
rect -1301 28714 -1203 28733
rect -1301 28650 -1284 28714
rect -1220 28650 -1203 28714
rect -1301 28635 -1203 28650
rect -913 28447 -815 28467
rect -913 28383 -896 28447
rect -832 28383 -815 28447
rect -913 28369 -815 28383
rect 685 28369 1079 28508
rect 1707 28369 1788 28370
rect 14601 28369 14875 28567
rect 21374 28376 21476 28547
rect 20802 28375 21476 28376
rect -91 28365 1788 28369
rect -91 28364 1716 28365
rect -91 28308 -78 28364
rect -22 28308 1716 28364
rect -91 28304 1716 28308
rect 1776 28304 1788 28365
rect -91 28300 1788 28304
rect -1540 27972 -1220 28197
rect -1800 27929 -1220 27972
rect -1800 27695 -1775 27929
rect -1541 27695 -1220 27929
rect -1800 27652 -1220 27695
rect -900 27972 -580 28204
rect -900 27929 -320 27972
rect -900 27695 -579 27929
rect -345 27695 -320 27929
rect -900 27652 -320 27695
rect 685 27689 1079 28300
rect 1707 28299 1788 28300
rect 13909 28364 15339 28369
rect 13909 28363 15274 28364
rect 13909 28305 13920 28363
rect 13977 28307 15274 28363
rect 15331 28307 15339 28364
rect 13977 28305 15339 28307
rect 13909 28297 15339 28305
rect 20802 28365 22191 28375
rect 20802 28306 20816 28365
rect 20877 28363 22191 28365
rect 20877 28307 22117 28363
rect 22174 28307 22191 28363
rect 20877 28306 22191 28307
rect 20802 28297 22191 28306
rect 14601 27728 14875 28297
rect 20802 27727 20911 28297
rect -1540 27609 -580 27652
rect -1540 27375 -1219 27609
rect -901 27375 -580 27609
rect -1540 27332 -580 27375
rect -1800 27289 -1220 27332
rect -1800 27055 -1775 27289
rect -1541 27055 -1220 27289
rect -1800 27012 -1220 27055
rect -900 27289 -320 27332
rect -900 27055 -579 27289
rect -345 27055 -320 27289
rect -900 27012 -320 27055
rect -1540 26969 -580 27012
rect -1540 26735 -1219 26969
rect -901 26735 -580 26969
rect -1540 26692 -580 26735
rect 13789 26725 14198 27045
rect -1800 26649 -1220 26692
rect -1800 26415 -1775 26649
rect -1541 26415 -1220 26649
rect -1800 26372 -1220 26415
rect -900 26649 -320 26692
rect -900 26415 -579 26649
rect -345 26415 -320 26649
rect -900 26372 -320 26415
rect -1540 26329 -580 26372
rect -1540 26095 -1219 26329
rect -901 26095 -580 26329
rect -1540 26052 -580 26095
rect -1800 26009 -1220 26052
rect -1800 25775 -1775 26009
rect -1541 25775 -1220 26009
rect -1800 25732 -1220 25775
rect -900 26009 2 26052
rect -900 25775 -579 26009
rect -345 25775 2 26009
rect 13798 25875 14207 26195
rect -900 25732 2 25775
rect -1540 25689 -580 25732
rect -1540 25455 -1219 25689
rect -901 25455 -580 25689
rect -1540 25412 -580 25455
rect -1800 25369 -1220 25412
rect -1800 25135 -1775 25369
rect -1541 25135 -1220 25369
rect -1800 25092 -1220 25135
rect -900 25369 -320 25412
rect -900 25135 -579 25369
rect -345 25135 -320 25369
rect -900 25092 -320 25135
rect -1540 25049 -580 25092
rect -1540 24815 -1219 25049
rect -901 24815 -580 25049
rect 13790 25023 14199 25343
rect -1540 24772 -580 24815
rect -1800 24729 -1220 24772
rect -1800 24495 -1775 24729
rect -1541 24495 -1220 24729
rect -1800 24452 -1220 24495
rect -900 24729 2 24772
rect -900 24495 -579 24729
rect -345 24495 2 24729
rect -900 24452 2 24495
rect -1540 24409 -580 24452
rect -1540 24175 -1219 24409
rect -901 24175 -580 24409
rect -1540 24132 -580 24175
rect -1800 24089 -1220 24132
rect -1800 23855 -1775 24089
rect -1541 23855 -1220 24089
rect -1800 23812 -1220 23855
rect -900 24089 -320 24132
rect -900 23855 -579 24089
rect -345 23855 -320 24089
rect -900 23812 -320 23855
rect -1540 23769 -580 23812
rect -1540 23535 -1219 23769
rect -901 23535 -580 23769
rect -1540 23492 -580 23535
rect -1800 23449 -1220 23492
rect -1800 23215 -1775 23449
rect -1541 23215 -1220 23449
rect -1800 23172 -1220 23215
rect -900 23449 2 23492
rect -900 23215 -579 23449
rect -345 23215 2 23449
rect 13785 23322 14194 23642
rect -900 23172 2 23215
rect -1540 23129 -580 23172
rect -1540 22895 -1219 23129
rect -901 22895 -580 23129
rect -1540 22852 -580 22895
rect -1800 22809 -1220 22852
rect -1800 22575 -1775 22809
rect -1541 22575 -1220 22809
rect -1800 22532 -1220 22575
rect -900 22809 -320 22852
rect -900 22575 -579 22809
rect -345 22575 -320 22809
rect -900 22532 -320 22575
rect -1540 22489 -580 22532
rect -1540 22255 -1219 22489
rect -901 22255 -580 22489
rect 13795 22427 14204 22747
rect -1540 22212 -580 22255
rect -1800 22169 -1220 22212
rect -1800 21935 -1775 22169
rect -1541 21935 -1220 22169
rect -1800 21892 -1220 21935
rect -900 22169 2 22212
rect -900 21935 -579 22169
rect -345 21935 2 22169
rect -900 21892 2 21935
rect -1540 21849 -580 21892
rect -1540 21615 -1219 21849
rect -901 21615 -580 21849
rect -1540 21572 -580 21615
rect -1800 21529 -1220 21572
rect -1800 21295 -1775 21529
rect -1541 21295 -1220 21529
rect -1800 21252 -1220 21295
rect -900 21529 -320 21572
rect 13786 21544 14195 21864
rect -900 21295 -579 21529
rect -345 21295 -320 21529
rect -900 21252 -320 21295
rect -1540 21209 -580 21252
rect -1540 20975 -1219 21209
rect -901 20975 -580 21209
rect -1540 20932 -580 20975
rect -1800 20889 -1220 20932
rect -1800 20655 -1775 20889
rect -1541 20655 -1220 20889
rect -1800 20612 -1220 20655
rect -900 20889 2 20932
rect -900 20655 -579 20889
rect -345 20655 2 20889
rect -900 20612 2 20655
rect -1540 20569 -580 20612
rect -1540 20335 -1219 20569
rect -901 20335 -580 20569
rect -1540 20292 -580 20335
rect -1800 20249 -1220 20292
rect -1800 20015 -1775 20249
rect -1541 20015 -1220 20249
rect -1800 19972 -1220 20015
rect -900 20249 -320 20292
rect -900 20015 -579 20249
rect -345 20015 -320 20249
rect -900 19972 -320 20015
rect -1540 19929 -580 19972
rect -1540 19695 -1219 19929
rect -901 19695 -580 19929
rect 13805 19840 14214 20160
rect -1540 19652 -580 19695
rect -1800 19609 -1220 19652
rect -1800 19375 -1775 19609
rect -1541 19375 -1220 19609
rect -1800 19332 -1220 19375
rect -900 19609 2 19652
rect -900 19375 -579 19609
rect -345 19375 2 19609
rect -900 19332 2 19375
rect -1540 19289 -580 19332
rect -1540 19055 -1219 19289
rect -901 19055 -580 19289
rect -1540 19012 -580 19055
rect -1800 18969 -1220 19012
rect -1800 18735 -1775 18969
rect -1541 18735 -1220 18969
rect -1800 18692 -1220 18735
rect -900 18969 -320 19012
rect -900 18735 -579 18969
rect -345 18735 -320 18969
rect 13800 18958 14209 19278
rect -900 18692 -320 18735
rect -1540 18649 -580 18692
rect -1540 18415 -1219 18649
rect -901 18415 -580 18649
rect -1540 18372 -580 18415
rect -1800 18329 -1220 18372
rect -1800 18095 -1775 18329
rect -1541 18095 -1220 18329
rect -1800 18052 -1220 18095
rect -900 18329 2 18372
rect -900 18095 -579 18329
rect -345 18095 2 18329
rect -900 18052 2 18095
rect 13811 18061 14220 18381
rect -1540 18009 -580 18052
rect -1540 17775 -1219 18009
rect -901 17775 -580 18009
rect -1540 17732 -580 17775
rect -1800 17689 -1220 17732
rect -1800 17455 -1775 17689
rect -1541 17455 -1220 17689
rect -1800 17412 -1220 17455
rect -900 17689 -320 17732
rect -900 17455 -579 17689
rect -345 17455 -320 17689
rect -900 17412 -320 17455
rect -1540 17369 -580 17412
rect -1540 17135 -1219 17369
rect -901 17135 -580 17369
rect -1540 17092 -580 17135
rect -1800 17049 -1220 17092
rect -1800 16815 -1775 17049
rect -1541 16815 -1220 17049
rect -1800 16772 -1220 16815
rect -900 17049 2 17092
rect -900 16815 -579 17049
rect -345 16815 2 17049
rect -900 16772 2 16815
rect -1540 16729 -580 16772
rect -1540 16495 -1219 16729
rect -901 16495 -580 16729
rect -1540 16452 -580 16495
rect -1800 16409 -1220 16452
rect -1800 16175 -1775 16409
rect -1541 16175 -1220 16409
rect -1800 16132 -1220 16175
rect -900 16409 -320 16452
rect -900 16175 -579 16409
rect -345 16175 -320 16409
rect 13800 16368 14209 16688
rect -900 16132 -320 16175
rect -1540 16089 -580 16132
rect -1540 15855 -1219 16089
rect -901 15855 -580 16089
rect -1540 15812 -580 15855
rect -1800 15769 -1220 15812
rect -1800 15535 -1775 15769
rect -1541 15535 -1220 15769
rect -1800 15492 -1220 15535
rect -900 15769 2 15812
rect -900 15535 -579 15769
rect -345 15535 2 15769
rect -900 15492 2 15535
rect -1540 15449 -580 15492
rect 13806 15470 14215 15790
rect -1540 15215 -1219 15449
rect -901 15215 -580 15449
rect -1540 15172 -580 15215
rect -1800 15129 -1220 15172
rect -1800 14895 -1775 15129
rect -1541 14895 -1220 15129
rect -1800 14852 -1220 14895
rect -900 15129 -320 15172
rect -900 14895 -579 15129
rect -345 14895 -320 15129
rect -900 14852 -320 14895
rect -1540 14809 -580 14852
rect -1540 14575 -1219 14809
rect -901 14575 -580 14809
rect 13809 14577 14218 14897
rect -1540 14532 -580 14575
rect -1800 14489 -1220 14532
rect -1800 14255 -1775 14489
rect -1541 14255 -1220 14489
rect -1800 14212 -1220 14255
rect -900 14489 2 14532
rect -900 14255 -579 14489
rect -345 14255 2 14489
rect -900 14212 2 14255
rect -1540 14169 -580 14212
rect -1540 13935 -1219 14169
rect -901 13935 -580 14169
rect -1540 13892 -580 13935
rect -1800 13849 -1220 13892
rect -1800 13615 -1775 13849
rect -1541 13615 -1220 13849
rect -1800 13572 -1220 13615
rect -900 13849 -320 13892
rect -900 13615 -579 13849
rect -345 13615 -320 13849
rect -900 13572 -320 13615
rect -1540 13529 -580 13572
rect -1540 13295 -1219 13529
rect -901 13295 -580 13529
rect -1540 13252 -580 13295
rect -1800 13209 -1220 13252
rect -1800 12975 -1775 13209
rect -1541 12975 -1220 13209
rect -1800 12932 -1220 12975
rect -900 13209 2 13252
rect -900 12975 -579 13209
rect -345 12975 2 13209
rect -900 12932 2 12975
rect -1540 12889 -580 12932
rect -1540 12655 -1219 12889
rect -901 12655 -580 12889
rect 13814 12881 14223 13201
rect -1540 12612 -580 12655
rect -1800 12569 -1220 12612
rect -1800 12335 -1775 12569
rect -1541 12335 -1220 12569
rect -1800 12292 -1220 12335
rect -900 12569 -320 12612
rect -900 12335 -579 12569
rect -345 12335 -320 12569
rect -900 12292 -320 12335
rect -1540 12249 -580 12292
rect -1540 12015 -1219 12249
rect -901 12015 -580 12249
rect -1540 11972 -580 12015
rect 13809 11988 14218 12308
rect -1800 11929 -1220 11972
rect -1800 11695 -1775 11929
rect -1541 11695 -1220 11929
rect -1800 11652 -1220 11695
rect -900 11929 2 11972
rect -900 11695 -579 11929
rect -345 11695 2 11929
rect -900 11652 2 11695
rect -1540 11609 -580 11652
rect -1540 11375 -1219 11609
rect -901 11375 -580 11609
rect -1540 11332 -580 11375
rect -1800 11289 -1220 11332
rect -1800 11055 -1775 11289
rect -1541 11055 -1220 11289
rect -1800 11012 -1220 11055
rect -900 11289 -320 11332
rect -900 11055 -579 11289
rect -345 11055 -320 11289
rect 13815 11093 14224 11413
rect -900 11012 -320 11055
rect -1540 10969 -580 11012
rect -1540 10735 -1219 10969
rect -901 10735 -580 10969
rect -1540 10692 -580 10735
rect -1800 10649 -1220 10692
rect -1800 10415 -1775 10649
rect -1541 10415 -1220 10649
rect -1800 10372 -1220 10415
rect -900 10649 2 10692
rect -900 10415 -579 10649
rect -345 10415 2 10649
rect -900 10372 2 10415
rect -1540 10329 -580 10372
rect -1540 10095 -1219 10329
rect -901 10095 -580 10329
rect -1540 10052 -580 10095
rect -1800 10009 -1220 10052
rect -1800 9775 -1775 10009
rect -1541 9775 -1220 10009
rect -1800 9732 -1220 9775
rect -900 10009 -320 10052
rect -900 9775 -579 10009
rect -345 9775 -320 10009
rect -900 9732 -320 9775
rect -1540 9689 -580 9732
rect -1540 9455 -1219 9689
rect -901 9455 -580 9689
rect -1540 9412 -580 9455
rect -1800 9369 -1220 9412
rect -1800 9135 -1775 9369
rect -1541 9135 -1220 9369
rect -1800 9092 -1220 9135
rect -900 9369 2 9412
rect 13813 9395 14222 9715
rect -900 9135 -579 9369
rect -345 9135 2 9369
rect -900 9092 2 9135
rect -1540 9049 -580 9092
rect -1540 8815 -1219 9049
rect -901 8815 -580 9049
rect -1540 8772 -580 8815
rect -1800 8729 -1220 8772
rect -1800 8495 -1775 8729
rect -1541 8495 -1220 8729
rect -1800 8452 -1220 8495
rect -900 8729 -320 8772
rect -900 8495 -579 8729
rect -345 8495 -320 8729
rect 13810 8502 14219 8822
rect -900 8452 -320 8495
rect -1540 8409 -580 8452
rect -1540 8175 -1219 8409
rect -901 8175 -580 8409
rect -1540 8132 -580 8175
rect -1800 8089 -1220 8132
rect -1800 7855 -1775 8089
rect -1541 7855 -1220 8089
rect -1800 7812 -1220 7855
rect -900 8089 2 8132
rect -900 7855 -579 8089
rect -345 7855 2 8089
rect -900 7812 2 7855
rect -1540 7769 -580 7812
rect -1540 7535 -1219 7769
rect -901 7535 -580 7769
rect 13806 7610 14208 7930
rect -1540 7492 -580 7535
rect -1800 7449 -1220 7492
rect -1800 7215 -1775 7449
rect -1541 7215 -1220 7449
rect -1800 7172 -1220 7215
rect -900 7449 -320 7492
rect -900 7215 -579 7449
rect -345 7215 -320 7449
rect -900 7172 -320 7215
rect -1540 7129 -580 7172
rect -1540 6895 -1219 7129
rect -901 6895 -580 7129
rect -1540 6852 -580 6895
rect -1800 6809 -1220 6852
rect -1800 6575 -1775 6809
rect -1541 6575 -1220 6809
rect -1800 6532 -1220 6575
rect -900 6809 2 6852
rect -900 6575 -579 6809
rect -345 6575 2 6809
rect -900 6532 2 6575
rect -1540 6489 -580 6532
rect -1540 6255 -1219 6489
rect -901 6255 -580 6489
rect -1540 6212 -580 6255
rect -1800 6169 -1220 6212
rect -1800 5935 -1775 6169
rect -1541 5935 -1220 6169
rect -1800 5892 -1220 5935
rect -900 6169 -320 6212
rect -900 5935 -579 6169
rect -345 5935 -320 6169
rect -900 5892 -320 5935
rect 13808 5914 14210 6234
rect -1540 5849 -580 5892
rect -1540 5615 -1219 5849
rect -901 5615 -580 5849
rect -1540 5572 -580 5615
rect -1800 5529 -1220 5572
rect -1800 5295 -1775 5529
rect -1541 5295 -1220 5529
rect -1800 5252 -1220 5295
rect -900 5529 2 5572
rect -900 5295 -579 5529
rect -345 5295 2 5529
rect -900 5252 2 5295
rect -1540 5209 -580 5252
rect -1540 4975 -1219 5209
rect -901 4975 -580 5209
rect 13812 5020 14214 5340
rect -1540 4932 -580 4975
rect -1800 4889 -1220 4932
rect -1800 4655 -1775 4889
rect -1541 4655 -1220 4889
rect -1800 4612 -1220 4655
rect -900 4889 -320 4932
rect -900 4655 -579 4889
rect -345 4655 -320 4889
rect -900 4612 -320 4655
rect -1540 4569 -580 4612
rect -1540 4335 -1219 4569
rect -901 4335 -580 4569
rect -1540 4292 -580 4335
rect -1800 4249 -1220 4292
rect -1800 4015 -1775 4249
rect -1541 4015 -1220 4249
rect -1800 3972 -1220 4015
rect -900 4249 2 4292
rect -900 4015 -579 4249
rect -345 4015 2 4249
rect 13804 4126 14206 4446
rect -900 3972 2 4015
rect -1540 3929 -580 3972
rect -1540 3695 -1219 3929
rect -901 3695 -580 3929
rect -1540 3652 -580 3695
rect -1800 3609 -1220 3652
rect -1800 3375 -1775 3609
rect -1541 3375 -1220 3609
rect -1800 3332 -1220 3375
rect -900 3609 -320 3652
rect -900 3375 -579 3609
rect -345 3375 -320 3609
rect -900 3332 -320 3375
rect -1540 3289 -580 3332
rect -1540 3055 -1219 3289
rect -901 3055 -580 3289
rect -1540 3012 -580 3055
rect -1800 2969 -1220 3012
rect -1800 2735 -1775 2969
rect -1541 2735 -1220 2969
rect -1800 2692 -1220 2735
rect -900 2969 2 3012
rect -900 2735 -579 2969
rect -345 2735 2 2969
rect -900 2692 2 2735
rect -1540 2649 -580 2692
rect -1540 2415 -1219 2649
rect -901 2415 -580 2649
rect 13812 2430 14214 2750
rect -1540 2372 -580 2415
rect -1800 2329 -1220 2372
rect -1800 2095 -1775 2329
rect -1541 2095 -1220 2329
rect -1800 2052 -1220 2095
rect -900 2329 -320 2372
rect -900 2095 -579 2329
rect -345 2095 -320 2329
rect -900 2052 -320 2095
rect -1540 2009 -580 2052
rect -1540 1775 -1219 2009
rect -901 1775 -580 2009
rect -1540 1732 -580 1775
rect -1800 1689 -1220 1732
rect -1800 1455 -1775 1689
rect -1541 1455 -1220 1689
rect -1800 1412 -1220 1455
rect -1540 372 -1220 1412
rect -900 1689 2 1732
rect -900 1455 -579 1689
rect -345 1455 2 1689
rect 13803 1541 14212 1861
rect -900 1412 2 1455
rect -900 372 -580 1412
rect 13794 676 14203 996
rect -1485 301 -1276 307
rect -1485 112 -1479 301
rect -1282 112 -1276 301
rect -1485 -1285 -1276 112
rect -844 301 -635 307
rect -844 112 -838 301
rect -641 112 -635 301
rect -844 -644 -635 112
rect 2 -343 322 13
rect 2 -577 45 -343
rect 279 -577 322 -343
rect 2 -578 322 -577
rect 642 -343 962 -318
rect 642 -577 685 -343
rect 919 -577 962 -343
rect 642 -578 962 -577
rect 1282 -343 1602 2
rect 1282 -577 1325 -343
rect 1559 -577 1602 -343
rect 1282 -578 1602 -577
rect 1922 -343 2242 -318
rect 1922 -577 1965 -343
rect 2199 -577 2242 -343
rect 1922 -578 2242 -577
rect 2562 -343 2882 2
rect 2562 -577 2605 -343
rect 2839 -577 2882 -343
rect 2562 -578 2882 -577
rect 3202 -343 3522 -318
rect 3202 -577 3245 -343
rect 3479 -577 3522 -343
rect 3202 -578 3522 -577
rect 3842 -343 4162 2
rect 3842 -577 3885 -343
rect 4119 -577 4162 -343
rect 3842 -578 4162 -577
rect 4482 -343 4802 -318
rect 4482 -577 4525 -343
rect 4759 -577 4802 -343
rect 4482 -578 4802 -577
rect 5122 -343 5442 2
rect 5122 -577 5165 -343
rect 5399 -577 5442 -343
rect 5122 -578 5442 -577
rect 5762 -343 6082 -318
rect 5762 -577 5805 -343
rect 6039 -577 6082 -343
rect 5762 -578 6082 -577
rect 6402 -343 6722 2
rect 6402 -577 6445 -343
rect 6679 -577 6722 -343
rect 6402 -578 6722 -577
rect 7042 -343 7362 -318
rect 7042 -577 7085 -343
rect 7319 -577 7362 -343
rect 7042 -578 7362 -577
rect 7682 -343 8002 2
rect 7682 -577 7725 -343
rect 7959 -577 8002 -343
rect 7682 -578 8002 -577
rect 8322 -343 8642 -318
rect 8322 -577 8365 -343
rect 8599 -577 8642 -343
rect 8322 -578 8642 -577
rect 8962 -343 9282 2
rect 8962 -577 9005 -343
rect 9239 -577 9282 -343
rect 8962 -578 9282 -577
rect 9602 -343 9922 -318
rect 9602 -577 9645 -343
rect 9879 -577 9922 -343
rect 9602 -578 9922 -577
rect 10242 -343 10562 2
rect 10242 -577 10285 -343
rect 10519 -577 10562 -343
rect 10242 -578 10562 -577
rect 10882 -343 11202 -318
rect 10882 -577 10925 -343
rect 11159 -577 11202 -343
rect 10882 -578 11202 -577
rect 11522 -343 11842 2
rect 11522 -577 11565 -343
rect 11799 -577 11842 -343
rect 11522 -578 11842 -577
rect 12162 -343 12482 -318
rect 12162 -577 12205 -343
rect 12439 -577 12482 -343
rect 12162 -578 12482 -577
rect 12802 -343 13122 2
rect 12802 -577 12845 -343
rect 13079 -577 13122 -343
rect 12802 -578 13122 -577
rect 13442 -343 13762 -318
rect 13442 -577 13485 -343
rect 13719 -577 13762 -343
rect 13442 -578 13762 -577
rect 14082 -343 14402 -318
rect 14082 -577 14125 -343
rect 14359 -577 14402 -343
rect 14082 -578 14402 -577
rect 14722 -343 15042 -318
rect 14722 -577 14765 -343
rect 14999 -577 15042 -343
rect 14722 -578 15042 -577
rect 15362 -343 15682 2
rect 15362 -577 15405 -343
rect 15639 -577 15682 -343
rect 15362 -578 15682 -577
rect 16002 -343 16322 -318
rect 16002 -577 16045 -343
rect 16279 -577 16322 -343
rect 16002 -578 16322 -577
rect 16642 -343 16962 2
rect 16642 -577 16685 -343
rect 16919 -577 16962 -343
rect 16642 -578 16962 -577
rect 17282 -343 17602 -318
rect 17282 -577 17325 -343
rect 17559 -577 17602 -343
rect 17282 -578 17602 -577
rect 17922 -343 18242 2
rect 17922 -577 17965 -343
rect 18199 -577 18242 -343
rect 17922 -578 18242 -577
rect 18562 -343 18882 -318
rect 18562 -577 18605 -343
rect 18839 -577 18882 -343
rect 18562 -578 18882 -577
rect 19202 -343 19522 2
rect 19202 -577 19245 -343
rect 19479 -577 19522 -343
rect 19202 -578 19522 -577
rect 19842 -343 20162 -318
rect 19842 -577 19885 -343
rect 20119 -577 20162 -343
rect 19842 -578 20162 -577
rect 20482 -343 20802 2
rect 20482 -577 20525 -343
rect 20759 -577 20802 -343
rect 20482 -578 20802 -577
rect 21122 -343 21442 -318
rect 21122 -577 21165 -343
rect 21399 -577 21442 -343
rect 21122 -578 21442 -577
rect 21762 -343 22082 -318
rect 21762 -577 21805 -343
rect 22039 -577 22082 -343
rect 21762 -578 22082 -577
rect 22402 -343 22722 -318
rect 22402 -577 22445 -343
rect 22679 -577 22722 -343
rect 22402 -578 22722 -577
rect 23042 -343 23362 -318
rect 23042 -577 23085 -343
rect 23319 -577 23362 -343
rect 23042 -578 23362 -577
rect 23682 -343 24002 -318
rect 23682 -577 23725 -343
rect 23959 -577 24002 -343
rect 23682 -578 24002 -577
rect 24322 -343 24642 -318
rect 24322 -577 24365 -343
rect 24599 -577 24642 -343
rect 24322 -578 24642 -577
rect 24962 -343 25282 -318
rect 24962 -577 25005 -343
rect 25239 -577 25282 -343
rect 24962 -578 25282 -577
rect -844 -833 -838 -644
rect -641 -833 -635 -644
rect -844 -837 -635 -833
rect -570 -898 25922 -578
rect 322 -899 642 -898
rect 322 -1217 365 -899
rect 599 -1217 642 -899
rect 322 -1218 642 -1217
rect 962 -899 1282 -898
rect 962 -1217 1005 -899
rect 1239 -1217 1282 -899
rect 962 -1218 1282 -1217
rect 1602 -899 1922 -898
rect 1602 -1217 1645 -899
rect 1879 -1217 1922 -899
rect 1602 -1218 1922 -1217
rect 2242 -899 2562 -898
rect 2242 -1217 2285 -899
rect 2519 -1217 2562 -899
rect 2242 -1218 2562 -1217
rect 2882 -899 3202 -898
rect 2882 -1217 2925 -899
rect 3159 -1217 3202 -899
rect 2882 -1218 3202 -1217
rect 3522 -899 3842 -898
rect 3522 -1217 3565 -899
rect 3799 -1217 3842 -899
rect 3522 -1218 3842 -1217
rect 4162 -899 4482 -898
rect 4162 -1217 4205 -899
rect 4439 -1217 4482 -899
rect 4162 -1218 4482 -1217
rect 4802 -899 5122 -898
rect 4802 -1217 4845 -899
rect 5079 -1217 5122 -899
rect 4802 -1218 5122 -1217
rect 5442 -899 5762 -898
rect 5442 -1217 5485 -899
rect 5719 -1217 5762 -899
rect 5442 -1218 5762 -1217
rect 6082 -899 6402 -898
rect 6082 -1217 6125 -899
rect 6359 -1217 6402 -899
rect 6082 -1218 6402 -1217
rect 6722 -899 7042 -898
rect 6722 -1217 6765 -899
rect 6999 -1217 7042 -899
rect 6722 -1218 7042 -1217
rect 7362 -899 7682 -898
rect 7362 -1217 7405 -899
rect 7639 -1217 7682 -899
rect 7362 -1218 7682 -1217
rect 8002 -899 8322 -898
rect 8002 -1217 8045 -899
rect 8279 -1217 8322 -899
rect 8002 -1218 8322 -1217
rect 8642 -899 8962 -898
rect 8642 -1217 8685 -899
rect 8919 -1217 8962 -899
rect 8642 -1218 8962 -1217
rect 9282 -899 9602 -898
rect 9282 -1217 9325 -899
rect 9559 -1217 9602 -899
rect 9282 -1218 9602 -1217
rect 9922 -899 10242 -898
rect 9922 -1217 9965 -899
rect 10199 -1217 10242 -899
rect 9922 -1218 10242 -1217
rect 10562 -899 10882 -898
rect 10562 -1217 10605 -899
rect 10839 -1217 10882 -899
rect 10562 -1218 10882 -1217
rect 11202 -899 11522 -898
rect 11202 -1217 11245 -899
rect 11479 -1217 11522 -899
rect 11202 -1218 11522 -1217
rect 11842 -899 12162 -898
rect 11842 -1217 11885 -899
rect 12119 -1217 12162 -899
rect 11842 -1218 12162 -1217
rect 12482 -899 12802 -898
rect 12482 -1217 12525 -899
rect 12759 -1217 12802 -899
rect 12482 -1218 12802 -1217
rect 13122 -899 13442 -898
rect 13122 -1217 13165 -899
rect 13399 -1217 13442 -899
rect 13122 -1218 13442 -1217
rect 13762 -899 14082 -898
rect 13762 -1217 13805 -899
rect 14039 -1217 14082 -899
rect 13762 -1218 14082 -1217
rect 14402 -899 14722 -898
rect 14402 -1217 14445 -899
rect 14679 -1217 14722 -899
rect 14402 -1218 14722 -1217
rect 15042 -899 15362 -898
rect 15042 -1217 15085 -899
rect 15319 -1217 15362 -899
rect 15042 -1218 15362 -1217
rect 15682 -899 16002 -898
rect 15682 -1217 15725 -899
rect 15959 -1217 16002 -899
rect 15682 -1218 16002 -1217
rect 16322 -899 16642 -898
rect 16322 -1217 16365 -899
rect 16599 -1217 16642 -899
rect 16322 -1218 16642 -1217
rect 16962 -899 17282 -898
rect 16962 -1217 17005 -899
rect 17239 -1217 17282 -899
rect 16962 -1218 17282 -1217
rect 17602 -899 17922 -898
rect 17602 -1217 17645 -899
rect 17879 -1217 17922 -899
rect 17602 -1218 17922 -1217
rect 18242 -899 18562 -898
rect 18242 -1217 18285 -899
rect 18519 -1217 18562 -899
rect 18242 -1218 18562 -1217
rect 18882 -899 19202 -898
rect 18882 -1217 18925 -899
rect 19159 -1217 19202 -899
rect 18882 -1218 19202 -1217
rect 19522 -899 19842 -898
rect 19522 -1217 19565 -899
rect 19799 -1217 19842 -899
rect 19522 -1218 19842 -1217
rect 20162 -899 20482 -898
rect 20162 -1217 20205 -899
rect 20439 -1217 20482 -899
rect 20162 -1218 20482 -1217
rect 20802 -899 21122 -898
rect 20802 -1217 20845 -899
rect 21079 -1217 21122 -899
rect 20802 -1218 21122 -1217
rect 21442 -899 21762 -898
rect 21442 -1217 21485 -899
rect 21719 -1217 21762 -899
rect 21442 -1218 21762 -1217
rect 22082 -899 22402 -898
rect 22082 -1217 22125 -899
rect 22359 -1217 22402 -899
rect 22082 -1218 22402 -1217
rect 22722 -899 23042 -898
rect 22722 -1217 22765 -899
rect 22999 -1217 23042 -899
rect 22722 -1218 23042 -1217
rect 23362 -899 23682 -898
rect 23362 -1217 23405 -899
rect 23639 -1217 23682 -899
rect 23362 -1218 23682 -1217
rect 24002 -899 24322 -898
rect 24002 -1217 24045 -899
rect 24279 -1217 24322 -899
rect 24002 -1218 24322 -1217
rect 24642 -899 24962 -898
rect 24642 -1217 24685 -899
rect 24919 -1217 24962 -899
rect 24642 -1218 24962 -1217
rect -1485 -1474 -1479 -1285
rect -1282 -1474 -1276 -1285
rect -1485 -1478 -1276 -1474
rect -1211 -1538 25922 -1218
rect 2 -1539 322 -1538
rect 2 -1773 45 -1539
rect 279 -1773 322 -1539
rect 2 -1798 322 -1773
rect 642 -1539 962 -1538
rect 642 -1773 685 -1539
rect 919 -1773 962 -1539
rect 642 -1798 962 -1773
rect 1282 -1539 1602 -1538
rect 1282 -1773 1325 -1539
rect 1559 -1773 1602 -1539
rect 1282 -1798 1602 -1773
rect 1922 -1539 2242 -1538
rect 1922 -1773 1965 -1539
rect 2199 -1773 2242 -1539
rect 1922 -1798 2242 -1773
rect 2562 -1539 2882 -1538
rect 2562 -1773 2605 -1539
rect 2839 -1773 2882 -1539
rect 2562 -1798 2882 -1773
rect 3202 -1539 3522 -1538
rect 3202 -1773 3245 -1539
rect 3479 -1773 3522 -1539
rect 3202 -1798 3522 -1773
rect 3842 -1539 4162 -1538
rect 3842 -1773 3885 -1539
rect 4119 -1773 4162 -1539
rect 3842 -1798 4162 -1773
rect 4482 -1539 4802 -1538
rect 4482 -1773 4525 -1539
rect 4759 -1773 4802 -1539
rect 4482 -1798 4802 -1773
rect 5122 -1539 5442 -1538
rect 5122 -1773 5165 -1539
rect 5399 -1773 5442 -1539
rect 5122 -1798 5442 -1773
rect 5762 -1539 6082 -1538
rect 5762 -1773 5805 -1539
rect 6039 -1773 6082 -1539
rect 5762 -1798 6082 -1773
rect 6402 -1539 6722 -1538
rect 6402 -1773 6445 -1539
rect 6679 -1773 6722 -1539
rect 6402 -1798 6722 -1773
rect 7042 -1539 7362 -1538
rect 7042 -1773 7085 -1539
rect 7319 -1773 7362 -1539
rect 7042 -1798 7362 -1773
rect 7682 -1539 8002 -1538
rect 7682 -1773 7725 -1539
rect 7959 -1773 8002 -1539
rect 7682 -1798 8002 -1773
rect 8322 -1539 8642 -1538
rect 8322 -1773 8365 -1539
rect 8599 -1773 8642 -1539
rect 8322 -1798 8642 -1773
rect 8962 -1539 9282 -1538
rect 8962 -1773 9005 -1539
rect 9239 -1773 9282 -1539
rect 8962 -1798 9282 -1773
rect 9602 -1539 9922 -1538
rect 9602 -1773 9645 -1539
rect 9879 -1773 9922 -1539
rect 9602 -1798 9922 -1773
rect 10242 -1539 10562 -1538
rect 10242 -1773 10285 -1539
rect 10519 -1773 10562 -1539
rect 10242 -1798 10562 -1773
rect 10882 -1539 11202 -1538
rect 10882 -1773 10925 -1539
rect 11159 -1773 11202 -1539
rect 10882 -1798 11202 -1773
rect 11522 -1539 11842 -1538
rect 11522 -1773 11565 -1539
rect 11799 -1773 11842 -1539
rect 11522 -1798 11842 -1773
rect 12162 -1539 12482 -1538
rect 12162 -1773 12205 -1539
rect 12439 -1773 12482 -1539
rect 12162 -1798 12482 -1773
rect 12802 -1539 13122 -1538
rect 12802 -1773 12845 -1539
rect 13079 -1773 13122 -1539
rect 12802 -1798 13122 -1773
rect 13442 -1539 13762 -1538
rect 13442 -1773 13485 -1539
rect 13719 -1773 13762 -1539
rect 13442 -1798 13762 -1773
rect 14082 -1539 14402 -1538
rect 14082 -1773 14125 -1539
rect 14359 -1773 14402 -1539
rect 14082 -1798 14402 -1773
rect 14722 -1539 15042 -1538
rect 14722 -1773 14765 -1539
rect 14999 -1773 15042 -1539
rect 14722 -1798 15042 -1773
rect 15362 -1539 15682 -1538
rect 15362 -1773 15405 -1539
rect 15639 -1773 15682 -1539
rect 15362 -1798 15682 -1773
rect 16002 -1539 16322 -1538
rect 16002 -1773 16045 -1539
rect 16279 -1773 16322 -1539
rect 16002 -1798 16322 -1773
rect 16642 -1539 16962 -1538
rect 16642 -1773 16685 -1539
rect 16919 -1773 16962 -1539
rect 16642 -1798 16962 -1773
rect 17282 -1539 17602 -1538
rect 17282 -1773 17325 -1539
rect 17559 -1773 17602 -1539
rect 17282 -1798 17602 -1773
rect 17922 -1539 18242 -1538
rect 17922 -1773 17965 -1539
rect 18199 -1773 18242 -1539
rect 17922 -1798 18242 -1773
rect 18562 -1539 18882 -1538
rect 18562 -1773 18605 -1539
rect 18839 -1773 18882 -1539
rect 18562 -1798 18882 -1773
rect 19202 -1539 19522 -1538
rect 19202 -1773 19245 -1539
rect 19479 -1773 19522 -1539
rect 19202 -1798 19522 -1773
rect 19842 -1539 20162 -1538
rect 19842 -1773 19885 -1539
rect 20119 -1773 20162 -1539
rect 19842 -1798 20162 -1773
rect 20482 -1539 20802 -1538
rect 20482 -1773 20525 -1539
rect 20759 -1773 20802 -1539
rect 20482 -1798 20802 -1773
rect 21122 -1539 21442 -1538
rect 21122 -1773 21165 -1539
rect 21399 -1773 21442 -1539
rect 21122 -1798 21442 -1773
rect 21762 -1539 22082 -1538
rect 21762 -1773 21805 -1539
rect 22039 -1773 22082 -1539
rect 21762 -1798 22082 -1773
rect 22402 -1539 22722 -1538
rect 22402 -1773 22445 -1539
rect 22679 -1773 22722 -1539
rect 22402 -1798 22722 -1773
rect 23042 -1539 23362 -1538
rect 23042 -1773 23085 -1539
rect 23319 -1773 23362 -1539
rect 23042 -1798 23362 -1773
rect 23682 -1539 24002 -1538
rect 23682 -1773 23725 -1539
rect 23959 -1773 24002 -1539
rect 23682 -1798 24002 -1773
rect 24322 -1539 24642 -1538
rect 24322 -1773 24365 -1539
rect 24599 -1773 24642 -1539
rect 24322 -1798 24642 -1773
rect 24962 -1539 25282 -1538
rect 24962 -1773 25005 -1539
rect 25239 -1773 25282 -1539
rect 24962 -1798 25282 -1773
<< via3 >>
rect -1284 28710 -1220 28714
rect -1284 28654 -1280 28710
rect -1280 28654 -1224 28710
rect -1224 28654 -1220 28710
rect -1284 28650 -1220 28654
rect -896 28443 -832 28447
rect -896 28387 -892 28443
rect -892 28387 -836 28443
rect -836 28387 -832 28443
rect -896 28383 -832 28387
rect -1775 27695 -1541 27929
rect -579 27695 -345 27929
rect -1219 27375 -901 27609
rect -1775 27055 -1541 27289
rect -579 27055 -345 27289
rect -1219 26735 -901 26969
rect -1775 26415 -1541 26649
rect -579 26415 -345 26649
rect -1219 26095 -901 26329
rect -1775 25775 -1541 26009
rect -579 25775 -345 26009
rect -1219 25455 -901 25689
rect -1775 25135 -1541 25369
rect -579 25135 -345 25369
rect -1219 24815 -901 25049
rect -1775 24495 -1541 24729
rect -579 24495 -345 24729
rect -1219 24175 -901 24409
rect -1775 23855 -1541 24089
rect -579 23855 -345 24089
rect -1219 23535 -901 23769
rect -1775 23215 -1541 23449
rect -579 23215 -345 23449
rect -1219 22895 -901 23129
rect -1775 22575 -1541 22809
rect -579 22575 -345 22809
rect -1219 22255 -901 22489
rect -1775 21935 -1541 22169
rect -579 21935 -345 22169
rect -1219 21615 -901 21849
rect -1775 21295 -1541 21529
rect -579 21295 -345 21529
rect -1219 20975 -901 21209
rect -1775 20655 -1541 20889
rect -579 20655 -345 20889
rect -1219 20335 -901 20569
rect -1775 20015 -1541 20249
rect -579 20015 -345 20249
rect -1219 19695 -901 19929
rect -1775 19375 -1541 19609
rect -579 19375 -345 19609
rect -1219 19055 -901 19289
rect -1775 18735 -1541 18969
rect -579 18735 -345 18969
rect -1219 18415 -901 18649
rect -1775 18095 -1541 18329
rect -579 18095 -345 18329
rect -1219 17775 -901 18009
rect -1775 17455 -1541 17689
rect -579 17455 -345 17689
rect -1219 17135 -901 17369
rect -1775 16815 -1541 17049
rect -579 16815 -345 17049
rect -1219 16495 -901 16729
rect -1775 16175 -1541 16409
rect -579 16175 -345 16409
rect -1219 15855 -901 16089
rect -1775 15535 -1541 15769
rect -579 15535 -345 15769
rect -1219 15215 -901 15449
rect -1775 14895 -1541 15129
rect -579 14895 -345 15129
rect -1219 14575 -901 14809
rect -1775 14255 -1541 14489
rect -579 14255 -345 14489
rect -1219 13935 -901 14169
rect -1775 13615 -1541 13849
rect -579 13615 -345 13849
rect -1219 13295 -901 13529
rect -1775 12975 -1541 13209
rect -579 12975 -345 13209
rect -1219 12655 -901 12889
rect -1775 12335 -1541 12569
rect -579 12335 -345 12569
rect -1219 12015 -901 12249
rect -1775 11695 -1541 11929
rect -579 11695 -345 11929
rect -1219 11375 -901 11609
rect -1775 11055 -1541 11289
rect -579 11055 -345 11289
rect -1219 10735 -901 10969
rect -1775 10415 -1541 10649
rect -579 10415 -345 10649
rect -1219 10095 -901 10329
rect -1775 9775 -1541 10009
rect -579 9775 -345 10009
rect -1219 9455 -901 9689
rect -1775 9135 -1541 9369
rect -579 9135 -345 9369
rect -1219 8815 -901 9049
rect -1775 8495 -1541 8729
rect -579 8495 -345 8729
rect -1219 8175 -901 8409
rect -1775 7855 -1541 8089
rect -579 7855 -345 8089
rect -1219 7535 -901 7769
rect -1775 7215 -1541 7449
rect -579 7215 -345 7449
rect -1219 6895 -901 7129
rect -1775 6575 -1541 6809
rect -579 6575 -345 6809
rect -1219 6255 -901 6489
rect -1775 5935 -1541 6169
rect -579 5935 -345 6169
rect -1219 5615 -901 5849
rect -1775 5295 -1541 5529
rect -579 5295 -345 5529
rect -1219 4975 -901 5209
rect -1775 4655 -1541 4889
rect -579 4655 -345 4889
rect -1219 4335 -901 4569
rect -1775 4015 -1541 4249
rect -579 4015 -345 4249
rect -1219 3695 -901 3929
rect -1775 3375 -1541 3609
rect -579 3375 -345 3609
rect -1219 3055 -901 3289
rect -1775 2735 -1541 2969
rect -579 2735 -345 2969
rect -1219 2415 -901 2649
rect -1775 2095 -1541 2329
rect -579 2095 -345 2329
rect -1219 1775 -901 2009
rect -1775 1455 -1541 1689
rect -579 1455 -345 1689
rect -1479 112 -1282 301
rect -838 112 -641 301
rect 45 -577 279 -343
rect 685 -577 919 -343
rect 1325 -577 1559 -343
rect 1965 -577 2199 -343
rect 2605 -577 2839 -343
rect 3245 -577 3479 -343
rect 3885 -577 4119 -343
rect 4525 -577 4759 -343
rect 5165 -577 5399 -343
rect 5805 -577 6039 -343
rect 6445 -577 6679 -343
rect 7085 -577 7319 -343
rect 7725 -577 7959 -343
rect 8365 -577 8599 -343
rect 9005 -577 9239 -343
rect 9645 -577 9879 -343
rect 10285 -577 10519 -343
rect 10925 -577 11159 -343
rect 11565 -577 11799 -343
rect 12205 -577 12439 -343
rect 12845 -577 13079 -343
rect 13485 -577 13719 -343
rect 14125 -577 14359 -343
rect 14765 -577 14999 -343
rect 15405 -577 15639 -343
rect 16045 -577 16279 -343
rect 16685 -577 16919 -343
rect 17325 -577 17559 -343
rect 17965 -577 18199 -343
rect 18605 -577 18839 -343
rect 19245 -577 19479 -343
rect 19885 -577 20119 -343
rect 20525 -577 20759 -343
rect 21165 -577 21399 -343
rect 21805 -577 22039 -343
rect 22445 -577 22679 -343
rect 23085 -577 23319 -343
rect 23725 -577 23959 -343
rect 24365 -577 24599 -343
rect 25005 -577 25239 -343
rect -838 -833 -641 -644
rect 365 -1217 599 -899
rect 1005 -1217 1239 -899
rect 1645 -1217 1879 -899
rect 2285 -1217 2519 -899
rect 2925 -1217 3159 -899
rect 3565 -1217 3799 -899
rect 4205 -1217 4439 -899
rect 4845 -1217 5079 -899
rect 5485 -1217 5719 -899
rect 6125 -1217 6359 -899
rect 6765 -1217 6999 -899
rect 7405 -1217 7639 -899
rect 8045 -1217 8279 -899
rect 8685 -1217 8919 -899
rect 9325 -1217 9559 -899
rect 9965 -1217 10199 -899
rect 10605 -1217 10839 -899
rect 11245 -1217 11479 -899
rect 11885 -1217 12119 -899
rect 12525 -1217 12759 -899
rect 13165 -1217 13399 -899
rect 13805 -1217 14039 -899
rect 14445 -1217 14679 -899
rect 15085 -1217 15319 -899
rect 15725 -1217 15959 -899
rect 16365 -1217 16599 -899
rect 17005 -1217 17239 -899
rect 17645 -1217 17879 -899
rect 18285 -1217 18519 -899
rect 18925 -1217 19159 -899
rect 19565 -1217 19799 -899
rect 20205 -1217 20439 -899
rect 20845 -1217 21079 -899
rect 21485 -1217 21719 -899
rect 22125 -1217 22359 -899
rect 22765 -1217 22999 -899
rect 23405 -1217 23639 -899
rect 24045 -1217 24279 -899
rect 24685 -1217 24919 -899
rect -1479 -1474 -1282 -1285
rect 45 -1773 279 -1539
rect 685 -1773 919 -1539
rect 1325 -1773 1559 -1539
rect 1965 -1773 2199 -1539
rect 2605 -1773 2839 -1539
rect 3245 -1773 3479 -1539
rect 3885 -1773 4119 -1539
rect 4525 -1773 4759 -1539
rect 5165 -1773 5399 -1539
rect 5805 -1773 6039 -1539
rect 6445 -1773 6679 -1539
rect 7085 -1773 7319 -1539
rect 7725 -1773 7959 -1539
rect 8365 -1773 8599 -1539
rect 9005 -1773 9239 -1539
rect 9645 -1773 9879 -1539
rect 10285 -1773 10519 -1539
rect 10925 -1773 11159 -1539
rect 11565 -1773 11799 -1539
rect 12205 -1773 12439 -1539
rect 12845 -1773 13079 -1539
rect 13485 -1773 13719 -1539
rect 14125 -1773 14359 -1539
rect 14765 -1773 14999 -1539
rect 15405 -1773 15639 -1539
rect 16045 -1773 16279 -1539
rect 16685 -1773 16919 -1539
rect 17325 -1773 17559 -1539
rect 17965 -1773 18199 -1539
rect 18605 -1773 18839 -1539
rect 19245 -1773 19479 -1539
rect 19885 -1773 20119 -1539
rect 20525 -1773 20759 -1539
rect 21165 -1773 21399 -1539
rect 21805 -1773 22039 -1539
rect 22445 -1773 22679 -1539
rect 23085 -1773 23319 -1539
rect 23725 -1773 23959 -1539
rect 24365 -1773 24599 -1539
rect 25005 -1773 25239 -1539
<< metal4 >>
rect -1480 28714 -1217 28721
rect -1480 28650 -1284 28714
rect -1220 28650 -1217 28714
rect -1480 28648 -1217 28650
rect -1480 301 -1281 28648
rect 51 28500 175 28600
rect 1462 28515 1655 28587
rect 2048 28515 2207 28587
rect 5050 28515 5139 28587
rect 5872 28515 5961 28587
rect 6347 28515 6986 28587
rect -913 28447 -640 28462
rect -913 28383 -896 28447
rect -832 28383 -640 28447
rect -913 28369 -640 28383
rect -1480 112 -1479 301
rect -1282 112 -1281 301
rect -1480 111 -1281 112
rect -839 301 -640 28369
rect 2099 27080 2207 28515
rect 6859 27015 6986 28515
rect 12486 28515 13665 28587
rect 14049 28515 14285 28587
rect 15106 28515 15226 28587
rect 15597 28515 16330 28587
rect 12486 27082 12673 28515
rect 16196 27096 16330 28515
rect 19693 28515 20564 28587
rect 20947 28515 21254 28587
rect 19693 27095 19870 28515
rect 21109 28510 21254 28515
rect 21736 28515 22085 28587
rect 22452 28515 22578 28587
rect 21736 28512 21845 28515
rect 22453 27054 22578 28515
rect 13789 26725 14198 27045
rect 13798 25875 14207 26195
rect 13790 25023 14199 25343
rect 13785 23322 14194 23642
rect 13795 22427 14204 22747
rect 13786 21544 14195 21864
rect 13805 19840 14214 20160
rect 13800 18958 14209 19278
rect 13811 18061 14220 18381
rect 13800 16368 14209 16688
rect 13806 15470 14215 15790
rect 13809 14577 14218 14897
rect 13814 12881 14223 13201
rect 13809 11988 14218 12308
rect 13815 11093 14224 11413
rect 13813 9395 14222 9715
rect 13810 8502 14219 8822
rect 13806 7610 14208 7930
rect 13808 5914 14210 6234
rect 13812 5020 14214 5340
rect 13804 4126 14206 4446
rect 13812 2430 14214 2750
rect 13803 1541 14212 1861
rect 13794 676 14203 996
rect -839 112 -838 301
rect -641 112 -640 301
rect -839 111 -640 112
rect -1540 -644 25922 -638
rect -1540 -833 -838 -644
rect -641 -833 25922 -644
rect -1540 -837 25922 -833
rect -1540 -1285 25922 -1279
rect -1540 -1474 -1479 -1285
rect -1282 -1474 25922 -1285
rect -1540 -1478 25922 -1474
<< via4 >>
rect -1776 27929 -1540 27930
rect -1776 27695 -1775 27929
rect -1775 27695 -1541 27929
rect -1541 27695 -1540 27929
rect -1776 27694 -1540 27695
rect -1776 27289 -1540 27290
rect -1776 27055 -1775 27289
rect -1775 27055 -1541 27289
rect -1541 27055 -1540 27289
rect -1776 27054 -1540 27055
rect -1776 26649 -1540 26650
rect -1776 26415 -1775 26649
rect -1775 26415 -1541 26649
rect -1541 26415 -1540 26649
rect -1776 26414 -1540 26415
rect -1776 26009 -1540 26010
rect -1776 25775 -1775 26009
rect -1775 25775 -1541 26009
rect -1541 25775 -1540 26009
rect -1776 25774 -1540 25775
rect -1776 25369 -1540 25370
rect -1776 25135 -1775 25369
rect -1775 25135 -1541 25369
rect -1541 25135 -1540 25369
rect -1776 25134 -1540 25135
rect -1776 24729 -1540 24730
rect -1776 24495 -1775 24729
rect -1775 24495 -1541 24729
rect -1541 24495 -1540 24729
rect -1776 24494 -1540 24495
rect -1776 24089 -1540 24090
rect -1776 23855 -1775 24089
rect -1775 23855 -1541 24089
rect -1541 23855 -1540 24089
rect -1776 23854 -1540 23855
rect -1776 23449 -1540 23450
rect -1776 23215 -1775 23449
rect -1775 23215 -1541 23449
rect -1541 23215 -1540 23449
rect -1776 23214 -1540 23215
rect -1776 22809 -1540 22810
rect -1776 22575 -1775 22809
rect -1775 22575 -1541 22809
rect -1541 22575 -1540 22809
rect -1776 22574 -1540 22575
rect -1776 22169 -1540 22170
rect -1776 21935 -1775 22169
rect -1775 21935 -1541 22169
rect -1541 21935 -1540 22169
rect -1776 21934 -1540 21935
rect -1776 21529 -1540 21530
rect -1776 21295 -1775 21529
rect -1775 21295 -1541 21529
rect -1541 21295 -1540 21529
rect -1776 21294 -1540 21295
rect -1776 20889 -1540 20890
rect -1776 20655 -1775 20889
rect -1775 20655 -1541 20889
rect -1541 20655 -1540 20889
rect -1776 20654 -1540 20655
rect -1776 20249 -1540 20250
rect -1776 20015 -1775 20249
rect -1775 20015 -1541 20249
rect -1541 20015 -1540 20249
rect -1776 20014 -1540 20015
rect -1776 19609 -1540 19610
rect -1776 19375 -1775 19609
rect -1775 19375 -1541 19609
rect -1541 19375 -1540 19609
rect -1776 19374 -1540 19375
rect -1776 18969 -1540 18970
rect -1776 18735 -1775 18969
rect -1775 18735 -1541 18969
rect -1541 18735 -1540 18969
rect -1776 18734 -1540 18735
rect -1776 18329 -1540 18330
rect -1776 18095 -1775 18329
rect -1775 18095 -1541 18329
rect -1541 18095 -1540 18329
rect -1776 18094 -1540 18095
rect -1776 17689 -1540 17690
rect -1776 17455 -1775 17689
rect -1775 17455 -1541 17689
rect -1541 17455 -1540 17689
rect -1776 17454 -1540 17455
rect -1776 17049 -1540 17050
rect -1776 16815 -1775 17049
rect -1775 16815 -1541 17049
rect -1541 16815 -1540 17049
rect -1776 16814 -1540 16815
rect -1776 16409 -1540 16410
rect -1776 16175 -1775 16409
rect -1775 16175 -1541 16409
rect -1541 16175 -1540 16409
rect -1776 16174 -1540 16175
rect -1776 15769 -1540 15770
rect -1776 15535 -1775 15769
rect -1775 15535 -1541 15769
rect -1541 15535 -1540 15769
rect -1776 15534 -1540 15535
rect -1776 15129 -1540 15130
rect -1776 14895 -1775 15129
rect -1775 14895 -1541 15129
rect -1541 14895 -1540 15129
rect -1776 14894 -1540 14895
rect -1776 14489 -1540 14490
rect -1776 14255 -1775 14489
rect -1775 14255 -1541 14489
rect -1541 14255 -1540 14489
rect -1776 14254 -1540 14255
rect -1776 13849 -1540 13850
rect -1776 13615 -1775 13849
rect -1775 13615 -1541 13849
rect -1541 13615 -1540 13849
rect -1776 13614 -1540 13615
rect -1776 13209 -1540 13210
rect -1776 12975 -1775 13209
rect -1775 12975 -1541 13209
rect -1541 12975 -1540 13209
rect -1776 12974 -1540 12975
rect -1776 12569 -1540 12570
rect -1776 12335 -1775 12569
rect -1775 12335 -1541 12569
rect -1541 12335 -1540 12569
rect -1776 12334 -1540 12335
rect -1776 11929 -1540 11930
rect -1776 11695 -1775 11929
rect -1775 11695 -1541 11929
rect -1541 11695 -1540 11929
rect -1776 11694 -1540 11695
rect -1776 11289 -1540 11290
rect -1776 11055 -1775 11289
rect -1775 11055 -1541 11289
rect -1541 11055 -1540 11289
rect -1776 11054 -1540 11055
rect -1776 10649 -1540 10650
rect -1776 10415 -1775 10649
rect -1775 10415 -1541 10649
rect -1541 10415 -1540 10649
rect -1776 10414 -1540 10415
rect -1776 10009 -1540 10010
rect -1776 9775 -1775 10009
rect -1775 9775 -1541 10009
rect -1541 9775 -1540 10009
rect -1776 9774 -1540 9775
rect -1776 9369 -1540 9370
rect -1776 9135 -1775 9369
rect -1775 9135 -1541 9369
rect -1541 9135 -1540 9369
rect -1776 9134 -1540 9135
rect -1776 8729 -1540 8730
rect -1776 8495 -1775 8729
rect -1775 8495 -1541 8729
rect -1541 8495 -1540 8729
rect -1776 8494 -1540 8495
rect -1776 8089 -1540 8090
rect -1776 7855 -1775 8089
rect -1775 7855 -1541 8089
rect -1541 7855 -1540 8089
rect -1776 7854 -1540 7855
rect -1776 7449 -1540 7450
rect -1776 7215 -1775 7449
rect -1775 7215 -1541 7449
rect -1541 7215 -1540 7449
rect -1776 7214 -1540 7215
rect -1776 6809 -1540 6810
rect -1776 6575 -1775 6809
rect -1775 6575 -1541 6809
rect -1541 6575 -1540 6809
rect -1776 6574 -1540 6575
rect -1776 6169 -1540 6170
rect -1776 5935 -1775 6169
rect -1775 5935 -1541 6169
rect -1541 5935 -1540 6169
rect -1776 5934 -1540 5935
rect -1776 5529 -1540 5530
rect -1776 5295 -1775 5529
rect -1775 5295 -1541 5529
rect -1541 5295 -1540 5529
rect -1776 5294 -1540 5295
rect -1776 4889 -1540 4890
rect -1776 4655 -1775 4889
rect -1775 4655 -1541 4889
rect -1541 4655 -1540 4889
rect -1776 4654 -1540 4655
rect -1776 4249 -1540 4250
rect -1776 4015 -1775 4249
rect -1775 4015 -1541 4249
rect -1541 4015 -1540 4249
rect -1776 4014 -1540 4015
rect -1776 3609 -1540 3610
rect -1776 3375 -1775 3609
rect -1775 3375 -1541 3609
rect -1541 3375 -1540 3609
rect -1776 3374 -1540 3375
rect -1776 2969 -1540 2970
rect -1776 2735 -1775 2969
rect -1775 2735 -1541 2969
rect -1541 2735 -1540 2969
rect -1776 2734 -1540 2735
rect -1776 2329 -1540 2330
rect -1776 2095 -1775 2329
rect -1775 2095 -1541 2329
rect -1541 2095 -1540 2329
rect -1776 2094 -1540 2095
rect -1776 1689 -1540 1690
rect -1776 1455 -1775 1689
rect -1775 1455 -1541 1689
rect -1541 1455 -1540 1689
rect -1776 1454 -1540 1455
rect -1220 27609 -900 27610
rect -1220 27375 -1219 27609
rect -1219 27375 -901 27609
rect -901 27375 -900 27609
rect -1220 27374 -900 27375
rect -1220 26969 -900 26970
rect -1220 26735 -1219 26969
rect -1219 26735 -901 26969
rect -901 26735 -900 26969
rect -1220 26734 -900 26735
rect -1220 26329 -900 26330
rect -1220 26095 -1219 26329
rect -1219 26095 -901 26329
rect -901 26095 -900 26329
rect -1220 26094 -900 26095
rect -1220 25689 -900 25690
rect -1220 25455 -1219 25689
rect -1219 25455 -901 25689
rect -901 25455 -900 25689
rect -1220 25454 -900 25455
rect -1220 25049 -900 25050
rect -1220 24815 -1219 25049
rect -1219 24815 -901 25049
rect -901 24815 -900 25049
rect -1220 24814 -900 24815
rect -1220 24409 -900 24410
rect -1220 24175 -1219 24409
rect -1219 24175 -901 24409
rect -901 24175 -900 24409
rect -1220 24174 -900 24175
rect -1220 23769 -900 23770
rect -1220 23535 -1219 23769
rect -1219 23535 -901 23769
rect -901 23535 -900 23769
rect -1220 23534 -900 23535
rect -1220 23129 -900 23130
rect -1220 22895 -1219 23129
rect -1219 22895 -901 23129
rect -901 22895 -900 23129
rect -1220 22894 -900 22895
rect -1220 22489 -900 22490
rect -1220 22255 -1219 22489
rect -1219 22255 -901 22489
rect -901 22255 -900 22489
rect -1220 22254 -900 22255
rect -1220 21849 -900 21850
rect -1220 21615 -1219 21849
rect -1219 21615 -901 21849
rect -901 21615 -900 21849
rect -1220 21614 -900 21615
rect -1220 21209 -900 21210
rect -1220 20975 -1219 21209
rect -1219 20975 -901 21209
rect -901 20975 -900 21209
rect -1220 20974 -900 20975
rect -1220 20569 -900 20570
rect -1220 20335 -1219 20569
rect -1219 20335 -901 20569
rect -901 20335 -900 20569
rect -1220 20334 -900 20335
rect -1220 19929 -900 19930
rect -1220 19695 -1219 19929
rect -1219 19695 -901 19929
rect -901 19695 -900 19929
rect -1220 19694 -900 19695
rect -1220 19289 -900 19290
rect -1220 19055 -1219 19289
rect -1219 19055 -901 19289
rect -901 19055 -900 19289
rect -1220 19054 -900 19055
rect -1220 18649 -900 18650
rect -1220 18415 -1219 18649
rect -1219 18415 -901 18649
rect -901 18415 -900 18649
rect -1220 18414 -900 18415
rect -1220 18009 -900 18010
rect -1220 17775 -1219 18009
rect -1219 17775 -901 18009
rect -901 17775 -900 18009
rect -1220 17774 -900 17775
rect -1220 17369 -900 17370
rect -1220 17135 -1219 17369
rect -1219 17135 -901 17369
rect -901 17135 -900 17369
rect -1220 17134 -900 17135
rect -1220 16729 -900 16730
rect -1220 16495 -1219 16729
rect -1219 16495 -901 16729
rect -901 16495 -900 16729
rect -1220 16494 -900 16495
rect -1220 16089 -900 16090
rect -1220 15855 -1219 16089
rect -1219 15855 -901 16089
rect -901 15855 -900 16089
rect -1220 15854 -900 15855
rect -1220 15449 -900 15450
rect -1220 15215 -1219 15449
rect -1219 15215 -901 15449
rect -901 15215 -900 15449
rect -1220 15214 -900 15215
rect -1220 14809 -900 14810
rect -1220 14575 -1219 14809
rect -1219 14575 -901 14809
rect -901 14575 -900 14809
rect -1220 14574 -900 14575
rect -1220 14169 -900 14170
rect -1220 13935 -1219 14169
rect -1219 13935 -901 14169
rect -901 13935 -900 14169
rect -1220 13934 -900 13935
rect -1220 13529 -900 13530
rect -1220 13295 -1219 13529
rect -1219 13295 -901 13529
rect -901 13295 -900 13529
rect -1220 13294 -900 13295
rect -1220 12889 -900 12890
rect -1220 12655 -1219 12889
rect -1219 12655 -901 12889
rect -901 12655 -900 12889
rect -1220 12654 -900 12655
rect -1220 12249 -900 12250
rect -1220 12015 -1219 12249
rect -1219 12015 -901 12249
rect -901 12015 -900 12249
rect -1220 12014 -900 12015
rect -1220 11609 -900 11610
rect -1220 11375 -1219 11609
rect -1219 11375 -901 11609
rect -901 11375 -900 11609
rect -1220 11374 -900 11375
rect -1220 10969 -900 10970
rect -1220 10735 -1219 10969
rect -1219 10735 -901 10969
rect -901 10735 -900 10969
rect -1220 10734 -900 10735
rect -1220 10329 -900 10330
rect -1220 10095 -1219 10329
rect -1219 10095 -901 10329
rect -901 10095 -900 10329
rect -1220 10094 -900 10095
rect -1220 9689 -900 9690
rect -1220 9455 -1219 9689
rect -1219 9455 -901 9689
rect -901 9455 -900 9689
rect -1220 9454 -900 9455
rect -1220 9049 -900 9050
rect -1220 8815 -1219 9049
rect -1219 8815 -901 9049
rect -901 8815 -900 9049
rect -1220 8814 -900 8815
rect -1220 8409 -900 8410
rect -1220 8175 -1219 8409
rect -1219 8175 -901 8409
rect -901 8175 -900 8409
rect -1220 8174 -900 8175
rect -1220 7769 -900 7770
rect -1220 7535 -1219 7769
rect -1219 7535 -901 7769
rect -901 7535 -900 7769
rect -1220 7534 -900 7535
rect -1220 7129 -900 7130
rect -1220 6895 -1219 7129
rect -1219 6895 -901 7129
rect -901 6895 -900 7129
rect -1220 6894 -900 6895
rect -1220 6489 -900 6490
rect -1220 6255 -1219 6489
rect -1219 6255 -901 6489
rect -901 6255 -900 6489
rect -1220 6254 -900 6255
rect -1220 5849 -900 5850
rect -1220 5615 -1219 5849
rect -1219 5615 -901 5849
rect -901 5615 -900 5849
rect -1220 5614 -900 5615
rect -1220 5209 -900 5210
rect -1220 4975 -1219 5209
rect -1219 4975 -901 5209
rect -901 4975 -900 5209
rect -1220 4974 -900 4975
rect -1220 4569 -900 4570
rect -1220 4335 -1219 4569
rect -1219 4335 -901 4569
rect -901 4335 -900 4569
rect -1220 4334 -900 4335
rect -1220 3929 -900 3930
rect -1220 3695 -1219 3929
rect -1219 3695 -901 3929
rect -901 3695 -900 3929
rect -1220 3694 -900 3695
rect -1220 3289 -900 3290
rect -1220 3055 -1219 3289
rect -1219 3055 -901 3289
rect -901 3055 -900 3289
rect -1220 3054 -900 3055
rect -1220 2649 -900 2650
rect -1220 2415 -1219 2649
rect -1219 2415 -901 2649
rect -901 2415 -900 2649
rect -1220 2414 -900 2415
rect -1220 2009 -900 2010
rect -1220 1775 -1219 2009
rect -1219 1775 -901 2009
rect -901 1775 -900 2009
rect -1220 1774 -900 1775
rect -580 27929 -344 27930
rect -580 27695 -579 27929
rect -579 27695 -345 27929
rect -345 27695 -344 27929
rect -580 27694 -344 27695
rect -580 27289 -344 27290
rect -580 27055 -579 27289
rect -579 27055 -345 27289
rect -345 27055 -344 27289
rect -580 27054 -344 27055
rect -580 26649 -344 26650
rect -580 26415 -579 26649
rect -579 26415 -345 26649
rect -345 26415 -344 26649
rect -580 26414 -344 26415
rect -580 26009 -344 26010
rect -580 25775 -579 26009
rect -579 25775 -345 26009
rect -345 25775 -344 26009
rect -580 25774 -344 25775
rect -580 25369 -344 25370
rect -580 25135 -579 25369
rect -579 25135 -345 25369
rect -345 25135 -344 25369
rect -580 25134 -344 25135
rect -580 24729 -344 24730
rect -580 24495 -579 24729
rect -579 24495 -345 24729
rect -345 24495 -344 24729
rect -580 24494 -344 24495
rect -580 24089 -344 24090
rect -580 23855 -579 24089
rect -579 23855 -345 24089
rect -345 23855 -344 24089
rect -580 23854 -344 23855
rect -580 23449 -344 23450
rect -580 23215 -579 23449
rect -579 23215 -345 23449
rect -345 23215 -344 23449
rect -580 23214 -344 23215
rect -580 22809 -344 22810
rect -580 22575 -579 22809
rect -579 22575 -345 22809
rect -345 22575 -344 22809
rect -580 22574 -344 22575
rect -580 22169 -344 22170
rect -580 21935 -579 22169
rect -579 21935 -345 22169
rect -345 21935 -344 22169
rect -580 21934 -344 21935
rect -580 21529 -344 21530
rect -580 21295 -579 21529
rect -579 21295 -345 21529
rect -345 21295 -344 21529
rect -580 21294 -344 21295
rect -580 20889 -344 20890
rect -580 20655 -579 20889
rect -579 20655 -345 20889
rect -345 20655 -344 20889
rect -580 20654 -344 20655
rect -580 20249 -344 20250
rect -580 20015 -579 20249
rect -579 20015 -345 20249
rect -345 20015 -344 20249
rect -580 20014 -344 20015
rect -580 19609 -344 19610
rect -580 19375 -579 19609
rect -579 19375 -345 19609
rect -345 19375 -344 19609
rect -580 19374 -344 19375
rect -580 18969 -344 18970
rect -580 18735 -579 18969
rect -579 18735 -345 18969
rect -345 18735 -344 18969
rect -580 18734 -344 18735
rect -580 18329 -344 18330
rect -580 18095 -579 18329
rect -579 18095 -345 18329
rect -345 18095 -344 18329
rect -580 18094 -344 18095
rect -580 17689 -344 17690
rect -580 17455 -579 17689
rect -579 17455 -345 17689
rect -345 17455 -344 17689
rect -580 17454 -344 17455
rect -580 17049 -344 17050
rect -580 16815 -579 17049
rect -579 16815 -345 17049
rect -345 16815 -344 17049
rect -580 16814 -344 16815
rect -580 16409 -344 16410
rect -580 16175 -579 16409
rect -579 16175 -345 16409
rect -345 16175 -344 16409
rect -580 16174 -344 16175
rect -580 15769 -344 15770
rect -580 15535 -579 15769
rect -579 15535 -345 15769
rect -345 15535 -344 15769
rect -580 15534 -344 15535
rect -580 15129 -344 15130
rect -580 14895 -579 15129
rect -579 14895 -345 15129
rect -345 14895 -344 15129
rect -580 14894 -344 14895
rect -580 14489 -344 14490
rect -580 14255 -579 14489
rect -579 14255 -345 14489
rect -345 14255 -344 14489
rect -580 14254 -344 14255
rect -580 13849 -344 13850
rect -580 13615 -579 13849
rect -579 13615 -345 13849
rect -345 13615 -344 13849
rect -580 13614 -344 13615
rect -580 13209 -344 13210
rect -580 12975 -579 13209
rect -579 12975 -345 13209
rect -345 12975 -344 13209
rect -580 12974 -344 12975
rect -580 12569 -344 12570
rect -580 12335 -579 12569
rect -579 12335 -345 12569
rect -345 12335 -344 12569
rect -580 12334 -344 12335
rect -580 11929 -344 11930
rect -580 11695 -579 11929
rect -579 11695 -345 11929
rect -345 11695 -344 11929
rect -580 11694 -344 11695
rect -580 11289 -344 11290
rect -580 11055 -579 11289
rect -579 11055 -345 11289
rect -345 11055 -344 11289
rect -580 11054 -344 11055
rect -580 10649 -344 10650
rect -580 10415 -579 10649
rect -579 10415 -345 10649
rect -345 10415 -344 10649
rect -580 10414 -344 10415
rect -580 10009 -344 10010
rect -580 9775 -579 10009
rect -579 9775 -345 10009
rect -345 9775 -344 10009
rect -580 9774 -344 9775
rect -580 9369 -344 9370
rect -580 9135 -579 9369
rect -579 9135 -345 9369
rect -345 9135 -344 9369
rect -580 9134 -344 9135
rect -580 8729 -344 8730
rect -580 8495 -579 8729
rect -579 8495 -345 8729
rect -345 8495 -344 8729
rect -580 8494 -344 8495
rect -580 8089 -344 8090
rect -580 7855 -579 8089
rect -579 7855 -345 8089
rect -345 7855 -344 8089
rect -580 7854 -344 7855
rect -580 7449 -344 7450
rect -580 7215 -579 7449
rect -579 7215 -345 7449
rect -345 7215 -344 7449
rect -580 7214 -344 7215
rect -580 6809 -344 6810
rect -580 6575 -579 6809
rect -579 6575 -345 6809
rect -345 6575 -344 6809
rect -580 6574 -344 6575
rect -580 6169 -344 6170
rect -580 5935 -579 6169
rect -579 5935 -345 6169
rect -345 5935 -344 6169
rect -580 5934 -344 5935
rect -580 5529 -344 5530
rect -580 5295 -579 5529
rect -579 5295 -345 5529
rect -345 5295 -344 5529
rect -580 5294 -344 5295
rect -580 4889 -344 4890
rect -580 4655 -579 4889
rect -579 4655 -345 4889
rect -345 4655 -344 4889
rect -580 4654 -344 4655
rect -580 4249 -344 4250
rect -580 4015 -579 4249
rect -579 4015 -345 4249
rect -345 4015 -344 4249
rect -580 4014 -344 4015
rect -580 3609 -344 3610
rect -580 3375 -579 3609
rect -579 3375 -345 3609
rect -345 3375 -344 3609
rect -580 3374 -344 3375
rect -580 2969 -344 2970
rect -580 2735 -579 2969
rect -579 2735 -345 2969
rect -345 2735 -344 2969
rect -580 2734 -344 2735
rect -580 2329 -344 2330
rect -580 2095 -579 2329
rect -579 2095 -345 2329
rect -345 2095 -344 2329
rect -580 2094 -344 2095
rect -580 1689 -344 1690
rect -580 1455 -579 1689
rect -579 1455 -345 1689
rect -345 1455 -344 1689
rect -580 1454 -344 1455
rect 44 -343 280 -342
rect 44 -577 45 -343
rect 45 -577 279 -343
rect 279 -577 280 -343
rect 44 -578 280 -577
rect 684 -343 920 -342
rect 684 -577 685 -343
rect 685 -577 919 -343
rect 919 -577 920 -343
rect 684 -578 920 -577
rect 1324 -343 1560 -342
rect 1324 -577 1325 -343
rect 1325 -577 1559 -343
rect 1559 -577 1560 -343
rect 1324 -578 1560 -577
rect 1964 -343 2200 -342
rect 1964 -577 1965 -343
rect 1965 -577 2199 -343
rect 2199 -577 2200 -343
rect 1964 -578 2200 -577
rect 2604 -343 2840 -342
rect 2604 -577 2605 -343
rect 2605 -577 2839 -343
rect 2839 -577 2840 -343
rect 2604 -578 2840 -577
rect 3244 -343 3480 -342
rect 3244 -577 3245 -343
rect 3245 -577 3479 -343
rect 3479 -577 3480 -343
rect 3244 -578 3480 -577
rect 3884 -343 4120 -342
rect 3884 -577 3885 -343
rect 3885 -577 4119 -343
rect 4119 -577 4120 -343
rect 3884 -578 4120 -577
rect 4524 -343 4760 -342
rect 4524 -577 4525 -343
rect 4525 -577 4759 -343
rect 4759 -577 4760 -343
rect 4524 -578 4760 -577
rect 5164 -343 5400 -342
rect 5164 -577 5165 -343
rect 5165 -577 5399 -343
rect 5399 -577 5400 -343
rect 5164 -578 5400 -577
rect 5804 -343 6040 -342
rect 5804 -577 5805 -343
rect 5805 -577 6039 -343
rect 6039 -577 6040 -343
rect 5804 -578 6040 -577
rect 6444 -343 6680 -342
rect 6444 -577 6445 -343
rect 6445 -577 6679 -343
rect 6679 -577 6680 -343
rect 6444 -578 6680 -577
rect 7084 -343 7320 -342
rect 7084 -577 7085 -343
rect 7085 -577 7319 -343
rect 7319 -577 7320 -343
rect 7084 -578 7320 -577
rect 7724 -343 7960 -342
rect 7724 -577 7725 -343
rect 7725 -577 7959 -343
rect 7959 -577 7960 -343
rect 7724 -578 7960 -577
rect 8364 -343 8600 -342
rect 8364 -577 8365 -343
rect 8365 -577 8599 -343
rect 8599 -577 8600 -343
rect 8364 -578 8600 -577
rect 9004 -343 9240 -342
rect 9004 -577 9005 -343
rect 9005 -577 9239 -343
rect 9239 -577 9240 -343
rect 9004 -578 9240 -577
rect 9644 -343 9880 -342
rect 9644 -577 9645 -343
rect 9645 -577 9879 -343
rect 9879 -577 9880 -343
rect 9644 -578 9880 -577
rect 10284 -343 10520 -342
rect 10284 -577 10285 -343
rect 10285 -577 10519 -343
rect 10519 -577 10520 -343
rect 10284 -578 10520 -577
rect 10924 -343 11160 -342
rect 10924 -577 10925 -343
rect 10925 -577 11159 -343
rect 11159 -577 11160 -343
rect 10924 -578 11160 -577
rect 11564 -343 11800 -342
rect 11564 -577 11565 -343
rect 11565 -577 11799 -343
rect 11799 -577 11800 -343
rect 11564 -578 11800 -577
rect 12204 -343 12440 -342
rect 12204 -577 12205 -343
rect 12205 -577 12439 -343
rect 12439 -577 12440 -343
rect 12204 -578 12440 -577
rect 12844 -343 13080 -342
rect 12844 -577 12845 -343
rect 12845 -577 13079 -343
rect 13079 -577 13080 -343
rect 12844 -578 13080 -577
rect 13484 -343 13720 -342
rect 13484 -577 13485 -343
rect 13485 -577 13719 -343
rect 13719 -577 13720 -343
rect 13484 -578 13720 -577
rect 14124 -343 14360 -342
rect 14124 -577 14125 -343
rect 14125 -577 14359 -343
rect 14359 -577 14360 -343
rect 14124 -578 14360 -577
rect 14764 -343 15000 -342
rect 14764 -577 14765 -343
rect 14765 -577 14999 -343
rect 14999 -577 15000 -343
rect 14764 -578 15000 -577
rect 15404 -343 15640 -342
rect 15404 -577 15405 -343
rect 15405 -577 15639 -343
rect 15639 -577 15640 -343
rect 15404 -578 15640 -577
rect 16044 -343 16280 -342
rect 16044 -577 16045 -343
rect 16045 -577 16279 -343
rect 16279 -577 16280 -343
rect 16044 -578 16280 -577
rect 16684 -343 16920 -342
rect 16684 -577 16685 -343
rect 16685 -577 16919 -343
rect 16919 -577 16920 -343
rect 16684 -578 16920 -577
rect 17324 -343 17560 -342
rect 17324 -577 17325 -343
rect 17325 -577 17559 -343
rect 17559 -577 17560 -343
rect 17324 -578 17560 -577
rect 17964 -343 18200 -342
rect 17964 -577 17965 -343
rect 17965 -577 18199 -343
rect 18199 -577 18200 -343
rect 17964 -578 18200 -577
rect 18604 -343 18840 -342
rect 18604 -577 18605 -343
rect 18605 -577 18839 -343
rect 18839 -577 18840 -343
rect 18604 -578 18840 -577
rect 19244 -343 19480 -342
rect 19244 -577 19245 -343
rect 19245 -577 19479 -343
rect 19479 -577 19480 -343
rect 19244 -578 19480 -577
rect 19884 -343 20120 -342
rect 19884 -577 19885 -343
rect 19885 -577 20119 -343
rect 20119 -577 20120 -343
rect 19884 -578 20120 -577
rect 20524 -343 20760 -342
rect 20524 -577 20525 -343
rect 20525 -577 20759 -343
rect 20759 -577 20760 -343
rect 20524 -578 20760 -577
rect 21164 -343 21400 -342
rect 21164 -577 21165 -343
rect 21165 -577 21399 -343
rect 21399 -577 21400 -343
rect 21164 -578 21400 -577
rect 21804 -343 22040 -342
rect 21804 -577 21805 -343
rect 21805 -577 22039 -343
rect 22039 -577 22040 -343
rect 21804 -578 22040 -577
rect 22444 -343 22680 -342
rect 22444 -577 22445 -343
rect 22445 -577 22679 -343
rect 22679 -577 22680 -343
rect 22444 -578 22680 -577
rect 23084 -343 23320 -342
rect 23084 -577 23085 -343
rect 23085 -577 23319 -343
rect 23319 -577 23320 -343
rect 23084 -578 23320 -577
rect 23724 -343 23960 -342
rect 23724 -577 23725 -343
rect 23725 -577 23959 -343
rect 23959 -577 23960 -343
rect 23724 -578 23960 -577
rect 24364 -343 24600 -342
rect 24364 -577 24365 -343
rect 24365 -577 24599 -343
rect 24599 -577 24600 -343
rect 24364 -578 24600 -577
rect 25004 -343 25240 -342
rect 25004 -577 25005 -343
rect 25005 -577 25239 -343
rect 25239 -577 25240 -343
rect 25004 -578 25240 -577
rect 364 -899 600 -898
rect 364 -1217 365 -899
rect 365 -1217 599 -899
rect 599 -1217 600 -899
rect 364 -1218 600 -1217
rect 1004 -899 1240 -898
rect 1004 -1217 1005 -899
rect 1005 -1217 1239 -899
rect 1239 -1217 1240 -899
rect 1004 -1218 1240 -1217
rect 1644 -899 1880 -898
rect 1644 -1217 1645 -899
rect 1645 -1217 1879 -899
rect 1879 -1217 1880 -899
rect 1644 -1218 1880 -1217
rect 2284 -899 2520 -898
rect 2284 -1217 2285 -899
rect 2285 -1217 2519 -899
rect 2519 -1217 2520 -899
rect 2284 -1218 2520 -1217
rect 2924 -899 3160 -898
rect 2924 -1217 2925 -899
rect 2925 -1217 3159 -899
rect 3159 -1217 3160 -899
rect 2924 -1218 3160 -1217
rect 3564 -899 3800 -898
rect 3564 -1217 3565 -899
rect 3565 -1217 3799 -899
rect 3799 -1217 3800 -899
rect 3564 -1218 3800 -1217
rect 4204 -899 4440 -898
rect 4204 -1217 4205 -899
rect 4205 -1217 4439 -899
rect 4439 -1217 4440 -899
rect 4204 -1218 4440 -1217
rect 4844 -899 5080 -898
rect 4844 -1217 4845 -899
rect 4845 -1217 5079 -899
rect 5079 -1217 5080 -899
rect 4844 -1218 5080 -1217
rect 5484 -899 5720 -898
rect 5484 -1217 5485 -899
rect 5485 -1217 5719 -899
rect 5719 -1217 5720 -899
rect 5484 -1218 5720 -1217
rect 6124 -899 6360 -898
rect 6124 -1217 6125 -899
rect 6125 -1217 6359 -899
rect 6359 -1217 6360 -899
rect 6124 -1218 6360 -1217
rect 6764 -899 7000 -898
rect 6764 -1217 6765 -899
rect 6765 -1217 6999 -899
rect 6999 -1217 7000 -899
rect 6764 -1218 7000 -1217
rect 7404 -899 7640 -898
rect 7404 -1217 7405 -899
rect 7405 -1217 7639 -899
rect 7639 -1217 7640 -899
rect 7404 -1218 7640 -1217
rect 8044 -899 8280 -898
rect 8044 -1217 8045 -899
rect 8045 -1217 8279 -899
rect 8279 -1217 8280 -899
rect 8044 -1218 8280 -1217
rect 8684 -899 8920 -898
rect 8684 -1217 8685 -899
rect 8685 -1217 8919 -899
rect 8919 -1217 8920 -899
rect 8684 -1218 8920 -1217
rect 9324 -899 9560 -898
rect 9324 -1217 9325 -899
rect 9325 -1217 9559 -899
rect 9559 -1217 9560 -899
rect 9324 -1218 9560 -1217
rect 9964 -899 10200 -898
rect 9964 -1217 9965 -899
rect 9965 -1217 10199 -899
rect 10199 -1217 10200 -899
rect 9964 -1218 10200 -1217
rect 10604 -899 10840 -898
rect 10604 -1217 10605 -899
rect 10605 -1217 10839 -899
rect 10839 -1217 10840 -899
rect 10604 -1218 10840 -1217
rect 11244 -899 11480 -898
rect 11244 -1217 11245 -899
rect 11245 -1217 11479 -899
rect 11479 -1217 11480 -899
rect 11244 -1218 11480 -1217
rect 11884 -899 12120 -898
rect 11884 -1217 11885 -899
rect 11885 -1217 12119 -899
rect 12119 -1217 12120 -899
rect 11884 -1218 12120 -1217
rect 12524 -899 12760 -898
rect 12524 -1217 12525 -899
rect 12525 -1217 12759 -899
rect 12759 -1217 12760 -899
rect 12524 -1218 12760 -1217
rect 13164 -899 13400 -898
rect 13164 -1217 13165 -899
rect 13165 -1217 13399 -899
rect 13399 -1217 13400 -899
rect 13164 -1218 13400 -1217
rect 13804 -899 14040 -898
rect 13804 -1217 13805 -899
rect 13805 -1217 14039 -899
rect 14039 -1217 14040 -899
rect 13804 -1218 14040 -1217
rect 14444 -899 14680 -898
rect 14444 -1217 14445 -899
rect 14445 -1217 14679 -899
rect 14679 -1217 14680 -899
rect 14444 -1218 14680 -1217
rect 15084 -899 15320 -898
rect 15084 -1217 15085 -899
rect 15085 -1217 15319 -899
rect 15319 -1217 15320 -899
rect 15084 -1218 15320 -1217
rect 15724 -899 15960 -898
rect 15724 -1217 15725 -899
rect 15725 -1217 15959 -899
rect 15959 -1217 15960 -899
rect 15724 -1218 15960 -1217
rect 16364 -899 16600 -898
rect 16364 -1217 16365 -899
rect 16365 -1217 16599 -899
rect 16599 -1217 16600 -899
rect 16364 -1218 16600 -1217
rect 17004 -899 17240 -898
rect 17004 -1217 17005 -899
rect 17005 -1217 17239 -899
rect 17239 -1217 17240 -899
rect 17004 -1218 17240 -1217
rect 17644 -899 17880 -898
rect 17644 -1217 17645 -899
rect 17645 -1217 17879 -899
rect 17879 -1217 17880 -899
rect 17644 -1218 17880 -1217
rect 18284 -899 18520 -898
rect 18284 -1217 18285 -899
rect 18285 -1217 18519 -899
rect 18519 -1217 18520 -899
rect 18284 -1218 18520 -1217
rect 18924 -899 19160 -898
rect 18924 -1217 18925 -899
rect 18925 -1217 19159 -899
rect 19159 -1217 19160 -899
rect 18924 -1218 19160 -1217
rect 19564 -899 19800 -898
rect 19564 -1217 19565 -899
rect 19565 -1217 19799 -899
rect 19799 -1217 19800 -899
rect 19564 -1218 19800 -1217
rect 20204 -899 20440 -898
rect 20204 -1217 20205 -899
rect 20205 -1217 20439 -899
rect 20439 -1217 20440 -899
rect 20204 -1218 20440 -1217
rect 20844 -899 21080 -898
rect 20844 -1217 20845 -899
rect 20845 -1217 21079 -899
rect 21079 -1217 21080 -899
rect 20844 -1218 21080 -1217
rect 21484 -899 21720 -898
rect 21484 -1217 21485 -899
rect 21485 -1217 21719 -899
rect 21719 -1217 21720 -899
rect 21484 -1218 21720 -1217
rect 22124 -899 22360 -898
rect 22124 -1217 22125 -899
rect 22125 -1217 22359 -899
rect 22359 -1217 22360 -899
rect 22124 -1218 22360 -1217
rect 22764 -899 23000 -898
rect 22764 -1217 22765 -899
rect 22765 -1217 22999 -899
rect 22999 -1217 23000 -899
rect 22764 -1218 23000 -1217
rect 23404 -899 23640 -898
rect 23404 -1217 23405 -899
rect 23405 -1217 23639 -899
rect 23639 -1217 23640 -899
rect 23404 -1218 23640 -1217
rect 24044 -899 24280 -898
rect 24044 -1217 24045 -899
rect 24045 -1217 24279 -899
rect 24279 -1217 24280 -899
rect 24044 -1218 24280 -1217
rect 24684 -899 24920 -898
rect 24684 -1217 24685 -899
rect 24685 -1217 24919 -899
rect 24919 -1217 24920 -899
rect 24684 -1218 24920 -1217
rect 44 -1539 280 -1538
rect 44 -1773 45 -1539
rect 45 -1773 279 -1539
rect 279 -1773 280 -1539
rect 44 -1774 280 -1773
rect 684 -1539 920 -1538
rect 684 -1773 685 -1539
rect 685 -1773 919 -1539
rect 919 -1773 920 -1539
rect 684 -1774 920 -1773
rect 1324 -1539 1560 -1538
rect 1324 -1773 1325 -1539
rect 1325 -1773 1559 -1539
rect 1559 -1773 1560 -1539
rect 1324 -1774 1560 -1773
rect 1964 -1539 2200 -1538
rect 1964 -1773 1965 -1539
rect 1965 -1773 2199 -1539
rect 2199 -1773 2200 -1539
rect 1964 -1774 2200 -1773
rect 2604 -1539 2840 -1538
rect 2604 -1773 2605 -1539
rect 2605 -1773 2839 -1539
rect 2839 -1773 2840 -1539
rect 2604 -1774 2840 -1773
rect 3244 -1539 3480 -1538
rect 3244 -1773 3245 -1539
rect 3245 -1773 3479 -1539
rect 3479 -1773 3480 -1539
rect 3244 -1774 3480 -1773
rect 3884 -1539 4120 -1538
rect 3884 -1773 3885 -1539
rect 3885 -1773 4119 -1539
rect 4119 -1773 4120 -1539
rect 3884 -1774 4120 -1773
rect 4524 -1539 4760 -1538
rect 4524 -1773 4525 -1539
rect 4525 -1773 4759 -1539
rect 4759 -1773 4760 -1539
rect 4524 -1774 4760 -1773
rect 5164 -1539 5400 -1538
rect 5164 -1773 5165 -1539
rect 5165 -1773 5399 -1539
rect 5399 -1773 5400 -1539
rect 5164 -1774 5400 -1773
rect 5804 -1539 6040 -1538
rect 5804 -1773 5805 -1539
rect 5805 -1773 6039 -1539
rect 6039 -1773 6040 -1539
rect 5804 -1774 6040 -1773
rect 6444 -1539 6680 -1538
rect 6444 -1773 6445 -1539
rect 6445 -1773 6679 -1539
rect 6679 -1773 6680 -1539
rect 6444 -1774 6680 -1773
rect 7084 -1539 7320 -1538
rect 7084 -1773 7085 -1539
rect 7085 -1773 7319 -1539
rect 7319 -1773 7320 -1539
rect 7084 -1774 7320 -1773
rect 7724 -1539 7960 -1538
rect 7724 -1773 7725 -1539
rect 7725 -1773 7959 -1539
rect 7959 -1773 7960 -1539
rect 7724 -1774 7960 -1773
rect 8364 -1539 8600 -1538
rect 8364 -1773 8365 -1539
rect 8365 -1773 8599 -1539
rect 8599 -1773 8600 -1539
rect 8364 -1774 8600 -1773
rect 9004 -1539 9240 -1538
rect 9004 -1773 9005 -1539
rect 9005 -1773 9239 -1539
rect 9239 -1773 9240 -1539
rect 9004 -1774 9240 -1773
rect 9644 -1539 9880 -1538
rect 9644 -1773 9645 -1539
rect 9645 -1773 9879 -1539
rect 9879 -1773 9880 -1539
rect 9644 -1774 9880 -1773
rect 10284 -1539 10520 -1538
rect 10284 -1773 10285 -1539
rect 10285 -1773 10519 -1539
rect 10519 -1773 10520 -1539
rect 10284 -1774 10520 -1773
rect 10924 -1539 11160 -1538
rect 10924 -1773 10925 -1539
rect 10925 -1773 11159 -1539
rect 11159 -1773 11160 -1539
rect 10924 -1774 11160 -1773
rect 11564 -1539 11800 -1538
rect 11564 -1773 11565 -1539
rect 11565 -1773 11799 -1539
rect 11799 -1773 11800 -1539
rect 11564 -1774 11800 -1773
rect 12204 -1539 12440 -1538
rect 12204 -1773 12205 -1539
rect 12205 -1773 12439 -1539
rect 12439 -1773 12440 -1539
rect 12204 -1774 12440 -1773
rect 12844 -1539 13080 -1538
rect 12844 -1773 12845 -1539
rect 12845 -1773 13079 -1539
rect 13079 -1773 13080 -1539
rect 12844 -1774 13080 -1773
rect 13484 -1539 13720 -1538
rect 13484 -1773 13485 -1539
rect 13485 -1773 13719 -1539
rect 13719 -1773 13720 -1539
rect 13484 -1774 13720 -1773
rect 14124 -1539 14360 -1538
rect 14124 -1773 14125 -1539
rect 14125 -1773 14359 -1539
rect 14359 -1773 14360 -1539
rect 14124 -1774 14360 -1773
rect 14764 -1539 15000 -1538
rect 14764 -1773 14765 -1539
rect 14765 -1773 14999 -1539
rect 14999 -1773 15000 -1539
rect 14764 -1774 15000 -1773
rect 15404 -1539 15640 -1538
rect 15404 -1773 15405 -1539
rect 15405 -1773 15639 -1539
rect 15639 -1773 15640 -1539
rect 15404 -1774 15640 -1773
rect 16044 -1539 16280 -1538
rect 16044 -1773 16045 -1539
rect 16045 -1773 16279 -1539
rect 16279 -1773 16280 -1539
rect 16044 -1774 16280 -1773
rect 16684 -1539 16920 -1538
rect 16684 -1773 16685 -1539
rect 16685 -1773 16919 -1539
rect 16919 -1773 16920 -1539
rect 16684 -1774 16920 -1773
rect 17324 -1539 17560 -1538
rect 17324 -1773 17325 -1539
rect 17325 -1773 17559 -1539
rect 17559 -1773 17560 -1539
rect 17324 -1774 17560 -1773
rect 17964 -1539 18200 -1538
rect 17964 -1773 17965 -1539
rect 17965 -1773 18199 -1539
rect 18199 -1773 18200 -1539
rect 17964 -1774 18200 -1773
rect 18604 -1539 18840 -1538
rect 18604 -1773 18605 -1539
rect 18605 -1773 18839 -1539
rect 18839 -1773 18840 -1539
rect 18604 -1774 18840 -1773
rect 19244 -1539 19480 -1538
rect 19244 -1773 19245 -1539
rect 19245 -1773 19479 -1539
rect 19479 -1773 19480 -1539
rect 19244 -1774 19480 -1773
rect 19884 -1539 20120 -1538
rect 19884 -1773 19885 -1539
rect 19885 -1773 20119 -1539
rect 20119 -1773 20120 -1539
rect 19884 -1774 20120 -1773
rect 20524 -1539 20760 -1538
rect 20524 -1773 20525 -1539
rect 20525 -1773 20759 -1539
rect 20759 -1773 20760 -1539
rect 20524 -1774 20760 -1773
rect 21164 -1539 21400 -1538
rect 21164 -1773 21165 -1539
rect 21165 -1773 21399 -1539
rect 21399 -1773 21400 -1539
rect 21164 -1774 21400 -1773
rect 21804 -1539 22040 -1538
rect 21804 -1773 21805 -1539
rect 21805 -1773 22039 -1539
rect 22039 -1773 22040 -1539
rect 21804 -1774 22040 -1773
rect 22444 -1539 22680 -1538
rect 22444 -1773 22445 -1539
rect 22445 -1773 22679 -1539
rect 22679 -1773 22680 -1539
rect 22444 -1774 22680 -1773
rect 23084 -1539 23320 -1538
rect 23084 -1773 23085 -1539
rect 23085 -1773 23319 -1539
rect 23319 -1773 23320 -1539
rect 23084 -1774 23320 -1773
rect 23724 -1539 23960 -1538
rect 23724 -1773 23725 -1539
rect 23725 -1773 23959 -1539
rect 23959 -1773 23960 -1539
rect 23724 -1774 23960 -1773
rect 24364 -1539 24600 -1538
rect 24364 -1773 24365 -1539
rect 24365 -1773 24599 -1539
rect 24599 -1773 24600 -1539
rect 24364 -1774 24600 -1773
rect 25004 -1539 25240 -1538
rect 25004 -1773 25005 -1539
rect 25005 -1773 25239 -1539
rect 25239 -1773 25240 -1539
rect 25004 -1774 25240 -1773
<< metal5 >>
rect -1540 27972 -1220 28197
rect -1800 27930 -1220 27972
rect -1800 27694 -1776 27930
rect -1540 27694 -1220 27930
rect -1800 27652 -1220 27694
rect -900 27972 -580 28204
rect -900 27930 -320 27972
rect -900 27694 -580 27930
rect -344 27694 -320 27930
rect -900 27652 -320 27694
rect -1540 27610 -580 27652
rect -1540 27374 -1220 27610
rect -900 27374 -580 27610
rect -1540 27332 -580 27374
rect -1800 27290 -1220 27332
rect -1800 27054 -1776 27290
rect -1540 27054 -1220 27290
rect -1800 27012 -1220 27054
rect -900 27290 -320 27332
rect -900 27054 -580 27290
rect -344 27054 -320 27290
rect -900 27012 -320 27054
rect -1540 26970 -580 27012
rect -1540 26734 -1220 26970
rect -900 26734 -580 26970
rect -1540 26692 -580 26734
rect 13789 26725 14198 27045
rect -1800 26650 -1220 26692
rect -1800 26414 -1776 26650
rect -1540 26414 -1220 26650
rect -1800 26372 -1220 26414
rect -900 26650 -320 26692
rect -900 26414 -580 26650
rect -344 26414 -320 26650
rect -900 26372 -320 26414
rect -1540 26330 -580 26372
rect -1540 26094 -1220 26330
rect -900 26094 -580 26330
rect -1540 26052 -580 26094
rect -1800 26010 -1220 26052
rect -1800 25774 -1776 26010
rect -1540 25774 -1220 26010
rect -1800 25732 -1220 25774
rect -900 26010 2 26052
rect -900 25774 -580 26010
rect -344 25774 2 26010
rect 13798 25875 14207 26195
rect -900 25732 2 25774
rect -1540 25690 -580 25732
rect -1540 25454 -1220 25690
rect -900 25454 -580 25690
rect -1540 25412 -580 25454
rect -1800 25370 -1220 25412
rect -1800 25134 -1776 25370
rect -1540 25134 -1220 25370
rect -1800 25092 -1220 25134
rect -900 25370 -320 25412
rect -900 25134 -580 25370
rect -344 25134 -320 25370
rect -900 25092 -320 25134
rect -1540 25050 -580 25092
rect -1540 24814 -1220 25050
rect -900 24814 -580 25050
rect 13790 25023 14199 25343
rect -1540 24772 -580 24814
rect -1800 24730 -1220 24772
rect -1800 24494 -1776 24730
rect -1540 24494 -1220 24730
rect -1800 24452 -1220 24494
rect -900 24730 2 24772
rect -900 24494 -580 24730
rect -344 24494 2 24730
rect -900 24452 2 24494
rect -1540 24410 -580 24452
rect -1540 24174 -1220 24410
rect -900 24174 -580 24410
rect -1540 24132 -580 24174
rect -1800 24090 -1220 24132
rect -1800 23854 -1776 24090
rect -1540 23854 -1220 24090
rect -1800 23812 -1220 23854
rect -900 24090 -320 24132
rect -900 23854 -580 24090
rect -344 23854 -320 24090
rect -900 23812 -320 23854
rect -1540 23770 -580 23812
rect -1540 23534 -1220 23770
rect -900 23534 -580 23770
rect -1540 23492 -580 23534
rect -1800 23450 -1220 23492
rect -1800 23214 -1776 23450
rect -1540 23214 -1220 23450
rect -1800 23172 -1220 23214
rect -900 23450 2 23492
rect -900 23214 -580 23450
rect -344 23214 2 23450
rect 13785 23322 14194 23642
rect -900 23172 2 23214
rect -1540 23130 -580 23172
rect -1540 22894 -1220 23130
rect -900 22894 -580 23130
rect -1540 22852 -580 22894
rect -1800 22810 -1220 22852
rect -1800 22574 -1776 22810
rect -1540 22574 -1220 22810
rect -1800 22532 -1220 22574
rect -900 22810 -320 22852
rect -900 22574 -580 22810
rect -344 22574 -320 22810
rect -900 22532 -320 22574
rect -1540 22490 -580 22532
rect -1540 22254 -1220 22490
rect -900 22254 -580 22490
rect 13795 22427 14204 22747
rect -1540 22212 -580 22254
rect -1800 22170 -1220 22212
rect -1800 21934 -1776 22170
rect -1540 21934 -1220 22170
rect -1800 21892 -1220 21934
rect -900 22170 2 22212
rect -900 21934 -580 22170
rect -344 21934 2 22170
rect -900 21892 2 21934
rect -1540 21850 -580 21892
rect -1540 21614 -1220 21850
rect -900 21614 -580 21850
rect -1540 21572 -580 21614
rect -1800 21530 -1220 21572
rect -1800 21294 -1776 21530
rect -1540 21294 -1220 21530
rect -1800 21252 -1220 21294
rect -900 21530 -320 21572
rect 13786 21544 14195 21864
rect -900 21294 -580 21530
rect -344 21294 -320 21530
rect -900 21252 -320 21294
rect -1540 21210 -580 21252
rect -1540 20974 -1220 21210
rect -900 20974 -580 21210
rect -1540 20932 -580 20974
rect -1800 20890 -1220 20932
rect -1800 20654 -1776 20890
rect -1540 20654 -1220 20890
rect -1800 20612 -1220 20654
rect -900 20890 2 20932
rect -900 20654 -580 20890
rect -344 20654 2 20890
rect -900 20612 2 20654
rect -1540 20570 -580 20612
rect -1540 20334 -1220 20570
rect -900 20334 -580 20570
rect -1540 20292 -580 20334
rect -1800 20250 -1220 20292
rect -1800 20014 -1776 20250
rect -1540 20014 -1220 20250
rect -1800 19972 -1220 20014
rect -900 20250 -320 20292
rect -900 20014 -580 20250
rect -344 20014 -320 20250
rect -900 19972 -320 20014
rect -1540 19930 -580 19972
rect -1540 19694 -1220 19930
rect -900 19694 -580 19930
rect 13805 19840 14214 20160
rect -1540 19652 -580 19694
rect -1800 19610 -1220 19652
rect -1800 19374 -1776 19610
rect -1540 19374 -1220 19610
rect -1800 19332 -1220 19374
rect -900 19610 2 19652
rect -900 19374 -580 19610
rect -344 19374 2 19610
rect -900 19332 2 19374
rect -1540 19290 -580 19332
rect -1540 19054 -1220 19290
rect -900 19054 -580 19290
rect -1540 19012 -580 19054
rect -1800 18970 -1220 19012
rect -1800 18734 -1776 18970
rect -1540 18734 -1220 18970
rect -1800 18692 -1220 18734
rect -900 18970 -320 19012
rect -900 18734 -580 18970
rect -344 18734 -320 18970
rect 13800 18958 14209 19278
rect -900 18692 -320 18734
rect -1540 18650 -580 18692
rect -1540 18414 -1220 18650
rect -900 18414 -580 18650
rect -1540 18372 -580 18414
rect -1800 18330 -1220 18372
rect -1800 18094 -1776 18330
rect -1540 18094 -1220 18330
rect -1800 18052 -1220 18094
rect -900 18330 2 18372
rect -900 18094 -580 18330
rect -344 18094 2 18330
rect -900 18052 2 18094
rect 13811 18061 14220 18381
rect -1540 18010 -580 18052
rect -1540 17774 -1220 18010
rect -900 17774 -580 18010
rect -1540 17732 -580 17774
rect -1800 17690 -1220 17732
rect -1800 17454 -1776 17690
rect -1540 17454 -1220 17690
rect -1800 17412 -1220 17454
rect -900 17690 -320 17732
rect -900 17454 -580 17690
rect -344 17454 -320 17690
rect -900 17412 -320 17454
rect -1540 17370 -580 17412
rect -1540 17134 -1220 17370
rect -900 17134 -580 17370
rect -1540 17092 -580 17134
rect -1800 17050 -1220 17092
rect -1800 16814 -1776 17050
rect -1540 16814 -1220 17050
rect -1800 16772 -1220 16814
rect -900 17050 2 17092
rect -900 16814 -580 17050
rect -344 16814 2 17050
rect -900 16772 2 16814
rect -1540 16730 -580 16772
rect -1540 16494 -1220 16730
rect -900 16494 -580 16730
rect -1540 16452 -580 16494
rect -1800 16410 -1220 16452
rect -1800 16174 -1776 16410
rect -1540 16174 -1220 16410
rect -1800 16132 -1220 16174
rect -900 16410 -320 16452
rect -900 16174 -580 16410
rect -344 16174 -320 16410
rect 13800 16368 14209 16688
rect -900 16132 -320 16174
rect -1540 16090 -580 16132
rect -1540 15854 -1220 16090
rect -900 15854 -580 16090
rect -1540 15812 -580 15854
rect -1800 15770 -1220 15812
rect -1800 15534 -1776 15770
rect -1540 15534 -1220 15770
rect -1800 15492 -1220 15534
rect -900 15770 2 15812
rect -900 15534 -580 15770
rect -344 15534 2 15770
rect -900 15492 2 15534
rect -1540 15450 -580 15492
rect 13806 15470 14215 15790
rect -1540 15214 -1220 15450
rect -900 15214 -580 15450
rect -1540 15172 -580 15214
rect -1800 15130 -1220 15172
rect -1800 14894 -1776 15130
rect -1540 14894 -1220 15130
rect -1800 14852 -1220 14894
rect -900 15130 -320 15172
rect -900 14894 -580 15130
rect -344 14894 -320 15130
rect -900 14852 -320 14894
rect -1540 14810 -580 14852
rect -1540 14574 -1220 14810
rect -900 14574 -580 14810
rect 13809 14577 14218 14897
rect -1540 14532 -580 14574
rect -1800 14490 -1220 14532
rect -1800 14254 -1776 14490
rect -1540 14254 -1220 14490
rect -1800 14212 -1220 14254
rect -900 14490 2 14532
rect -900 14254 -580 14490
rect -344 14254 2 14490
rect -900 14212 2 14254
rect -1540 14170 -580 14212
rect -1540 13934 -1220 14170
rect -900 13934 -580 14170
rect -1540 13892 -580 13934
rect -1800 13850 -1220 13892
rect -1800 13614 -1776 13850
rect -1540 13614 -1220 13850
rect -1800 13572 -1220 13614
rect -900 13850 -320 13892
rect -900 13614 -580 13850
rect -344 13614 -320 13850
rect -900 13572 -320 13614
rect -1540 13530 -580 13572
rect -1540 13294 -1220 13530
rect -900 13294 -580 13530
rect -1540 13252 -580 13294
rect -1800 13210 -1220 13252
rect -1800 12974 -1776 13210
rect -1540 12974 -1220 13210
rect -1800 12932 -1220 12974
rect -900 13210 2 13252
rect -900 12974 -580 13210
rect -344 12974 2 13210
rect -900 12932 2 12974
rect -1540 12890 -580 12932
rect -1540 12654 -1220 12890
rect -900 12654 -580 12890
rect 13814 12881 14223 13201
rect -1540 12612 -580 12654
rect -1800 12570 -1220 12612
rect -1800 12334 -1776 12570
rect -1540 12334 -1220 12570
rect -1800 12292 -1220 12334
rect -900 12570 -320 12612
rect -900 12334 -580 12570
rect -344 12334 -320 12570
rect -900 12292 -320 12334
rect -1540 12250 -580 12292
rect -1540 12014 -1220 12250
rect -900 12014 -580 12250
rect -1540 11972 -580 12014
rect 13809 11988 14218 12308
rect -1800 11930 -1220 11972
rect -1800 11694 -1776 11930
rect -1540 11694 -1220 11930
rect -1800 11652 -1220 11694
rect -900 11930 2 11972
rect -900 11694 -580 11930
rect -344 11694 2 11930
rect -900 11652 2 11694
rect -1540 11610 -580 11652
rect -1540 11374 -1220 11610
rect -900 11374 -580 11610
rect -1540 11332 -580 11374
rect -1800 11290 -1220 11332
rect -1800 11054 -1776 11290
rect -1540 11054 -1220 11290
rect -1800 11012 -1220 11054
rect -900 11290 -320 11332
rect -900 11054 -580 11290
rect -344 11054 -320 11290
rect 13815 11093 14224 11413
rect -900 11012 -320 11054
rect -1540 10970 -580 11012
rect -1540 10734 -1220 10970
rect -900 10734 -580 10970
rect -1540 10692 -580 10734
rect -1800 10650 -1220 10692
rect -1800 10414 -1776 10650
rect -1540 10414 -1220 10650
rect -1800 10372 -1220 10414
rect -900 10650 2 10692
rect -900 10414 -580 10650
rect -344 10414 2 10650
rect -900 10372 2 10414
rect -1540 10330 -580 10372
rect -1540 10094 -1220 10330
rect -900 10094 -580 10330
rect -1540 10052 -580 10094
rect -1800 10010 -1220 10052
rect -1800 9774 -1776 10010
rect -1540 9774 -1220 10010
rect -1800 9732 -1220 9774
rect -900 10010 -320 10052
rect -900 9774 -580 10010
rect -344 9774 -320 10010
rect -900 9732 -320 9774
rect -1540 9690 -580 9732
rect -1540 9454 -1220 9690
rect -900 9454 -580 9690
rect -1540 9412 -580 9454
rect -1800 9370 -1220 9412
rect -1800 9134 -1776 9370
rect -1540 9134 -1220 9370
rect -1800 9092 -1220 9134
rect -900 9370 2 9412
rect 13813 9395 14222 9715
rect -900 9134 -580 9370
rect -344 9134 2 9370
rect -900 9092 2 9134
rect -1540 9050 -580 9092
rect -1540 8814 -1220 9050
rect -900 8814 -580 9050
rect -1540 8772 -580 8814
rect -1800 8730 -1220 8772
rect -1800 8494 -1776 8730
rect -1540 8494 -1220 8730
rect -1800 8452 -1220 8494
rect -900 8730 -320 8772
rect -900 8494 -580 8730
rect -344 8494 -320 8730
rect 13810 8502 14219 8822
rect -900 8452 -320 8494
rect -1540 8410 -580 8452
rect -1540 8174 -1220 8410
rect -900 8174 -580 8410
rect -1540 8132 -580 8174
rect -1800 8090 -1220 8132
rect -1800 7854 -1776 8090
rect -1540 7854 -1220 8090
rect -1800 7812 -1220 7854
rect -900 8090 2 8132
rect -900 7854 -580 8090
rect -344 7854 2 8090
rect -900 7812 2 7854
rect -1540 7770 -580 7812
rect -1540 7534 -1220 7770
rect -900 7534 -580 7770
rect 13806 7610 14208 7930
rect -1540 7492 -580 7534
rect -1800 7450 -1220 7492
rect -1800 7214 -1776 7450
rect -1540 7214 -1220 7450
rect -1800 7172 -1220 7214
rect -900 7450 -320 7492
rect -900 7214 -580 7450
rect -344 7214 -320 7450
rect -900 7172 -320 7214
rect -1540 7130 -580 7172
rect -1540 6894 -1220 7130
rect -900 6894 -580 7130
rect -1540 6852 -580 6894
rect -1800 6810 -1220 6852
rect -1800 6574 -1776 6810
rect -1540 6574 -1220 6810
rect -1800 6532 -1220 6574
rect -900 6810 2 6852
rect -900 6574 -580 6810
rect -344 6574 2 6810
rect -900 6532 2 6574
rect -1540 6490 -580 6532
rect -1540 6254 -1220 6490
rect -900 6254 -580 6490
rect -1540 6212 -580 6254
rect -1800 6170 -1220 6212
rect -1800 5934 -1776 6170
rect -1540 5934 -1220 6170
rect -1800 5892 -1220 5934
rect -900 6170 -320 6212
rect -900 5934 -580 6170
rect -344 5934 -320 6170
rect -900 5892 -320 5934
rect 13808 5914 14210 6234
rect -1540 5850 -580 5892
rect -1540 5614 -1220 5850
rect -900 5614 -580 5850
rect -1540 5572 -580 5614
rect -1800 5530 -1220 5572
rect -1800 5294 -1776 5530
rect -1540 5294 -1220 5530
rect -1800 5252 -1220 5294
rect -900 5530 2 5572
rect -900 5294 -580 5530
rect -344 5294 2 5530
rect -900 5252 2 5294
rect -1540 5210 -580 5252
rect -1540 4974 -1220 5210
rect -900 4974 -580 5210
rect 13812 5020 14214 5340
rect -1540 4932 -580 4974
rect -1800 4890 -1220 4932
rect -1800 4654 -1776 4890
rect -1540 4654 -1220 4890
rect -1800 4612 -1220 4654
rect -900 4890 -320 4932
rect -900 4654 -580 4890
rect -344 4654 -320 4890
rect -900 4612 -320 4654
rect -1540 4570 -580 4612
rect -1540 4334 -1220 4570
rect -900 4334 -580 4570
rect -1540 4292 -580 4334
rect -1800 4250 -1220 4292
rect -1800 4014 -1776 4250
rect -1540 4014 -1220 4250
rect -1800 3972 -1220 4014
rect -900 4250 2 4292
rect -900 4014 -580 4250
rect -344 4014 2 4250
rect 13804 4126 14206 4446
rect -900 3972 2 4014
rect -1540 3930 -580 3972
rect -1540 3694 -1220 3930
rect -900 3694 -580 3930
rect -1540 3652 -580 3694
rect -1800 3610 -1220 3652
rect -1800 3374 -1776 3610
rect -1540 3374 -1220 3610
rect -1800 3332 -1220 3374
rect -900 3610 -320 3652
rect -900 3374 -580 3610
rect -344 3374 -320 3610
rect -900 3332 -320 3374
rect -1540 3290 -580 3332
rect -1540 3054 -1220 3290
rect -900 3054 -580 3290
rect -1540 3012 -580 3054
rect -1800 2970 -1220 3012
rect -1800 2734 -1776 2970
rect -1540 2734 -1220 2970
rect -1800 2692 -1220 2734
rect -900 2970 2 3012
rect -900 2734 -580 2970
rect -344 2734 2 2970
rect -900 2692 2 2734
rect -1540 2650 -580 2692
rect -1540 2414 -1220 2650
rect -900 2414 -580 2650
rect 13812 2430 14214 2750
rect -1540 2372 -580 2414
rect -1800 2330 -1220 2372
rect -1800 2094 -1776 2330
rect -1540 2094 -1220 2330
rect -1800 2052 -1220 2094
rect -900 2330 -320 2372
rect -900 2094 -580 2330
rect -344 2094 -320 2330
rect -900 2052 -320 2094
rect -1540 2010 -580 2052
rect -1540 1774 -1220 2010
rect -900 1774 -580 2010
rect -1540 1732 -580 1774
rect -1800 1690 -1220 1732
rect -1800 1454 -1776 1690
rect -1540 1454 -1220 1690
rect -1800 1412 -1220 1454
rect -1540 -578 -1220 1412
rect -900 1690 2 1732
rect -900 1454 -580 1690
rect -344 1454 2 1690
rect 13803 1541 14212 1861
rect -900 1412 2 1454
rect -900 -578 -580 1412
rect 13794 676 14203 996
rect 2 -342 322 13
rect 2 -578 44 -342
rect 280 -578 322 -342
rect 642 -342 962 -318
rect 642 -578 684 -342
rect 920 -578 962 -342
rect 1282 -342 1602 2
rect 1282 -578 1324 -342
rect 1560 -578 1602 -342
rect 1922 -342 2242 -318
rect 1922 -578 1964 -342
rect 2200 -578 2242 -342
rect 2562 -342 2882 2
rect 2562 -578 2604 -342
rect 2840 -578 2882 -342
rect 3202 -342 3522 -318
rect 3202 -578 3244 -342
rect 3480 -578 3522 -342
rect 3842 -342 4162 2
rect 3842 -578 3884 -342
rect 4120 -578 4162 -342
rect 4482 -342 4802 -318
rect 4482 -578 4524 -342
rect 4760 -578 4802 -342
rect 5122 -342 5442 2
rect 5122 -578 5164 -342
rect 5400 -578 5442 -342
rect 5762 -342 6082 -318
rect 5762 -578 5804 -342
rect 6040 -578 6082 -342
rect 6402 -342 6722 2
rect 6402 -578 6444 -342
rect 6680 -578 6722 -342
rect 7042 -342 7362 -318
rect 7042 -578 7084 -342
rect 7320 -578 7362 -342
rect 7682 -342 8002 2
rect 7682 -578 7724 -342
rect 7960 -578 8002 -342
rect 8322 -342 8642 -318
rect 8322 -578 8364 -342
rect 8600 -578 8642 -342
rect 8962 -342 9282 2
rect 8962 -578 9004 -342
rect 9240 -578 9282 -342
rect 9602 -342 9922 -318
rect 9602 -578 9644 -342
rect 9880 -578 9922 -342
rect 10242 -342 10562 2
rect 10242 -578 10284 -342
rect 10520 -578 10562 -342
rect 10882 -342 11202 -318
rect 10882 -578 10924 -342
rect 11160 -578 11202 -342
rect 11522 -342 11842 2
rect 11522 -578 11564 -342
rect 11800 -578 11842 -342
rect 12162 -342 12482 -318
rect 12162 -578 12204 -342
rect 12440 -578 12482 -342
rect 12802 -342 13122 2
rect 12802 -578 12844 -342
rect 13080 -578 13122 -342
rect 13442 -342 13762 -318
rect 13442 -578 13484 -342
rect 13720 -578 13762 -342
rect 14082 -342 14402 -318
rect 14082 -578 14124 -342
rect 14360 -578 14402 -342
rect 14722 -342 15042 -318
rect 14722 -578 14764 -342
rect 15000 -578 15042 -342
rect 15362 -342 15682 2
rect 15362 -578 15404 -342
rect 15640 -578 15682 -342
rect 16002 -342 16322 -318
rect 16002 -578 16044 -342
rect 16280 -578 16322 -342
rect 16642 -342 16962 2
rect 16642 -578 16684 -342
rect 16920 -578 16962 -342
rect 17282 -342 17602 -318
rect 17282 -578 17324 -342
rect 17560 -578 17602 -342
rect 17922 -342 18242 2
rect 17922 -578 17964 -342
rect 18200 -578 18242 -342
rect 18562 -342 18882 -318
rect 18562 -578 18604 -342
rect 18840 -578 18882 -342
rect 19202 -342 19522 2
rect 19202 -578 19244 -342
rect 19480 -578 19522 -342
rect 19842 -342 20162 -318
rect 19842 -578 19884 -342
rect 20120 -578 20162 -342
rect 20482 -342 20802 2
rect 20482 -578 20524 -342
rect 20760 -578 20802 -342
rect 21122 -342 21442 -318
rect 21122 -578 21164 -342
rect 21400 -578 21442 -342
rect 21762 -342 22082 -318
rect 21762 -578 21804 -342
rect 22040 -578 22082 -342
rect 22402 -342 22722 -318
rect 22402 -578 22444 -342
rect 22680 -578 22722 -342
rect 23042 -342 23362 -318
rect 23042 -578 23084 -342
rect 23320 -578 23362 -342
rect 23682 -342 24002 -318
rect 23682 -578 23724 -342
rect 23960 -578 24002 -342
rect 24322 -342 24642 -318
rect 24322 -578 24364 -342
rect 24600 -578 24642 -342
rect 24962 -342 25282 -318
rect 24962 -578 25004 -342
rect 25240 -578 25282 -342
rect -1540 -898 25922 -578
rect -1540 -1218 -1220 -898
rect 322 -1218 364 -898
rect 600 -1218 642 -898
rect 962 -1218 1004 -898
rect 1240 -1218 1282 -898
rect 1602 -1218 1644 -898
rect 1880 -1218 1922 -898
rect 2242 -1218 2284 -898
rect 2520 -1218 2562 -898
rect 2882 -1218 2924 -898
rect 3160 -1218 3202 -898
rect 3522 -1218 3564 -898
rect 3800 -1218 3842 -898
rect 4162 -1218 4204 -898
rect 4440 -1218 4482 -898
rect 4802 -1218 4844 -898
rect 5080 -1218 5122 -898
rect 5442 -1218 5484 -898
rect 5720 -1218 5762 -898
rect 6082 -1218 6124 -898
rect 6360 -1218 6402 -898
rect 6722 -1218 6764 -898
rect 7000 -1218 7042 -898
rect 7362 -1218 7404 -898
rect 7640 -1218 7682 -898
rect 8002 -1218 8044 -898
rect 8280 -1218 8322 -898
rect 8642 -1218 8684 -898
rect 8920 -1218 8962 -898
rect 9282 -1218 9324 -898
rect 9560 -1218 9602 -898
rect 9922 -1218 9964 -898
rect 10200 -1218 10242 -898
rect 10562 -1218 10604 -898
rect 10840 -1218 10882 -898
rect 11202 -1218 11244 -898
rect 11480 -1218 11522 -898
rect 11842 -1218 11884 -898
rect 12120 -1218 12162 -898
rect 12482 -1218 12524 -898
rect 12760 -1218 12802 -898
rect 13122 -1218 13164 -898
rect 13400 -1218 13442 -898
rect 13762 -1218 13804 -898
rect 14040 -1218 14082 -898
rect 14402 -1218 14444 -898
rect 14680 -1218 14722 -898
rect 15042 -1218 15084 -898
rect 15320 -1218 15362 -898
rect 15682 -1218 15724 -898
rect 15960 -1218 16002 -898
rect 16322 -1218 16364 -898
rect 16600 -1218 16642 -898
rect 16962 -1218 17004 -898
rect 17240 -1218 17282 -898
rect 17602 -1218 17644 -898
rect 17880 -1218 17922 -898
rect 18242 -1218 18284 -898
rect 18520 -1218 18562 -898
rect 18882 -1218 18924 -898
rect 19160 -1218 19202 -898
rect 19522 -1218 19564 -898
rect 19800 -1218 19842 -898
rect 20162 -1218 20204 -898
rect 20440 -1218 20482 -898
rect 20802 -1218 20844 -898
rect 21080 -1218 21122 -898
rect 21442 -1218 21484 -898
rect 21720 -1218 21762 -898
rect 22082 -1218 22124 -898
rect 22360 -1218 22402 -898
rect 22722 -1218 22764 -898
rect 23000 -1218 23042 -898
rect 23362 -1218 23404 -898
rect 23640 -1218 23682 -898
rect 24002 -1218 24044 -898
rect 24280 -1218 24322 -898
rect 24642 -1218 24684 -898
rect 24920 -1218 24962 -898
rect -1540 -1538 25922 -1218
rect 2 -1774 44 -1538
rect 280 -1774 322 -1538
rect 2 -1798 322 -1774
rect 642 -1774 684 -1538
rect 920 -1774 962 -1538
rect 642 -1798 962 -1774
rect 1282 -1774 1324 -1538
rect 1560 -1774 1602 -1538
rect 1282 -1798 1602 -1774
rect 1922 -1774 1964 -1538
rect 2200 -1774 2242 -1538
rect 1922 -1798 2242 -1774
rect 2562 -1774 2604 -1538
rect 2840 -1774 2882 -1538
rect 2562 -1798 2882 -1774
rect 3202 -1774 3244 -1538
rect 3480 -1774 3522 -1538
rect 3202 -1798 3522 -1774
rect 3842 -1774 3884 -1538
rect 4120 -1774 4162 -1538
rect 3842 -1798 4162 -1774
rect 4482 -1774 4524 -1538
rect 4760 -1774 4802 -1538
rect 4482 -1798 4802 -1774
rect 5122 -1774 5164 -1538
rect 5400 -1774 5442 -1538
rect 5122 -1798 5442 -1774
rect 5762 -1774 5804 -1538
rect 6040 -1774 6082 -1538
rect 5762 -1798 6082 -1774
rect 6402 -1774 6444 -1538
rect 6680 -1774 6722 -1538
rect 6402 -1798 6722 -1774
rect 7042 -1774 7084 -1538
rect 7320 -1774 7362 -1538
rect 7042 -1798 7362 -1774
rect 7682 -1774 7724 -1538
rect 7960 -1774 8002 -1538
rect 7682 -1798 8002 -1774
rect 8322 -1774 8364 -1538
rect 8600 -1774 8642 -1538
rect 8322 -1798 8642 -1774
rect 8962 -1774 9004 -1538
rect 9240 -1774 9282 -1538
rect 8962 -1798 9282 -1774
rect 9602 -1774 9644 -1538
rect 9880 -1774 9922 -1538
rect 9602 -1798 9922 -1774
rect 10242 -1774 10284 -1538
rect 10520 -1774 10562 -1538
rect 10242 -1798 10562 -1774
rect 10882 -1774 10924 -1538
rect 11160 -1774 11202 -1538
rect 10882 -1798 11202 -1774
rect 11522 -1774 11564 -1538
rect 11800 -1774 11842 -1538
rect 11522 -1798 11842 -1774
rect 12162 -1774 12204 -1538
rect 12440 -1774 12482 -1538
rect 12162 -1798 12482 -1774
rect 12802 -1774 12844 -1538
rect 13080 -1774 13122 -1538
rect 12802 -1798 13122 -1774
rect 13442 -1774 13484 -1538
rect 13720 -1774 13762 -1538
rect 13442 -1798 13762 -1774
rect 14082 -1774 14124 -1538
rect 14360 -1774 14402 -1538
rect 14082 -1798 14402 -1774
rect 14722 -1774 14764 -1538
rect 15000 -1774 15042 -1538
rect 14722 -1798 15042 -1774
rect 15362 -1774 15404 -1538
rect 15640 -1774 15682 -1538
rect 15362 -1798 15682 -1774
rect 16002 -1774 16044 -1538
rect 16280 -1774 16322 -1538
rect 16002 -1798 16322 -1774
rect 16642 -1774 16684 -1538
rect 16920 -1774 16962 -1538
rect 16642 -1798 16962 -1774
rect 17282 -1774 17324 -1538
rect 17560 -1774 17602 -1538
rect 17282 -1798 17602 -1774
rect 17922 -1774 17964 -1538
rect 18200 -1774 18242 -1538
rect 17922 -1798 18242 -1774
rect 18562 -1774 18604 -1538
rect 18840 -1774 18882 -1538
rect 18562 -1798 18882 -1774
rect 19202 -1774 19244 -1538
rect 19480 -1774 19522 -1538
rect 19202 -1798 19522 -1774
rect 19842 -1774 19884 -1538
rect 20120 -1774 20162 -1538
rect 19842 -1798 20162 -1774
rect 20482 -1774 20524 -1538
rect 20760 -1774 20802 -1538
rect 20482 -1798 20802 -1774
rect 21122 -1774 21164 -1538
rect 21400 -1774 21442 -1538
rect 21122 -1798 21442 -1774
rect 21762 -1774 21804 -1538
rect 22040 -1774 22082 -1538
rect 21762 -1798 22082 -1774
rect 22402 -1774 22444 -1538
rect 22680 -1774 22722 -1538
rect 22402 -1798 22722 -1774
rect 23042 -1774 23084 -1538
rect 23320 -1774 23362 -1538
rect 23042 -1798 23362 -1774
rect 23682 -1774 23724 -1538
rect 23960 -1774 24002 -1538
rect 23682 -1798 24002 -1774
rect 24322 -1774 24364 -1538
rect 24600 -1774 24642 -1538
rect 24322 -1798 24642 -1774
rect 24962 -1774 25004 -1538
rect 25240 -1774 25282 -1538
rect 24962 -1798 25282 -1774
use cap_3pF  cap_3pF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654658877
transform 0 1 19258 -1 0 21107
box -6669 2096 15759 5484
use cap_6pF  cap_6pF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654658794
transform 0 1 17599 -1 0 24342
box -2674 -2673 19758 3439
use cap_10fF  cap_10fF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654307754
transform 1 0 21137 0 1 28534
box -28 -28 708 628
use cap_10fF  cap_10fF_1
timestamp 1654307754
transform 1 0 5164 0 1 28515
box -28 -28 708 628
use cap_12pF  cap_12pF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654658794
transform 0 1 3438 -1 0 24342
box -2674 -2674 19758 8878
use cap_20fF  cap_20fF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654307754
transform 1 0 14293 0 1 28538
box -28 -28 828 1028
use cap_40fF  cap_40fF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654602114
transform 1 0 159 0 1 28488
box -28 -28 1368 1228
use cmos_switch  cmos_switch_0 ~/Documents/fossi_cochlea/mag/final_designs/switch
timestamp 1654602114
transform 1 0 -183 0 1 28398
box -175 -95 235 381
use cmos_switch  cmos_switch_1
timestamp 1654602114
transform -1 0 1877 0 1 28398
box -175 -95 235 381
use cmos_switch  cmos_switch_2
timestamp 1654602114
transform 1 0 13817 0 1 28398
box -175 -95 235 381
use cmos_switch  cmos_switch_3
timestamp 1654602114
transform -1 0 15435 0 1 28398
box -175 -95 235 381
use cmos_switch  cmos_switch_4
timestamp 1654602114
transform 1 0 20717 0 1 28398
box -175 -95 235 381
use cmos_switch  cmos_switch_5
timestamp 1654602114
transform -1 0 22277 0 1 28398
box -175 -95 235 381
use cmos_switch  cmos_switch_6
timestamp 1654602114
transform 1 0 4817 0 1 28398
box -175 -95 235 381
use cmos_switch  cmos_switch_7
timestamp 1654602114
transform -1 0 6187 0 1 28398
box -175 -95 235 381
use mux  mux_0 ~/Documents/fossi_cochlea/mag/final_designs/mux
timestamp 1654652041
transform 0 -1 -744 1 0 28489
box -224 -79 685 681
<< end >>
