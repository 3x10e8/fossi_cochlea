magic
tech sky130A
magscale 1 2
timestamp 1654748317
<< nwell >>
rect 987 322 1294 630
<< nmos >>
rect 1108 96 1138 180
<< pmos >>
rect 1106 466 1136 550
<< ndiff >>
rect 1034 168 1108 180
rect 1034 110 1054 168
rect 1088 110 1108 168
rect 1034 96 1108 110
rect 1138 168 1212 180
rect 1138 110 1158 168
rect 1192 110 1212 168
rect 1138 96 1212 110
<< pdiff >>
rect 1032 538 1106 550
rect 1032 480 1052 538
rect 1086 480 1106 538
rect 1032 466 1106 480
rect 1136 538 1210 550
rect 1136 480 1156 538
rect 1190 480 1210 538
rect 1136 466 1210 480
<< ndiffc >>
rect 1054 110 1088 168
rect 1158 110 1192 168
<< pdiffc >>
rect 1052 480 1086 538
rect 1156 480 1190 538
<< poly >>
rect 1106 550 1136 576
rect 1106 400 1136 466
rect 1090 388 1156 400
rect 1090 354 1106 388
rect 1140 354 1156 388
rect 1090 340 1156 354
rect 1090 258 1156 270
rect 1090 224 1106 258
rect 1140 224 1156 258
rect 1090 212 1156 224
rect 1108 180 1138 212
rect 1108 70 1138 96
<< polycont >>
rect 1106 354 1140 388
rect 1106 224 1140 258
<< locali >>
rect 1036 538 1102 546
rect 1036 480 1052 538
rect 1086 480 1102 538
rect 1036 470 1102 480
rect 1140 538 1210 546
rect 1140 480 1156 538
rect 1190 480 1210 538
rect 1140 470 1210 480
rect 1090 388 1156 400
rect 1090 354 1106 388
rect 1140 354 1156 388
rect 1090 340 1156 354
rect 1106 270 1140 340
rect 1090 260 1156 270
rect 1090 258 1203 260
rect 1090 224 1106 258
rect 1140 224 1203 258
rect 1241 224 1245 260
rect 1090 212 1156 224
rect 1038 168 1104 176
rect 1038 110 1054 168
rect 1088 110 1104 168
rect 1038 100 1104 110
rect 1142 168 1212 176
rect 1142 110 1158 168
rect 1192 110 1212 168
rect 1142 100 1212 110
<< viali >>
rect 1052 480 1086 538
rect 1156 480 1190 538
rect 1203 224 1241 260
rect 1054 110 1088 168
rect 1158 110 1192 168
<< metal1 >>
rect 1140 584 1210 652
rect 1156 546 1190 584
rect 1040 538 1098 546
rect 1040 480 1052 538
rect 1086 480 1098 538
rect 1040 470 1098 480
rect 1144 538 1202 546
rect 1144 480 1156 538
rect 1190 480 1202 538
rect 1144 470 1202 480
rect 1042 176 1076 470
rect 1189 260 1255 274
rect 1189 224 1203 260
rect 1241 224 1255 260
rect 1189 210 1255 224
rect 1042 168 1100 176
rect 1042 110 1054 168
rect 1088 110 1100 168
rect 1042 100 1100 110
rect 1146 168 1204 176
rect 1146 110 1158 168
rect 1192 110 1204 168
rect 1146 92 1204 110
rect 1144 32 1208 92
<< labels >>
rlabel viali 1221 244 1221 244 3 A
port 3 e
<< end >>
