magic
tech sky130A
magscale 1 2
timestamp 1654749871
use unison_side_1  unison_side_1_0
timestamp 1654749871
transform 1 0 -22 0 1 -14
box 0 0 443111 35463
use unison_side_1  unison_side_1_1
timestamp 1654749871
transform 1 0 -22 0 -1 152912
box 0 0 443111 35463
<< end >>
