magic
tech sky130A
magscale 1 2
timestamp 1654479361
<< error_s >>
rect -40 433 -39 517
rect -8 450 45 503
rect 125 450 178 502
rect 258 450 312 503
rect 392 450 445 502
rect 525 450 578 503
rect 609 433 610 517
rect 56 362 91 386
rect -133 355 97 362
rect 43 352 97 355
rect 212 352 247 386
rect 323 352 358 386
rect 479 362 514 386
rect 473 355 703 362
rect 473 352 527 355
rect 50 346 96 352
rect 474 346 520 352
rect 50 338 90 346
rect 480 338 520 346
rect -161 327 125 334
rect 15 324 125 327
rect 445 327 731 334
rect 445 324 555 327
rect 22 318 124 324
rect 446 318 548 324
rect 22 310 118 318
rect 452 310 548 318
rect 56 172 91 206
rect 212 172 247 206
rect 258 202 312 254
rect 323 172 358 206
rect 479 172 514 206
rect -40 48 -39 132
rect -9 63 45 115
rect 125 63 178 115
rect 258 63 312 115
rect 392 63 445 115
rect 525 63 579 115
rect 609 48 610 132
<< nwell >>
rect 258 450 312 503
<< pdiff >>
rect 258 450 312 503
<< locali >>
rect 258 450 312 503
rect 242 352 328 386
rect 242 172 328 206
rect -8 14 43 55
rect 527 14 578 52
rect -8 -20 578 14
<< via1 >>
rect 258 450 312 503
<< metal2 >>
rect 258 503 312 509
rect 258 444 312 450
use mux  mux_0
timestamp 1654479361
transform 1 0 91 0 1 -31
box -224 -79 685 681
use mux  mux_1
timestamp 1654479361
transform -1 0 479 0 1 -31
box -224 -79 685 681
<< end >>
