magic
tech sky130B
magscale 1 2
timestamp 1663464516
use filter_p_m  filter_p_m_0
array 0 7 50784 0 0 13945
timestamp 1663464270
transform 1 0 26 0 1 0
box -26 0 51192 35689
<< end >>
