magic
tech sky130A
timestamp 1647809156
<< nwell >>
rect -191 -3 226 82
rect 383 -4 923 81
<< pmos >>
rect -144 17 -129 59
rect -100 17 -85 59
rect 0 17 15 59
rect 44 17 59 59
rect 88 17 103 59
rect 132 17 147 59
rect 431 16 446 58
rect 476 16 491 58
rect 622 16 637 58
rect 669 16 684 58
rect 815 16 830 58
rect 860 16 875 58
<< nmoslvt >>
rect -199 -133 -184 -91
rect -152 -133 -137 -91
rect -52 -133 -37 -91
rect 0 -133 15 -91
rect 44 -133 59 -91
rect 88 -133 103 -91
rect 132 -133 147 -91
rect 477 -188 492 -146
rect 521 -188 536 -146
rect 622 -158 637 -116
rect 669 -158 684 -116
rect 770 -188 785 -146
rect 814 -188 829 -146
rect 633 -235 675 -220
<< ndiff >>
rect -228 -102 -199 -91
rect -228 -119 -222 -102
rect -205 -119 -199 -102
rect -228 -133 -199 -119
rect -184 -102 -152 -91
rect -184 -119 -175 -102
rect -158 -119 -152 -102
rect -184 -133 -152 -119
rect -137 -102 -110 -91
rect -137 -119 -131 -102
rect -114 -119 -110 -102
rect -137 -133 -110 -119
rect -79 -102 -52 -91
rect -79 -119 -75 -102
rect -58 -119 -52 -102
rect -79 -133 -52 -119
rect -37 -108 0 -91
rect -37 -125 -30 -108
rect -13 -125 0 -108
rect -37 -133 0 -125
rect 15 -102 44 -91
rect 15 -119 21 -102
rect 38 -119 44 -102
rect 15 -133 44 -119
rect 59 -102 88 -91
rect 59 -119 65 -102
rect 82 -119 88 -102
rect 59 -133 88 -119
rect 103 -102 132 -91
rect 103 -119 109 -102
rect 126 -119 132 -102
rect 103 -133 132 -119
rect 147 -102 177 -91
rect 147 -119 153 -102
rect 170 -119 177 -102
rect 147 -133 177 -119
rect 593 -127 622 -116
rect 593 -144 599 -127
rect 616 -144 622 -127
rect 450 -158 477 -146
rect 450 -175 454 -158
rect 471 -175 477 -158
rect 450 -188 477 -175
rect 492 -158 521 -146
rect 492 -175 498 -158
rect 515 -175 521 -158
rect 492 -188 521 -175
rect 536 -158 564 -146
rect 593 -158 622 -144
rect 637 -127 669 -116
rect 637 -144 646 -127
rect 663 -144 669 -127
rect 637 -158 669 -144
rect 684 -125 713 -116
rect 684 -142 690 -125
rect 707 -142 713 -125
rect 684 -158 713 -142
rect 742 -158 770 -146
rect 536 -175 542 -158
rect 559 -175 564 -158
rect 536 -188 564 -175
rect 742 -175 747 -158
rect 764 -175 770 -158
rect 742 -188 770 -175
rect 785 -158 814 -146
rect 785 -175 791 -158
rect 808 -175 814 -158
rect 785 -188 814 -175
rect 829 -158 856 -146
rect 829 -175 835 -158
rect 852 -175 856 -158
rect 829 -188 856 -175
rect 633 -197 675 -192
rect 633 -214 646 -197
rect 663 -214 675 -197
rect 633 -220 675 -214
rect 633 -241 675 -235
rect 633 -258 646 -241
rect 663 -258 675 -241
rect 633 -264 675 -258
<< pdiff >>
rect -173 48 -144 59
rect -173 31 -167 48
rect -150 31 -144 48
rect -173 17 -144 31
rect -129 48 -100 59
rect -129 31 -123 48
rect -106 31 -100 48
rect -129 17 -100 31
rect -85 48 -58 59
rect -85 31 -79 48
rect -62 31 -58 48
rect -85 17 -58 31
rect -27 48 0 59
rect -27 31 -23 48
rect -6 31 0 48
rect -27 17 0 31
rect 15 48 44 59
rect 15 31 21 48
rect 38 31 44 48
rect 15 17 44 31
rect 59 48 88 59
rect 59 31 65 48
rect 82 31 88 48
rect 59 17 88 31
rect 103 48 132 59
rect 103 31 109 48
rect 126 31 132 48
rect 103 17 132 31
rect 147 48 177 59
rect 147 31 153 48
rect 170 31 177 48
rect 147 17 177 31
rect 404 46 431 58
rect 404 29 408 46
rect 425 29 431 46
rect 404 16 431 29
rect 446 46 476 58
rect 446 29 453 46
rect 470 29 476 46
rect 446 16 476 29
rect 491 46 519 58
rect 491 29 498 46
rect 515 29 519 46
rect 491 16 519 29
rect 593 47 622 58
rect 593 30 599 47
rect 616 30 622 47
rect 593 16 622 30
rect 637 47 669 58
rect 637 30 644 47
rect 661 30 669 47
rect 637 16 669 30
rect 684 47 713 58
rect 684 30 690 47
rect 707 30 713 47
rect 684 16 713 30
rect 787 46 815 58
rect 787 29 791 46
rect 808 29 815 46
rect 787 16 815 29
rect 830 46 860 58
rect 830 29 836 46
rect 853 29 860 46
rect 830 16 860 29
rect 875 46 902 58
rect 875 29 881 46
rect 898 29 902 46
rect 875 16 902 29
<< ndiffc >>
rect -222 -119 -205 -102
rect -175 -119 -158 -102
rect -131 -119 -114 -102
rect -75 -119 -58 -102
rect -30 -125 -13 -108
rect 21 -119 38 -102
rect 65 -119 82 -102
rect 109 -119 126 -102
rect 153 -119 170 -102
rect 599 -144 616 -127
rect 454 -175 471 -158
rect 498 -175 515 -158
rect 646 -144 663 -127
rect 690 -142 707 -125
rect 542 -175 559 -158
rect 747 -175 764 -158
rect 791 -175 808 -158
rect 835 -175 852 -158
rect 646 -214 663 -197
rect 646 -258 663 -241
<< pdiffc >>
rect -167 31 -150 48
rect -123 31 -106 48
rect -79 31 -62 48
rect -23 31 -6 48
rect 21 31 38 48
rect 65 31 82 48
rect 109 31 126 48
rect 153 31 170 48
rect 408 29 425 46
rect 453 29 470 46
rect 498 29 515 46
rect 599 30 616 47
rect 644 30 661 47
rect 690 30 707 47
rect 791 29 808 46
rect 836 29 853 46
rect 881 29 898 46
<< psubdiff >>
rect 177 -103 208 -91
rect 177 -120 191 -103
rect 177 -133 208 -120
<< nsubdiff >>
rect 177 46 208 59
rect 177 29 191 46
rect 177 17 208 29
<< psubdiffcont >>
rect 191 -120 208 -103
<< nsubdiffcont >>
rect 191 29 208 46
<< poly >>
rect 21 115 54 123
rect -219 108 -186 110
rect -219 105 -35 108
rect -219 88 -211 105
rect -194 93 -35 105
rect 21 98 29 115
rect 46 113 54 115
rect 476 114 509 119
rect 46 98 147 113
rect 21 93 54 98
rect -194 88 -186 93
rect -219 83 -186 88
rect -144 59 -129 72
rect -100 59 -85 72
rect -144 7 -129 17
rect -100 7 -85 17
rect -144 -8 -85 7
rect -245 -17 -213 -8
rect -245 -34 -238 -17
rect -221 -34 -213 -17
rect -102 -30 -85 -8
rect -50 6 -35 93
rect 0 59 15 72
rect 44 59 59 72
rect 88 59 103 72
rect 132 59 147 98
rect 476 97 484 114
rect 501 97 509 114
rect 476 92 509 97
rect 797 114 830 119
rect 797 97 805 114
rect 822 97 830 114
rect 797 92 830 97
rect 431 58 446 71
rect 476 58 491 92
rect 622 58 637 71
rect 669 58 684 71
rect 815 58 830 92
rect 860 58 875 71
rect 0 6 15 17
rect -50 -9 15 6
rect -245 -42 -213 -34
rect -163 -35 -130 -30
rect -237 -65 -222 -42
rect -163 -52 -155 -35
rect -138 -52 -130 -35
rect -163 -57 -130 -52
rect -102 -35 -50 -30
rect -102 -52 -76 -35
rect -59 -52 -50 -35
rect 44 -39 59 17
rect 88 1 103 17
rect 132 4 147 17
rect 84 -7 111 1
rect 84 -24 89 -7
rect 106 -24 111 -7
rect 84 -32 111 -24
rect -102 -57 -50 -52
rect 36 -42 59 -39
rect 36 -50 63 -42
rect -237 -80 -184 -65
rect -199 -91 -184 -80
rect -152 -91 -137 -57
rect -199 -146 -184 -133
rect -152 -146 -137 -133
rect -102 -141 -87 -57
rect 36 -67 41 -50
rect 58 -67 63 -50
rect 36 -75 63 -67
rect -52 -91 -37 -78
rect 0 -91 15 -78
rect 44 -91 59 -75
rect 88 -91 103 -32
rect 152 -47 179 -39
rect 152 -57 157 -47
rect 132 -64 157 -57
rect 174 -64 179 -47
rect 132 -72 179 -64
rect 132 -91 147 -72
rect 431 -101 446 16
rect 476 3 491 16
rect 622 3 637 16
rect 669 3 684 16
rect 815 3 830 16
rect 622 -8 684 3
rect 622 -12 646 -8
rect 641 -25 646 -12
rect 663 -12 684 -8
rect 860 0 875 16
rect 860 -8 887 0
rect 663 -25 668 -12
rect 641 -33 668 -25
rect 860 -25 865 -8
rect 882 -25 887 -8
rect 860 -33 887 -25
rect 604 -60 637 -55
rect 604 -77 612 -60
rect 629 -77 637 -60
rect 604 -82 637 -77
rect 426 -106 456 -101
rect 423 -123 431 -106
rect 448 -123 456 -106
rect 622 -116 637 -82
rect 669 -60 702 -55
rect 669 -77 677 -60
rect 694 -77 702 -60
rect 669 -82 702 -77
rect 669 -116 684 -82
rect 426 -128 492 -123
rect -52 -141 -37 -133
rect -102 -156 -37 -141
rect 0 -167 15 -133
rect 44 -146 59 -133
rect 88 -146 103 -133
rect 132 -167 147 -133
rect 431 -138 492 -128
rect 477 -146 492 -138
rect 521 -146 536 -133
rect 0 -182 147 -167
rect 860 -123 875 -33
rect 770 -146 785 -133
rect 814 -138 875 -123
rect 814 -146 829 -138
rect 622 -171 637 -158
rect 669 -171 684 -158
rect 477 -201 492 -188
rect 521 -222 536 -188
rect 503 -230 536 -222
rect 503 -247 508 -230
rect 525 -247 536 -230
rect 588 -219 621 -214
rect 588 -236 596 -219
rect 613 -220 621 -219
rect 688 -219 721 -214
rect 688 -220 696 -219
rect 613 -235 633 -220
rect 675 -235 696 -220
rect 613 -236 621 -235
rect 588 -241 621 -236
rect 688 -236 696 -235
rect 713 -236 721 -219
rect 688 -241 721 -236
rect 770 -222 785 -188
rect 814 -201 829 -188
rect 770 -230 803 -222
rect 503 -255 536 -247
rect 770 -247 781 -230
rect 798 -247 803 -230
rect 770 -255 803 -247
<< polycont >>
rect -211 88 -194 105
rect 29 98 46 115
rect -238 -34 -221 -17
rect 484 97 501 114
rect 805 97 822 114
rect -155 -52 -138 -35
rect -76 -52 -59 -35
rect 89 -24 106 -7
rect 41 -67 58 -50
rect 157 -64 174 -47
rect 646 -25 663 -8
rect 865 -25 882 -8
rect 612 -77 629 -60
rect 431 -123 448 -106
rect 677 -77 694 -60
rect 508 -247 525 -230
rect 596 -236 613 -219
rect 696 -236 713 -219
rect 781 -247 798 -230
<< locali >>
rect -286 134 -268 151
rect -251 134 -232 151
rect -215 134 -196 151
rect -179 134 -160 151
rect -143 134 -124 151
rect -107 134 -88 151
rect -71 134 -52 151
rect -35 134 -16 151
rect 1 134 20 151
rect 37 134 56 151
rect 73 134 92 151
rect 109 134 128 151
rect 145 134 164 151
rect 181 134 200 151
rect 217 134 236 151
rect 253 134 268 151
rect 372 134 377 151
rect 394 134 425 151
rect 442 134 473 151
rect 490 134 521 151
rect 538 134 569 151
rect 586 134 617 151
rect 634 134 665 151
rect 682 134 713 151
rect 730 134 761 151
rect 778 134 809 151
rect 826 134 857 151
rect 874 134 905 151
rect 922 134 953 151
rect -219 105 -186 108
rect -219 88 -211 105
rect -194 88 -186 105
rect -219 85 -186 88
rect -215 40 -198 85
rect -123 56 -106 134
rect -75 115 54 117
rect -75 100 29 115
rect -75 56 -58 100
rect 21 98 29 100
rect 46 98 54 115
rect 21 90 54 98
rect 76 101 98 134
rect 76 90 93 101
rect 71 73 93 90
rect 71 56 88 73
rect -171 48 -146 56
rect -171 40 -167 48
rect -215 31 -167 40
rect -150 31 -146 48
rect -215 23 -146 31
rect -127 48 -102 56
rect -127 31 -123 48
rect -106 31 -102 48
rect -127 23 -102 31
rect -83 48 -58 56
rect -83 31 -79 48
rect -62 31 -58 48
rect -83 23 -58 31
rect -215 11 -182 23
rect -238 -17 -221 -8
rect -238 -43 -221 -34
rect -201 -60 -182 11
rect -75 6 -58 23
rect -119 -11 -58 6
rect -27 48 -2 56
rect -27 31 -23 48
rect -6 31 -2 48
rect -27 23 -2 31
rect 17 48 42 56
rect 17 31 21 48
rect 38 31 42 48
rect 17 23 42 31
rect 61 48 88 56
rect 61 31 65 48
rect 82 31 88 48
rect 61 23 88 31
rect 105 48 130 56
rect 105 31 109 48
rect 126 31 130 48
rect 105 23 130 31
rect 149 48 174 56
rect 149 31 153 48
rect 170 31 174 48
rect 149 23 174 31
rect 191 46 208 134
rect -27 -7 -10 23
rect 89 -7 106 1
rect 153 -2 170 23
rect 191 21 208 29
rect 408 46 425 134
rect 476 97 484 114
rect 501 97 595 114
rect 578 55 595 97
rect 643 55 662 134
rect 711 97 805 114
rect 822 97 830 114
rect 711 55 728 97
rect 408 21 425 29
rect 453 46 470 54
rect 453 21 470 29
rect 498 46 515 54
rect -155 -35 -138 -27
rect -155 -60 -138 -52
rect -218 -77 -182 -60
rect -119 -77 -102 -11
rect -27 -24 89 -7
rect -84 -52 -76 -35
rect -59 -52 -51 -35
rect -218 -94 -201 -77
rect -127 -94 -102 -77
rect 7 -94 24 -24
rect 89 -32 106 -24
rect 123 -19 170 -2
rect 498 -7 515 29
rect 41 -50 58 -42
rect 123 -50 140 -19
rect 58 -67 140 -50
rect 41 -75 58 -67
rect 110 -74 140 -67
rect 157 -47 174 -39
rect 157 -72 174 -64
rect 110 -94 127 -74
rect -226 -102 -201 -94
rect -226 -119 -222 -102
rect -205 -119 -201 -102
rect -226 -127 -201 -119
rect -179 -102 -154 -94
rect -179 -119 -175 -102
rect -158 -119 -154 -102
rect -179 -127 -154 -119
rect -135 -102 -110 -94
rect -135 -119 -131 -102
rect -114 -119 -110 -102
rect -135 -127 -110 -119
rect -78 -102 -54 -94
rect -78 -119 -75 -102
rect -58 -119 -54 -102
rect -78 -127 -54 -119
rect -33 -108 -10 -100
rect -33 -125 -30 -108
rect -13 -125 -10 -108
rect 7 -102 42 -94
rect 7 -111 21 -102
rect -174 -145 -157 -127
rect -78 -145 -61 -127
rect -33 -133 -10 -125
rect 17 -119 21 -111
rect 38 -119 42 -102
rect 17 -127 42 -119
rect 61 -102 86 -94
rect 61 -119 65 -102
rect 82 -119 86 -102
rect 61 -127 86 -119
rect 105 -102 130 -94
rect 105 -119 109 -102
rect 126 -119 130 -102
rect 105 -127 130 -119
rect 149 -102 174 -94
rect 149 -119 153 -102
rect 170 -119 174 -102
rect 149 -127 174 -119
rect 191 -103 208 -94
rect -174 -162 -61 -145
rect -27 -182 -10 -133
rect 66 -182 83 -127
rect 154 -182 171 -127
rect 191 -182 208 -120
rect 423 -123 431 -106
rect 448 -123 456 -106
rect 454 -158 471 -150
rect -286 -199 -196 -182
rect -179 -199 -160 -182
rect -143 -199 -124 -182
rect -107 -199 -88 -182
rect -71 -199 -52 -182
rect -35 -199 -16 -182
rect 1 -199 20 -182
rect 37 -199 56 -182
rect 73 -199 92 -182
rect 109 -199 128 -182
rect 145 -199 164 -182
rect 181 -199 200 -182
rect 217 -199 236 -182
rect 253 -199 268 -182
rect 454 -282 471 -175
rect 498 -158 515 -24
rect 578 47 620 55
rect 578 30 599 47
rect 616 30 620 47
rect 578 22 620 30
rect 640 47 665 55
rect 640 30 644 47
rect 661 30 665 47
rect 640 22 665 30
rect 686 47 728 55
rect 686 30 690 47
rect 707 30 728 47
rect 686 22 728 30
rect 578 -119 595 22
rect 638 -25 646 -8
rect 663 -25 671 -8
rect 612 -60 629 -52
rect 612 -85 629 -77
rect 677 -60 694 -52
rect 677 -85 694 -77
rect 711 -117 728 22
rect 578 -127 620 -119
rect 578 -144 599 -127
rect 616 -144 620 -127
rect 498 -183 515 -175
rect 542 -158 559 -149
rect 578 -152 620 -144
rect 642 -127 667 -119
rect 642 -144 646 -127
rect 663 -144 667 -127
rect 642 -152 667 -144
rect 686 -125 728 -117
rect 686 -142 690 -125
rect 707 -142 728 -125
rect 686 -151 728 -142
rect 791 46 808 54
rect 791 -106 808 29
rect 836 46 853 54
rect 836 21 853 29
rect 881 46 898 134
rect 881 21 898 29
rect 857 -25 865 -8
rect 882 -25 890 -8
rect 508 -229 525 -222
rect 508 -255 525 -247
rect 542 -282 559 -175
rect 646 -197 663 -152
rect 747 -158 764 -149
rect 596 -219 613 -211
rect 638 -214 646 -197
rect 663 -214 672 -197
rect 596 -244 613 -236
rect 696 -219 713 -211
rect 638 -258 646 -241
rect 663 -258 671 -241
rect 696 -244 713 -236
rect 646 -282 663 -258
rect 747 -282 764 -175
rect 791 -158 808 -123
rect 791 -183 808 -175
rect 835 -158 852 -150
rect 781 -229 798 -222
rect 781 -255 798 -247
rect 835 -282 852 -175
rect 372 -299 377 -282
rect 394 -299 425 -282
rect 442 -299 473 -282
rect 490 -299 521 -282
rect 538 -299 569 -282
rect 586 -299 617 -282
rect 634 -299 665 -282
rect 682 -299 713 -282
rect 730 -299 761 -282
rect 778 -299 809 -282
rect 826 -299 857 -282
rect 874 -299 905 -282
rect 922 -299 953 -282
<< viali >>
rect -268 134 -251 151
rect -232 134 -215 151
rect -196 134 -179 151
rect -160 134 -143 151
rect -124 134 -107 151
rect -88 134 -71 151
rect -52 134 -35 151
rect -16 134 1 151
rect 20 134 37 151
rect 56 134 73 151
rect 92 134 109 151
rect 128 134 145 151
rect 164 134 181 151
rect 200 134 217 151
rect 236 134 253 151
rect 377 134 394 151
rect 425 134 442 151
rect 473 134 490 151
rect 521 134 538 151
rect 569 134 586 151
rect 617 134 634 151
rect 665 134 682 151
rect 713 134 730 151
rect 761 134 778 151
rect 809 134 826 151
rect 857 134 874 151
rect 905 134 922 151
rect 498 -24 515 -7
rect 431 -123 448 -106
rect -196 -199 -179 -182
rect -160 -199 -143 -182
rect -124 -199 -107 -182
rect -88 -199 -71 -182
rect -52 -199 -35 -182
rect -16 -199 1 -182
rect 20 -199 37 -182
rect 56 -199 73 -182
rect 92 -199 109 -182
rect 128 -199 145 -182
rect 164 -199 181 -182
rect 200 -199 217 -182
rect 236 -199 253 -182
rect 646 -25 663 -8
rect 865 -25 882 -8
rect 791 -123 808 -106
rect 508 -230 525 -229
rect 508 -246 525 -230
rect 596 -236 613 -219
rect 696 -236 713 -219
rect 781 -230 798 -229
rect 781 -246 798 -230
rect 377 -299 394 -282
rect 425 -299 442 -282
rect 473 -299 490 -282
rect 521 -299 538 -282
rect 569 -299 586 -282
rect 617 -299 634 -282
rect 665 -299 682 -282
rect 713 -299 730 -282
rect 761 -299 778 -282
rect 809 -299 826 -282
rect 857 -299 874 -282
rect 905 -299 922 -282
<< metal1 >>
rect -286 151 268 167
rect -286 134 -268 151
rect -251 134 -232 151
rect -215 134 -196 151
rect -179 134 -160 151
rect -143 134 -124 151
rect -107 134 -88 151
rect -71 134 -52 151
rect -35 134 -16 151
rect 1 134 20 151
rect 37 134 56 151
rect 73 134 92 151
rect 109 134 128 151
rect 145 134 164 151
rect 181 134 200 151
rect 217 134 236 151
rect 253 134 268 151
rect -286 118 268 134
rect 372 151 953 167
rect 372 134 377 151
rect 394 134 425 151
rect 442 134 473 151
rect 490 134 521 151
rect 538 134 569 151
rect 586 134 617 151
rect 634 134 665 151
rect 682 134 713 151
rect 730 134 761 151
rect 778 134 809 151
rect 826 134 857 151
rect 874 134 905 151
rect 922 134 953 151
rect 372 118 953 134
rect 609 14 882 31
rect 492 -7 521 -1
rect 609 -7 626 14
rect 492 -24 498 -7
rect 515 -24 626 -7
rect 642 -3 668 0
rect 865 -5 882 14
rect 492 -30 521 -24
rect 642 -32 668 -29
rect 861 -8 885 -5
rect 861 -25 865 -8
rect 882 -25 885 -8
rect 861 -31 885 -25
rect 425 -106 455 -102
rect 788 -106 814 -100
rect 425 -123 431 -106
rect 448 -123 791 -106
rect 808 -123 814 -106
rect 425 -128 455 -123
rect 788 -130 814 -123
rect -286 -182 268 -166
rect -286 -199 -196 -182
rect -179 -199 -160 -182
rect -143 -199 -124 -182
rect -107 -199 -88 -182
rect -71 -199 -52 -182
rect -35 -199 -16 -182
rect 1 -199 20 -182
rect 37 -199 56 -182
rect 73 -199 92 -182
rect 109 -199 128 -182
rect 145 -199 164 -182
rect 181 -199 200 -182
rect 217 -199 236 -182
rect 253 -199 268 -182
rect -286 -215 268 -199
rect 508 -175 798 -158
rect 508 -226 525 -175
rect 590 -219 616 -216
rect 638 -219 641 -215
rect 503 -229 530 -226
rect 503 -246 508 -229
rect 525 -246 530 -229
rect 590 -236 596 -219
rect 613 -236 641 -219
rect 590 -239 616 -236
rect 638 -241 641 -236
rect 667 -219 670 -215
rect 693 -219 719 -216
rect 667 -236 696 -219
rect 713 -236 719 -219
rect 781 -225 798 -175
rect 667 -241 670 -236
rect 693 -239 719 -236
rect 775 -229 804 -225
rect 503 -252 530 -246
rect 775 -246 781 -229
rect 798 -246 804 -229
rect 775 -252 804 -246
rect 372 -282 953 -266
rect 372 -299 377 -282
rect 394 -299 425 -282
rect 442 -299 473 -282
rect 490 -299 521 -282
rect 538 -299 569 -282
rect 586 -299 617 -282
rect 634 -299 665 -282
rect 682 -299 713 -282
rect 730 -299 761 -282
rect 778 -299 809 -282
rect 826 -299 857 -282
rect 874 -299 905 -282
rect 922 -299 953 -282
rect 372 -315 953 -299
<< via1 >>
rect 642 -8 668 -3
rect 642 -25 646 -8
rect 646 -25 663 -8
rect 663 -25 668 -8
rect 642 -29 668 -25
rect 641 -241 667 -215
<< metal2 >>
rect 642 -3 668 0
rect 642 -32 668 -29
rect 646 -215 663 -32
rect 638 -241 641 -215
rect 667 -241 670 -215
<< labels >>
rlabel locali 728 -97 728 -97 3 FN
rlabel locali 578 -94 578 -94 7 FP
flabel polycont 612 -77 629 -60 0 FreeSans 80 0 0 0 inp
flabel polycont 677 -77 694 -60 0 FreeSans 80 0 0 0 inm
flabel metal2 646 -25 663 -8 0 FreeSans 80 0 0 0 phi1
rlabel locali 515 -130 515 -130 3 high
rlabel locali 791 -125 791 -125 7 low
rlabel locali 461 21 461 21 5 pfetw
rlabel locali 845 21 845 21 5 pfete
flabel metal1 508 -246 525 -229 0 FreeSans 80 0 0 0 phi1b
flabel metal1 781 -246 798 -229 0 FreeSans 80 0 0 0 phi1b
flabel viali 498 -24 515 -7 0 FreeSans 80 0 0 0 high
flabel viali 791 -123 808 -106 0 FreeSans 80 0 0 0 low
rlabel locali -102 -51 -102 -51 3 FN
rlabel locali -104 -145 -104 -145 1 tail
rlabel locali 165 -39 165 -39 1 phi1b
rlabel locali 30 -94 30 -94 1 high
rlabel locali 118 -94 118 -94 1 low
rlabel locali 30 56 30 56 1 pfetw
rlabel locali 118 56 118 56 1 pfete
rlabel locali -51 -44 -51 -44 3 phi1
flabel polycont -76 -52 -59 -35 0 FreeSans 56 0 0 0 phi1
flabel polycont 157 -64 174 -47 0 FreeSans 56 0 0 0 phi1b
flabel polycont 41 -67 58 -50 0 FreeSans 56 0 0 0 low
flabel polycont 89 -24 106 -7 0 FreeSans 56 0 0 0 high
flabel polycont -238 -34 -221 -17 0 FreeSans 56 0 0 0 inp
flabel polycont -155 -52 -138 -35 0 FreeSans 56 0 0 0 inm
rlabel locali -229 -8 -229 -8 1 inp
rlabel locali -147 -27 -147 -27 1 inm
rlabel locali 268 142 268 142 3 VDD
rlabel locali 268 -189 268 -189 3 GND
rlabel locali -198 -54 -198 -54 3 FP
<< end >>
