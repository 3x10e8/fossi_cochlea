magic
tech sky130A
magscale 1 2
timestamp 1654749026
<< obsli1 >>
rect 1104 2159 96876 77809
<< obsm1 >>
rect 1104 2128 97230 78736
<< metal2 >>
rect 2686 79200 2742 80000
rect 8114 79200 8170 80000
rect 13542 79200 13598 80000
rect 18970 79200 19026 80000
rect 24398 79200 24454 80000
rect 29826 79200 29882 80000
rect 35346 79200 35402 80000
rect 40774 79200 40830 80000
rect 46202 79200 46258 80000
rect 51630 79200 51686 80000
rect 57058 79200 57114 80000
rect 62486 79200 62542 80000
rect 68006 79200 68062 80000
rect 73434 79200 73490 80000
rect 78862 79200 78918 80000
rect 84290 79200 84346 80000
rect 89718 79200 89774 80000
rect 95146 79200 95202 80000
rect 7010 0 7066 800
rect 20994 0 21050 800
rect 34978 0 35034 800
rect 48962 0 49018 800
rect 62946 0 63002 800
rect 76930 0 76986 800
rect 90914 0 90970 800
<< obsm2 >>
rect 1398 79144 2630 79393
rect 2798 79144 8058 79393
rect 8226 79144 13486 79393
rect 13654 79144 18914 79393
rect 19082 79144 24342 79393
rect 24510 79144 29770 79393
rect 29938 79144 35290 79393
rect 35458 79144 40718 79393
rect 40886 79144 46146 79393
rect 46314 79144 51574 79393
rect 51742 79144 57002 79393
rect 57170 79144 62430 79393
rect 62598 79144 67950 79393
rect 68118 79144 73378 79393
rect 73546 79144 78806 79393
rect 78974 79144 84234 79393
rect 84402 79144 89662 79393
rect 89830 79144 95090 79393
rect 95258 79144 97224 79393
rect 1398 856 97224 79144
rect 1398 734 6954 856
rect 7122 734 20938 856
rect 21106 734 34922 856
rect 35090 734 48906 856
rect 49074 734 62890 856
rect 63058 734 76874 856
rect 77042 734 90858 856
rect 91026 734 97224 856
<< metal3 >>
rect 0 77528 800 77648
rect 97200 77664 98000 77784
rect 97200 73176 98000 73296
rect 0 72768 800 72888
rect 97200 68824 98000 68944
rect 0 68144 800 68264
rect 97200 64336 98000 64456
rect 0 63384 800 63504
rect 97200 59848 98000 59968
rect 0 58760 800 58880
rect 97200 55496 98000 55616
rect 0 54000 800 54120
rect 97200 51008 98000 51128
rect 0 49240 800 49360
rect 97200 46520 98000 46640
rect 0 44616 800 44736
rect 97200 42168 98000 42288
rect 0 39856 800 39976
rect 97200 37680 98000 37800
rect 0 35232 800 35352
rect 97200 33192 98000 33312
rect 0 30472 800 30592
rect 97200 28840 98000 28960
rect 0 25712 800 25832
rect 97200 24352 98000 24472
rect 0 21088 800 21208
rect 97200 19864 98000 19984
rect 0 16328 800 16448
rect 97200 15512 98000 15632
rect 0 11704 800 11824
rect 97200 11024 98000 11144
rect 0 6944 800 7064
rect 97200 6536 98000 6656
rect 0 2320 800 2440
rect 97200 2184 98000 2304
<< obsm3 >>
rect 800 77864 97200 79389
rect 800 77728 97120 77864
rect 880 77584 97120 77728
rect 880 77448 97200 77584
rect 800 73376 97200 77448
rect 800 73096 97120 73376
rect 800 72968 97200 73096
rect 880 72688 97200 72968
rect 800 69024 97200 72688
rect 800 68744 97120 69024
rect 800 68344 97200 68744
rect 880 68064 97200 68344
rect 800 64536 97200 68064
rect 800 64256 97120 64536
rect 800 63584 97200 64256
rect 880 63304 97200 63584
rect 800 60048 97200 63304
rect 800 59768 97120 60048
rect 800 58960 97200 59768
rect 880 58680 97200 58960
rect 800 55696 97200 58680
rect 800 55416 97120 55696
rect 800 54200 97200 55416
rect 880 53920 97200 54200
rect 800 51208 97200 53920
rect 800 50928 97120 51208
rect 800 49440 97200 50928
rect 880 49160 97200 49440
rect 800 46720 97200 49160
rect 800 46440 97120 46720
rect 800 44816 97200 46440
rect 880 44536 97200 44816
rect 800 42368 97200 44536
rect 800 42088 97120 42368
rect 800 40056 97200 42088
rect 880 39776 97200 40056
rect 800 37880 97200 39776
rect 800 37600 97120 37880
rect 800 35432 97200 37600
rect 880 35152 97200 35432
rect 800 33392 97200 35152
rect 800 33112 97120 33392
rect 800 30672 97200 33112
rect 880 30392 97200 30672
rect 800 29040 97200 30392
rect 800 28760 97120 29040
rect 800 25912 97200 28760
rect 880 25632 97200 25912
rect 800 24552 97200 25632
rect 800 24272 97120 24552
rect 800 21288 97200 24272
rect 880 21008 97200 21288
rect 800 20064 97200 21008
rect 800 19784 97120 20064
rect 800 16528 97200 19784
rect 880 16248 97200 16528
rect 800 15712 97200 16248
rect 800 15432 97120 15712
rect 800 11904 97200 15432
rect 880 11624 97200 11904
rect 800 11224 97200 11624
rect 800 10944 97120 11224
rect 800 7144 97200 10944
rect 880 6864 97200 7144
rect 800 6736 97200 6864
rect 800 6456 97120 6736
rect 800 2520 97200 6456
rect 880 2384 97200 2520
rect 880 2240 97120 2384
rect 800 2143 97120 2240
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
rect 65648 2128 65968 77840
rect 81008 2128 81328 77840
rect 96368 2128 96688 77840
<< obsm4 >>
rect 13675 77920 93965 79389
rect 13675 13227 19488 77920
rect 19968 13227 34848 77920
rect 35328 13227 50208 77920
rect 50688 13227 65568 77920
rect 66048 13227 80928 77920
rect 81408 13227 93965 77920
<< labels >>
rlabel metal3 s 0 25712 800 25832 6 cclk_I[0]
port 1 nsew signal output
rlabel metal3 s 0 58760 800 58880 6 cclk_I[1]
port 2 nsew signal output
rlabel metal3 s 97200 6536 98000 6656 6 cclk_Q[0]
port 3 nsew signal output
rlabel metal3 s 97200 37680 98000 37800 6 cclk_Q[1]
port 4 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 clk_master
port 5 nsew signal input
rlabel metal2 s 8114 79200 8170 80000 6 clk_master_out
port 6 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 clkdiv2_I[0]
port 7 nsew signal output
rlabel metal3 s 0 54000 800 54120 6 clkdiv2_I[1]
port 8 nsew signal output
rlabel metal3 s 97200 11024 98000 11144 6 clkdiv2_Q[0]
port 9 nsew signal output
rlabel metal3 s 97200 42168 98000 42288 6 clkdiv2_Q[1]
port 10 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 comp_high_I[0]
port 11 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 comp_high_I[1]
port 12 nsew signal input
rlabel metal3 s 97200 15512 98000 15632 6 comp_high_Q[0]
port 13 nsew signal input
rlabel metal3 s 97200 46520 98000 46640 6 comp_high_Q[1]
port 14 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 cos_out[0]
port 15 nsew signal output
rlabel metal3 s 0 63384 800 63504 6 cos_out[1]
port 16 nsew signal output
rlabel metal3 s 0 2320 800 2440 6 cos_outb[0]
port 17 nsew signal output
rlabel metal3 s 0 35232 800 35352 6 cos_outb[1]
port 18 nsew signal output
rlabel metal2 s 18970 79200 19026 80000 6 div2out
port 19 nsew signal output
rlabel metal3 s 0 6944 800 7064 6 fb1_I[0]
port 20 nsew signal output
rlabel metal3 s 0 39856 800 39976 6 fb1_I[1]
port 21 nsew signal output
rlabel metal3 s 97200 24352 98000 24472 6 fb1_Q[0]
port 22 nsew signal output
rlabel metal3 s 97200 55496 98000 55616 6 fb1_Q[1]
port 23 nsew signal output
rlabel metal2 s 95146 79200 95202 80000 6 fb2_I[0]
port 24 nsew signal output
rlabel metal3 s 97200 77664 98000 77784 6 fb2_I[1]
port 25 nsew signal output
rlabel metal3 s 97200 73176 98000 73296 6 fb2_Q[0]
port 26 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 fb2_Q[1]
port 27 nsew signal output
rlabel metal2 s 73434 79200 73490 80000 6 gray_clk_out[10]
port 28 nsew signal output
rlabel metal2 s 24398 79200 24454 80000 6 gray_clk_out[1]
port 29 nsew signal output
rlabel metal2 s 29826 79200 29882 80000 6 gray_clk_out[2]
port 30 nsew signal output
rlabel metal2 s 35346 79200 35402 80000 6 gray_clk_out[3]
port 31 nsew signal output
rlabel metal2 s 40774 79200 40830 80000 6 gray_clk_out[4]
port 32 nsew signal output
rlabel metal2 s 46202 79200 46258 80000 6 gray_clk_out[5]
port 33 nsew signal output
rlabel metal2 s 51630 79200 51686 80000 6 gray_clk_out[6]
port 34 nsew signal output
rlabel metal2 s 57058 79200 57114 80000 6 gray_clk_out[7]
port 35 nsew signal output
rlabel metal2 s 62486 79200 62542 80000 6 gray_clk_out[8]
port 36 nsew signal output
rlabel metal2 s 68006 79200 68062 80000 6 gray_clk_out[9]
port 37 nsew signal output
rlabel metal2 s 78862 79200 78918 80000 6 no_ones_below_out[0]
port 38 nsew signal output
rlabel metal2 s 84290 79200 84346 80000 6 no_ones_below_out[1]
port 39 nsew signal output
rlabel metal2 s 89718 79200 89774 80000 6 no_ones_below_out[2]
port 40 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 phi1b_dig_I[0]
port 41 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 phi1b_dig_I[1]
port 42 nsew signal input
rlabel metal3 s 97200 19864 98000 19984 6 phi1b_dig_Q[0]
port 43 nsew signal input
rlabel metal3 s 97200 51008 98000 51128 6 phi1b_dig_Q[1]
port 44 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 read_out_I[0]
port 45 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 read_out_I[1]
port 46 nsew signal output
rlabel metal3 s 0 68144 800 68264 6 read_out_I_top[0]
port 47 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 read_out_I_top[1]
port 48 nsew signal output
rlabel metal2 s 90914 0 90970 800 6 read_out_Q[0]
port 49 nsew signal output
rlabel metal2 s 76930 0 76986 800 6 read_out_Q[1]
port 50 nsew signal output
rlabel metal3 s 97200 64336 98000 64456 6 read_out_Q_top[0]
port 51 nsew signal output
rlabel metal3 s 97200 68824 98000 68944 6 read_out_Q_top[1]
port 52 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 rstb
port 53 nsew signal input
rlabel metal2 s 2686 79200 2742 80000 6 rstb_out
port 54 nsew signal output
rlabel metal3 s 97200 2184 98000 2304 6 sin_out[0]
port 55 nsew signal output
rlabel metal3 s 97200 33192 98000 33312 6 sin_out[1]
port 56 nsew signal output
rlabel metal3 s 97200 28840 98000 28960 6 sin_outb[0]
port 57 nsew signal output
rlabel metal3 s 97200 59848 98000 59968 6 sin_outb[1]
port 58 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 ud_en
port 59 nsew signal input
rlabel metal2 s 13542 79200 13598 80000 6 ud_en_out
port 60 nsew signal output
rlabel metal4 s 4208 2128 4528 77840 6 vccd1
port 61 nsew power input
rlabel metal4 s 34928 2128 35248 77840 6 vccd1
port 61 nsew power input
rlabel metal4 s 65648 2128 65968 77840 6 vccd1
port 61 nsew power input
rlabel metal4 s 96368 2128 96688 77840 6 vccd1
port 61 nsew power input
rlabel metal4 s 19568 2128 19888 77840 6 vssd1
port 62 nsew ground input
rlabel metal4 s 50288 2128 50608 77840 6 vssd1
port 62 nsew ground input
rlabel metal4 s 81008 2128 81328 77840 6 vssd1
port 62 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 98000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9269336
string GDS_FILE /Volumes/export/isn/abhinav/fossi_cochlea/openlane/first_dual_core/runs/first_dual_core/results/finishing/first_dual_core.magic.gds
string GDS_START 447134
<< end >>

