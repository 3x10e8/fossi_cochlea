magic
tech sky130A
timestamp 1654156239
<< metal3 >>
rect 56 1011 216 1046
rect 412 1011 572 1046
rect 762 1011 922 1046
rect -22 927 1006 1011
rect -57 767 1041 927
rect -22 577 1006 767
rect -57 417 1041 577
rect -22 221 1006 417
rect -57 61 1041 221
rect -22 -17 1006 61
rect 56 -52 216 -17
rect 412 -52 572 -17
rect 762 -52 922 -17
<< mimcap >>
rect -8 897 992 997
rect -8 97 92 897
rect 193 547 441 797
rect 542 547 791 797
rect 193 197 441 447
rect 542 197 791 447
rect 892 97 992 897
rect -8 -3 992 97
<< mimcapcontact >>
rect 92 797 892 897
rect 92 547 193 797
rect 441 547 542 797
rect 791 547 892 797
rect 92 447 892 547
rect 92 197 193 447
rect 441 197 542 447
rect 791 197 892 447
rect 92 97 892 197
<< metal4 >>
rect 56 1011 216 1046
rect 412 1011 572 1046
rect 762 1011 922 1046
rect -22 927 1006 1011
rect -57 897 1041 927
rect -57 767 92 897
rect -22 577 92 767
rect -57 417 92 577
rect 193 547 441 797
rect 542 547 791 797
rect 892 767 1041 897
rect 892 577 1006 767
rect -22 221 92 417
rect -57 97 92 221
rect 193 197 441 447
rect 542 197 791 447
rect 892 417 1041 577
rect 892 221 1006 417
rect 892 97 1041 221
rect -57 61 1041 97
rect -22 -17 1006 61
rect 56 -52 216 -17
rect 412 -52 572 -17
rect 762 -52 922 -17
<< mimcap2 >>
rect -8 906 992 997
rect -8 88 83 906
rect 201 556 433 788
rect 551 556 783 788
rect 201 206 433 438
rect 551 206 783 438
rect 901 88 992 906
rect -8 -3 992 88
<< mimcap2contact >>
rect 83 788 901 906
rect 83 556 201 788
rect 433 556 551 788
rect 783 556 901 788
rect 83 438 901 556
rect 83 206 201 438
rect 433 206 551 438
rect 783 206 901 438
rect 83 88 901 206
<< metal5 >>
rect 56 927 216 1046
rect 412 927 572 1046
rect 762 927 922 1046
rect -57 906 1041 927
rect -57 767 83 906
rect 56 577 83 767
rect -57 417 83 577
rect 201 767 433 788
rect 201 577 216 767
rect 412 577 433 767
rect 201 556 433 577
rect 551 767 783 788
rect 551 577 572 767
rect 762 577 783 767
rect 551 556 783 577
rect 901 767 1041 906
rect 901 577 922 767
rect 56 221 83 417
rect -57 88 83 221
rect 201 417 433 438
rect 201 221 216 417
rect 412 221 433 417
rect 201 206 433 221
rect 551 417 783 438
rect 551 221 572 417
rect 762 221 783 417
rect 551 206 783 221
rect 901 417 1041 577
rect 901 221 922 417
rect 901 88 1041 221
rect -57 61 1041 88
rect 56 -52 216 61
rect 412 -52 572 61
rect 762 -52 922 61
<< end >>
