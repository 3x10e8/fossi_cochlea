magic
tech sky130A
timestamp 1654307754
use cap_10_10__side_x2  cap_10_10__side_x2_0
array 0 0 1397 0 5 -1742
timestamp 1654307754
transform 0 -1 1368 1 0 34
box -34 -374 1363 1368
use cap_10_10__side_x2  cap_10_10__side_x2_1
array 0 0 1397 0 5 -1742
timestamp 1654307754
transform 0 1 9084 -1 0 2760
box -34 -374 1363 1368
use cap_10_10_edge_x2  cap_10_10_edge_x2_0
timestamp 1654307754
transform 1 0 -1363 0 1 29
box -34 -29 1363 1368
use cap_10_10_edge_x2  cap_10_10_edge_x2_1
timestamp 1654307754
transform 0 1 -1368 -1 0 2760
box -34 -29 1363 1368
use cap_10_10_edge_x2  cap_10_10_edge_x2_2
timestamp 1654307754
transform -1 0 11815 0 -1 2765
box -34 -29 1363 1368
use cap_10_10_edge_x2  cap_10_10_edge_x2_3
timestamp 1654307754
transform 0 -1 11820 1 0 34
box -34 -29 1363 1368
<< end >>
