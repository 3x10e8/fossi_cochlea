** sch_path:
*+ /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/archive/mux/multiplier_differential.sch
**.subckt multiplier_differential inp inm outp outm ctrl ctrlbar vdda vssa
*.ipin inp
*.ipin inm
*.opin outp
*.opin outm
*.ipin ctrl
*.ipin ctrlbar
*.ipin vdda
*.ipin vssa
x1 inm inp ctrlbar ctrl outp vssa vdda analogMux
x2 inp inm ctrlbar ctrl outm vssa vdda analogMux
**.ends

* expanding   symbol:  mux/analogMux.sym # of pins=7
** sym_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/mux/analogMux.sym
** sch_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/mux/analogMux.sch
.subckt analogMux  vref2 vref1 c cbar out vssa vdda
*.ipin vref1
*.opin out
*.ipin vref2
*.ipin c
*.ipin cbar
*.ipin vssa
*.ipin vdda
XM2 vref1 c out vssa sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 vref1 cbar out vdda sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 out cbar vref2 vssa sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 out c vref2 vdda sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
