magic
tech sky130A
magscale 1 2
timestamp 1654748254
<< locali >>
rect 22218 28813 22252 29386
rect 25824 28777 25858 29363
<< viali >>
rect 22218 29386 22252 29420
<< metal1 >>
rect 24646 34222 24698 34228
rect 23265 34172 24646 34216
rect 24646 34164 24698 34170
rect 24403 33734 24455 33740
rect 23252 33685 24403 33729
rect 24403 33676 24455 33682
rect 24210 33113 24262 33119
rect 23256 33065 24210 33109
rect 24210 33055 24262 33061
rect 23757 32641 23810 32647
rect 23250 32597 23757 32641
rect 23757 32583 23810 32589
rect 23593 32016 23646 32022
rect 23229 31959 23593 32016
rect 23645 31959 23646 32016
rect 23593 31953 23646 31959
rect 23225 31614 23277 31620
rect 23225 31447 23277 31453
rect 13786 30310 22323 30350
rect 25813 30311 25866 30350
rect 25881 30311 34418 30350
rect 25884 30310 34418 30311
rect 13796 30190 22333 30230
rect 22335 30190 22387 30230
rect 25686 30190 25738 30230
rect 25744 30190 34281 30230
rect 24402 30120 24456 30126
rect 24402 30068 24403 30120
rect 24455 30068 24456 30120
rect 24402 30062 24456 30068
rect 24645 29997 24697 30003
rect 24645 29939 24697 29945
rect 23758 29880 23810 29886
rect 23758 29822 23810 29828
rect 24209 29756 24261 29762
rect 24209 29698 24261 29704
rect 23593 28713 23645 28719
rect 22201 28666 23593 28711
rect 23645 28666 25876 28711
rect 23593 28654 23645 28661
rect 23224 28544 23276 28550
rect 22279 28496 23224 28541
rect 23276 28496 25793 28541
rect 23224 28486 23276 28492
rect 24645 28453 24697 28459
rect 23390 28447 23442 28453
rect 22206 28406 23390 28440
rect 23442 28406 24645 28440
rect 24697 28406 25871 28440
rect 24645 28395 24697 28401
rect 23390 28389 23442 28395
<< via1 >>
rect 24646 34170 24698 34222
rect 24403 33682 24455 33734
rect 24210 33061 24262 33113
rect 23757 32589 23810 32641
rect 23593 31959 23645 32016
rect 23225 31453 23277 31614
rect 24403 30068 24455 30120
rect 24645 29945 24697 29997
rect 23758 29828 23810 29880
rect 24209 29704 24261 29756
rect 23593 28661 23645 28713
rect 23224 28492 23276 28544
rect 23390 28395 23442 28447
rect 24645 28401 24697 28453
rect 24018 26706 24070 26758
<< metal2 >>
rect 24646 34222 24698 34228
rect 24646 34164 24698 34170
rect 24403 33734 24455 33740
rect 24403 33676 24455 33682
rect 24210 33113 24262 33119
rect 24210 33055 24262 33061
rect 23757 32641 23810 32647
rect 23757 32583 23810 32589
rect 23593 32016 23646 32022
rect 23645 31959 23646 32016
rect 23593 31953 23646 31959
rect 23225 31614 23277 31620
rect 23225 31447 23277 31453
rect 21701 30758 21757 30767
rect 21701 30693 21757 30702
rect 21714 30481 21748 30693
rect 22096 30579 22130 30580
rect 22085 30570 22141 30579
rect 22085 30505 22141 30514
rect 21713 28443 21749 30481
rect 21713 28405 21922 28443
rect 22095 28442 22131 30505
rect 22202 28666 22240 28717
rect 23227 28551 23275 31447
rect 23594 28719 23644 31953
rect 23758 29880 23810 32583
rect 23758 29809 23810 29828
rect 24009 30958 24080 30970
rect 24009 30902 24017 30958
rect 24073 30902 24080 30958
rect 23593 28713 23645 28719
rect 23593 28654 23645 28661
rect 23224 28544 23276 28551
rect 23224 28486 23276 28492
rect 23390 28447 23442 28453
rect 23390 28389 23442 28395
rect 23400 26902 23434 28389
rect 24009 26758 24080 30902
rect 24211 29762 24260 33055
rect 24404 30126 24454 33676
rect 24402 30120 24456 30126
rect 24402 30068 24403 30120
rect 24455 30068 24456 30120
rect 24402 30062 24456 30068
rect 24404 30060 24454 30062
rect 24647 30003 24696 34164
rect 25935 30765 25991 30774
rect 25935 30700 25991 30709
rect 24645 29997 24697 30003
rect 24645 29939 24697 29945
rect 24647 29925 24696 29939
rect 24209 29756 24261 29762
rect 24209 29698 24261 29704
rect 25820 28683 25861 28717
rect 24645 28453 24697 28459
rect 25946 28432 25980 30700
rect 26315 30568 26371 30578
rect 26315 30503 26371 30512
rect 26328 28440 26362 30503
rect 26152 28403 26362 28440
rect 24645 28395 24697 28401
rect 24656 26902 24690 28395
rect 24009 26706 24018 26758
rect 24070 26706 24080 26758
rect 24009 26700 24080 26706
rect 46310 26270 47033 26314
rect 46310 26064 46355 26270
rect 1063 26007 1751 26051
<< via2 >>
rect 21701 30702 21757 30758
rect 22085 30514 22141 30570
rect 24017 30902 24073 30958
rect 25935 30709 25991 30765
rect 26315 30512 26371 30568
<< metal3 >>
rect 21701 30758 21757 30767
rect 21701 30693 21757 30702
rect 25935 30765 25991 30774
rect 25935 30700 25991 30709
rect 22085 30570 22141 30579
rect 22085 30505 22141 30514
rect 26315 30568 26371 30578
rect 26315 30503 26371 30512
<< via3 >>
rect 18624 30895 18710 30971
rect 22940 29565 23014 29636
rect 22483 29373 22555 29445
<< metal4 >>
rect 18618 30971 18716 31605
rect 18618 30895 18624 30971
rect 18710 30895 18716 30971
rect 18618 30886 18716 30895
rect 22481 29445 22558 31276
rect 22933 29636 23019 31187
rect 22933 29565 22940 29636
rect 23014 29565 23019 29636
rect 22933 29532 23019 29565
rect 22481 29373 22483 29445
rect 22555 29373 22558 29445
rect 22481 29341 22558 29373
use comparator  comparator_0 ~/Documents/fossi_cochlea/mag/final_designs/comparator
timestamp 1654741520
transform 1 0 23898 0 1 26079
box -779 -1057 1059 897
use filter  filter_0
timestamp 1654748254
transform 1 0 1272 0 1 -2522
box -1575 2522 22766 33508
use filter  filter_1
timestamp 1654748254
transform -1 0 46804 0 1 -2522
box -1575 2522 22766 33508
use filter_clkgen  filter_clkgen_0 ~/Documents/fossi_cochlea/mag/final_designs/clkgen
timestamp 1654741520
transform 1 0 20194 0 1 33321
box -1661 -2136 3360 1229
<< end >>
