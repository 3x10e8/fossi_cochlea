magic
tech sky130A
timestamp 1647865954
<< nwell >>
rect -256 -3 562 82
<< pmos >>
rect -209 17 -194 59
rect -165 17 -150 59
rect 0 17 15 59
rect 44 17 59 59
rect 88 17 103 59
rect 132 17 147 59
rect 264 15 279 57
rect 309 15 324 57
rect 451 15 466 57
rect 496 15 511 57
<< nmoslvt >>
rect -215 -133 -200 -91
rect -162 -133 -147 -91
rect -52 -133 -37 -91
rect 0 -133 15 -91
rect 44 -133 59 -91
rect 88 -133 103 -91
rect 132 -133 147 -91
rect 264 -133 279 -91
rect 309 -133 324 -91
rect 451 -133 466 -91
rect 496 -133 511 -91
<< ndiff >>
rect -252 -102 -215 -91
rect -252 -119 -248 -102
rect -231 -119 -215 -102
rect -252 -133 -215 -119
rect -200 -102 -162 -91
rect -200 -119 -189 -102
rect -172 -119 -162 -102
rect -200 -133 -162 -119
rect -147 -102 -110 -91
rect -147 -119 -131 -102
rect -114 -119 -110 -102
rect -147 -133 -110 -119
rect -79 -102 -52 -91
rect -79 -119 -75 -102
rect -58 -119 -52 -102
rect -79 -133 -52 -119
rect -37 -108 0 -91
rect -37 -125 -30 -108
rect -13 -125 0 -108
rect -37 -133 0 -125
rect 15 -102 44 -91
rect 15 -119 21 -102
rect 38 -119 44 -102
rect 15 -133 44 -119
rect 59 -102 88 -91
rect 59 -119 65 -102
rect 82 -119 88 -102
rect 59 -133 88 -119
rect 103 -102 132 -91
rect 103 -119 109 -102
rect 126 -119 132 -102
rect 103 -133 132 -119
rect 147 -102 177 -91
rect 147 -119 153 -102
rect 170 -119 177 -102
rect 147 -133 177 -119
rect 235 -102 264 -91
rect 235 -119 241 -102
rect 258 -119 264 -102
rect 235 -133 264 -119
rect 279 -102 309 -91
rect 279 -119 285 -102
rect 302 -119 309 -102
rect 279 -133 309 -119
rect 324 -102 354 -91
rect 324 -119 330 -102
rect 347 -119 354 -102
rect 421 -102 451 -91
rect 324 -133 354 -119
rect 421 -119 428 -102
rect 445 -119 451 -102
rect 421 -133 451 -119
rect 466 -102 496 -91
rect 466 -119 472 -102
rect 489 -119 496 -102
rect 466 -133 496 -119
rect 511 -102 540 -91
rect 511 -119 517 -102
rect 534 -119 540 -102
rect 511 -133 540 -119
<< pdiff >>
rect -238 48 -209 59
rect -238 31 -232 48
rect -215 31 -209 48
rect -238 17 -209 31
rect -194 48 -165 59
rect -194 31 -188 48
rect -171 31 -165 48
rect -194 17 -165 31
rect -150 48 -123 59
rect -150 31 -144 48
rect -127 31 -123 48
rect -150 17 -123 31
rect -27 48 0 59
rect -27 31 -23 48
rect -6 31 0 48
rect -27 17 0 31
rect 15 48 44 59
rect 15 31 21 48
rect 38 31 44 48
rect 15 17 44 31
rect 59 48 88 59
rect 59 31 65 48
rect 82 31 88 48
rect 59 17 88 31
rect 103 48 132 59
rect 103 31 109 48
rect 126 31 132 48
rect 103 17 132 31
rect 147 48 177 59
rect 147 31 153 48
rect 170 31 177 48
rect 147 17 177 31
rect 235 43 264 57
rect 235 26 241 43
rect 258 26 264 43
rect 235 15 264 26
rect 279 43 309 57
rect 279 26 286 43
rect 303 26 309 43
rect 279 15 309 26
rect 324 43 354 57
rect 324 26 330 43
rect 347 26 354 43
rect 421 43 451 57
rect 324 15 354 26
rect 421 26 428 43
rect 445 26 451 43
rect 421 15 451 26
rect 466 43 496 57
rect 466 26 473 43
rect 490 26 496 43
rect 466 15 496 26
rect 511 43 540 57
rect 511 26 517 43
rect 534 26 540 43
rect 511 15 540 26
<< ndiffc >>
rect -248 -119 -231 -102
rect -189 -119 -172 -102
rect -131 -119 -114 -102
rect -75 -119 -58 -102
rect -30 -125 -13 -108
rect 21 -119 38 -102
rect 65 -119 82 -102
rect 109 -119 126 -102
rect 153 -119 170 -102
rect 241 -119 258 -102
rect 285 -119 302 -102
rect 330 -119 347 -102
rect 428 -119 445 -102
rect 472 -119 489 -102
rect 517 -119 534 -102
<< pdiffc >>
rect -232 31 -215 48
rect -188 31 -171 48
rect -144 31 -127 48
rect -23 31 -6 48
rect 21 31 38 48
rect 65 31 82 48
rect 109 31 126 48
rect 153 31 170 48
rect 241 26 258 43
rect 286 26 303 43
rect 330 26 347 43
rect 428 26 445 43
rect 473 26 490 43
rect 517 26 534 43
<< psubdiff >>
rect 177 -103 208 -91
rect 177 -120 191 -103
rect 177 -133 208 -120
rect 354 -114 421 -91
rect 354 -131 385 -114
rect 402 -131 421 -114
rect 354 -133 421 -131
<< nsubdiff >>
rect 177 46 208 59
rect 177 29 191 46
rect 177 17 208 29
rect 354 55 421 57
rect 354 38 391 55
rect 408 38 421 55
rect 354 15 421 38
<< psubdiffcont >>
rect 191 -120 208 -103
rect 385 -131 402 -114
<< nsubdiffcont >>
rect 191 29 208 46
rect 391 38 408 55
<< poly >>
rect 75 115 108 123
rect 75 98 83 115
rect 100 113 108 115
rect 100 98 147 113
rect 75 93 108 98
rect -209 59 -194 72
rect -165 59 -150 72
rect 0 59 15 72
rect 44 59 59 72
rect 88 59 103 72
rect 132 59 147 98
rect -77 42 -35 50
rect -77 25 -72 42
rect -55 25 -35 42
rect -77 17 -35 25
rect 264 57 279 70
rect 309 57 324 70
rect 451 57 466 70
rect 496 57 511 70
rect -209 7 -194 17
rect -165 7 -150 17
rect -209 -8 -102 7
rect -50 6 -35 17
rect 0 6 15 17
rect -123 -13 -86 -8
rect -50 -9 15 6
rect -123 -15 -85 -13
rect -118 -23 -85 -15
rect -102 -30 -85 -23
rect -102 -35 -50 -30
rect -223 -45 -191 -36
rect -223 -62 -216 -45
rect -199 -62 -191 -45
rect -223 -70 -191 -62
rect -170 -45 -139 -36
rect -170 -62 -163 -45
rect -146 -62 -139 -45
rect -170 -70 -139 -62
rect -102 -52 -76 -35
rect -59 -52 -50 -35
rect 44 -39 59 17
rect 88 1 103 17
rect 132 4 147 17
rect 84 -7 111 1
rect 84 -24 89 -7
rect 106 -24 111 -7
rect 84 -32 111 -24
rect 206 -18 233 -10
rect -102 -57 -50 -52
rect 36 -42 59 -39
rect 36 -50 63 -42
rect -215 -91 -200 -70
rect -162 -91 -147 -70
rect -215 -146 -200 -133
rect -162 -146 -147 -133
rect -102 -141 -87 -57
rect 36 -67 41 -50
rect 58 -67 63 -50
rect 36 -75 63 -67
rect -52 -91 -37 -78
rect 0 -91 15 -78
rect 44 -91 59 -75
rect 88 -91 103 -32
rect 206 -35 211 -18
rect 228 -19 233 -18
rect 264 -19 279 15
rect 228 -34 279 -19
rect 309 -29 324 15
rect 393 -18 420 -10
rect 228 -35 233 -34
rect 152 -47 179 -39
rect 206 -43 233 -35
rect 152 -57 157 -47
rect 132 -64 157 -57
rect 174 -64 179 -47
rect 132 -72 179 -64
rect 132 -91 147 -72
rect 264 -91 279 -34
rect 303 -37 330 -29
rect 303 -54 308 -37
rect 325 -54 330 -37
rect 393 -35 398 -18
rect 415 -19 420 -18
rect 451 -19 466 15
rect 415 -34 466 -19
rect 496 -29 511 15
rect 415 -35 420 -34
rect 393 -43 420 -35
rect 303 -62 330 -54
rect 309 -91 324 -62
rect 451 -91 466 -34
rect 490 -37 517 -29
rect 490 -54 495 -37
rect 512 -54 517 -37
rect 490 -62 517 -54
rect 496 -91 511 -62
rect -52 -141 -37 -133
rect -102 -156 -37 -141
rect 0 -167 15 -133
rect 44 -146 59 -133
rect 88 -146 103 -133
rect 132 -167 147 -133
rect 264 -146 279 -133
rect 309 -146 324 -133
rect 451 -146 466 -133
rect 496 -146 511 -133
rect 0 -182 147 -167
<< polycont >>
rect 83 98 100 115
rect -72 25 -55 42
rect -216 -62 -199 -45
rect -163 -62 -146 -45
rect -76 -52 -59 -35
rect 89 -24 106 -7
rect 41 -67 58 -50
rect 211 -35 228 -18
rect 157 -64 174 -47
rect 308 -54 325 -37
rect 398 -35 415 -18
rect 495 -54 512 -37
<< locali >>
rect -286 134 -255 151
rect -238 134 -207 151
rect -190 134 -159 151
rect -142 134 -111 151
rect -94 134 -63 151
rect -46 134 -15 151
rect 2 134 33 151
rect 50 134 81 151
rect 98 134 129 151
rect 146 134 177 151
rect 194 134 225 151
rect 242 134 273 151
rect 290 134 321 151
rect 338 134 369 151
rect 386 134 417 151
rect 434 134 465 151
rect 482 134 513 151
rect 530 134 561 151
rect 578 134 609 151
rect -188 56 -171 134
rect -140 115 108 117
rect -140 100 83 115
rect -140 56 -123 100
rect 75 98 83 100
rect 100 98 108 115
rect 75 90 108 98
rect -252 48 -211 56
rect -252 31 -232 48
rect -215 31 -211 48
rect -252 23 -211 31
rect -192 48 -167 56
rect -192 31 -188 48
rect -171 31 -167 48
rect -192 23 -167 31
rect -148 55 -123 56
rect -148 48 -109 55
rect -148 31 -144 48
rect -127 31 -109 48
rect -148 23 -109 31
rect -252 -94 -235 23
rect -216 -45 -199 -36
rect -216 -70 -199 -62
rect -163 -45 -146 -36
rect -163 -70 -146 -62
rect -126 -94 -109 23
rect -75 42 -52 50
rect -75 25 -72 42
rect -55 25 -52 42
rect -75 17 -52 25
rect -27 48 -2 56
rect -27 31 -23 48
rect -6 31 -2 48
rect -27 23 -2 31
rect 17 48 42 56
rect 17 31 21 48
rect 38 31 42 48
rect 17 23 42 31
rect 61 48 88 56
rect 61 31 65 48
rect 82 31 88 48
rect 61 23 88 31
rect 105 48 130 56
rect 105 31 109 48
rect 126 31 130 48
rect 105 23 130 31
rect 149 48 174 56
rect 149 31 153 48
rect 170 31 174 48
rect 149 23 174 31
rect 191 46 208 134
rect 285 51 302 134
rect 391 55 408 134
rect -27 -7 -10 23
rect 89 -7 106 1
rect 153 -2 170 23
rect 191 21 208 29
rect 241 43 262 51
rect 258 26 262 43
rect 241 18 262 26
rect 282 43 307 51
rect 282 26 286 43
rect 303 26 307 43
rect 282 18 307 26
rect 326 43 368 51
rect 326 26 330 43
rect 347 26 368 43
rect 472 51 489 134
rect 391 30 408 38
rect 428 43 449 51
rect 326 18 368 26
rect 445 26 449 43
rect 428 18 449 26
rect 469 43 494 51
rect 469 26 473 43
rect 490 26 494 43
rect 469 18 494 26
rect 513 43 555 51
rect 513 26 517 43
rect 534 26 555 43
rect 513 18 555 26
rect -27 -24 89 -7
rect -84 -52 -76 -35
rect -59 -52 -51 -35
rect 7 -94 24 -24
rect 89 -32 106 -24
rect 123 -19 170 -2
rect 211 -18 228 -10
rect 41 -50 58 -42
rect 123 -50 140 -19
rect 58 -67 140 -50
rect 41 -75 58 -67
rect 110 -74 140 -67
rect 157 -47 174 -39
rect 211 -43 228 -35
rect 245 -37 262 18
rect 308 -37 325 -29
rect 157 -72 174 -64
rect 245 -54 308 -37
rect 110 -94 127 -74
rect 245 -94 262 -54
rect 308 -62 325 -54
rect 351 -94 368 18
rect 398 -18 415 -10
rect 398 -43 415 -35
rect 432 -37 449 18
rect 495 -37 512 -29
rect 432 -54 495 -37
rect 432 -94 449 -54
rect 495 -62 512 -54
rect 538 -94 555 18
rect -252 -102 -227 -94
rect -252 -119 -248 -102
rect -231 -119 -227 -102
rect -252 -127 -227 -119
rect -193 -102 -168 -94
rect -193 -119 -189 -102
rect -172 -119 -168 -102
rect -193 -127 -168 -119
rect -135 -102 -109 -94
rect -135 -119 -131 -102
rect -114 -111 -109 -102
rect -78 -102 -54 -94
rect -114 -119 -110 -111
rect -135 -127 -110 -119
rect -78 -119 -75 -102
rect -58 -119 -54 -102
rect -78 -127 -54 -119
rect -33 -108 -10 -100
rect -33 -125 -30 -108
rect -13 -125 -10 -108
rect 7 -102 42 -94
rect 7 -111 21 -102
rect -190 -145 -173 -127
rect -78 -145 -61 -127
rect -33 -133 -10 -125
rect 17 -119 21 -111
rect 38 -119 42 -102
rect 17 -127 42 -119
rect 61 -102 86 -94
rect 61 -119 65 -102
rect 82 -119 86 -102
rect 61 -127 86 -119
rect 105 -102 130 -94
rect 105 -119 109 -102
rect 126 -119 130 -102
rect 105 -127 130 -119
rect 149 -102 174 -94
rect 149 -119 153 -102
rect 170 -119 174 -102
rect 149 -127 174 -119
rect 191 -103 208 -94
rect -190 -162 -61 -145
rect -27 -182 -10 -133
rect 66 -182 83 -127
rect 154 -182 171 -127
rect 191 -182 208 -120
rect 241 -102 262 -94
rect 258 -119 262 -102
rect 241 -127 262 -119
rect 281 -102 306 -94
rect 281 -119 285 -102
rect 302 -119 306 -102
rect 281 -127 306 -119
rect 326 -102 368 -94
rect 326 -119 330 -102
rect 347 -119 368 -102
rect 428 -102 449 -94
rect 326 -127 368 -119
rect 385 -114 402 -106
rect 286 -182 303 -127
rect 445 -119 449 -102
rect 428 -127 449 -119
rect 468 -102 493 -94
rect 468 -119 472 -102
rect 489 -119 493 -102
rect 468 -127 493 -119
rect 513 -102 555 -94
rect 513 -119 517 -102
rect 534 -119 555 -102
rect 513 -127 555 -119
rect 385 -182 402 -131
rect 473 -182 490 -127
rect -286 -199 -255 -182
rect -238 -199 -207 -182
rect -190 -199 -159 -182
rect -142 -199 -111 -182
rect -94 -199 -63 -182
rect -46 -199 -15 -182
rect 2 -199 33 -182
rect 50 -199 81 -182
rect 98 -199 129 -182
rect 146 -199 177 -182
rect 194 -199 225 -182
rect 242 -199 273 -182
rect 290 -199 321 -182
rect 338 -199 369 -182
rect 386 -199 417 -182
rect 434 -199 465 -182
rect 482 -199 513 -182
rect 530 -199 561 -182
rect 578 -199 609 -182
<< viali >>
rect -255 134 -238 151
rect -207 134 -190 151
rect -159 134 -142 151
rect -111 134 -94 151
rect -63 134 -46 151
rect -15 134 2 151
rect 33 134 50 151
rect 81 134 98 151
rect 129 134 146 151
rect 177 134 194 151
rect 225 134 242 151
rect 273 134 290 151
rect 321 134 338 151
rect 369 134 386 151
rect 417 134 434 151
rect 465 134 482 151
rect 513 134 530 151
rect 561 134 578 151
rect -232 31 -215 48
rect -72 25 -55 42
rect 65 31 82 48
rect 89 -24 106 -7
rect 211 -35 228 -18
rect 41 -67 58 -50
rect 398 -35 415 -18
rect -255 -199 -238 -182
rect -207 -199 -190 -182
rect -159 -199 -142 -182
rect -111 -199 -94 -182
rect -63 -199 -46 -182
rect -15 -199 2 -182
rect 33 -199 50 -182
rect 81 -199 98 -182
rect 129 -199 146 -182
rect 177 -199 194 -182
rect 225 -199 242 -182
rect 273 -199 290 -182
rect 321 -199 338 -182
rect 369 -199 386 -182
rect 417 -199 434 -182
rect 465 -199 482 -182
rect 513 -199 530 -182
rect 561 -199 578 -182
<< metal1 >>
rect -286 151 609 167
rect -286 134 -255 151
rect -238 134 -207 151
rect -190 134 -159 151
rect -142 134 -111 151
rect -94 134 -63 151
rect -46 134 -15 151
rect 2 134 33 151
rect 50 134 81 151
rect 98 134 129 151
rect 146 134 177 151
rect 194 134 225 151
rect 242 134 273 151
rect 290 134 321 151
rect 338 134 369 151
rect 386 134 417 151
rect 434 134 465 151
rect 482 134 513 151
rect 530 134 561 151
rect 578 134 609 151
rect -286 118 609 134
rect -238 49 -211 52
rect 65 51 82 118
rect -238 48 -52 49
rect -238 31 -232 48
rect -215 42 -52 48
rect -215 31 -72 42
rect -238 30 -72 31
rect -238 27 -211 30
rect -75 25 -72 30
rect -55 25 -52 42
rect 62 48 85 51
rect 62 31 65 48
rect 82 31 85 48
rect 62 25 85 31
rect -75 18 -52 25
rect 84 -7 111 1
rect 84 -24 89 -7
rect 106 -18 233 -7
rect 106 -24 211 -18
rect 84 -32 111 -24
rect 206 -35 211 -24
rect 228 -35 233 -18
rect 36 -50 63 -41
rect 206 -43 233 -35
rect 395 -18 420 -7
rect 395 -35 398 -18
rect 415 -35 420 -18
rect 395 -43 420 -35
rect 36 -67 41 -50
rect 58 -67 63 -50
rect 36 -75 63 -67
rect 41 -102 58 -75
rect 398 -102 415 -43
rect 41 -119 415 -102
rect -286 -182 609 -166
rect -286 -199 -255 -182
rect -238 -199 -207 -182
rect -190 -199 -159 -182
rect -142 -199 -111 -182
rect -94 -199 -63 -182
rect -46 -199 -15 -182
rect 2 -199 33 -182
rect 50 -199 81 -182
rect 98 -199 129 -182
rect 146 -199 177 -182
rect 194 -199 225 -182
rect 242 -199 273 -182
rect 290 -199 321 -182
rect 338 -199 369 -182
rect 386 -199 417 -182
rect 434 -199 465 -182
rect 482 -199 513 -182
rect 530 -199 561 -182
rect 578 -199 609 -182
rect -286 -215 609 -199
<< labels >>
flabel polycont 89 -24 106 -7 0 FreeSans 56 0 0 0 high
flabel polycont 41 -67 58 -50 0 FreeSans 56 0 0 0 low
flabel polycont 157 -64 174 -47 0 FreeSans 56 0 0 0 phi1b
flabel polycont -76 -52 -59 -35 0 FreeSans 56 0 0 0 phi1
rlabel locali -51 -44 -51 -44 3 phi1
rlabel locali 118 56 118 56 1 pfete
rlabel locali 30 56 30 56 1 pfetw
rlabel locali 118 -94 118 -94 1 low
rlabel locali 30 -94 30 -94 1 high
rlabel locali 165 -39 165 -39 1 phi1b
rlabel locali -104 -145 -104 -145 1 tail
rlabel locali -155 -37 -155 -37 1 inm
flabel polycont -163 -62 -146 -45 0 FreeSans 56 0 0 0 inm
flabel polycont -216 -62 -199 -45 0 FreeSans 56 0 0 0 inp
rlabel locali -207 -36 -207 -36 1 inp
rlabel locali -235 -20 -235 -20 3 FP
rlabel locali -126 -23 -126 -23 7 FN
rlabel locali 273 144 273 144 3 VDD
rlabel locali 273 -191 273 -191 3 GND
flabel pdiffc 330 26 347 43 0 FreeSans 56 0 0 0 high_buffered
flabel ndiffc 517 -119 534 -102 0 FreeSans 56 0 0 0 low_buffered
<< end >>
