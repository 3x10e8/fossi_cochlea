** sch_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/tryandtest/for_lvs.sch
**.subckt for_lvs
x1 cc phi2b phi2 phi1b phi1 cclkb cclk vpb vnb vdda GND vccd div2 filter_clkgen_balanced_clks
XC1 net1 GND sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=32 m=32
XC2 GND net1 sky130_fd_pr__cap_mim_m3_2 W=10 L=10 VM=32 m=32
XC3 net2 GND sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=16 m=16
XC4 GND net2 sky130_fd_pr__cap_mim_m3_2 W=10 L=10 VM=16 m=16
XC5 net3 net4 sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=8 m=8
XC6 net4 net3 sky130_fd_pr__cap_mim_m3_2 W=10 L=10 VM=8 m=8
XC7 net5 GND sky130_fd_pr__cap_mim_m3_1 W=6 L=6.7 MF=1 m=1
XC8 net8 GND sky130_fd_pr__cap_mim_m3_1 W=3.4 L=3 MF=1 m=1
XC9 net6 GND sky130_fd_pr__cap_mim_m3_1 W=4 L=5 MF=1 m=1
XC10 net7 GND sky130_fd_pr__cap_mim_m3_1 W=3.4 L=3 MF=1 m=1
x2 th2 th1 cclk cclkb net4 GND vdda analogMux
x3 net3 net11 net19 phi1_ana phi1b_ana net20 vdda GND comparator_single_tail Wplus=0.42 Lplus=0.42
+ Wminus=0.42 Lminus=0.15
XC11 net9 GND sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=32 m=32
XC12 GND net9 sky130_fd_pr__cap_mim_m3_2 W=10 L=10 VM=32 m=32
XC13 net10 GND sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=16 m=16
XC14 GND net10 sky130_fd_pr__cap_mim_m3_2 W=10 L=10 VM=16 m=16
XC15 net11 net12 sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=8 m=8
XC16 net12 net11 sky130_fd_pr__cap_mim_m3_2 W=10 L=10 VM=8 m=8
XC17 net13 GND sky130_fd_pr__cap_mim_m3_1 W=6 L=6.7 MF=1 m=1
XC18 net16 GND sky130_fd_pr__cap_mim_m3_1 W=3.4 L=3 MF=1 m=1
XC19 net14 GND sky130_fd_pr__cap_mim_m3_1 W=4 L=5 MF=1 m=1
XC20 net15 GND sky130_fd_pr__cap_mim_m3_1 W=3.4 L=3 MF=1 m=1
x4 th1 th2 cclk cclkb net12 GND vdda analogMux
x5 inm inp sin sinb net17 GND vdda analogMux
x6 inp inm sin sinb x GND vdda analogMux
x7 inm inp cos cosb y GND vdda analogMux
x8 inp inm cos cosb net18 GND vdda analogMux
x9 net19 GND GND vdda VPWR net21 sky130_fd_sc_hd__buf_1
x10 net21 GND GND vdda VPWR high sky130_fd_sc_hd__buf_1
x11 net20 GND GND vdda VPWR net22 sky130_fd_sc_hd__buf_1
x12 net22 GND GND vdda VPWR low sky130_fd_sc_hd__buf_1
x13 fb net8 phi1b phi1 vdda GND tg Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x14 net8 net1 phi2b phi2 vdda GND tg Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x15 net17 net5 phi1b phi1 vdda GND tg Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x16 net5 net1 phi2b phi2 vdda GND tg Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x17 net1 net6 phi1b phi1 vdda GND tg Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x18 net6 net2 phi2b phi2 vdda GND tg Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x19 net2 net7 phi1b phi1 vdda GND tg Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x20 net7 net3 phi2b phi2 vdda GND tg Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x21 net15 net11 phi2b phi2 vdda GND tg Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x22 net10 net15 phi1b phi1 vdda GND tg Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x23 net14 net10 phi2b phi2 vdda GND tg Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x24 net9 net14 phi1b phi1 vdda GND tg Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x25 net13 net9 phi2b phi2 vdda GND tg Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x26 net18 net13 phi1b phi1 vdda GND tg Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x27 fb_inv net16 phi1b phi1 vdda GND tg Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x28 net16 net9 phi2b phi2 vdda GND tg Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
**.ends

* expanding   symbol:  clkgen/filter_clkgen_balanced_clks.sym # of pins=13
** sym_path:
*+ /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/clkgen/filter_clkgen_balanced_clks.sym
** sch_path:
*+ /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/clkgen/filter_clkgen_balanced_clks.sch
.subckt filter_clkgen_balanced_clks  cclk phi2b phi2 phi1b phi1 cclkb_ana cclk_ana vpb vnb vdda vssd
+ vccd div2
*.ipin div2
*.opin phi2
*.opin phi2b
*.opin phi1
*.opin phi1b
*.opin cclk_ana
*.opin cclkb_ana
*.ipin vpb
*.ipin vnb
*.ipin cclk
*.iopin vdda
*.iopin vccd
*.iopin vssd
X4 phi2dd phi2 phi2b vdda vssd comp_clks Wpmos=1.26 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
X7 phi1dd phi1 phi1b vdda vssd comp_clks Wpmos=1.26 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
X10 div2dd cclk_ana cclkb_ana vdda vssd comp_clks Wpmos=1.26 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
X1 div2 net3 net7 vccd vssd comp_clks_1stage Wpmos=1.26 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
X2 net1 phi2d vnb vdda vssd inv_weak_pulldown Wpmos=1.26 Lpmos= Wnmos= Lnmos=0.54
X5 net2 phi1d vnb vdda vssd inv_weak_pulldown Wpmos=1.26 Lpmos= Wnmos= Lnmos=0.54
X8 net5 div2d vnb vdda vssd inv_weak_pulldown Wpmos=1.26 Lpmos= Wnmos= Lnmos=0.54
X9 div2d div2dd vnb vdda vssd inv_weak_pulldown Wpmos=1.26 Lpmos= Wnmos= Lnmos=0.54
X3 phi2d phi2dd vpb vdda vssd inv_weak_pullup Wpmos=1.26 Lpmos=0.54 Wnmos= Lnmos=
X6 phi1d phi1dd vpb vdda vssd inv_weak_pullup Wpmos=1.26 Lpmos=0.54 Wnmos= Lnmos=
X11 cclk net4 net6 vccd vssd comp_clks_1stage Wpmos=1.26 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
x15 vdda vccd net3 net2 net1 vssd net7 level_up_shifter_no_inv
X14 vdda vccd net4 outb_alone net5 vssd net6 level_up_shifter_no_inv
.ends


* expanding   symbol:  mux/analogMux.sym # of pins=7
** sym_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/mux/analogMux.sym
** sch_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/mux/analogMux.sch
.subckt analogMux  vref2 vref1 c cbar out vssa vdda
*.ipin vref1
*.opin out
*.ipin vref2
*.ipin c
*.ipin cbar
*.ipin vssa
*.ipin vdda
XM2 vref1 c out vssa sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 vref1 cbar out vdda sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 out cbar vref2 vssa sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 out c vref2 vdda sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  comparator_latest/comparator_single_tail.sym # of pins=8
** sym_path:
*+ /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/comparator_latest/comparator_single_tail.sym
** sch_path:
*+ /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/comparator_latest/comparator_single_tail.sch
.subckt comparator_single_tail  inp inm high phi1 phi1b low vccd vssd   Wplus=0.42 Lplus=0.15
+ Wminus=0.42 Lminus=0.15
*.ipin phi1
*.opin high
*.ipin phi1b
*.ipin inp
*.ipin inm
*.opin low
*.iopin vccd
*.iopin vssd
XM12 FP inp tail GND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM13 FN inm tail GND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM14 pfetw low VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 high FP pfetw VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 pfete FN low VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 VDD high pfete VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 GND phi1b low GND sky130_fd_pr__nfet_01v8_lvt L=2 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 GND phi1b high GND sky130_fd_pr__nfet_01v8_lvt L=2 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 low high GND GND sky130_fd_pr__nfet_01v8_lvt L=2 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 high low GND GND sky130_fd_pr__nfet_01v8_lvt L=2 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 tail phi1 GND GND sky130_fd_pr__nfet_01v8_lvt L=2 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 VDD phi1 FP VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 FN phi1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  transmission_gate/tg.sym # of pins=6
** sym_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/transmission_gate/tg.sym
** sch_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/transmission_gate/tg.sch
.subckt tg  in out ctrl_ ctrl vdda vssa   Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
*.iopin in
*.iopin out
*.ipin ctrl_
*.ipin ctrl
*.ipin vdda
*.ipin vssa
XM1 out ctrl in vssa sky130_fd_pr__nfet_01v8 L=Lnmos W=Wnmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out ctrl_ in vdda sky130_fd_pr__pfet_01v8 L=Lpmos W=Wpmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
.ends


* expanding   symbol:  clkgen/comp_clks.sym # of pins=5
** sym_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/clkgen/comp_clks.sym
** sch_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/clkgen/comp_clks.sch
.subckt comp_clks  clk clka clkb vdda vssa   Wpmos=1.26 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
*.ipin clk
*.opin clka
*.opin clkb
*.ipin vdda
*.ipin vssa
X3 clk clkt vssa vdda vdda vssa transmission_gate Wpmos=Wpmos Lpmos=Lpmos Wnmos=Wnmos Lnmos=Lnmos
X1 clk clki vdda vssa inv Wpmos=Wpmos Lpmos=Lpmos Wnmos=Wnmos Lnmos=Lnmos
X2 clki clka vdda vssa inv Wpmos=Wpmos Lpmos=Lpmos Wnmos=Wnmos Lnmos=Lnmos
X4 clkt clkb vdda vssa inv Wpmos=Wpmos Lpmos=Lpmos Wnmos=Wnmos Lnmos=Lnmos
.ends


* expanding   symbol:  clkgen/comp_clks_1stage.sym # of pins=5
** sym_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/clkgen/comp_clks_1stage.sym
** sch_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/clkgen/comp_clks_1stage.sch
.subckt comp_clks_1stage  clk clka clkb vdda vssa   Wpmos=1.26 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
*.ipin clk
*.opin clka
*.opin clkb
*.ipin vdda
*.ipin vssa
X3 clk clkb vssa vdda vdda vssa transmission_gate Wpmos=Wpmos Lpmos=Lpmos Wnmos=Wnmos Lnmos=Lnmos
X1 clk clka vdda vssa inv Wpmos=Wpmos Lpmos=Lpmos Wnmos=Wnmos Lnmos=Lnmos
.ends


* expanding   symbol:  inv/inv_weak_pulldown.sym # of pins=5
** sym_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/inv/inv_weak_pulldown.sym
** sch_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/inv/inv_weak_pulldown.sch
.subckt inv_weak_pulldown  in out Vnb vdda vssa   Wpmos=1.26 Lmin=0.18 Wmin=0.42 Lnmos=0.54
*.ipin in
*.iopin out
*.ipin Vnb
*.ipin vdda
*.ipin vssa
XM1 net1 in vssa vssa sky130_fd_pr__nfet_01v8 L=Lmin W=Wmin nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 out Vnb net1 vssa sky130_fd_pr__nfet_01v8 L=Lnmos W=Wmin nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 out in vdda vdda sky130_fd_pr__pfet_01v8 L=Lmin W=Wpmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  inv/inv_weak_pullup.sym # of pins=5
** sym_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/inv/inv_weak_pullup.sym
** sch_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/inv/inv_weak_pullup.sch
.subckt inv_weak_pullup  in out Vpb vdda vssa   Wpmos=1.26 Lpmos=0.54 Wmin=0.42 Lmin=0.18
*.ipin in
*.iopin out
*.ipin Vpb
*.ipin vdda
*.ipin vssa
XM1 out in vssa vssa sky130_fd_pr__nfet_01v8 L=Lmin W=Wmin nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 out Vpb net1 vdda sky130_fd_pr__pfet_01v8 L=Lmin W=Wpmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net1 in vdda vdda sky130_fd_pr__pfet_01v8 L=Lmin W=Wpmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  level_shifter/level_up_shifter_no_inv.sym # of pins=7
** sym_path:
*+ /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/level_shifter/level_up_shifter_no_inv.sym
** sch_path:
*+ /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/level_shifter/level_up_shifter_no_inv.sch
.subckt level_up_shifter_no_inv  vdda1 vccd1 in outb out vssd1 inb
*.ipin in
*.iopin vdda1
*.opin out
*.opin outb
*.ipin inb
*.iopin vssd1
*.iopin vccd1
XM7 outb out vdda1 vdda1 sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 out outb vdda1 vdda1 sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 outb inb vdda1 vssd1 sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM3 outb in vssd1 vssd1 sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM4 vssd1 in outb vssd1 sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM5 out inb vssd1 vssd1 sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM6 vssd1 inb out vssd1 sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM9 vdda1 in out vssd1 sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM10 out in vdda1 vssd1 sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM11 vdda1 inb outb vssd1 sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
.ends


* expanding   symbol:  transmission_gate/transmission_gate.sym # of pins=6
** sym_path:
*+ /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/transmission_gate/transmission_gate.sym
** sch_path:
*+ /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/transmission_gate/transmission_gate.sch
.subckt transmission_gate  in out ctrl_ ctrl vdda vssa   Wpmos=0.42 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
*.iopin in
*.iopin out
*.ipin ctrl_
*.ipin ctrl
*.ipin vdda
*.ipin vssa
XM1 out ctrl in vssa sky130_fd_pr__nfet_01v8 L=Lnmos W=Wnmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out ctrl_ in vdda sky130_fd_pr__pfet_01v8 L=Lpmos W=Wpmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM3 in ctrl_ out vdda sky130_fd_pr__pfet_01v8 L=Lpmos W=Wpmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
.ends


* expanding   symbol:  inv/inv.sym # of pins=4
** sym_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/inv/inv.sym
** sch_path: /Volumes/export/isn/ankur/Documents/fossi_cochlea/xschem/inv/inv.sch
.subckt inv  in out vdda vssa   Wpmos=3 Lpmos=0.18 Wnmos=1 Lnmos=0.18
*.ipin in
*.iopin out
*.ipin vdda
*.ipin vssa
XM1 vssa in out vssa sky130_fd_pr__nfet_01v8 L=Lnmos W=Wnmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 vdda in out vdda sky130_fd_pr__pfet_01v8 L=Lpmos W=Wpmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 out in vdda vdda sky130_fd_pr__pfet_01v8 L=Lpmos W=Wpmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
