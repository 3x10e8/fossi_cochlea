magic
tech sky130B
magscale 1 2
timestamp 1663635562
use analog_core_Q  analog_core_Q_0 final_designs
timestamp 1663635562
transform 1 0 0 0 1 -35689
box 0 0 406272 35689
use digital_unison  digital_unison_0
timestamp 1663374934
transform 1 0 0 0 1 0
box 0 0 406984 24000
<< end >>
