magic
tech sky130B
magscale 1 2
timestamp 1662946268
<< nwell >>
rect 1715 1303 2125 1535
<< nmos >>
rect 1230 1060 1260 1180
rect 1316 1060 1346 1180
rect 1403 1060 1433 1180
rect 1489 1060 1519 1180
rect 1576 1060 1606 1180
rect 1662 1060 1692 1180
rect 1749 1060 1779 1180
rect 1835 1060 1865 1180
rect 1922 1060 1952 1180
rect 2008 1060 2038 1180
rect 2095 1060 2125 1180
rect 2181 1060 2211 1180
rect 2268 1060 2298 1180
rect 2354 1060 2384 1180
rect 2441 1060 2471 1180
rect 2527 1060 2557 1180
rect 1230 620 1260 740
rect 1316 620 1346 740
rect 1403 620 1433 740
rect 1489 620 1519 740
rect 1576 620 1606 740
rect 1662 620 1692 740
rect 1749 620 1779 740
rect 1835 620 1865 740
rect 1922 620 1952 740
rect 2008 620 2038 740
rect 2095 620 2125 740
rect 2181 620 2211 740
rect 2268 620 2298 740
rect 2354 620 2384 740
rect 2441 620 2471 740
rect 2527 620 2557 740
<< pmos >>
rect 1829 1375 1859 1459
rect 1930 1375 1960 1459
<< ndiff >>
rect 1173 1168 1230 1180
rect 1173 1134 1185 1168
rect 1219 1134 1230 1168
rect 1173 1060 1230 1134
rect 1260 1106 1316 1180
rect 1260 1072 1271 1106
rect 1305 1072 1316 1106
rect 1260 1060 1316 1072
rect 1346 1168 1403 1180
rect 1346 1134 1358 1168
rect 1392 1134 1403 1168
rect 1346 1060 1403 1134
rect 1433 1106 1489 1180
rect 1433 1072 1444 1106
rect 1478 1072 1489 1106
rect 1433 1060 1489 1072
rect 1519 1168 1576 1180
rect 1519 1134 1531 1168
rect 1565 1134 1576 1168
rect 1519 1060 1576 1134
rect 1606 1106 1662 1180
rect 1606 1072 1617 1106
rect 1651 1072 1662 1106
rect 1606 1060 1662 1072
rect 1692 1168 1749 1180
rect 1692 1134 1704 1168
rect 1738 1134 1749 1168
rect 1692 1060 1749 1134
rect 1779 1106 1835 1180
rect 1779 1072 1790 1106
rect 1824 1072 1835 1106
rect 1779 1060 1835 1072
rect 1865 1168 1922 1180
rect 1865 1134 1877 1168
rect 1911 1134 1922 1168
rect 1865 1060 1922 1134
rect 1952 1106 2008 1180
rect 1952 1072 1963 1106
rect 1997 1072 2008 1106
rect 1952 1060 2008 1072
rect 2038 1168 2095 1180
rect 2038 1134 2050 1168
rect 2084 1134 2095 1168
rect 2038 1060 2095 1134
rect 2125 1106 2181 1180
rect 2125 1072 2136 1106
rect 2170 1072 2181 1106
rect 2125 1060 2181 1072
rect 2211 1168 2268 1180
rect 2211 1134 2223 1168
rect 2257 1134 2268 1168
rect 2211 1060 2268 1134
rect 2298 1106 2354 1180
rect 2298 1072 2309 1106
rect 2343 1072 2354 1106
rect 2298 1060 2354 1072
rect 2384 1168 2441 1180
rect 2384 1134 2396 1168
rect 2430 1134 2441 1168
rect 2384 1060 2441 1134
rect 2471 1106 2527 1180
rect 2471 1072 2482 1106
rect 2516 1072 2527 1106
rect 2471 1060 2527 1072
rect 2557 1168 2614 1180
rect 2557 1134 2569 1168
rect 2603 1134 2614 1168
rect 2557 1060 2614 1134
rect 1170 728 1230 740
rect 1170 694 1185 728
rect 1219 694 1230 728
rect 1170 620 1230 694
rect 1260 666 1316 740
rect 1260 632 1271 666
rect 1305 632 1316 666
rect 1260 620 1316 632
rect 1346 728 1403 740
rect 1346 694 1358 728
rect 1392 694 1403 728
rect 1346 620 1403 694
rect 1433 666 1489 740
rect 1433 632 1444 666
rect 1478 632 1489 666
rect 1433 620 1489 632
rect 1519 728 1576 740
rect 1519 694 1531 728
rect 1565 694 1576 728
rect 1519 620 1576 694
rect 1606 667 1662 740
rect 1606 633 1617 667
rect 1651 633 1662 667
rect 1606 620 1662 633
rect 1692 728 1749 740
rect 1692 694 1704 728
rect 1738 694 1749 728
rect 1692 620 1749 694
rect 1779 666 1835 740
rect 1779 632 1790 666
rect 1824 632 1835 666
rect 1779 620 1835 632
rect 1865 728 1922 740
rect 1865 694 1877 728
rect 1911 694 1922 728
rect 1865 620 1922 694
rect 1952 666 2008 740
rect 1952 632 1963 666
rect 1997 632 2008 666
rect 1952 620 2008 632
rect 2038 728 2095 740
rect 2038 694 2050 728
rect 2084 694 2095 728
rect 2038 620 2095 694
rect 2125 666 2181 740
rect 2125 632 2136 666
rect 2170 632 2181 666
rect 2125 620 2181 632
rect 2211 728 2268 740
rect 2211 694 2223 728
rect 2257 694 2268 728
rect 2211 620 2268 694
rect 2298 666 2354 740
rect 2298 632 2309 666
rect 2343 632 2354 666
rect 2298 620 2354 632
rect 2384 728 2441 740
rect 2384 694 2396 728
rect 2430 694 2441 728
rect 2384 620 2441 694
rect 2471 666 2527 740
rect 2471 632 2482 666
rect 2516 632 2527 666
rect 2471 620 2527 632
rect 2557 728 2618 740
rect 2557 694 2569 728
rect 2603 694 2618 728
rect 2557 620 2618 694
<< pdiff >>
rect 1763 1435 1829 1459
rect 1763 1401 1783 1435
rect 1817 1401 1829 1435
rect 1763 1375 1829 1401
rect 1859 1435 1930 1459
rect 1859 1401 1877 1435
rect 1911 1401 1930 1435
rect 1859 1375 1930 1401
rect 1960 1435 2020 1459
rect 1960 1401 1975 1435
rect 2009 1401 2020 1435
rect 1960 1375 2020 1401
<< ndiffc >>
rect 1185 1134 1219 1168
rect 1271 1072 1305 1106
rect 1358 1134 1392 1168
rect 1444 1072 1478 1106
rect 1531 1134 1565 1168
rect 1617 1072 1651 1106
rect 1704 1134 1738 1168
rect 1790 1072 1824 1106
rect 1877 1134 1911 1168
rect 1963 1072 1997 1106
rect 2050 1134 2084 1168
rect 2136 1072 2170 1106
rect 2223 1134 2257 1168
rect 2309 1072 2343 1106
rect 2396 1134 2430 1168
rect 2482 1072 2516 1106
rect 2569 1134 2603 1168
rect 1185 694 1219 728
rect 1271 632 1305 666
rect 1358 694 1392 728
rect 1444 632 1478 666
rect 1531 694 1565 728
rect 1617 633 1651 667
rect 1704 694 1738 728
rect 1790 632 1824 666
rect 1877 694 1911 728
rect 1963 632 1997 666
rect 2050 694 2084 728
rect 2136 632 2170 666
rect 2223 694 2257 728
rect 2309 632 2343 666
rect 2396 694 2430 728
rect 2482 632 2516 666
rect 2569 694 2603 728
<< pdiffc >>
rect 1783 1401 1817 1435
rect 1877 1401 1911 1435
rect 1975 1401 2009 1435
<< psubdiff >>
rect 1112 707 1170 740
rect 1112 673 1113 707
rect 1147 673 1170 707
rect 1112 620 1170 673
rect 2618 713 2691 740
rect 2618 679 2647 713
rect 2681 679 2691 713
rect 2618 620 2691 679
<< nsubdiff >>
rect 2020 1435 2089 1459
rect 2020 1401 2043 1435
rect 2077 1401 2089 1435
rect 2020 1375 2089 1401
<< psubdiffcont >>
rect 1113 673 1147 707
rect 2647 679 2681 713
<< nsubdiffcont >>
rect 2043 1401 2077 1435
<< poly >>
rect 1817 1540 1871 1550
rect 1811 1506 1827 1540
rect 1861 1506 1877 1540
rect 1817 1496 1871 1506
rect 1829 1459 1859 1496
rect 1930 1459 1960 1485
rect 1829 1349 1859 1375
rect 1930 1338 1960 1375
rect 1918 1328 1972 1338
rect 1912 1294 1928 1328
rect 1962 1294 1978 1328
rect 1918 1284 1972 1294
rect 1203 1253 1269 1269
rect 1203 1219 1219 1253
rect 1254 1219 1269 1253
rect 1209 1209 1264 1219
rect 1230 1180 1260 1209
rect 1316 1180 1346 1206
rect 1403 1180 1433 1206
rect 1489 1180 1519 1206
rect 1576 1180 1606 1206
rect 1662 1180 1692 1206
rect 1749 1180 1779 1206
rect 1835 1180 1865 1206
rect 1922 1180 1952 1206
rect 2008 1180 2038 1206
rect 2095 1180 2125 1206
rect 2181 1180 2211 1206
rect 2268 1180 2298 1206
rect 2354 1180 2384 1206
rect 2441 1180 2471 1206
rect 2527 1180 2557 1206
rect 1230 1034 1260 1060
rect 1316 1034 1346 1060
rect 1403 1034 1433 1060
rect 1489 1034 1519 1060
rect 1576 1034 1606 1060
rect 1662 1034 1692 1060
rect 1749 1034 1779 1060
rect 1835 1034 1865 1060
rect 1230 1004 1865 1034
rect 1922 1034 1952 1060
rect 2008 1034 2038 1060
rect 2095 1034 2125 1060
rect 2181 1034 2211 1060
rect 2268 1034 2298 1060
rect 2354 1034 2384 1060
rect 2441 1034 2471 1060
rect 2527 1034 2557 1060
rect 1922 1004 2557 1034
rect 1778 970 1788 1004
rect 1823 970 1833 1004
rect 1778 954 1833 970
rect 1922 912 1952 1004
rect 1785 882 1952 912
rect 1235 820 1290 836
rect 1235 796 1245 820
rect 1230 786 1245 796
rect 1280 796 1290 820
rect 1785 796 1815 882
rect 1977 830 2032 846
rect 1977 796 1987 830
rect 2022 796 2032 830
rect 1280 786 1865 796
rect 1230 766 1865 786
rect 1230 740 1260 766
rect 1316 740 1346 766
rect 1403 740 1433 766
rect 1489 740 1519 766
rect 1576 740 1606 766
rect 1662 740 1692 766
rect 1749 740 1779 766
rect 1835 740 1865 766
rect 1922 766 2557 796
rect 1922 740 1952 766
rect 2008 740 2038 766
rect 2095 740 2125 766
rect 2181 740 2211 766
rect 2268 740 2298 766
rect 2354 740 2384 766
rect 2441 740 2471 766
rect 2527 740 2557 766
rect 1230 594 1260 620
rect 1316 594 1346 620
rect 1403 594 1433 620
rect 1489 594 1519 620
rect 1576 594 1606 620
rect 1662 594 1692 620
rect 1749 594 1779 620
rect 1835 594 1865 620
rect 1922 594 1952 620
rect 2008 594 2038 620
rect 2095 594 2125 620
rect 2181 594 2211 620
rect 2268 594 2298 620
rect 2354 594 2384 620
rect 2441 594 2471 620
rect 2527 594 2557 620
<< polycont >>
rect 1827 1506 1861 1540
rect 1928 1294 1962 1328
rect 1219 1219 1254 1253
rect 1788 970 1823 1004
rect 1245 786 1280 820
rect 1987 796 2022 830
<< locali >>
rect 1506 1617 1535 1651
rect 1569 1617 1627 1651
rect 1661 1617 1719 1651
rect 1753 1617 1811 1651
rect 1845 1617 1903 1651
rect 1937 1617 1995 1651
rect 2029 1617 2087 1651
rect 2121 1617 2179 1651
rect 2213 1617 2271 1651
rect 2305 1617 2363 1651
rect 2397 1617 2455 1651
rect 2489 1617 2547 1651
rect 2581 1617 2639 1651
rect 2673 1617 2731 1651
rect 2765 1617 2794 1651
rect 1811 1506 1827 1540
rect 1861 1506 2170 1540
rect 1783 1435 1817 1451
rect 1783 1328 1817 1401
rect 1877 1435 1911 1451
rect 1877 1385 1911 1401
rect 1975 1435 2009 1506
rect 1975 1385 2009 1401
rect 2043 1435 2077 1451
rect 2043 1385 2077 1401
rect 1783 1294 1928 1328
rect 1962 1294 1978 1328
rect 934 1219 1219 1253
rect 1254 1219 1270 1253
rect 1185 1168 1219 1184
rect 1185 1118 1219 1134
rect 1358 1168 1392 1184
rect 1271 1106 1305 1122
rect 1358 1118 1392 1134
rect 1531 1168 1565 1184
rect 1271 1056 1305 1072
rect 1444 1106 1478 1122
rect 1531 1118 1565 1134
rect 1704 1168 1738 1184
rect 1444 1056 1478 1072
rect 1617 1106 1651 1122
rect 1704 1118 1738 1134
rect 1617 1056 1651 1072
rect 1790 1106 1824 1294
rect 1877 1168 1911 1184
rect 1877 1118 1911 1134
rect 2050 1168 2084 1184
rect 1790 1056 1824 1072
rect 1963 1106 1997 1122
rect 2050 1118 2084 1134
rect 1963 1056 1997 1072
rect 2136 1106 2170 1506
rect 2223 1168 2257 1184
rect 2223 1118 2257 1134
rect 2396 1168 2430 1184
rect 2136 1056 2170 1072
rect 2309 1106 2343 1122
rect 2396 1118 2430 1134
rect 2569 1168 2603 1184
rect 2309 1056 2343 1072
rect 2482 1106 2516 1122
rect 2569 1118 2603 1134
rect 2482 1056 2516 1072
rect 1772 970 1788 1004
rect 1823 970 1839 1004
rect 759 851 1280 886
rect 1245 820 1280 851
rect 1788 830 1823 970
rect 1788 796 1987 830
rect 2022 796 2038 830
rect 1245 770 1280 786
rect 1185 728 1219 744
rect 1113 707 1147 723
rect 1185 678 1219 694
rect 1358 728 1392 744
rect 1113 657 1147 673
rect 1271 666 1305 682
rect 1358 678 1392 694
rect 1531 728 1565 744
rect 1271 616 1305 632
rect 1444 666 1478 682
rect 1531 678 1565 694
rect 1704 728 1738 744
rect 1444 616 1478 632
rect 1617 667 1651 683
rect 1704 678 1738 694
rect 1877 728 1911 744
rect 1617 616 1651 633
rect 1790 666 1824 682
rect 1877 678 1911 694
rect 2050 728 2084 744
rect 1790 616 1824 632
rect 1963 666 1997 682
rect 2050 678 2084 694
rect 2223 728 2257 744
rect 1963 616 1997 632
rect 2136 666 2170 682
rect 2223 678 2257 694
rect 2396 728 2430 744
rect 2136 616 2170 632
rect 2309 666 2343 682
rect 2396 678 2430 694
rect 2569 728 2603 744
rect 2309 616 2343 632
rect 2482 666 2516 682
rect 2569 678 2603 694
rect 2647 713 2681 729
rect 2482 616 2516 632
rect 2647 563 2681 679
rect 1596 529 1627 563
rect 1663 529 1719 563
rect 1753 529 1811 563
rect 1845 529 1903 563
rect 1937 529 1995 563
rect 2029 529 2087 563
rect 2121 529 2179 563
rect 2213 529 2271 563
rect 2305 529 2363 563
rect 2397 529 2455 563
rect 2489 529 2547 563
rect 2581 529 2639 563
rect 2673 529 2731 563
rect 2765 529 2794 563
<< viali >>
rect 1535 1617 1569 1651
rect 1627 1617 1661 1651
rect 1719 1617 1753 1651
rect 1811 1617 1845 1651
rect 1903 1617 1937 1651
rect 1995 1617 2029 1651
rect 2087 1617 2121 1651
rect 2179 1617 2213 1651
rect 2271 1617 2305 1651
rect 2363 1617 2397 1651
rect 2455 1617 2489 1651
rect 2547 1617 2581 1651
rect 2639 1617 2673 1651
rect 2731 1617 2765 1651
rect 1877 1401 1911 1435
rect 2043 1401 2077 1435
rect 1185 1134 1219 1168
rect 1358 1134 1392 1168
rect 1531 1134 1565 1168
rect 1271 1072 1305 1106
rect 1704 1134 1738 1168
rect 1444 1072 1478 1106
rect 1617 1072 1651 1106
rect 1877 1134 1911 1168
rect 2050 1134 2084 1168
rect 1790 1072 1824 1106
rect 1963 1072 1997 1106
rect 2223 1134 2257 1168
rect 2396 1134 2430 1168
rect 2136 1072 2170 1106
rect 2569 1134 2603 1168
rect 2309 1072 2343 1106
rect 2482 1072 2516 1106
rect 1113 673 1147 707
rect 1185 694 1219 728
rect 1358 694 1392 728
rect 1531 694 1565 728
rect 1271 632 1305 666
rect 1704 694 1738 728
rect 1444 632 1478 666
rect 1877 694 1911 728
rect 1617 633 1651 667
rect 2050 694 2084 728
rect 1790 632 1824 666
rect 2223 694 2257 728
rect 1963 632 1997 666
rect 2396 694 2430 728
rect 2136 632 2170 666
rect 2569 694 2603 728
rect 2309 632 2343 666
rect 2647 679 2681 713
rect 2482 632 2516 666
rect 1627 529 1663 563
rect 1719 529 1753 563
rect 1811 529 1845 563
rect 1903 529 1937 563
rect 1995 529 2029 563
rect 2087 529 2121 563
rect 2179 529 2213 563
rect 2271 529 2305 563
rect 2363 529 2397 563
rect 2455 529 2489 563
rect 2547 529 2581 563
rect 2639 529 2673 563
rect 2731 529 2765 563
<< metal1 >>
rect 427 1321 681 1361
rect 985 1329 1029 1683
rect 1506 1651 2794 1682
rect 1506 1617 1535 1651
rect 1569 1617 1627 1651
rect 1661 1617 1719 1651
rect 1753 1617 1811 1651
rect 1845 1617 1903 1651
rect 1937 1617 1995 1651
rect 2029 1617 2087 1651
rect 2121 1617 2179 1651
rect 2213 1617 2271 1651
rect 2305 1617 2363 1651
rect 2397 1617 2455 1651
rect 2489 1617 2547 1651
rect 2581 1617 2639 1651
rect 2673 1617 2731 1651
rect 2765 1617 2794 1651
rect 1506 1586 2794 1617
rect 1910 1447 1998 1586
rect 1871 1435 1998 1447
rect 2037 1435 2083 1441
rect 1871 1401 1877 1435
rect 1911 1401 2043 1435
rect 2077 1401 2089 1435
rect 1871 1395 1917 1401
rect 2037 1395 2083 1401
rect 427 1042 471 1321
rect 837 1289 1029 1329
rect 1877 1174 1911 1395
rect 1173 1168 2615 1174
rect 1173 1134 1185 1168
rect 1219 1142 1358 1168
rect 1219 1134 1231 1142
rect 1173 1128 1231 1134
rect 1346 1134 1358 1142
rect 1392 1142 1531 1168
rect 1392 1134 1404 1142
rect 1346 1128 1404 1134
rect 1519 1134 1531 1142
rect 1565 1142 1704 1168
rect 1565 1134 1577 1142
rect 1519 1128 1577 1134
rect 1692 1134 1704 1142
rect 1738 1142 1877 1168
rect 1738 1134 1750 1142
rect 1692 1128 1750 1134
rect 1865 1134 1877 1142
rect 1911 1142 2050 1168
rect 1911 1134 1923 1142
rect 1865 1128 1923 1134
rect 2038 1134 2050 1142
rect 2084 1142 2223 1168
rect 2084 1134 2096 1142
rect 2038 1128 2096 1134
rect 2211 1134 2223 1142
rect 2257 1142 2396 1168
rect 2257 1134 2269 1142
rect 2211 1128 2269 1134
rect 2384 1134 2396 1142
rect 2430 1142 2569 1168
rect 2430 1134 2442 1142
rect 2384 1128 2442 1134
rect 2557 1134 2569 1142
rect 2603 1134 2615 1168
rect 2557 1128 2615 1134
rect 1259 1106 1320 1114
rect 1259 1072 1271 1106
rect 1305 1097 1320 1106
rect 1432 1106 1493 1114
rect 1432 1097 1444 1106
rect 1305 1072 1444 1097
rect 1478 1097 1493 1106
rect 1603 1097 1609 1114
rect 1478 1072 1609 1097
rect 1661 1097 1667 1114
rect 1778 1106 1839 1114
rect 1778 1097 1790 1106
rect 1661 1072 1790 1097
rect 1824 1072 1839 1106
rect 1951 1106 2012 1114
rect 1951 1097 1963 1106
rect 1259 1066 1609 1072
rect 1603 1062 1609 1066
rect 1661 1066 1839 1072
rect 1950 1072 1963 1097
rect 1997 1097 2012 1106
rect 2121 1097 2127 1114
rect 1997 1072 2127 1097
rect 2179 1097 2185 1114
rect 2297 1106 2358 1114
rect 2297 1097 2309 1106
rect 2179 1072 2309 1097
rect 2343 1097 2358 1106
rect 2470 1106 2531 1114
rect 2470 1097 2482 1106
rect 2343 1072 2482 1097
rect 2516 1097 2531 1106
rect 2516 1072 2614 1097
rect 1950 1066 2127 1072
rect 1661 1062 1667 1066
rect 2121 1062 2127 1066
rect 2179 1066 2614 1072
rect 2179 1062 2185 1066
rect 1603 1061 1667 1062
rect 1107 728 2687 734
rect 1107 707 1185 728
rect 1107 673 1113 707
rect 1147 694 1185 707
rect 1219 702 1358 728
rect 1219 694 1231 702
rect 1147 688 1231 694
rect 1346 694 1358 702
rect 1392 702 1531 728
rect 1392 694 1404 702
rect 1346 688 1404 694
rect 1519 694 1531 702
rect 1565 703 1704 728
rect 1565 694 1577 703
rect 1519 688 1577 694
rect 1692 694 1704 703
rect 1738 702 1877 728
rect 1738 694 1750 702
rect 1692 688 1750 694
rect 1865 694 1877 702
rect 1911 702 2050 728
rect 1911 694 1923 702
rect 1865 688 1923 694
rect 2038 694 2050 702
rect 2084 704 2223 728
rect 2084 694 2096 704
rect 2211 694 2223 704
rect 2257 702 2396 728
rect 2257 694 2269 702
rect 2038 688 2096 694
rect 2215 688 2269 694
rect 2384 694 2396 702
rect 2430 702 2569 728
rect 2430 694 2442 702
rect 2384 688 2442 694
rect 2557 694 2569 702
rect 2603 713 2687 728
rect 2603 694 2647 713
rect 2557 688 2647 694
rect 1147 673 1157 688
rect 1107 661 1157 673
rect 1259 666 1320 674
rect 1259 632 1271 666
rect 1305 657 1320 666
rect 1432 666 1493 674
rect 1432 657 1444 666
rect 1305 632 1444 657
rect 1478 657 1493 666
rect 1603 657 1609 675
rect 1478 632 1609 657
rect 1661 657 1667 675
rect 1778 666 1839 674
rect 1778 657 1790 666
rect 1259 626 1609 632
rect 1603 623 1609 626
rect 1661 632 1790 657
rect 1824 632 1839 666
rect 1661 626 1839 632
rect 1661 623 1667 626
rect 1603 622 1667 623
rect 1877 594 1911 688
rect 2639 679 2647 688
rect 2681 679 2687 713
rect 1951 666 2012 674
rect 1951 657 1963 666
rect 1950 632 1963 657
rect 1997 657 2012 666
rect 2123 657 2129 674
rect 1997 632 2129 657
rect 2181 657 2187 674
rect 2297 666 2358 674
rect 2297 657 2309 666
rect 2181 632 2309 657
rect 2343 657 2358 666
rect 2470 666 2531 674
rect 2639 667 2687 679
rect 2470 657 2482 666
rect 2343 632 2482 657
rect 2516 632 2531 666
rect 1950 626 2129 632
rect 2123 622 2129 626
rect 2181 626 2531 632
rect 2181 622 2187 626
rect 1571 572 2794 594
rect 1571 520 1617 572
rect 1670 563 2794 572
rect 1670 529 1719 563
rect 1753 529 1811 563
rect 1845 529 1903 563
rect 1937 529 1995 563
rect 2029 529 2087 563
rect 2121 529 2179 563
rect 2213 529 2271 563
rect 2305 529 2363 563
rect 2397 529 2455 563
rect 2489 529 2547 563
rect 2581 529 2639 563
rect 2673 529 2731 563
rect 2765 529 2794 563
rect 1670 520 2794 529
rect 1571 498 2794 520
<< via1 >>
rect 1609 1106 1661 1114
rect 1609 1072 1617 1106
rect 1617 1072 1651 1106
rect 1651 1072 1661 1106
rect 1609 1062 1661 1072
rect 2127 1106 2179 1114
rect 2127 1072 2136 1106
rect 2136 1072 2170 1106
rect 2170 1072 2179 1106
rect 2127 1062 2179 1072
rect 1609 667 1661 675
rect 1609 633 1617 667
rect 1617 633 1651 667
rect 1651 633 1661 667
rect 1609 623 1661 633
rect 2129 666 2181 674
rect 2129 632 2136 666
rect 2136 632 2170 666
rect 2170 632 2181 666
rect 2129 622 2181 632
rect 1617 563 1670 572
rect 1617 529 1627 563
rect 1627 529 1663 563
rect 1663 529 1670 563
rect 1617 520 1670 529
<< metal2 >>
rect 1603 1062 1609 1114
rect 1661 1062 1667 1114
rect 2121 1062 2127 1114
rect 2179 1062 2185 1114
rect 1617 675 1651 1062
rect 1603 623 1609 675
rect 1661 623 1667 675
rect 2136 674 2170 1062
rect 1603 622 1667 623
rect 2123 622 2129 674
rect 2181 622 2187 674
rect 2123 620 2187 622
rect 1607 572 1681 574
rect 1607 520 1617 572
rect 1670 520 1681 572
rect 1607 518 1681 520
use comp_clks_stg1  comp_clks_stg1_0 clkgen
timestamp 1662946268
transform 1 0 402 0 -1 1138
box 0 -547 644 640
<< end >>
