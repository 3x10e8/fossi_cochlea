magic
tech sky130B
magscale 1 2
timestamp 1654756118
<< viali >>
rect -9808 42802 -9634 43538
<< metal1 >>
rect -9846 43538 -9590 43598
rect -9846 42802 -9808 43538
rect -9634 42802 -9590 43538
rect -9846 42746 -9590 42802
rect -9733 37898 -9671 42746
rect -22638 37836 -9671 37898
rect -19438 34012 -6846 34030
rect -19438 33954 -19418 34012
rect -19366 33954 -6846 34012
rect -19438 33938 -6846 33954
rect -19010 32590 -18874 32596
rect -19010 32546 -19004 32590
rect -26706 32540 -19004 32546
rect -26710 32470 -19004 32540
rect -18882 32524 -18874 32590
rect -18882 32470 -18872 32524
rect -26710 32422 -18872 32470
rect -26710 31910 -26674 32422
rect -6956 31274 -6864 33938
<< via1 >>
rect -9808 42802 -9634 43538
rect -19418 33954 -19366 34012
rect -19004 32470 -18882 32590
<< metal2 >>
rect -9846 43538 -9590 43598
rect -16028 43328 -15818 43354
rect -16028 42794 -15982 43328
rect -15842 42794 -15818 43328
rect -16028 42780 -15818 42794
rect -9846 42802 -9808 43538
rect -9634 42802 -9590 43538
rect -15987 42731 -15861 42780
rect -9846 42746 -9590 42802
rect -19008 42605 -15861 42731
rect -26160 42242 -26108 42272
rect -35742 42190 -26108 42242
rect -35742 36712 -35690 42190
rect -26160 41392 -26108 42190
rect -26856 41224 -26778 41234
rect -26856 41216 -26848 41224
rect -27750 41166 -26848 41216
rect -26788 41166 -26778 41224
rect -26856 41160 -26778 41166
rect -26818 40948 -26638 41000
rect -26818 40378 -26774 40948
rect -26818 40334 -19370 40378
rect -30362 38244 -30272 38254
rect -30362 38182 -30352 38244
rect -30282 38182 -30272 38244
rect -30362 38172 -30272 38182
rect -30360 37638 -30278 37648
rect -30360 37578 -30350 37638
rect -30288 37578 -30278 37638
rect -30360 37568 -30278 37578
rect -43040 36660 -35690 36712
rect -43040 36376 -42988 36660
rect -43040 31302 -42986 36376
rect -19414 34022 -19370 40334
rect -19424 34012 -19360 34022
rect -19424 33954 -19418 34012
rect -19366 33954 -19360 34012
rect -19424 33944 -19360 33954
rect -19008 32596 -18882 42605
rect -19010 32590 -18874 32596
rect -19010 32470 -19004 32590
rect -18882 32470 -18874 32590
rect -19010 32464 -18874 32470
<< via2 >>
rect -15982 42794 -15842 43328
rect -9808 42802 -9634 43538
rect -26848 41166 -26788 41224
rect -30352 38182 -30282 38244
rect -30350 37578 -30288 37638
<< metal3 >>
rect -28384 43127 -28044 43602
rect -9846 43538 -9590 43598
rect -31098 42941 -28044 43127
rect -31098 41582 -30912 42941
rect -28384 42788 -28044 42941
rect -22424 42535 -21460 43508
rect -16028 43328 -15818 43354
rect -16028 42794 -15982 43328
rect -15842 42794 -15818 43328
rect -16028 42780 -15818 42794
rect -9846 42802 -9808 43538
rect -9634 42802 -9590 43538
rect -9846 42746 -9590 42802
rect -30758 42456 -21460 42535
rect -30758 42436 -21927 42456
rect -31098 37650 -30916 41582
rect -30758 38252 -30659 42436
rect -22081 42408 -21927 42436
rect -26876 41234 -26770 41268
rect -26876 41160 -26856 41234
rect -26778 41160 -26770 41234
rect -26876 41136 -26770 41160
rect -30366 38252 -30272 38254
rect -30758 38244 -30272 38252
rect -30758 38182 -30352 38244
rect -30282 38182 -30272 38244
rect -30758 38172 -30272 38182
rect -30758 38170 -30274 38172
rect -30366 38168 -30274 38170
rect -31098 37638 -30278 37650
rect -31098 37578 -30350 37638
rect -30288 37578 -30278 37638
rect -31098 37568 -30278 37578
<< via3 >>
rect -3708 42866 -3600 43434
rect -26856 41224 -26778 41234
rect -26856 41166 -26848 41224
rect -26848 41166 -26788 41224
rect -26788 41166 -26778 41224
rect -26856 41160 -26778 41166
<< metal4 >>
rect -3730 43434 -3554 43600
rect -3730 42866 -3708 43434
rect -3600 42866 -3554 43434
rect -26876 41234 -26770 41268
rect -26876 41160 -26856 41234
rect -26778 41232 -26770 41234
rect -3730 41232 -3554 42866
rect -26778 41160 -3507 41232
rect -26876 41150 -3507 41160
rect -26876 41136 -26770 41150
rect -3730 41134 -3554 41150
use filter_p_m  filter_p_m_0
array 0 1 -48682 0 0 34550
timestamp 1654754989
transform 1 0 -321 0 1 5258
box -303 0 48379 37136
use filter_p_m  filter_p_m_1
array 0 1 -48682 0 0 34550
timestamp 1654754989
transform -1 0 -927 0 -1 159808
box -303 0 48379 37136
use first_dual_core  first_dual_core_0 ../digital
timestamp 1654751233
transform 0 -1 48362 1 0 42794
box 0 0 80000 98000
<< end >>
