VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO comparator_final
  CLASS BLOCK ;
  FOREIGN comparator_final ;
  ORIGIN 2.870 2.150 ;
  SIZE 51.080 BY 4.155 ;
  OBS
      LAYER nwell ;
        RECT 5.745 0.820 47.885 1.615 ;
        RECT -2.560 -0.030 47.885 0.820 ;
        RECT 5.745 -0.250 47.885 -0.030 ;
      LAYER pwell ;
        RECT 9.940 -0.760 10.900 -0.540 ;
        RECT 13.170 -0.760 14.540 -0.540 ;
        RECT 18.580 -0.760 19.540 -0.540 ;
        RECT 21.810 -0.760 23.180 -0.540 ;
        RECT 27.220 -0.760 28.180 -0.540 ;
        RECT 30.450 -0.760 31.820 -0.540 ;
        RECT 35.860 -0.760 36.820 -0.540 ;
        RECT 39.090 -0.760 40.460 -0.540 ;
        RECT 7.100 -1.045 14.540 -0.760 ;
        RECT 15.740 -0.765 23.180 -0.760 ;
        RECT 15.740 -1.045 23.295 -0.765 ;
        RECT 24.380 -0.780 31.820 -0.760 ;
        RECT 24.380 -1.045 31.945 -0.780 ;
        RECT 33.020 -0.795 40.460 -0.760 ;
        RECT 33.020 -1.045 40.540 -0.795 ;
        RECT 5.940 -1.050 14.540 -1.045 ;
        RECT 14.580 -1.050 40.540 -1.045 ;
        RECT 5.940 -1.645 40.540 -1.050 ;
        RECT 5.940 -1.660 23.180 -1.645 ;
        RECT 23.220 -1.660 40.540 -1.645 ;
        RECT 40.575 -1.660 43.800 -0.590 ;
        RECT 44.185 -1.660 46.055 -0.700 ;
        RECT 46.260 -1.660 47.690 -0.700 ;
        RECT 5.935 -1.905 47.695 -1.660 ;
        RECT 44.455 -1.940 44.795 -1.905 ;
      LAYER li1 ;
        RECT -2.860 1.340 47.695 1.510 ;
        RECT -1.880 0.560 -1.710 1.340 ;
        RECT -1.400 1.000 1.080 1.170 ;
        RECT -1.400 0.560 -1.230 1.000 ;
        RECT 0.750 0.900 1.080 1.000 ;
        RECT -2.520 0.230 -2.110 0.560 ;
        RECT -1.920 0.230 -1.670 0.560 ;
        RECT -1.480 0.550 -1.230 0.560 ;
        RECT -1.480 0.230 -1.090 0.550 ;
        RECT -2.520 -0.940 -2.350 0.230 ;
        RECT -2.160 -0.700 -1.990 -0.360 ;
        RECT -1.630 -0.700 -1.460 -0.360 ;
        RECT -1.260 -0.940 -1.090 0.230 ;
        RECT -0.750 0.170 -0.520 0.500 ;
        RECT -0.270 0.230 -0.020 0.560 ;
        RECT 0.170 0.230 0.420 0.560 ;
        RECT 0.610 0.230 0.880 0.560 ;
        RECT 1.050 0.230 1.300 0.560 ;
        RECT 1.490 0.230 1.740 0.560 ;
        RECT -0.270 -0.070 -0.100 0.230 ;
        RECT 0.890 -0.070 1.060 0.010 ;
        RECT 1.530 -0.020 1.700 0.230 ;
        RECT 1.910 0.210 2.080 1.340 ;
        RECT 2.850 0.510 3.020 1.340 ;
        RECT 2.410 0.180 2.620 0.510 ;
        RECT 2.820 0.180 3.070 0.510 ;
        RECT 3.260 0.180 3.680 0.510 ;
        RECT 3.910 0.300 4.080 1.340 ;
        RECT 4.720 0.510 4.890 1.340 ;
        RECT 6.030 0.755 6.360 1.340 ;
        RECT 4.280 0.180 4.490 0.510 ;
        RECT 4.690 0.180 4.940 0.510 ;
        RECT 5.130 0.180 5.550 0.510 ;
        RECT -0.270 -0.240 1.060 -0.070 ;
        RECT -0.840 -0.520 -0.510 -0.350 ;
        RECT 0.070 -0.940 0.240 -0.240 ;
        RECT 0.890 -0.320 1.060 -0.240 ;
        RECT 1.230 -0.190 1.700 -0.020 ;
        RECT 0.410 -0.500 0.580 -0.420 ;
        RECT 1.230 -0.500 1.400 -0.190 ;
        RECT 0.410 -0.670 1.400 -0.500 ;
        RECT 0.410 -0.750 0.580 -0.670 ;
        RECT 1.100 -0.740 1.400 -0.670 ;
        RECT 1.570 -0.720 1.740 -0.390 ;
        RECT 2.110 -0.430 2.280 -0.100 ;
        RECT 2.450 -0.370 2.620 0.180 ;
        RECT 3.080 -0.370 3.250 -0.290 ;
        RECT 2.450 -0.540 3.250 -0.370 ;
        RECT 1.100 -0.940 1.270 -0.740 ;
        RECT 2.450 -0.940 2.620 -0.540 ;
        RECT 3.080 -0.620 3.250 -0.540 ;
        RECT 3.510 -0.940 3.680 0.180 ;
        RECT 3.980 -0.430 4.150 -0.100 ;
        RECT 4.320 -0.370 4.490 0.180 ;
        RECT 4.950 -0.370 5.120 -0.290 ;
        RECT 4.320 -0.540 5.120 -0.370 ;
        RECT 4.320 -0.940 4.490 -0.540 ;
        RECT 4.950 -0.620 5.120 -0.540 ;
        RECT 5.380 -0.940 5.550 0.180 ;
        RECT -2.520 -1.270 -2.270 -0.940 ;
        RECT -1.930 -1.270 -1.680 -0.940 ;
        RECT -1.350 -1.110 -1.090 -0.940 ;
        RECT -1.350 -1.270 -1.100 -1.110 ;
        RECT -0.780 -1.270 -0.540 -0.940 ;
        RECT -1.900 -1.450 -1.730 -1.270 ;
        RECT -0.780 -1.450 -0.610 -1.270 ;
        RECT -0.330 -1.330 -0.100 -1.000 ;
        RECT 0.070 -1.110 0.420 -0.940 ;
        RECT 0.170 -1.270 0.420 -1.110 ;
        RECT 0.610 -1.270 0.860 -0.940 ;
        RECT 1.050 -1.270 1.300 -0.940 ;
        RECT 1.490 -1.270 1.740 -0.940 ;
        RECT -1.900 -1.620 -0.610 -1.450 ;
        RECT -0.270 -1.820 -0.100 -1.330 ;
        RECT 0.660 -1.820 0.830 -1.270 ;
        RECT 1.540 -1.820 1.710 -1.270 ;
        RECT 1.910 -1.820 2.080 -0.940 ;
        RECT 2.410 -1.270 2.620 -0.940 ;
        RECT 2.810 -1.270 3.060 -0.940 ;
        RECT 3.260 -1.270 3.680 -0.940 ;
        RECT 2.860 -1.820 3.030 -1.270 ;
        RECT 3.850 -1.820 4.020 -1.060 ;
        RECT 4.280 -1.270 4.490 -0.940 ;
        RECT 4.680 -1.270 4.930 -0.940 ;
        RECT 5.130 -1.270 5.550 -0.940 ;
        RECT 6.020 -1.065 6.360 0.585 ;
        RECT 4.730 -1.820 4.900 -1.270 ;
        RECT 6.030 -1.820 6.360 -1.235 ;
        RECT 6.530 -1.575 6.975 1.145 ;
        RECT 7.145 0.200 7.355 0.960 ;
        RECT 7.525 0.380 7.855 1.340 ;
        RECT 8.025 0.855 9.625 1.035 ;
        RECT 8.025 0.200 8.205 0.855 ;
        RECT 7.145 0.030 8.205 0.200 ;
        RECT 7.145 -1.265 7.520 0.030 ;
        RECT 7.875 -0.765 8.205 -0.140 ;
        RECT 8.375 -0.685 8.565 0.685 ;
        RECT 8.735 -0.520 8.905 0.855 ;
        RECT 9.075 -0.680 9.285 0.685 ;
        RECT 9.455 0.550 9.625 0.855 ;
        RECT 9.910 0.720 10.240 1.340 ;
        RECT 9.455 0.380 11.100 0.550 ;
        RECT 9.540 0.010 10.750 0.210 ;
        RECT 9.540 -0.500 9.870 0.010 ;
        RECT 10.110 -0.680 10.360 -0.230 ;
        RECT 8.375 -0.935 8.555 -0.685 ;
        RECT 9.075 -0.850 10.360 -0.680 ;
        RECT 9.075 -0.870 9.275 -0.850 ;
        RECT 7.690 -1.820 7.970 -0.935 ;
        RECT 8.160 -1.265 8.555 -0.935 ;
        RECT 8.725 -1.040 9.275 -0.870 ;
        RECT 8.725 -1.265 8.995 -1.040 ;
        RECT 9.455 -1.820 10.360 -1.020 ;
        RECT 10.530 -1.320 10.740 0.010 ;
        RECT 10.920 -0.350 11.100 0.380 ;
        RECT 11.270 -0.030 11.590 0.850 ;
        RECT 12.085 0.070 12.465 1.340 ;
        RECT 10.920 -0.430 11.240 -0.350 ;
        RECT 10.910 -0.610 11.240 -0.430 ;
        RECT 11.420 -0.610 11.590 -0.030 ;
        RECT 12.685 -0.100 13.100 0.850 ;
        RECT 13.270 -0.090 13.550 1.340 ;
        RECT 11.960 -0.260 13.100 -0.100 ;
        RECT 11.960 -0.270 13.370 -0.260 ;
        RECT 11.960 -0.440 12.290 -0.270 ;
        RECT 12.500 -0.610 12.760 -0.450 ;
        RECT 11.420 -0.780 12.760 -0.610 ;
        RECT 12.930 -0.480 13.370 -0.270 ;
        RECT 11.080 -1.260 11.590 -0.780 ;
        RECT 12.930 -0.960 13.100 -0.480 ;
        RECT 11.935 -1.820 12.455 -0.960 ;
        RECT 12.625 -1.490 13.100 -0.960 ;
        RECT 13.270 -1.820 13.550 -0.650 ;
        RECT 13.720 -1.530 13.985 1.170 ;
        RECT 14.155 -0.090 14.390 1.340 ;
        RECT 14.670 0.755 15.000 1.340 ;
        RECT 14.155 -1.820 14.390 -0.650 ;
        RECT 14.660 -1.065 15.000 0.585 ;
        RECT 14.670 -1.820 15.000 -1.235 ;
        RECT 15.170 -1.575 15.615 1.145 ;
        RECT 15.785 0.200 15.995 0.960 ;
        RECT 16.165 0.380 16.495 1.340 ;
        RECT 16.665 0.855 18.265 1.035 ;
        RECT 16.665 0.200 16.845 0.855 ;
        RECT 15.785 0.030 16.845 0.200 ;
        RECT 15.785 -1.265 16.160 0.030 ;
        RECT 16.515 -0.765 16.845 -0.140 ;
        RECT 17.015 -0.685 17.205 0.685 ;
        RECT 17.375 -0.520 17.545 0.855 ;
        RECT 17.715 -0.680 17.925 0.685 ;
        RECT 18.095 0.550 18.265 0.855 ;
        RECT 18.550 0.720 18.880 1.340 ;
        RECT 18.095 0.380 19.740 0.550 ;
        RECT 18.180 0.010 19.390 0.210 ;
        RECT 18.180 -0.500 18.510 0.010 ;
        RECT 18.750 -0.680 19.000 -0.230 ;
        RECT 17.015 -0.935 17.195 -0.685 ;
        RECT 17.715 -0.850 19.000 -0.680 ;
        RECT 17.715 -0.870 17.915 -0.850 ;
        RECT 16.330 -1.820 16.610 -0.935 ;
        RECT 16.800 -1.265 17.195 -0.935 ;
        RECT 17.365 -1.040 17.915 -0.870 ;
        RECT 17.365 -1.265 17.635 -1.040 ;
        RECT 18.095 -1.820 19.000 -1.020 ;
        RECT 19.170 -1.320 19.380 0.010 ;
        RECT 19.560 -0.350 19.740 0.380 ;
        RECT 19.910 -0.030 20.230 0.850 ;
        RECT 20.725 0.070 21.105 1.340 ;
        RECT 19.560 -0.430 19.880 -0.350 ;
        RECT 19.550 -0.610 19.880 -0.430 ;
        RECT 20.060 -0.610 20.230 -0.030 ;
        RECT 21.325 -0.100 21.740 0.850 ;
        RECT 21.910 -0.090 22.190 1.340 ;
        RECT 20.600 -0.260 21.740 -0.100 ;
        RECT 20.600 -0.270 22.010 -0.260 ;
        RECT 20.600 -0.440 20.930 -0.270 ;
        RECT 21.140 -0.610 21.400 -0.450 ;
        RECT 20.060 -0.780 21.400 -0.610 ;
        RECT 21.570 -0.480 22.010 -0.270 ;
        RECT 19.720 -1.260 20.230 -0.780 ;
        RECT 21.570 -0.960 21.740 -0.480 ;
        RECT 20.575 -1.820 21.095 -0.960 ;
        RECT 21.265 -1.490 21.740 -0.960 ;
        RECT 21.910 -1.820 22.190 -0.650 ;
        RECT 22.360 -1.530 22.625 1.170 ;
        RECT 22.795 -0.090 23.030 1.340 ;
        RECT 23.310 0.755 23.640 1.340 ;
        RECT 22.795 -1.820 23.030 -0.650 ;
        RECT 23.300 -1.065 23.640 0.585 ;
        RECT 23.310 -1.820 23.640 -1.235 ;
        RECT 23.810 -1.575 24.255 1.145 ;
        RECT 24.425 0.200 24.635 0.960 ;
        RECT 24.805 0.380 25.135 1.340 ;
        RECT 25.305 0.855 26.905 1.035 ;
        RECT 25.305 0.200 25.485 0.855 ;
        RECT 24.425 0.030 25.485 0.200 ;
        RECT 24.425 -1.265 24.800 0.030 ;
        RECT 25.155 -0.765 25.485 -0.140 ;
        RECT 25.655 -0.685 25.845 0.685 ;
        RECT 26.015 -0.520 26.185 0.855 ;
        RECT 26.355 -0.680 26.565 0.685 ;
        RECT 26.735 0.550 26.905 0.855 ;
        RECT 27.190 0.720 27.520 1.340 ;
        RECT 26.735 0.380 28.380 0.550 ;
        RECT 26.820 0.010 28.030 0.210 ;
        RECT 26.820 -0.500 27.150 0.010 ;
        RECT 27.390 -0.680 27.640 -0.230 ;
        RECT 25.655 -0.935 25.835 -0.685 ;
        RECT 26.355 -0.850 27.640 -0.680 ;
        RECT 26.355 -0.870 26.555 -0.850 ;
        RECT 24.970 -1.820 25.250 -0.935 ;
        RECT 25.440 -1.265 25.835 -0.935 ;
        RECT 26.005 -1.040 26.555 -0.870 ;
        RECT 26.005 -1.265 26.275 -1.040 ;
        RECT 26.735 -1.820 27.640 -1.020 ;
        RECT 27.810 -1.320 28.020 0.010 ;
        RECT 28.200 -0.350 28.380 0.380 ;
        RECT 28.550 -0.030 28.870 0.850 ;
        RECT 29.365 0.070 29.745 1.340 ;
        RECT 28.200 -0.430 28.520 -0.350 ;
        RECT 28.190 -0.610 28.520 -0.430 ;
        RECT 28.700 -0.610 28.870 -0.030 ;
        RECT 29.965 -0.100 30.380 0.850 ;
        RECT 30.550 -0.090 30.830 1.340 ;
        RECT 29.240 -0.260 30.380 -0.100 ;
        RECT 29.240 -0.270 30.650 -0.260 ;
        RECT 29.240 -0.440 29.570 -0.270 ;
        RECT 29.780 -0.610 30.040 -0.450 ;
        RECT 28.700 -0.780 30.040 -0.610 ;
        RECT 30.210 -0.480 30.650 -0.270 ;
        RECT 28.360 -1.260 28.870 -0.780 ;
        RECT 30.210 -0.960 30.380 -0.480 ;
        RECT 29.215 -1.820 29.735 -0.960 ;
        RECT 29.905 -1.490 30.380 -0.960 ;
        RECT 30.550 -1.820 30.830 -0.650 ;
        RECT 31.000 -1.530 31.265 1.170 ;
        RECT 31.435 -0.090 31.670 1.340 ;
        RECT 31.950 0.755 32.280 1.340 ;
        RECT 31.435 -1.820 31.670 -0.650 ;
        RECT 31.940 -1.065 32.280 0.585 ;
        RECT 31.950 -1.820 32.280 -1.235 ;
        RECT 32.450 -1.575 32.895 1.145 ;
        RECT 33.065 0.200 33.275 0.960 ;
        RECT 33.445 0.380 33.775 1.340 ;
        RECT 33.945 0.855 35.545 1.035 ;
        RECT 33.945 0.200 34.125 0.855 ;
        RECT 33.065 0.030 34.125 0.200 ;
        RECT 33.065 -1.265 33.440 0.030 ;
        RECT 33.795 -0.765 34.125 -0.140 ;
        RECT 34.295 -0.685 34.485 0.685 ;
        RECT 34.655 -0.520 34.825 0.855 ;
        RECT 34.995 -0.680 35.205 0.685 ;
        RECT 35.375 0.550 35.545 0.855 ;
        RECT 35.830 0.720 36.160 1.340 ;
        RECT 35.375 0.380 37.020 0.550 ;
        RECT 35.460 0.010 36.670 0.210 ;
        RECT 35.460 -0.500 35.790 0.010 ;
        RECT 36.030 -0.680 36.280 -0.230 ;
        RECT 34.295 -0.935 34.475 -0.685 ;
        RECT 34.995 -0.850 36.280 -0.680 ;
        RECT 34.995 -0.870 35.195 -0.850 ;
        RECT 33.610 -1.820 33.890 -0.935 ;
        RECT 34.080 -1.265 34.475 -0.935 ;
        RECT 34.645 -1.040 35.195 -0.870 ;
        RECT 34.645 -1.265 34.915 -1.040 ;
        RECT 35.375 -1.820 36.280 -1.020 ;
        RECT 36.450 -1.320 36.660 0.010 ;
        RECT 36.840 -0.350 37.020 0.380 ;
        RECT 37.190 -0.030 37.510 0.850 ;
        RECT 38.005 0.070 38.385 1.340 ;
        RECT 36.840 -0.430 37.160 -0.350 ;
        RECT 36.830 -0.610 37.160 -0.430 ;
        RECT 37.340 -0.610 37.510 -0.030 ;
        RECT 38.605 -0.100 39.020 0.850 ;
        RECT 39.190 -0.090 39.470 1.340 ;
        RECT 37.880 -0.260 39.020 -0.100 ;
        RECT 37.880 -0.270 39.290 -0.260 ;
        RECT 37.880 -0.440 38.210 -0.270 ;
        RECT 38.420 -0.610 38.680 -0.450 ;
        RECT 37.340 -0.780 38.680 -0.610 ;
        RECT 38.850 -0.480 39.290 -0.270 ;
        RECT 37.000 -1.260 37.510 -0.780 ;
        RECT 38.850 -0.960 39.020 -0.480 ;
        RECT 37.855 -1.820 38.375 -0.960 ;
        RECT 38.545 -1.490 39.020 -0.960 ;
        RECT 39.190 -1.820 39.470 -0.650 ;
        RECT 39.640 -1.530 39.905 1.170 ;
        RECT 40.075 -0.090 40.310 1.340 ;
        RECT 40.665 0.330 40.995 1.170 ;
        RECT 41.485 0.500 41.765 1.340 ;
        RECT 41.935 0.840 42.265 1.170 ;
        RECT 42.460 1.010 42.790 1.340 ;
        RECT 43.430 0.840 43.760 1.020 ;
        RECT 41.935 0.670 43.760 0.840 ;
        RECT 41.935 0.500 42.265 0.670 ;
        RECT 42.435 0.330 43.730 0.500 ;
        RECT 40.665 0.160 42.605 0.330 ;
        RECT 40.580 -0.180 42.610 -0.010 ;
        RECT 43.000 -0.110 43.330 0.160 ;
        RECT 43.000 -0.155 43.230 -0.110 ;
        RECT 40.075 -1.820 40.310 -0.650 ;
        RECT 40.580 -0.695 40.950 -0.180 ;
        RECT 41.120 -0.695 42.260 -0.350 ;
        RECT 42.430 -0.560 42.610 -0.180 ;
        RECT 42.780 -0.335 43.230 -0.155 ;
        RECT 43.560 -0.280 43.730 0.330 ;
        RECT 44.275 0.050 44.605 1.340 ;
        RECT 44.775 0.185 45.105 0.380 ;
        RECT 45.400 0.355 45.730 1.340 ;
        RECT 44.775 0.015 45.730 0.185 ;
        RECT 42.780 -0.740 42.950 -0.335 ;
        RECT 43.400 -0.505 43.730 -0.280 ;
        RECT 43.940 -0.415 44.720 -0.155 ;
        RECT 44.890 -0.415 45.290 -0.155 ;
        RECT 40.665 -1.820 40.925 -0.865 ;
        RECT 41.095 -1.035 42.365 -0.865 ;
        RECT 41.095 -1.570 41.355 -1.035 ;
        RECT 41.525 -1.820 41.855 -1.205 ;
        RECT 42.195 -1.480 42.365 -1.035 ;
        RECT 42.535 -1.310 42.950 -0.740 ;
        RECT 43.120 -0.675 43.730 -0.505 ;
        RECT 45.480 -0.585 45.730 0.015 ;
        RECT 43.120 -1.480 43.290 -0.675 ;
        RECT 44.275 -0.755 45.730 -0.585 ;
        RECT 42.195 -1.650 43.290 -1.480 ;
        RECT 43.460 -1.820 43.710 -0.845 ;
        RECT 44.275 -1.205 44.605 -0.755 ;
        RECT 45.900 -0.925 46.170 1.170 ;
        RECT 46.350 -0.130 46.670 0.580 ;
        RECT 46.840 0.040 47.170 1.340 ;
        RECT 47.340 -0.040 47.610 1.170 ;
        RECT 46.350 -0.200 47.190 -0.130 ;
        RECT 46.350 -0.300 47.265 -0.200 ;
        RECT 46.340 -0.715 46.690 -0.470 ;
        RECT 47.000 -0.720 47.265 -0.300 ;
        RECT 47.000 -0.885 47.170 -0.720 ;
        RECT 47.435 -0.875 47.610 -0.040 ;
        RECT 44.520 -1.820 44.730 -1.555 ;
        RECT 45.065 -1.820 45.435 -0.925 ;
        RECT 45.605 -1.650 46.170 -0.925 ;
        RECT 46.350 -1.055 47.170 -0.885 ;
        RECT 46.350 -1.215 46.670 -1.055 ;
        RECT 46.840 -1.820 47.170 -1.225 ;
        RECT 47.340 -1.650 47.610 -0.875 ;
        RECT -2.860 -1.990 47.695 -1.820 ;
      LAYER mcon ;
        RECT -2.550 1.340 -2.380 1.510 ;
        RECT -2.070 1.340 -1.900 1.510 ;
        RECT -1.590 1.340 -1.420 1.510 ;
        RECT -1.110 1.340 -0.940 1.510 ;
        RECT -0.630 1.340 -0.460 1.510 ;
        RECT -0.150 1.340 0.020 1.510 ;
        RECT 0.330 1.340 0.500 1.510 ;
        RECT 0.810 1.340 0.980 1.510 ;
        RECT 1.290 1.340 1.460 1.510 ;
        RECT 1.770 1.340 1.940 1.510 ;
        RECT 2.250 1.340 2.420 1.510 ;
        RECT 2.730 1.340 2.900 1.510 ;
        RECT 3.210 1.340 3.380 1.510 ;
        RECT 3.690 1.340 3.860 1.510 ;
        RECT 4.170 1.340 4.340 1.510 ;
        RECT 4.650 1.340 4.820 1.510 ;
        RECT 5.130 1.340 5.300 1.510 ;
        RECT 5.610 1.340 5.780 1.510 ;
        RECT 6.090 1.340 6.260 1.510 ;
        RECT 6.570 1.340 6.740 1.510 ;
        RECT 7.050 1.340 7.220 1.510 ;
        RECT 7.530 1.340 7.700 1.510 ;
        RECT 8.010 1.340 8.180 1.510 ;
        RECT 8.490 1.340 8.660 1.510 ;
        RECT 8.970 1.340 9.140 1.510 ;
        RECT 9.450 1.340 9.620 1.510 ;
        RECT 9.930 1.340 10.100 1.510 ;
        RECT 10.410 1.340 10.580 1.510 ;
        RECT 10.890 1.340 11.060 1.510 ;
        RECT 11.370 1.340 11.540 1.510 ;
        RECT 11.850 1.340 12.020 1.510 ;
        RECT 12.330 1.340 12.500 1.510 ;
        RECT 12.810 1.340 12.980 1.510 ;
        RECT 13.290 1.340 13.460 1.510 ;
        RECT 13.770 1.340 13.940 1.510 ;
        RECT 14.250 1.340 14.420 1.510 ;
        RECT 14.730 1.340 14.900 1.510 ;
        RECT 15.210 1.340 15.380 1.510 ;
        RECT 15.690 1.340 15.860 1.510 ;
        RECT 16.170 1.340 16.340 1.510 ;
        RECT 16.650 1.340 16.820 1.510 ;
        RECT 17.130 1.340 17.300 1.510 ;
        RECT 17.610 1.340 17.780 1.510 ;
        RECT 18.090 1.340 18.260 1.510 ;
        RECT 18.570 1.340 18.740 1.510 ;
        RECT 19.050 1.340 19.220 1.510 ;
        RECT 19.530 1.340 19.700 1.510 ;
        RECT 20.010 1.340 20.180 1.510 ;
        RECT 20.490 1.340 20.660 1.510 ;
        RECT 20.970 1.340 21.140 1.510 ;
        RECT 21.450 1.340 21.620 1.510 ;
        RECT 21.930 1.340 22.100 1.510 ;
        RECT 22.410 1.340 22.580 1.510 ;
        RECT 22.890 1.340 23.060 1.510 ;
        RECT 23.370 1.340 23.540 1.510 ;
        RECT 23.850 1.340 24.020 1.510 ;
        RECT 24.330 1.340 24.500 1.510 ;
        RECT 24.810 1.340 24.980 1.510 ;
        RECT 25.290 1.340 25.460 1.510 ;
        RECT 25.770 1.340 25.940 1.510 ;
        RECT 26.250 1.340 26.420 1.510 ;
        RECT 26.730 1.340 26.900 1.510 ;
        RECT 27.210 1.340 27.380 1.510 ;
        RECT 27.690 1.340 27.860 1.510 ;
        RECT 28.170 1.340 28.340 1.510 ;
        RECT 28.650 1.340 28.820 1.510 ;
        RECT 29.130 1.340 29.300 1.510 ;
        RECT 29.610 1.340 29.780 1.510 ;
        RECT 30.090 1.340 30.260 1.510 ;
        RECT 30.570 1.340 30.740 1.510 ;
        RECT 31.050 1.340 31.220 1.510 ;
        RECT 31.530 1.340 31.700 1.510 ;
        RECT 32.010 1.340 32.180 1.510 ;
        RECT 32.490 1.340 32.660 1.510 ;
        RECT 32.970 1.340 33.140 1.510 ;
        RECT 33.450 1.340 33.620 1.510 ;
        RECT 33.930 1.340 34.100 1.510 ;
        RECT 34.410 1.340 34.580 1.510 ;
        RECT 34.890 1.340 35.060 1.510 ;
        RECT 35.370 1.340 35.540 1.510 ;
        RECT 35.850 1.340 36.020 1.510 ;
        RECT 36.330 1.340 36.500 1.510 ;
        RECT 36.810 1.340 36.980 1.510 ;
        RECT 37.290 1.340 37.460 1.510 ;
        RECT 37.770 1.340 37.940 1.510 ;
        RECT 38.250 1.340 38.420 1.510 ;
        RECT 38.730 1.340 38.900 1.510 ;
        RECT 39.210 1.340 39.380 1.510 ;
        RECT 39.690 1.340 39.860 1.510 ;
        RECT 40.170 1.340 40.340 1.510 ;
        RECT 40.650 1.340 40.820 1.510 ;
        RECT 41.130 1.340 41.300 1.510 ;
        RECT 41.610 1.340 41.780 1.510 ;
        RECT 42.090 1.340 42.260 1.510 ;
        RECT 42.570 1.340 42.740 1.510 ;
        RECT 43.050 1.340 43.220 1.510 ;
        RECT 43.530 1.340 43.700 1.510 ;
        RECT 44.010 1.340 44.180 1.510 ;
        RECT 44.490 1.340 44.660 1.510 ;
        RECT 44.970 1.340 45.140 1.510 ;
        RECT 45.450 1.340 45.620 1.510 ;
        RECT 45.930 1.340 46.100 1.510 ;
        RECT 46.410 1.340 46.580 1.510 ;
        RECT 46.890 1.340 47.060 1.510 ;
        RECT 47.370 1.340 47.540 1.510 ;
        RECT -2.320 0.310 -2.150 0.480 ;
        RECT -2.160 -0.620 -1.990 -0.450 ;
        RECT -1.630 -0.620 -1.460 -0.450 ;
        RECT -0.720 0.250 -0.550 0.420 ;
        RECT 0.650 0.310 0.820 0.480 ;
        RECT 3.295 0.260 3.470 0.430 ;
        RECT 0.890 -0.240 1.060 -0.070 ;
        RECT -0.760 -0.520 -0.590 -0.350 ;
        RECT 2.110 -0.350 2.280 -0.180 ;
        RECT 1.570 -0.640 1.740 -0.470 ;
        RECT 3.980 -0.350 4.150 -0.180 ;
        RECT 6.170 -0.645 6.340 -0.475 ;
        RECT 7.955 -0.585 8.135 -0.395 ;
        RECT 13.770 0.025 13.940 0.195 ;
        RECT 14.810 -0.645 14.980 -0.475 ;
        RECT 16.595 -0.355 16.765 -0.185 ;
        RECT 22.410 0.430 22.580 0.600 ;
        RECT 23.450 -0.645 23.620 -0.475 ;
        RECT 25.235 -0.355 25.405 -0.185 ;
        RECT 31.060 -0.085 31.230 0.085 ;
        RECT 32.090 -0.645 32.260 -0.475 ;
        RECT 33.875 -0.355 34.045 -0.185 ;
        RECT 39.680 -0.660 39.870 -0.475 ;
        RECT 43.080 -0.030 43.250 0.140 ;
        RECT 40.675 -0.620 40.875 -0.450 ;
        RECT 41.550 -0.555 41.720 -0.385 ;
        RECT 45.910 0.455 46.080 0.625 ;
        RECT 44.130 -0.405 44.310 -0.225 ;
        RECT 45.005 -0.375 45.195 -0.205 ;
        RECT 42.615 -0.930 42.785 -0.760 ;
        RECT 46.465 -0.705 46.645 -0.515 ;
        RECT 47.350 -1.130 47.530 -0.940 ;
        RECT -2.550 -1.990 -2.380 -1.820 ;
        RECT -2.070 -1.990 -1.900 -1.820 ;
        RECT -1.590 -1.990 -1.420 -1.820 ;
        RECT -1.110 -1.990 -0.940 -1.820 ;
        RECT -0.630 -1.990 -0.460 -1.820 ;
        RECT -0.150 -1.990 0.020 -1.820 ;
        RECT 0.330 -1.990 0.500 -1.820 ;
        RECT 0.810 -1.990 0.980 -1.820 ;
        RECT 1.290 -1.990 1.460 -1.820 ;
        RECT 1.770 -1.990 1.940 -1.820 ;
        RECT 2.250 -1.990 2.420 -1.820 ;
        RECT 2.730 -1.990 2.900 -1.820 ;
        RECT 3.210 -1.990 3.380 -1.820 ;
        RECT 3.690 -1.990 3.860 -1.820 ;
        RECT 4.170 -1.990 4.340 -1.820 ;
        RECT 4.650 -1.990 4.820 -1.820 ;
        RECT 5.130 -1.990 5.300 -1.820 ;
        RECT 5.610 -1.990 5.780 -1.820 ;
        RECT 6.090 -1.990 6.260 -1.820 ;
        RECT 6.570 -1.990 6.740 -1.820 ;
        RECT 7.050 -1.990 7.220 -1.820 ;
        RECT 7.530 -1.990 7.700 -1.820 ;
        RECT 8.010 -1.990 8.180 -1.820 ;
        RECT 8.490 -1.990 8.660 -1.820 ;
        RECT 8.970 -1.990 9.140 -1.820 ;
        RECT 9.450 -1.990 9.620 -1.820 ;
        RECT 9.930 -1.990 10.100 -1.820 ;
        RECT 10.410 -1.990 10.580 -1.820 ;
        RECT 10.890 -1.990 11.060 -1.820 ;
        RECT 11.370 -1.990 11.540 -1.820 ;
        RECT 11.850 -1.990 12.020 -1.820 ;
        RECT 12.330 -1.990 12.500 -1.820 ;
        RECT 12.810 -1.990 12.980 -1.820 ;
        RECT 13.290 -1.990 13.460 -1.820 ;
        RECT 13.770 -1.990 13.940 -1.820 ;
        RECT 14.250 -1.990 14.420 -1.820 ;
        RECT 14.730 -1.990 14.900 -1.820 ;
        RECT 15.210 -1.990 15.380 -1.820 ;
        RECT 15.690 -1.990 15.860 -1.820 ;
        RECT 16.170 -1.990 16.340 -1.820 ;
        RECT 16.650 -1.990 16.820 -1.820 ;
        RECT 17.130 -1.990 17.300 -1.820 ;
        RECT 17.610 -1.990 17.780 -1.820 ;
        RECT 18.090 -1.990 18.260 -1.820 ;
        RECT 18.570 -1.990 18.740 -1.820 ;
        RECT 19.050 -1.990 19.220 -1.820 ;
        RECT 19.530 -1.990 19.700 -1.820 ;
        RECT 20.010 -1.990 20.180 -1.820 ;
        RECT 20.490 -1.990 20.660 -1.820 ;
        RECT 20.970 -1.990 21.140 -1.820 ;
        RECT 21.450 -1.990 21.620 -1.820 ;
        RECT 21.930 -1.990 22.100 -1.820 ;
        RECT 22.410 -1.990 22.580 -1.820 ;
        RECT 22.890 -1.990 23.060 -1.820 ;
        RECT 23.370 -1.990 23.540 -1.820 ;
        RECT 23.850 -1.990 24.020 -1.820 ;
        RECT 24.330 -1.990 24.500 -1.820 ;
        RECT 24.810 -1.990 24.980 -1.820 ;
        RECT 25.290 -1.990 25.460 -1.820 ;
        RECT 25.770 -1.990 25.940 -1.820 ;
        RECT 26.250 -1.990 26.420 -1.820 ;
        RECT 26.730 -1.990 26.900 -1.820 ;
        RECT 27.210 -1.990 27.380 -1.820 ;
        RECT 27.690 -1.990 27.860 -1.820 ;
        RECT 28.170 -1.990 28.340 -1.820 ;
        RECT 28.650 -1.990 28.820 -1.820 ;
        RECT 29.130 -1.990 29.300 -1.820 ;
        RECT 29.610 -1.990 29.780 -1.820 ;
        RECT 30.090 -1.990 30.260 -1.820 ;
        RECT 30.570 -1.990 30.740 -1.820 ;
        RECT 31.050 -1.990 31.220 -1.820 ;
        RECT 31.530 -1.990 31.700 -1.820 ;
        RECT 32.010 -1.990 32.180 -1.820 ;
        RECT 32.490 -1.990 32.660 -1.820 ;
        RECT 32.970 -1.990 33.140 -1.820 ;
        RECT 33.450 -1.990 33.620 -1.820 ;
        RECT 33.930 -1.990 34.100 -1.820 ;
        RECT 34.410 -1.990 34.580 -1.820 ;
        RECT 34.890 -1.990 35.060 -1.820 ;
        RECT 35.370 -1.990 35.540 -1.820 ;
        RECT 35.850 -1.990 36.020 -1.820 ;
        RECT 36.330 -1.990 36.500 -1.820 ;
        RECT 36.810 -1.990 36.980 -1.820 ;
        RECT 37.290 -1.990 37.460 -1.820 ;
        RECT 37.770 -1.990 37.940 -1.820 ;
        RECT 38.250 -1.990 38.420 -1.820 ;
        RECT 38.730 -1.990 38.900 -1.820 ;
        RECT 39.210 -1.990 39.380 -1.820 ;
        RECT 39.690 -1.990 39.860 -1.820 ;
        RECT 40.170 -1.990 40.340 -1.820 ;
        RECT 40.650 -1.990 40.820 -1.820 ;
        RECT 41.130 -1.990 41.300 -1.820 ;
        RECT 41.610 -1.990 41.780 -1.820 ;
        RECT 42.090 -1.990 42.260 -1.820 ;
        RECT 42.570 -1.990 42.740 -1.820 ;
        RECT 43.050 -1.990 43.220 -1.820 ;
        RECT 43.530 -1.990 43.700 -1.820 ;
        RECT 44.010 -1.990 44.180 -1.820 ;
        RECT 44.490 -1.990 44.660 -1.820 ;
        RECT 44.970 -1.990 45.140 -1.820 ;
        RECT 45.450 -1.990 45.620 -1.820 ;
        RECT 45.930 -1.990 46.100 -1.820 ;
        RECT 46.410 -1.990 46.580 -1.820 ;
        RECT 46.890 -1.990 47.060 -1.820 ;
        RECT 47.370 -1.990 47.540 -1.820 ;
      LAYER met1 ;
        RECT -2.860 1.180 47.695 1.670 ;
        RECT -2.380 0.490 -2.110 0.520 ;
        RECT 0.650 0.510 0.820 1.180 ;
        RECT 22.350 0.585 22.640 0.660 ;
        RECT 45.845 0.625 46.160 0.685 ;
        RECT 25.175 0.585 41.610 0.595 ;
        RECT -2.380 0.300 -0.520 0.490 ;
        RECT -2.380 0.270 -2.110 0.300 ;
        RECT -0.750 0.180 -0.520 0.300 ;
        RECT 0.620 0.250 0.850 0.510 ;
        RECT 3.240 0.430 3.535 0.500 ;
        RECT 3.240 0.260 8.145 0.430 ;
        RECT 22.350 0.425 41.610 0.585 ;
        RECT 22.350 0.370 22.640 0.425 ;
        RECT 3.240 0.195 3.535 0.260 ;
        RECT 0.840 -0.070 1.110 0.010 ;
        RECT 0.840 -0.240 2.330 -0.070 ;
        RECT -2.250 -0.360 -1.990 -0.345 ;
        RECT -1.625 -0.355 -1.245 -0.325 ;
        RECT -2.250 -0.700 -1.910 -0.360 ;
        RECT -1.700 -0.700 -1.245 -0.355 ;
        RECT -0.875 -0.575 -0.480 -0.290 ;
        RECT 0.840 -0.320 1.110 -0.240 ;
        RECT -2.250 -0.715 -1.990 -0.700 ;
        RECT -1.625 -0.735 -1.245 -0.700 ;
        RECT 0.360 -0.750 0.630 -0.410 ;
        RECT 1.525 -0.735 1.800 -0.380 ;
        RECT 2.060 -0.430 2.330 -0.240 ;
        RECT 3.950 -0.430 4.200 -0.070 ;
        RECT 7.955 -0.350 8.145 0.260 ;
        RECT 13.710 0.195 14.005 0.230 ;
        RECT 13.710 0.025 16.845 0.195 ;
        RECT 13.710 -0.015 14.005 0.025 ;
        RECT 0.410 -1.020 0.580 -0.750 ;
        RECT 3.980 -1.020 4.150 -0.430 ;
        RECT 6.110 -0.735 6.400 -0.385 ;
        RECT 7.900 -0.625 8.185 -0.350 ;
        RECT 7.955 -0.695 8.145 -0.625 ;
        RECT 14.700 -0.760 15.105 -0.355 ;
        RECT 16.520 -0.385 16.845 0.025 ;
        RECT 25.230 -0.135 25.445 0.425 ;
        RECT 30.995 0.085 31.300 0.145 ;
        RECT 30.995 -0.085 34.075 0.085 ;
        RECT 23.355 -0.755 23.740 -0.360 ;
        RECT 25.175 -0.390 25.475 -0.135 ;
        RECT 30.995 -0.145 31.300 -0.085 ;
        RECT 31.970 -0.765 32.375 -0.370 ;
        RECT 33.815 -0.485 34.075 -0.085 ;
        RECT 41.425 -0.300 41.610 0.425 ;
        RECT 45.845 0.455 48.120 0.625 ;
        RECT 45.845 0.395 46.160 0.455 ;
        RECT 43.015 -0.005 45.270 0.185 ;
        RECT 43.015 -0.060 43.330 -0.005 ;
        RECT 41.275 -0.310 42.215 -0.300 ;
        RECT 43.940 -0.310 44.665 -0.160 ;
        RECT 39.650 -0.730 40.945 -0.405 ;
        RECT 41.275 -0.555 44.665 -0.310 ;
        RECT 44.895 -0.415 45.270 -0.005 ;
        RECT 41.275 -0.635 42.215 -0.555 ;
        RECT 42.545 -0.750 42.855 -0.705 ;
        RECT 46.405 -0.750 46.705 -0.430 ;
        RECT 42.545 -0.930 46.705 -0.750 ;
        RECT 42.545 -1.000 42.855 -0.930 ;
        RECT 47.290 -0.950 47.590 -0.880 ;
        RECT 0.410 -1.190 4.150 -1.020 ;
        RECT 47.290 -1.120 48.210 -0.950 ;
        RECT 47.290 -1.195 47.590 -1.120 ;
        RECT -2.860 -2.150 47.695 -1.660 ;
      LAYER via ;
        RECT -2.250 -0.650 -1.990 -0.390 ;
        RECT -1.630 -0.655 -1.370 -0.395 ;
        RECT -0.840 -0.575 -0.535 -0.290 ;
        RECT 1.540 -0.680 1.800 -0.415 ;
        RECT 6.110 -0.705 6.400 -0.415 ;
        RECT 14.775 -0.685 15.035 -0.425 ;
        RECT 23.415 -0.685 23.675 -0.425 ;
        RECT 32.045 -0.690 32.305 -0.425 ;
      LAYER met2 ;
        RECT -2.870 0.150 -2.720 2.005 ;
        RECT -1.820 1.095 -1.670 1.870 ;
        RECT -1.820 0.945 1.690 1.095 ;
        RECT -2.870 0.005 -0.495 0.150 ;
        RECT -0.730 -0.290 -0.495 0.005 ;
        RECT -2.320 -0.735 -1.990 -0.335 ;
        RECT -1.625 -0.365 -1.245 -0.325 ;
        RECT -1.630 -0.685 -1.245 -0.365 ;
        RECT -0.875 -0.575 -0.480 -0.290 ;
        RECT 1.525 -0.360 1.690 0.945 ;
        RECT -1.625 -0.735 -1.245 -0.685 ;
        RECT 1.520 -0.740 1.815 -0.360 ;
        RECT 6.080 -0.780 6.445 -0.340 ;
        RECT 14.700 -0.760 15.105 -0.355 ;
        RECT 23.355 -0.755 23.740 -0.360 ;
        RECT 31.970 -0.765 32.375 -0.370 ;
      LAYER via2 ;
        RECT -2.320 -0.690 -2.035 -0.380 ;
        RECT -1.575 -0.690 -1.295 -0.370 ;
        RECT 1.530 -0.695 1.810 -0.405 ;
        RECT 6.110 -0.735 6.400 -0.385 ;
        RECT 14.745 -0.715 15.060 -0.400 ;
        RECT 23.400 -0.710 23.695 -0.405 ;
        RECT 32.020 -0.720 32.325 -0.420 ;
      LAYER met3 ;
        RECT -2.775 -0.720 -1.990 -0.345 ;
        RECT -1.630 -0.720 -0.845 -0.345 ;
        RECT 1.500 -0.405 1.835 -0.360 ;
        RECT 6.080 -0.395 6.445 -0.340 ;
        RECT 14.700 -0.395 15.105 -0.355 ;
        RECT 23.355 -0.395 23.740 -0.360 ;
        RECT 31.970 -0.395 32.375 -0.370 ;
        RECT 5.865 -0.405 32.375 -0.395 ;
        RECT 1.500 -0.730 32.375 -0.405 ;
        RECT 1.500 -0.740 1.835 -0.730 ;
        RECT 6.080 -0.780 6.445 -0.730 ;
        RECT 14.700 -0.760 15.105 -0.730 ;
        RECT 23.355 -0.755 23.740 -0.730 ;
        RECT 31.970 -0.765 32.375 -0.730 ;
      LAYER via3 ;
        RECT -2.360 -0.700 -2.035 -0.365 ;
        RECT -1.575 -0.695 -1.255 -0.360 ;
      LAYER met4 ;
        RECT -1.370 -0.345 -0.980 -0.210 ;
        RECT -2.380 -0.370 -2.020 -0.355 ;
        RECT -2.775 -0.670 -2.020 -0.370 ;
        RECT -2.380 -0.710 -2.020 -0.670 ;
        RECT -1.590 -0.705 -0.980 -0.345 ;
  END
END comparator_final
MACRO fitler_cell
  CLASS BLOCK ;
  FOREIGN fitler_cell ;
  ORIGIN 26.440 48.250 ;
  SIZE 82.480 BY 79.280 ;
  OBS
      LAYER nwell ;
        RECT 8.410 -15.050 32.630 -14.210 ;
      LAYER li1 ;
        RECT 9.440 -13.670 9.720 -13.500 ;
        RECT 8.850 -14.200 9.180 -14.030 ;
        RECT 8.690 -15.990 8.860 -14.480 ;
        RECT 9.160 -15.200 9.330 -14.480 ;
        RECT 9.500 -14.810 9.670 -13.670 ;
        RECT 17.040 -14.030 17.210 -12.700 ;
        RECT 17.800 -14.030 17.970 -13.040 ;
        RECT 18.370 -13.500 18.540 -13.470 ;
        RECT 18.340 -13.670 18.570 -13.500 ;
        RECT 16.960 -14.200 17.290 -14.030 ;
        RECT 17.720 -14.200 18.050 -14.030 ;
        RECT 9.160 -15.370 9.410 -15.200 ;
        RECT 9.160 -15.990 9.330 -15.370 ;
        RECT 8.930 -16.240 9.100 -16.210 ;
        RECT 8.850 -16.410 9.180 -16.240 ;
        RECT 8.930 -16.440 9.100 -16.410 ;
        RECT 9.500 -17.000 9.670 -15.660 ;
        RECT 16.800 -15.990 16.970 -14.480 ;
        RECT 17.270 -15.990 17.730 -14.480 ;
        RECT 18.030 -15.200 18.200 -14.480 ;
        RECT 18.370 -14.810 18.540 -13.670 ;
        RECT 25.740 -14.030 25.910 -12.700 ;
        RECT 26.500 -14.030 26.670 -13.040 ;
        RECT 27.070 -13.500 27.240 -13.470 ;
        RECT 27.040 -13.670 27.270 -13.500 ;
        RECT 25.660 -14.200 25.990 -14.030 ;
        RECT 26.420 -14.200 26.750 -14.030 ;
        RECT 18.030 -15.370 18.280 -15.200 ;
        RECT 18.030 -15.990 18.200 -15.370 ;
        RECT 16.960 -16.410 17.290 -16.240 ;
        RECT 17.720 -16.410 18.050 -16.240 ;
        RECT 17.040 -17.820 17.210 -16.410 ;
        RECT 17.800 -17.480 17.970 -16.410 ;
        RECT 18.370 -17.000 18.540 -15.660 ;
        RECT 25.500 -15.990 25.670 -14.480 ;
        RECT 25.970 -15.990 26.430 -14.480 ;
        RECT 26.730 -15.200 26.900 -14.480 ;
        RECT 27.070 -14.810 27.240 -13.670 ;
        RECT 31.690 -14.030 31.860 -12.700 ;
        RECT 32.260 -13.500 32.430 -13.470 ;
        RECT 32.230 -13.670 32.460 -13.500 ;
        RECT 31.610 -14.200 31.940 -14.030 ;
        RECT 31.450 -15.190 31.620 -14.480 ;
        RECT 26.730 -15.370 26.980 -15.200 ;
        RECT 31.360 -15.360 31.620 -15.190 ;
        RECT 26.730 -15.990 26.900 -15.370 ;
        RECT 25.660 -16.410 25.990 -16.240 ;
        RECT 26.420 -16.410 26.750 -16.240 ;
        RECT 25.740 -17.820 25.910 -16.410 ;
        RECT 26.500 -17.480 26.670 -16.410 ;
        RECT 27.070 -16.830 27.240 -15.660 ;
        RECT 31.450 -15.990 31.620 -15.360 ;
        RECT 31.920 -15.200 32.090 -14.480 ;
        RECT 32.260 -14.810 32.430 -13.670 ;
        RECT 31.920 -15.370 32.170 -15.200 ;
        RECT 31.920 -15.990 32.090 -15.370 ;
        RECT 31.610 -16.410 31.940 -16.240 ;
        RECT 27.070 -17.000 27.300 -16.830 ;
        RECT 31.690 -17.820 31.860 -16.410 ;
        RECT 32.260 -17.000 32.430 -15.660 ;
      LAYER mcon ;
        RECT 17.040 -12.870 17.210 -12.700 ;
        RECT 9.500 -13.670 9.670 -13.500 ;
        RECT 8.930 -14.200 9.100 -14.030 ;
        RECT 8.690 -15.340 8.860 -15.170 ;
        RECT 25.740 -12.870 25.910 -12.700 ;
        RECT 17.800 -13.250 17.970 -13.080 ;
        RECT 18.370 -13.670 18.540 -13.500 ;
        RECT 9.240 -15.370 9.410 -15.200 ;
        RECT 16.800 -15.340 16.970 -15.170 ;
        RECT 8.930 -16.410 9.100 -16.240 ;
        RECT 17.270 -15.380 17.440 -15.210 ;
        RECT 31.690 -12.870 31.860 -12.700 ;
        RECT 26.500 -13.210 26.670 -13.040 ;
        RECT 27.070 -13.670 27.240 -13.500 ;
        RECT 18.110 -15.370 18.280 -15.200 ;
        RECT 25.500 -15.340 25.670 -15.170 ;
        RECT 25.970 -15.380 26.140 -15.210 ;
        RECT 32.260 -13.670 32.430 -13.500 ;
        RECT 26.810 -15.370 26.980 -15.200 ;
        RECT 17.800 -17.390 17.970 -17.220 ;
        RECT 32.000 -15.370 32.170 -15.200 ;
      LAYER met1 ;
        RECT 16.980 -12.730 17.270 -12.640 ;
        RECT 25.680 -12.730 25.970 -12.640 ;
        RECT 31.630 -12.730 31.920 -12.670 ;
        RECT 16.980 -12.870 55.960 -12.730 ;
        RECT 16.980 -12.900 17.270 -12.870 ;
        RECT 25.680 -12.900 25.970 -12.870 ;
        RECT 31.630 -12.900 31.920 -12.870 ;
        RECT 26.440 -13.040 26.720 -13.010 ;
        RECT 8.930 -13.180 55.960 -13.040 ;
        RECT 8.930 -13.970 9.100 -13.180 ;
        RECT 17.740 -13.300 18.030 -13.180 ;
        RECT 26.440 -13.270 26.720 -13.180 ;
        RECT 9.470 -13.500 9.700 -13.470 ;
        RECT 18.340 -13.500 18.570 -13.470 ;
        RECT 27.040 -13.500 27.270 -13.470 ;
        RECT 32.230 -13.500 32.460 -13.470 ;
        RECT 9.440 -13.670 55.960 -13.500 ;
        RECT 9.470 -13.700 9.700 -13.670 ;
        RECT 18.340 -13.700 18.570 -13.670 ;
        RECT 27.040 -13.700 27.270 -13.670 ;
        RECT 32.230 -13.700 32.460 -13.670 ;
        RECT 8.890 -14.260 9.140 -13.970 ;
        RECT 8.620 -15.120 8.920 -15.110 ;
        RECT 8.590 -15.490 9.020 -15.120 ;
        RECT 9.780 -15.160 10.080 -15.150 ;
        RECT 9.160 -15.400 10.110 -15.160 ;
        RECT 9.680 -15.530 10.110 -15.400 ;
        RECT 16.330 -15.460 17.000 -15.090 ;
        RECT 17.220 -15.160 17.560 -15.130 ;
        RECT 18.650 -15.160 18.950 -15.150 ;
        RECT 17.210 -15.460 17.560 -15.160 ;
        RECT 18.030 -15.400 18.980 -15.160 ;
        RECT 16.360 -15.470 16.660 -15.460 ;
        RECT 17.220 -15.490 17.560 -15.460 ;
        RECT 18.550 -15.530 18.980 -15.400 ;
        RECT 25.030 -15.460 25.700 -15.090 ;
        RECT 25.920 -15.160 26.260 -15.130 ;
        RECT 27.350 -15.160 27.650 -15.150 ;
        RECT 25.910 -15.460 26.260 -15.160 ;
        RECT 26.730 -15.400 27.680 -15.160 ;
        RECT 25.060 -15.470 25.360 -15.460 ;
        RECT 25.920 -15.490 26.260 -15.460 ;
        RECT 27.250 -15.530 27.680 -15.400 ;
        RECT 31.200 -15.460 31.630 -15.090 ;
        RECT 32.540 -15.160 32.840 -15.150 ;
        RECT 31.920 -15.400 32.870 -15.160 ;
        RECT 31.230 -15.470 31.530 -15.460 ;
        RECT 32.440 -15.530 32.870 -15.400 ;
        RECT 54.960 -15.850 55.230 -15.760 ;
        RECT 54.960 -15.990 55.960 -15.850 ;
        RECT 54.960 -16.080 55.230 -15.990 ;
        RECT 8.900 -16.440 9.130 -16.180 ;
        RECT 8.930 -17.340 9.100 -16.440 ;
        RECT 9.450 -16.770 9.720 -16.750 ;
        RECT 18.320 -16.770 18.590 -16.750 ;
        RECT 27.020 -16.770 27.290 -16.750 ;
        RECT 32.210 -16.770 32.480 -16.750 ;
        RECT 9.440 -17.060 9.730 -16.770 ;
        RECT 18.310 -17.060 18.600 -16.770 ;
        RECT 27.010 -17.060 27.300 -16.770 ;
        RECT 32.200 -17.060 32.490 -16.770 ;
        RECT 9.450 -17.080 9.720 -17.060 ;
        RECT 18.320 -17.080 18.590 -17.060 ;
        RECT 27.020 -17.080 27.290 -17.060 ;
        RECT 32.210 -17.080 32.480 -17.060 ;
        RECT 17.710 -17.340 18.030 -17.140 ;
        RECT 26.440 -17.340 26.730 -17.240 ;
        RECT 8.930 -17.480 55.960 -17.340 ;
        RECT 26.440 -17.520 26.730 -17.480 ;
        RECT 16.980 -17.660 17.270 -17.620 ;
        RECT 25.680 -17.660 25.980 -17.620 ;
        RECT 31.630 -17.660 31.920 -17.620 ;
        RECT 16.980 -17.800 55.960 -17.660 ;
        RECT 16.980 -17.880 17.270 -17.800 ;
        RECT 25.680 -17.910 25.980 -17.800 ;
        RECT 31.630 -17.880 31.920 -17.800 ;
      LAYER via ;
        RECT 8.640 -15.400 8.900 -15.140 ;
        RECT 9.800 -15.440 10.060 -15.180 ;
        RECT 16.380 -15.440 16.640 -15.180 ;
        RECT 17.240 -15.440 17.500 -15.180 ;
        RECT 18.670 -15.440 18.930 -15.180 ;
        RECT 25.080 -15.440 25.340 -15.180 ;
        RECT 25.940 -15.440 26.200 -15.180 ;
        RECT 27.370 -15.440 27.630 -15.180 ;
        RECT 31.250 -15.440 31.510 -15.180 ;
        RECT 32.560 -15.440 32.820 -15.180 ;
        RECT 54.960 -16.050 55.230 -15.790 ;
        RECT 9.450 -17.050 9.720 -16.780 ;
        RECT 18.320 -17.050 18.590 -16.780 ;
        RECT 27.020 -17.050 27.290 -16.780 ;
        RECT 32.210 -17.050 32.480 -16.780 ;
      LAYER met2 ;
        RECT 8.590 -15.460 8.950 -15.080 ;
        RECT 9.750 -15.500 10.110 -15.120 ;
        RECT 16.330 -15.500 16.690 -15.120 ;
        RECT 17.180 -15.490 17.560 -15.130 ;
        RECT 18.620 -15.500 18.980 -15.120 ;
        RECT 25.030 -15.500 25.390 -15.120 ;
        RECT 25.880 -15.490 26.260 -15.130 ;
        RECT 27.320 -15.500 27.680 -15.120 ;
        RECT 31.200 -15.500 31.560 -15.120 ;
        RECT 32.510 -15.500 32.870 -15.120 ;
        RECT 54.920 -16.140 55.260 -15.700 ;
        RECT 9.450 -16.780 9.720 -16.750 ;
        RECT 18.320 -16.780 18.590 -16.750 ;
        RECT 27.020 -16.780 27.290 -16.750 ;
        RECT 32.210 -16.780 32.480 -16.750 ;
        RECT 9.400 -17.060 9.780 -16.780 ;
        RECT 18.270 -17.060 18.650 -16.780 ;
        RECT 26.970 -17.060 27.350 -16.780 ;
        RECT 32.160 -17.060 32.540 -16.780 ;
        RECT 9.450 -17.080 9.720 -17.060 ;
        RECT 18.320 -17.080 18.590 -17.060 ;
        RECT 27.020 -17.080 27.290 -17.060 ;
        RECT 32.210 -17.080 32.480 -17.060 ;
      LAYER via2 ;
        RECT 8.630 -15.410 8.910 -15.130 ;
        RECT 9.790 -15.450 10.070 -15.170 ;
        RECT 16.370 -15.450 16.650 -15.170 ;
        RECT 17.230 -15.450 17.510 -15.170 ;
        RECT 18.660 -15.450 18.940 -15.170 ;
        RECT 25.070 -15.450 25.350 -15.170 ;
        RECT 25.930 -15.450 26.210 -15.170 ;
        RECT 27.360 -15.450 27.640 -15.170 ;
        RECT 31.240 -15.450 31.520 -15.170 ;
        RECT 32.550 -15.450 32.830 -15.170 ;
        RECT 54.920 -16.090 55.260 -15.750 ;
        RECT 9.450 -17.060 9.730 -16.780 ;
        RECT 18.320 -17.060 18.600 -16.780 ;
        RECT 27.020 -17.060 27.300 -16.780 ;
        RECT 32.210 -17.060 32.490 -16.780 ;
      LAYER met3 ;
        RECT -26.440 26.900 -23.150 28.530 ;
        RECT -24.830 25.270 -21.720 26.900 ;
        RECT -26.440 23.640 -23.150 25.270 ;
        RECT -24.830 22.010 -21.720 23.640 ;
        RECT -26.440 20.380 -23.150 22.010 ;
        RECT -24.830 18.750 -21.720 20.380 ;
        RECT -26.440 17.120 -23.150 18.750 ;
        RECT -24.830 15.490 -21.720 17.120 ;
        RECT -26.440 13.860 -23.150 15.490 ;
        RECT -24.830 12.230 -21.720 13.860 ;
        RECT -26.440 10.600 -23.150 12.230 ;
        RECT -24.830 8.970 -21.720 10.600 ;
        RECT -26.440 7.340 -23.150 8.970 ;
        RECT -24.830 5.710 -21.720 7.340 ;
        RECT -26.440 4.080 -23.150 5.710 ;
        RECT -24.830 2.450 -21.720 4.080 ;
        RECT -26.440 0.820 -23.150 2.450 ;
        RECT -24.830 -0.810 -21.720 0.820 ;
        RECT -26.440 -2.440 -23.150 -0.810 ;
        RECT -24.830 -4.070 -21.720 -2.440 ;
        RECT -26.440 -5.700 -23.150 -4.070 ;
        RECT -24.830 -7.330 -21.720 -5.700 ;
        RECT -26.440 -8.960 -23.150 -7.330 ;
        RECT -24.830 -8.970 -23.150 -8.960 ;
        RECT -24.830 -10.600 -21.720 -8.970 ;
        RECT -26.440 -12.230 -23.150 -10.600 ;
        RECT -24.830 -13.870 -23.150 -12.230 ;
        RECT -20.920 -12.500 56.040 28.620 ;
        RECT -26.440 -14.430 -23.150 -13.870 ;
        RECT 10.570 -13.060 11.490 -12.500 ;
        RECT -26.440 -15.500 7.820 -14.430 ;
        RECT 8.530 -15.490 9.020 -15.010 ;
        RECT -24.830 -15.790 7.820 -15.500 ;
        RECT 8.580 -15.530 9.020 -15.490 ;
        RECT 9.680 -15.570 10.170 -15.050 ;
        RECT -24.830 -15.830 8.280 -15.790 ;
        RECT -24.830 -16.090 8.390 -15.830 ;
        RECT 7.980 -16.670 8.390 -16.090 ;
        RECT 10.570 -16.670 15.850 -13.060 ;
        RECT 16.270 -15.570 16.760 -15.050 ;
        RECT 17.110 -15.560 17.630 -15.070 ;
        RECT 18.550 -15.570 19.040 -15.050 ;
        RECT 19.360 -16.670 24.640 -14.300 ;
        RECT 24.970 -15.570 25.460 -15.050 ;
        RECT 25.810 -15.560 26.330 -15.070 ;
        RECT 27.250 -15.570 27.740 -15.050 ;
        RECT 28.060 -16.670 30.840 -14.230 ;
        RECT 31.140 -15.570 31.630 -15.050 ;
        RECT 32.440 -15.510 32.930 -15.050 ;
        RECT 32.440 -15.570 32.860 -15.510 ;
        RECT 7.980 -17.160 32.550 -16.670 ;
        RECT 10.570 -17.340 15.850 -17.160 ;
        RECT 10.570 -17.970 11.510 -17.340 ;
        RECT 54.280 -17.970 55.920 -15.020 ;
        RECT -20.930 -48.250 30.190 -17.970 ;
        RECT 30.750 -48.250 56.040 -17.970 ;
      LAYER via3 ;
        RECT -25.800 27.580 -25.480 27.900 ;
        RECT -22.520 25.950 -22.200 26.270 ;
        RECT -25.800 24.320 -25.480 24.640 ;
        RECT -22.520 22.690 -22.200 23.010 ;
        RECT -25.800 21.060 -25.480 21.380 ;
        RECT -22.520 19.430 -22.200 19.750 ;
        RECT -25.800 17.800 -25.480 18.120 ;
        RECT -22.520 16.170 -22.200 16.490 ;
        RECT -25.800 14.540 -25.480 14.860 ;
        RECT -22.520 12.910 -22.200 13.230 ;
        RECT -25.800 11.280 -25.480 11.600 ;
        RECT -22.520 9.650 -22.200 9.970 ;
        RECT -25.800 8.020 -25.480 8.340 ;
        RECT -22.520 6.390 -22.200 6.710 ;
        RECT -25.800 4.760 -25.480 5.080 ;
        RECT -22.520 3.130 -22.200 3.450 ;
        RECT -25.800 1.500 -25.480 1.820 ;
        RECT -22.520 -0.130 -22.200 0.190 ;
        RECT -25.800 -1.760 -25.480 -1.440 ;
        RECT -22.520 -3.390 -22.200 -3.070 ;
        RECT -25.800 -5.020 -25.480 -4.700 ;
        RECT -22.520 -6.650 -22.200 -6.330 ;
        RECT -25.800 -8.280 -25.480 -7.960 ;
        RECT -22.520 -9.920 -22.200 -9.600 ;
        RECT -25.800 -11.550 -25.480 -11.230 ;
        RECT -25.800 -14.820 -25.480 -14.500 ;
        RECT 8.610 -15.430 8.930 -15.110 ;
        RECT 9.770 -15.470 10.090 -15.150 ;
        RECT 16.350 -15.470 16.670 -15.150 ;
        RECT 17.210 -15.470 17.530 -15.150 ;
        RECT 18.640 -15.470 18.960 -15.150 ;
        RECT 25.050 -15.470 25.370 -15.150 ;
        RECT 25.910 -15.470 26.230 -15.150 ;
        RECT 27.340 -15.470 27.660 -15.150 ;
        RECT 31.220 -15.470 31.540 -15.150 ;
        RECT 32.530 -15.470 32.850 -15.150 ;
        RECT 54.920 -16.090 55.260 -15.750 ;
      LAYER met4 ;
        RECT -26.440 26.900 -24.930 28.530 ;
        RECT -26.440 23.640 -24.930 25.270 ;
        RECT -26.440 20.380 -24.930 22.010 ;
        RECT -26.440 17.120 -24.930 18.750 ;
        RECT -26.440 13.860 -24.930 15.490 ;
        RECT -26.440 10.600 -24.930 12.230 ;
        RECT -26.440 7.340 -24.930 8.970 ;
        RECT -26.440 4.080 -24.930 5.710 ;
        RECT -26.440 0.820 -24.930 2.450 ;
        RECT -26.440 -2.440 -24.930 -0.810 ;
        RECT -26.440 -5.700 -24.930 -4.070 ;
        RECT -26.440 -8.960 -24.930 -7.330 ;
        RECT -26.440 -12.230 -24.930 -10.600 ;
        RECT -26.440 -15.500 -24.930 -13.870 ;
        RECT -24.140 -15.110 -23.840 31.030 ;
        RECT -23.090 25.270 -21.720 26.900 ;
        RECT -23.090 22.010 -21.720 23.640 ;
        RECT -23.090 18.750 -21.720 20.380 ;
        RECT -23.090 15.490 -21.720 17.120 ;
        RECT -23.090 12.230 -21.720 13.860 ;
        RECT -23.090 8.970 -21.720 10.600 ;
        RECT -23.090 5.710 -21.720 7.340 ;
        RECT -23.090 2.450 -21.720 4.080 ;
        RECT -23.090 -0.810 -21.720 0.820 ;
        RECT -23.090 -4.070 -21.720 -2.440 ;
        RECT -23.090 -7.330 -21.720 -5.700 ;
        RECT -23.090 -10.600 -21.720 -8.970 ;
        RECT -20.920 -12.500 56.040 28.620 ;
        RECT 8.510 -15.110 8.940 -15.080 ;
        RECT -24.140 -15.410 8.940 -15.110 ;
        RECT 8.510 -15.440 8.940 -15.410 ;
        RECT 9.760 -15.480 11.280 -15.120 ;
        RECT 10.900 -15.500 11.280 -15.480 ;
        RECT 15.180 -15.140 15.560 -15.130 ;
        RECT 15.180 -15.500 16.680 -15.140 ;
        RECT 17.180 -15.480 17.540 -12.500 ;
        RECT 18.630 -15.480 20.100 -15.120 ;
        RECT 24.040 -15.500 25.380 -15.140 ;
        RECT 25.880 -15.480 26.240 -15.130 ;
        RECT 27.330 -15.480 28.760 -15.120 ;
        RECT 15.180 -15.510 15.560 -15.500 ;
        RECT 25.910 -17.970 26.230 -15.480 ;
        RECT 30.240 -15.500 31.550 -15.140 ;
        RECT 32.480 -17.970 32.980 -15.090 ;
        RECT 54.540 -16.460 55.720 -15.280 ;
        RECT -20.930 -48.250 30.190 -17.970 ;
        RECT 30.750 -48.250 56.040 -17.970 ;
      LAYER via4 ;
        RECT -26.220 27.160 -25.040 28.340 ;
        RECT -26.220 23.900 -25.040 25.080 ;
        RECT -26.220 20.640 -25.040 21.820 ;
        RECT -26.220 17.380 -25.040 18.560 ;
        RECT -26.220 14.120 -25.040 15.300 ;
        RECT -26.220 10.860 -25.040 12.040 ;
        RECT -26.220 7.600 -25.040 8.780 ;
        RECT -26.220 4.340 -25.040 5.520 ;
        RECT -26.220 1.080 -25.040 2.260 ;
        RECT -26.220 -2.180 -25.040 -1.000 ;
        RECT -26.220 -5.440 -25.040 -4.260 ;
        RECT -26.220 -8.700 -25.040 -7.520 ;
        RECT -26.220 -11.970 -25.040 -10.790 ;
        RECT -26.220 -15.240 -25.040 -14.060 ;
        RECT -22.940 25.530 -21.760 26.710 ;
        RECT -22.940 22.270 -21.760 23.450 ;
        RECT -22.940 19.010 -21.760 20.190 ;
        RECT -22.940 15.750 -21.760 16.930 ;
        RECT -22.940 12.490 -21.760 13.670 ;
        RECT -22.940 9.230 -21.760 10.410 ;
        RECT -22.940 5.970 -21.760 7.150 ;
        RECT -22.940 2.710 -21.760 3.890 ;
        RECT -22.940 -0.550 -21.760 0.630 ;
        RECT -22.940 -3.810 -21.760 -2.630 ;
        RECT -22.940 -7.070 -21.760 -5.890 ;
        RECT -22.940 -10.340 -21.760 -9.160 ;
      LAYER met5 ;
        RECT -26.440 26.900 -23.150 28.530 ;
        RECT -24.830 25.270 -21.550 26.900 ;
        RECT -26.440 23.640 -23.150 25.270 ;
        RECT -24.830 22.010 -21.550 23.640 ;
        RECT -26.440 20.380 -23.150 22.010 ;
        RECT -24.830 18.750 -21.550 20.380 ;
        RECT -26.440 17.120 -23.150 18.750 ;
        RECT -24.830 15.490 -21.550 17.120 ;
        RECT -26.440 13.860 -23.150 15.490 ;
        RECT -24.830 12.230 -21.550 13.860 ;
        RECT -26.440 10.600 -23.150 12.230 ;
        RECT -24.830 8.970 -21.550 10.600 ;
        RECT -26.440 7.340 -23.150 8.970 ;
        RECT -24.830 5.710 -21.550 7.340 ;
        RECT 7.300 5.920 11.880 10.290 ;
        RECT -26.440 4.080 -23.150 5.710 ;
        RECT 38.090 5.690 42.660 10.130 ;
        RECT -24.830 2.450 -21.550 4.080 ;
        RECT -26.440 0.820 -23.150 2.450 ;
        RECT -24.830 -0.810 -21.550 0.820 ;
        RECT -26.440 -2.440 -23.150 -0.810 ;
        RECT -24.830 -4.070 -21.550 -2.440 ;
        RECT -26.440 -5.700 -23.150 -4.070 ;
        RECT -24.830 -7.330 -21.550 -5.700 ;
        RECT -26.440 -8.960 -23.150 -7.330 ;
        RECT -24.830 -8.970 -23.150 -8.960 ;
        RECT -24.830 -10.600 -21.550 -8.970 ;
        RECT -26.440 -12.230 -23.150 -10.600 ;
        RECT -24.830 -13.870 -23.150 -12.230 ;
        RECT -26.440 -14.430 -23.150 -13.870 ;
        RECT 6.390 -14.430 8.050 -10.730 ;
        RECT -26.440 -15.500 8.390 -14.430 ;
        RECT -24.830 -16.090 8.390 -15.500 ;
        RECT 5.560 -18.390 7.170 -16.090 ;
        RECT 2.180 -20.000 7.170 -18.390 ;
        RECT 54.280 -18.050 55.920 -15.020 ;
        RECT 54.280 -19.780 55.910 -18.050 ;
  END
END fitler_cell
MACRO filter_p_m_fin
  CLASS BLOCK ;
  FOREIGN filter_p_m_fin ;
  ORIGIN 26.420 52.755 ;
  SIZE 167.350 BY 89.955 ;
  PIN compout
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.252000 ;
    PORT
      LAYER li1 ;
        RECT 62.610 -50.010 63.030 -49.680 ;
        RECT 62.860 -51.130 63.030 -50.010 ;
        RECT 67.225 -50.955 67.555 -50.330 ;
        RECT 62.610 -51.460 63.030 -51.130 ;
      LAYER mcon ;
        RECT 62.645 -49.930 62.820 -49.760 ;
        RECT 67.305 -50.775 67.485 -50.585 ;
      LAYER met1 ;
        RECT 62.590 -49.760 62.885 -49.690 ;
        RECT 62.590 -49.930 67.495 -49.760 ;
        RECT 62.590 -49.995 62.885 -49.930 ;
        RECT 67.305 -50.505 67.495 -49.930 ;
        RECT 67.250 -50.910 67.540 -50.505 ;
      LAYER via ;
        RECT 67.265 -50.840 67.525 -50.580 ;
      LAYER met2 ;
        RECT 67.250 -52.755 67.540 -50.480 ;
    END
  END compout
  PIN vssa1
    ANTENNADIFFAREA 9.375800 ;
    PORT
      LAYER pwell ;
        RECT 69.290 -50.950 70.250 -50.730 ;
        RECT 72.520 -50.950 73.890 -50.730 ;
        RECT 77.930 -50.950 78.890 -50.730 ;
        RECT 81.160 -50.950 82.530 -50.730 ;
        RECT 86.570 -50.950 87.530 -50.730 ;
        RECT 89.800 -50.950 91.170 -50.730 ;
        RECT 95.210 -50.950 96.170 -50.730 ;
        RECT 98.440 -50.950 99.810 -50.730 ;
        RECT 66.450 -51.235 73.890 -50.950 ;
        RECT 75.090 -50.955 82.530 -50.950 ;
        RECT 75.090 -51.235 82.645 -50.955 ;
        RECT 83.730 -50.970 91.170 -50.950 ;
        RECT 83.730 -51.235 91.295 -50.970 ;
        RECT 92.370 -50.985 99.810 -50.950 ;
        RECT 92.370 -51.235 99.890 -50.985 ;
        RECT 65.290 -51.240 73.890 -51.235 ;
        RECT 73.930 -51.240 99.890 -51.235 ;
        RECT 65.290 -51.835 99.890 -51.240 ;
        RECT 65.290 -51.850 82.530 -51.835 ;
        RECT 82.570 -51.850 99.890 -51.835 ;
        RECT 99.925 -51.850 103.150 -50.780 ;
        RECT 103.535 -51.850 105.405 -50.890 ;
        RECT 105.610 -51.850 107.040 -50.890 ;
        RECT 65.285 -52.095 107.045 -51.850 ;
        RECT 103.805 -52.130 104.145 -52.095 ;
      LAYER li1 ;
        RECT 9.520 -17.000 9.690 -15.660 ;
        RECT 18.390 -17.000 18.560 -15.660 ;
        RECT 27.090 -16.830 27.260 -15.660 ;
        RECT 27.090 -17.000 27.320 -16.830 ;
        RECT 32.280 -17.000 32.450 -15.660 ;
        RECT 82.060 -17.000 82.230 -15.660 ;
        RECT 87.250 -16.830 87.420 -15.660 ;
        RECT 87.190 -17.000 87.420 -16.830 ;
        RECT 95.950 -17.000 96.120 -15.660 ;
        RECT 104.820 -17.000 104.990 -15.660 ;
        RECT 59.020 -51.520 59.250 -51.190 ;
        RECT 59.960 -51.460 60.210 -51.130 ;
        RECT 60.840 -51.460 61.090 -51.130 ;
        RECT 59.080 -52.010 59.250 -51.520 ;
        RECT 60.010 -52.010 60.180 -51.460 ;
        RECT 60.890 -52.010 61.060 -51.460 ;
        RECT 61.260 -52.010 61.430 -51.130 ;
        RECT 62.160 -51.460 62.410 -51.130 ;
        RECT 62.210 -52.010 62.380 -51.460 ;
        RECT 63.200 -52.010 63.370 -51.250 ;
        RECT 64.030 -51.460 64.280 -51.130 ;
        RECT 64.080 -52.010 64.250 -51.460 ;
        RECT 65.380 -52.010 65.710 -51.425 ;
        RECT 67.040 -52.010 67.320 -51.125 ;
        RECT 68.805 -52.010 69.710 -51.210 ;
        RECT 71.285 -52.010 71.805 -51.150 ;
        RECT 72.620 -52.010 72.900 -50.840 ;
        RECT 73.505 -52.010 73.740 -50.840 ;
        RECT 74.020 -52.010 74.350 -51.425 ;
        RECT 75.680 -52.010 75.960 -51.125 ;
        RECT 77.445 -52.010 78.350 -51.210 ;
        RECT 79.925 -52.010 80.445 -51.150 ;
        RECT 81.260 -52.010 81.540 -50.840 ;
        RECT 82.145 -52.010 82.380 -50.840 ;
        RECT 82.660 -52.010 82.990 -51.425 ;
        RECT 84.320 -52.010 84.600 -51.125 ;
        RECT 86.085 -52.010 86.990 -51.210 ;
        RECT 88.565 -52.010 89.085 -51.150 ;
        RECT 89.900 -52.010 90.180 -50.840 ;
        RECT 90.785 -52.010 91.020 -50.840 ;
        RECT 91.300 -52.010 91.630 -51.425 ;
        RECT 92.960 -52.010 93.240 -51.125 ;
        RECT 94.725 -52.010 95.630 -51.210 ;
        RECT 97.205 -52.010 97.725 -51.150 ;
        RECT 98.540 -52.010 98.820 -50.840 ;
        RECT 99.425 -52.010 99.660 -50.840 ;
        RECT 100.015 -52.010 100.275 -51.055 ;
        RECT 100.875 -52.010 101.205 -51.395 ;
        RECT 102.810 -52.010 103.060 -51.035 ;
        RECT 103.870 -52.010 104.080 -51.745 ;
        RECT 104.415 -52.010 104.785 -51.115 ;
        RECT 106.190 -52.010 106.520 -51.415 ;
        RECT 56.490 -52.180 107.045 -52.010 ;
      LAYER mcon ;
        RECT 87.250 -17.000 87.420 -16.830 ;
        RECT 56.800 -52.180 56.970 -52.010 ;
        RECT 57.280 -52.180 57.450 -52.010 ;
        RECT 57.760 -52.180 57.930 -52.010 ;
        RECT 58.240 -52.180 58.410 -52.010 ;
        RECT 58.720 -52.180 58.890 -52.010 ;
        RECT 59.200 -52.180 59.370 -52.010 ;
        RECT 59.680 -52.180 59.850 -52.010 ;
        RECT 60.160 -52.180 60.330 -52.010 ;
        RECT 60.640 -52.180 60.810 -52.010 ;
        RECT 61.120 -52.180 61.290 -52.010 ;
        RECT 61.600 -52.180 61.770 -52.010 ;
        RECT 62.080 -52.180 62.250 -52.010 ;
        RECT 62.560 -52.180 62.730 -52.010 ;
        RECT 63.040 -52.180 63.210 -52.010 ;
        RECT 63.520 -52.180 63.690 -52.010 ;
        RECT 64.000 -52.180 64.170 -52.010 ;
        RECT 64.480 -52.180 64.650 -52.010 ;
        RECT 64.960 -52.180 65.130 -52.010 ;
        RECT 65.440 -52.180 65.610 -52.010 ;
        RECT 65.920 -52.180 66.090 -52.010 ;
        RECT 66.400 -52.180 66.570 -52.010 ;
        RECT 66.880 -52.180 67.050 -52.010 ;
        RECT 67.360 -52.180 67.530 -52.010 ;
        RECT 67.840 -52.180 68.010 -52.010 ;
        RECT 68.320 -52.180 68.490 -52.010 ;
        RECT 68.800 -52.180 68.970 -52.010 ;
        RECT 69.280 -52.180 69.450 -52.010 ;
        RECT 69.760 -52.180 69.930 -52.010 ;
        RECT 70.240 -52.180 70.410 -52.010 ;
        RECT 70.720 -52.180 70.890 -52.010 ;
        RECT 71.200 -52.180 71.370 -52.010 ;
        RECT 71.680 -52.180 71.850 -52.010 ;
        RECT 72.160 -52.180 72.330 -52.010 ;
        RECT 72.640 -52.180 72.810 -52.010 ;
        RECT 73.120 -52.180 73.290 -52.010 ;
        RECT 73.600 -52.180 73.770 -52.010 ;
        RECT 74.080 -52.180 74.250 -52.010 ;
        RECT 74.560 -52.180 74.730 -52.010 ;
        RECT 75.040 -52.180 75.210 -52.010 ;
        RECT 75.520 -52.180 75.690 -52.010 ;
        RECT 76.000 -52.180 76.170 -52.010 ;
        RECT 76.480 -52.180 76.650 -52.010 ;
        RECT 76.960 -52.180 77.130 -52.010 ;
        RECT 77.440 -52.180 77.610 -52.010 ;
        RECT 77.920 -52.180 78.090 -52.010 ;
        RECT 78.400 -52.180 78.570 -52.010 ;
        RECT 78.880 -52.180 79.050 -52.010 ;
        RECT 79.360 -52.180 79.530 -52.010 ;
        RECT 79.840 -52.180 80.010 -52.010 ;
        RECT 80.320 -52.180 80.490 -52.010 ;
        RECT 80.800 -52.180 80.970 -52.010 ;
        RECT 81.280 -52.180 81.450 -52.010 ;
        RECT 81.760 -52.180 81.930 -52.010 ;
        RECT 82.240 -52.180 82.410 -52.010 ;
        RECT 82.720 -52.180 82.890 -52.010 ;
        RECT 83.200 -52.180 83.370 -52.010 ;
        RECT 83.680 -52.180 83.850 -52.010 ;
        RECT 84.160 -52.180 84.330 -52.010 ;
        RECT 84.640 -52.180 84.810 -52.010 ;
        RECT 85.120 -52.180 85.290 -52.010 ;
        RECT 85.600 -52.180 85.770 -52.010 ;
        RECT 86.080 -52.180 86.250 -52.010 ;
        RECT 86.560 -52.180 86.730 -52.010 ;
        RECT 87.040 -52.180 87.210 -52.010 ;
        RECT 87.520 -52.180 87.690 -52.010 ;
        RECT 88.000 -52.180 88.170 -52.010 ;
        RECT 88.480 -52.180 88.650 -52.010 ;
        RECT 88.960 -52.180 89.130 -52.010 ;
        RECT 89.440 -52.180 89.610 -52.010 ;
        RECT 89.920 -52.180 90.090 -52.010 ;
        RECT 90.400 -52.180 90.570 -52.010 ;
        RECT 90.880 -52.180 91.050 -52.010 ;
        RECT 91.360 -52.180 91.530 -52.010 ;
        RECT 91.840 -52.180 92.010 -52.010 ;
        RECT 92.320 -52.180 92.490 -52.010 ;
        RECT 92.800 -52.180 92.970 -52.010 ;
        RECT 93.280 -52.180 93.450 -52.010 ;
        RECT 93.760 -52.180 93.930 -52.010 ;
        RECT 94.240 -52.180 94.410 -52.010 ;
        RECT 94.720 -52.180 94.890 -52.010 ;
        RECT 95.200 -52.180 95.370 -52.010 ;
        RECT 95.680 -52.180 95.850 -52.010 ;
        RECT 96.160 -52.180 96.330 -52.010 ;
        RECT 96.640 -52.180 96.810 -52.010 ;
        RECT 97.120 -52.180 97.290 -52.010 ;
        RECT 97.600 -52.180 97.770 -52.010 ;
        RECT 98.080 -52.180 98.250 -52.010 ;
        RECT 98.560 -52.180 98.730 -52.010 ;
        RECT 99.040 -52.180 99.210 -52.010 ;
        RECT 99.520 -52.180 99.690 -52.010 ;
        RECT 100.000 -52.180 100.170 -52.010 ;
        RECT 100.480 -52.180 100.650 -52.010 ;
        RECT 100.960 -52.180 101.130 -52.010 ;
        RECT 101.440 -52.180 101.610 -52.010 ;
        RECT 101.920 -52.180 102.090 -52.010 ;
        RECT 102.400 -52.180 102.570 -52.010 ;
        RECT 102.880 -52.180 103.050 -52.010 ;
        RECT 103.360 -52.180 103.530 -52.010 ;
        RECT 103.840 -52.180 104.010 -52.010 ;
        RECT 104.320 -52.180 104.490 -52.010 ;
        RECT 104.800 -52.180 104.970 -52.010 ;
        RECT 105.280 -52.180 105.450 -52.010 ;
        RECT 105.760 -52.180 105.930 -52.010 ;
        RECT 106.240 -52.180 106.410 -52.010 ;
        RECT 106.720 -52.180 106.890 -52.010 ;
      LAYER met1 ;
        RECT 9.470 -16.770 9.740 -16.750 ;
        RECT 18.340 -16.770 18.610 -16.750 ;
        RECT 27.040 -16.770 27.310 -16.750 ;
        RECT 32.230 -16.770 32.500 -16.750 ;
        RECT 82.010 -16.770 82.280 -16.750 ;
        RECT 87.200 -16.770 87.470 -16.750 ;
        RECT 95.900 -16.770 96.170 -16.750 ;
        RECT 104.770 -16.770 105.040 -16.750 ;
        RECT 9.460 -17.060 9.750 -16.770 ;
        RECT 18.330 -17.060 18.620 -16.770 ;
        RECT 27.030 -17.060 27.320 -16.770 ;
        RECT 32.220 -17.060 32.510 -16.770 ;
        RECT 82.000 -17.060 82.290 -16.770 ;
        RECT 87.190 -17.060 87.480 -16.770 ;
        RECT 95.890 -17.060 96.180 -16.770 ;
        RECT 104.760 -17.060 105.050 -16.770 ;
        RECT 9.470 -17.080 9.740 -17.060 ;
        RECT 18.340 -17.080 18.610 -17.060 ;
        RECT 27.040 -17.080 27.310 -17.060 ;
        RECT 32.230 -17.080 32.500 -17.060 ;
        RECT 82.010 -17.080 82.280 -17.060 ;
        RECT 87.200 -17.080 87.470 -17.060 ;
        RECT 95.900 -17.080 96.170 -17.060 ;
        RECT 104.770 -17.080 105.040 -17.060 ;
        RECT 56.490 -52.340 107.045 -51.850 ;
      LAYER via ;
        RECT 9.470 -17.050 9.740 -16.780 ;
        RECT 18.340 -17.050 18.610 -16.780 ;
        RECT 27.040 -17.050 27.310 -16.780 ;
        RECT 32.230 -17.050 32.500 -16.780 ;
        RECT 82.010 -17.050 82.280 -16.780 ;
        RECT 87.200 -17.050 87.470 -16.780 ;
        RECT 95.900 -17.050 96.170 -16.780 ;
        RECT 104.770 -17.050 105.040 -16.780 ;
        RECT 97.360 -52.195 97.620 -51.935 ;
      LAYER met2 ;
        RECT 9.470 -16.780 9.740 -16.750 ;
        RECT 18.340 -16.780 18.610 -16.750 ;
        RECT 27.040 -16.780 27.310 -16.750 ;
        RECT 32.230 -16.780 32.500 -16.750 ;
        RECT 82.010 -16.780 82.280 -16.750 ;
        RECT 87.200 -16.780 87.470 -16.750 ;
        RECT 95.900 -16.780 96.170 -16.750 ;
        RECT 104.770 -16.780 105.040 -16.750 ;
        RECT 9.420 -17.060 9.800 -16.780 ;
        RECT 18.290 -17.060 18.670 -16.780 ;
        RECT 26.990 -17.060 27.370 -16.780 ;
        RECT 32.180 -17.060 32.560 -16.780 ;
        RECT 81.950 -17.060 82.330 -16.780 ;
        RECT 87.140 -17.060 87.520 -16.780 ;
        RECT 95.840 -17.060 96.220 -16.780 ;
        RECT 104.710 -17.060 105.090 -16.780 ;
        RECT 9.470 -17.080 9.740 -17.060 ;
        RECT 18.340 -17.080 18.610 -17.060 ;
        RECT 27.040 -17.080 27.310 -17.060 ;
        RECT 32.230 -17.080 32.500 -17.060 ;
        RECT 82.010 -17.080 82.280 -17.060 ;
        RECT 87.200 -17.080 87.470 -17.060 ;
        RECT 95.900 -17.080 96.170 -17.060 ;
        RECT 104.770 -17.080 105.040 -17.060 ;
        RECT 97.295 -52.265 97.680 -51.890 ;
      LAYER via2 ;
        RECT 9.470 -17.060 9.750 -16.780 ;
        RECT 18.340 -17.060 18.620 -16.780 ;
        RECT 27.040 -17.060 27.320 -16.780 ;
        RECT 32.230 -17.060 32.510 -16.780 ;
        RECT 82.000 -17.060 82.280 -16.780 ;
        RECT 87.190 -17.060 87.470 -16.780 ;
        RECT 95.890 -17.060 96.170 -16.780 ;
        RECT 104.760 -17.060 105.040 -16.780 ;
        RECT 97.345 -52.215 97.625 -51.935 ;
      LAYER met3 ;
        RECT -26.420 28.530 -25.480 30.060 ;
        RECT -26.420 26.900 -23.130 28.530 ;
        RECT -20.900 28.375 56.060 28.620 ;
        RECT 58.450 28.375 135.410 28.620 ;
        RECT -20.900 27.560 135.410 28.375 ;
        RECT -24.810 25.270 -21.700 26.900 ;
        RECT -26.420 23.640 -23.130 25.270 ;
        RECT -20.900 25.100 56.060 27.560 ;
        RECT 58.450 25.100 135.410 27.560 ;
        RECT 137.640 26.900 140.930 28.530 ;
        RECT 136.210 25.270 139.320 26.900 ;
        RECT -20.900 24.285 135.410 25.100 ;
        RECT -24.810 22.010 -21.700 23.640 ;
        RECT -26.420 20.380 -23.130 22.010 ;
        RECT -24.810 18.750 -21.700 20.380 ;
        RECT -26.420 17.120 -23.130 18.750 ;
        RECT -20.900 17.730 56.060 24.285 ;
        RECT 58.450 17.730 135.410 24.285 ;
        RECT 137.640 23.640 140.930 25.270 ;
        RECT 136.210 22.010 139.320 23.640 ;
        RECT 137.640 20.380 140.930 22.010 ;
        RECT 136.210 18.750 139.320 20.380 ;
        RECT -24.810 15.490 -21.700 17.120 ;
        RECT -20.900 16.365 135.410 17.730 ;
        RECT 137.640 17.120 140.930 18.750 ;
        RECT -26.420 13.860 -23.130 15.490 ;
        RECT -24.810 12.230 -21.700 13.860 ;
        RECT -26.420 10.600 -23.130 12.230 ;
        RECT -20.900 11.450 56.060 16.365 ;
        RECT 58.450 11.450 135.410 16.365 ;
        RECT 136.210 15.490 139.320 17.120 ;
        RECT 137.640 13.860 140.930 15.490 ;
        RECT 136.210 12.230 139.320 13.860 ;
        RECT -24.810 8.970 -21.700 10.600 ;
        RECT -20.900 10.085 135.410 11.450 ;
        RECT 137.640 10.600 140.930 12.230 ;
        RECT -26.420 7.340 -23.130 8.970 ;
        RECT -24.810 5.710 -21.700 7.340 ;
        RECT -26.420 4.080 -23.130 5.710 ;
        RECT -20.900 5.465 56.060 10.085 ;
        RECT 58.450 5.465 135.410 10.085 ;
        RECT 136.210 8.970 139.320 10.600 ;
        RECT 137.640 7.340 140.930 8.970 ;
        RECT 136.210 5.710 139.320 7.340 ;
        RECT -20.900 4.100 135.410 5.465 ;
        RECT -24.810 2.450 -21.700 4.080 ;
        RECT -26.420 0.820 -23.130 2.450 ;
        RECT -24.810 -0.810 -21.700 0.820 ;
        RECT -20.900 -0.175 56.060 4.100 ;
        RECT 58.450 -0.175 135.410 4.100 ;
        RECT 137.640 4.080 140.930 5.710 ;
        RECT 136.210 2.450 139.320 4.080 ;
        RECT 137.640 0.820 140.930 2.450 ;
        RECT -26.420 -2.440 -23.130 -0.810 ;
        RECT -20.900 -1.540 135.410 -0.175 ;
        RECT 136.210 -0.810 139.320 0.820 ;
        RECT -24.810 -4.070 -21.700 -2.440 ;
        RECT -26.420 -5.700 -23.130 -4.070 ;
        RECT -20.900 -5.670 56.060 -1.540 ;
        RECT 58.450 -5.670 135.410 -1.540 ;
        RECT 137.640 -2.440 140.930 -0.810 ;
        RECT 136.210 -4.070 139.320 -2.440 ;
        RECT -24.810 -7.330 -21.700 -5.700 ;
        RECT -20.900 -7.035 135.410 -5.670 ;
        RECT 137.640 -5.700 140.930 -4.070 ;
        RECT -26.420 -8.960 -23.130 -7.330 ;
        RECT -24.810 -8.970 -23.130 -8.960 ;
        RECT -24.810 -10.600 -21.700 -8.970 ;
        RECT -26.420 -12.230 -23.130 -10.600 ;
        RECT -24.810 -13.870 -23.130 -12.230 ;
        RECT -20.900 -12.500 56.060 -7.035 ;
        RECT 58.450 -12.500 135.410 -7.035 ;
        RECT 136.210 -7.330 139.320 -5.700 ;
        RECT 137.640 -8.960 140.930 -7.330 ;
        RECT 137.640 -8.970 139.320 -8.960 ;
        RECT 136.210 -10.600 139.320 -8.970 ;
        RECT 137.640 -12.230 140.930 -10.600 ;
        RECT -26.420 -14.430 -23.130 -13.870 ;
        RECT 10.590 -13.060 11.510 -12.500 ;
        RECT 103.000 -13.060 103.920 -12.500 ;
        RECT -26.420 -15.500 7.840 -14.430 ;
        RECT -24.810 -15.790 7.840 -15.500 ;
        RECT -24.810 -15.830 8.300 -15.790 ;
        RECT -24.810 -16.090 8.410 -15.830 ;
        RECT 8.000 -16.670 8.410 -16.090 ;
        RECT 10.590 -16.670 15.870 -13.060 ;
        RECT 19.380 -16.670 24.660 -14.300 ;
        RECT 28.080 -16.670 30.860 -14.230 ;
        RECT 83.650 -16.670 86.430 -14.230 ;
        RECT 89.850 -16.670 95.130 -14.300 ;
        RECT 98.640 -16.670 103.920 -13.060 ;
        RECT 137.640 -13.870 139.320 -12.230 ;
        RECT 137.640 -14.430 140.930 -13.870 ;
        RECT 106.670 -15.500 140.930 -14.430 ;
        RECT 106.670 -15.790 139.320 -15.500 ;
        RECT 106.210 -15.830 139.320 -15.790 ;
        RECT 106.100 -16.090 139.320 -15.830 ;
        RECT 106.100 -16.670 106.510 -16.090 ;
        RECT 8.000 -17.160 32.570 -16.670 ;
        RECT 81.940 -17.160 106.510 -16.670 ;
        RECT 10.590 -17.340 15.870 -17.160 ;
        RECT 98.640 -17.340 103.920 -17.160 ;
        RECT 10.590 -17.970 11.530 -17.340 ;
        RECT 102.980 -17.970 103.920 -17.340 ;
        RECT -20.910 -48.250 30.210 -17.970 ;
        RECT 84.300 -48.250 135.420 -17.970 ;
        RECT 97.075 -52.340 97.915 -48.250 ;
      LAYER via3 ;
        RECT -25.780 27.580 -25.460 27.900 ;
        RECT -22.500 25.950 -22.180 26.270 ;
        RECT -25.780 24.320 -25.460 24.640 ;
        RECT 139.970 27.580 140.290 27.900 ;
        RECT 136.690 25.950 137.010 26.270 ;
        RECT -22.500 22.690 -22.180 23.010 ;
        RECT -25.780 21.060 -25.460 21.380 ;
        RECT -22.500 19.430 -22.180 19.750 ;
        RECT -25.780 17.800 -25.460 18.120 ;
        RECT 139.970 24.320 140.290 24.640 ;
        RECT 136.690 22.690 137.010 23.010 ;
        RECT 139.970 21.060 140.290 21.380 ;
        RECT 136.690 19.430 137.010 19.750 ;
        RECT -22.500 16.170 -22.180 16.490 ;
        RECT 139.970 17.800 140.290 18.120 ;
        RECT -25.780 14.540 -25.460 14.860 ;
        RECT -22.500 12.910 -22.180 13.230 ;
        RECT -25.780 11.280 -25.460 11.600 ;
        RECT 136.690 16.170 137.010 16.490 ;
        RECT 139.970 14.540 140.290 14.860 ;
        RECT 136.690 12.910 137.010 13.230 ;
        RECT -22.500 9.650 -22.180 9.970 ;
        RECT 139.970 11.280 140.290 11.600 ;
        RECT -25.780 8.020 -25.460 8.340 ;
        RECT -22.500 6.390 -22.180 6.710 ;
        RECT -25.780 4.760 -25.460 5.080 ;
        RECT 136.690 9.650 137.010 9.970 ;
        RECT 139.970 8.020 140.290 8.340 ;
        RECT 136.690 6.390 137.010 6.710 ;
        RECT -22.500 3.130 -22.180 3.450 ;
        RECT -25.780 1.500 -25.460 1.820 ;
        RECT -22.500 -0.130 -22.180 0.190 ;
        RECT 139.970 4.760 140.290 5.080 ;
        RECT 136.690 3.130 137.010 3.450 ;
        RECT 139.970 1.500 140.290 1.820 ;
        RECT -25.780 -1.760 -25.460 -1.440 ;
        RECT 136.690 -0.130 137.010 0.190 ;
        RECT -22.500 -3.390 -22.180 -3.070 ;
        RECT -25.780 -5.020 -25.460 -4.700 ;
        RECT 139.970 -1.760 140.290 -1.440 ;
        RECT 136.690 -3.390 137.010 -3.070 ;
        RECT -22.500 -6.650 -22.180 -6.330 ;
        RECT 139.970 -5.020 140.290 -4.700 ;
        RECT -25.780 -8.280 -25.460 -7.960 ;
        RECT -22.500 -9.920 -22.180 -9.600 ;
        RECT -25.780 -11.550 -25.460 -11.230 ;
        RECT 136.690 -6.650 137.010 -6.330 ;
        RECT 139.970 -8.280 140.290 -7.960 ;
        RECT 136.690 -9.920 137.010 -9.600 ;
        RECT 139.970 -11.550 140.290 -11.230 ;
        RECT -25.780 -14.820 -25.460 -14.500 ;
        RECT 139.970 -14.820 140.290 -14.500 ;
      LAYER met4 ;
        RECT -26.420 26.900 -24.910 28.530 ;
        RECT 139.420 26.900 140.930 28.530 ;
        RECT -23.070 25.270 -21.700 26.900 ;
        RECT 136.210 25.270 137.580 26.900 ;
        RECT -26.420 23.640 -24.910 25.270 ;
        RECT 139.420 23.640 140.930 25.270 ;
        RECT -23.070 22.010 -21.700 23.640 ;
        RECT 136.210 22.010 137.580 23.640 ;
        RECT -26.420 20.380 -24.910 22.010 ;
        RECT 139.420 20.380 140.930 22.010 ;
        RECT -23.070 18.750 -21.700 20.380 ;
        RECT 136.210 18.750 137.580 20.380 ;
        RECT -26.420 17.120 -24.910 18.750 ;
        RECT 139.420 17.120 140.930 18.750 ;
        RECT -23.070 15.490 -21.700 17.120 ;
        RECT 136.210 15.490 137.580 17.120 ;
        RECT -26.420 13.860 -24.910 15.490 ;
        RECT 139.420 13.860 140.930 15.490 ;
        RECT -23.070 12.230 -21.700 13.860 ;
        RECT 136.210 12.230 137.580 13.860 ;
        RECT -26.420 10.600 -24.910 12.230 ;
        RECT 139.420 10.600 140.930 12.230 ;
        RECT -23.070 8.970 -21.700 10.600 ;
        RECT 136.210 8.970 137.580 10.600 ;
        RECT -26.420 7.340 -24.910 8.970 ;
        RECT 139.420 7.340 140.930 8.970 ;
        RECT -23.070 5.710 -21.700 7.340 ;
        RECT 136.210 5.710 137.580 7.340 ;
        RECT -26.420 4.080 -24.910 5.710 ;
        RECT 139.420 4.080 140.930 5.710 ;
        RECT -23.070 2.450 -21.700 4.080 ;
        RECT 136.210 2.450 137.580 4.080 ;
        RECT -26.420 0.820 -24.910 2.450 ;
        RECT 139.420 0.820 140.930 2.450 ;
        RECT -23.070 -0.810 -21.700 0.820 ;
        RECT 136.210 -0.810 137.580 0.820 ;
        RECT -26.420 -2.440 -24.910 -0.810 ;
        RECT 139.420 -2.440 140.930 -0.810 ;
        RECT -23.070 -4.070 -21.700 -2.440 ;
        RECT 136.210 -4.070 137.580 -2.440 ;
        RECT -26.420 -5.700 -24.910 -4.070 ;
        RECT 139.420 -5.700 140.930 -4.070 ;
        RECT -23.070 -7.330 -21.700 -5.700 ;
        RECT 136.210 -7.330 137.580 -5.700 ;
        RECT -26.420 -8.960 -24.910 -7.330 ;
        RECT 139.420 -8.960 140.930 -7.330 ;
        RECT -23.070 -10.600 -21.700 -8.970 ;
        RECT 136.210 -10.600 137.580 -8.970 ;
        RECT -26.420 -12.230 -24.910 -10.600 ;
        RECT 139.420 -12.230 140.930 -10.600 ;
        RECT -26.420 -15.500 -24.910 -13.870 ;
        RECT 139.420 -15.500 140.930 -13.870 ;
      LAYER via4 ;
        RECT -26.200 27.160 -25.020 28.340 ;
        RECT 139.530 27.160 140.710 28.340 ;
        RECT -22.920 25.530 -21.740 26.710 ;
        RECT 136.250 25.530 137.430 26.710 ;
        RECT -26.200 23.900 -25.020 25.080 ;
        RECT 139.530 23.900 140.710 25.080 ;
        RECT -22.920 22.270 -21.740 23.450 ;
        RECT 136.250 22.270 137.430 23.450 ;
        RECT -26.200 20.640 -25.020 21.820 ;
        RECT 139.530 20.640 140.710 21.820 ;
        RECT -22.920 19.010 -21.740 20.190 ;
        RECT 136.250 19.010 137.430 20.190 ;
        RECT -26.200 17.380 -25.020 18.560 ;
        RECT 139.530 17.380 140.710 18.560 ;
        RECT -22.920 15.750 -21.740 16.930 ;
        RECT 136.250 15.750 137.430 16.930 ;
        RECT -26.200 14.120 -25.020 15.300 ;
        RECT 139.530 14.120 140.710 15.300 ;
        RECT -22.920 12.490 -21.740 13.670 ;
        RECT 136.250 12.490 137.430 13.670 ;
        RECT -26.200 10.860 -25.020 12.040 ;
        RECT 139.530 10.860 140.710 12.040 ;
        RECT -22.920 9.230 -21.740 10.410 ;
        RECT 136.250 9.230 137.430 10.410 ;
        RECT -26.200 7.600 -25.020 8.780 ;
        RECT 139.530 7.600 140.710 8.780 ;
        RECT -22.920 5.970 -21.740 7.150 ;
        RECT 136.250 5.970 137.430 7.150 ;
        RECT -26.200 4.340 -25.020 5.520 ;
        RECT 139.530 4.340 140.710 5.520 ;
        RECT -22.920 2.710 -21.740 3.890 ;
        RECT 136.250 2.710 137.430 3.890 ;
        RECT -26.200 1.080 -25.020 2.260 ;
        RECT 139.530 1.080 140.710 2.260 ;
        RECT -22.920 -0.550 -21.740 0.630 ;
        RECT 136.250 -0.550 137.430 0.630 ;
        RECT -26.200 -2.180 -25.020 -1.000 ;
        RECT 139.530 -2.180 140.710 -1.000 ;
        RECT -22.920 -3.810 -21.740 -2.630 ;
        RECT 136.250 -3.810 137.430 -2.630 ;
        RECT -26.200 -5.440 -25.020 -4.260 ;
        RECT 139.530 -5.440 140.710 -4.260 ;
        RECT -22.920 -7.070 -21.740 -5.890 ;
        RECT 136.250 -7.070 137.430 -5.890 ;
        RECT -26.200 -8.700 -25.020 -7.520 ;
        RECT 139.530 -8.700 140.710 -7.520 ;
        RECT -22.920 -10.340 -21.740 -9.160 ;
        RECT 136.250 -10.340 137.430 -9.160 ;
        RECT -26.200 -11.970 -25.020 -10.790 ;
        RECT 139.530 -11.970 140.710 -10.790 ;
        RECT -26.200 -15.240 -25.020 -14.060 ;
        RECT 139.530 -15.240 140.710 -14.060 ;
      LAYER met5 ;
        RECT -26.420 26.900 -23.130 28.530 ;
        RECT 137.640 26.900 140.930 28.530 ;
        RECT -24.810 25.270 -21.530 26.900 ;
        RECT 136.040 25.270 139.320 26.900 ;
        RECT -26.420 23.640 -23.130 25.270 ;
        RECT 137.640 23.640 140.930 25.270 ;
        RECT -24.810 22.010 -21.530 23.640 ;
        RECT 136.040 22.010 139.320 23.640 ;
        RECT -26.420 20.380 -23.130 22.010 ;
        RECT 137.640 20.380 140.930 22.010 ;
        RECT -24.810 18.750 -21.530 20.380 ;
        RECT 136.040 18.750 139.320 20.380 ;
        RECT -26.420 17.120 -23.130 18.750 ;
        RECT 137.640 17.120 140.930 18.750 ;
        RECT -24.810 15.490 -21.530 17.120 ;
        RECT 136.040 15.490 139.320 17.120 ;
        RECT -26.420 13.860 -23.130 15.490 ;
        RECT 137.640 13.860 140.930 15.490 ;
        RECT -24.810 12.230 -21.530 13.860 ;
        RECT 136.040 12.230 139.320 13.860 ;
        RECT -26.420 10.600 -23.130 12.230 ;
        RECT 137.640 10.600 140.930 12.230 ;
        RECT -24.810 8.970 -21.530 10.600 ;
        RECT -26.420 7.340 -23.130 8.970 ;
        RECT -24.810 5.710 -21.530 7.340 ;
        RECT 7.320 5.920 11.900 10.290 ;
        RECT -26.420 4.080 -23.130 5.710 ;
        RECT 38.110 5.690 42.680 10.130 ;
        RECT 71.830 5.690 76.400 10.130 ;
        RECT 102.610 5.920 107.190 10.290 ;
        RECT 136.040 8.970 139.320 10.600 ;
        RECT 137.640 7.340 140.930 8.970 ;
        RECT 136.040 5.710 139.320 7.340 ;
        RECT 137.640 4.080 140.930 5.710 ;
        RECT -24.810 2.450 -21.530 4.080 ;
        RECT 136.040 2.450 139.320 4.080 ;
        RECT -26.420 0.820 -23.130 2.450 ;
        RECT 137.640 0.820 140.930 2.450 ;
        RECT -24.810 -0.810 -21.530 0.820 ;
        RECT 136.040 -0.810 139.320 0.820 ;
        RECT -26.420 -2.440 -23.130 -0.810 ;
        RECT 137.640 -2.440 140.930 -0.810 ;
        RECT -24.810 -4.070 -21.530 -2.440 ;
        RECT 136.040 -4.070 139.320 -2.440 ;
        RECT -26.420 -5.700 -23.130 -4.070 ;
        RECT 137.640 -5.700 140.930 -4.070 ;
        RECT -24.810 -7.330 -21.530 -5.700 ;
        RECT 136.040 -7.330 139.320 -5.700 ;
        RECT -26.420 -8.960 -23.130 -7.330 ;
        RECT -24.810 -8.970 -23.130 -8.960 ;
        RECT 137.640 -8.960 140.930 -7.330 ;
        RECT 137.640 -8.970 139.320 -8.960 ;
        RECT -24.810 -10.600 -21.530 -8.970 ;
        RECT 136.040 -10.600 139.320 -8.970 ;
        RECT -26.420 -12.230 -23.130 -10.600 ;
        RECT -24.810 -13.870 -23.130 -12.230 ;
        RECT -26.420 -14.430 -23.130 -13.870 ;
        RECT 6.410 -14.430 8.070 -10.730 ;
        RECT 106.440 -14.430 108.100 -10.730 ;
        RECT 137.640 -12.230 140.930 -10.600 ;
        RECT 137.640 -13.870 139.320 -12.230 ;
        RECT 137.640 -14.430 140.930 -13.870 ;
        RECT -26.420 -15.500 8.410 -14.430 ;
        RECT -24.810 -16.090 8.410 -15.500 ;
        RECT 106.100 -15.500 140.930 -14.430 ;
        RECT 106.100 -16.090 139.320 -15.500 ;
        RECT 5.580 -18.390 7.190 -16.090 ;
        RECT 2.200 -20.000 7.190 -18.390 ;
        RECT 107.320 -18.390 108.930 -16.090 ;
        RECT 107.320 -20.000 112.310 -18.390 ;
    END
  END vssa1
  PIN phi1b
    ANTENNAGATEAREA 1.140000 ;
    PORT
      LAYER li1 ;
        RECT 17.820 -14.030 17.990 -13.040 ;
        RECT 26.520 -14.030 26.690 -13.040 ;
        RECT 87.820 -14.030 87.990 -13.040 ;
        RECT 96.520 -14.030 96.690 -13.040 ;
        RECT 8.870 -14.200 9.200 -14.030 ;
        RECT 17.740 -14.200 18.070 -14.030 ;
        RECT 26.440 -14.200 26.770 -14.030 ;
        RECT 87.740 -14.200 88.070 -14.030 ;
        RECT 96.440 -14.200 96.770 -14.030 ;
        RECT 105.310 -14.200 105.640 -14.030 ;
        RECT 60.920 -50.910 61.090 -50.580 ;
        RECT 65.370 -51.255 65.710 -49.605 ;
        RECT 74.010 -51.255 74.350 -49.605 ;
        RECT 82.650 -51.255 82.990 -49.605 ;
        RECT 91.290 -51.255 91.630 -49.605 ;
      LAYER mcon ;
        RECT 17.820 -13.250 17.990 -13.080 ;
        RECT 26.520 -13.210 26.690 -13.040 ;
        RECT 87.820 -13.210 87.990 -13.040 ;
        RECT 96.520 -13.250 96.690 -13.080 ;
        RECT 8.950 -14.200 9.120 -14.030 ;
        RECT 105.390 -14.200 105.560 -14.030 ;
        RECT 60.920 -50.830 61.090 -50.660 ;
        RECT 65.520 -50.835 65.690 -50.665 ;
        RECT 74.160 -50.835 74.330 -50.665 ;
        RECT 82.800 -50.835 82.970 -50.665 ;
        RECT 91.440 -50.835 91.610 -50.665 ;
      LAYER met1 ;
        RECT 26.460 -13.040 26.740 -13.010 ;
        RECT 57.470 -13.040 57.730 -13.020 ;
        RECT 87.770 -13.040 88.050 -13.010 ;
        RECT 8.950 -13.180 105.560 -13.040 ;
        RECT 8.950 -13.970 9.120 -13.180 ;
        RECT 17.760 -13.300 18.050 -13.180 ;
        RECT 26.460 -13.270 26.740 -13.180 ;
        RECT 57.470 -13.340 57.730 -13.180 ;
        RECT 87.770 -13.270 88.050 -13.180 ;
        RECT 96.460 -13.300 96.750 -13.180 ;
        RECT 105.390 -13.970 105.560 -13.180 ;
        RECT 8.910 -14.260 9.160 -13.970 ;
        RECT 105.350 -14.260 105.600 -13.970 ;
        RECT 60.875 -50.925 61.150 -50.570 ;
        RECT 65.460 -50.925 65.750 -50.575 ;
        RECT 74.050 -50.950 74.455 -50.545 ;
        RECT 82.705 -50.945 83.090 -50.550 ;
        RECT 91.320 -50.955 91.725 -50.560 ;
      LAYER via ;
        RECT 57.470 -13.310 57.730 -13.050 ;
        RECT 60.890 -50.870 61.150 -50.605 ;
        RECT 65.460 -50.895 65.750 -50.605 ;
        RECT 74.125 -50.875 74.385 -50.615 ;
        RECT 82.765 -50.875 83.025 -50.615 ;
        RECT 91.395 -50.880 91.655 -50.615 ;
      LAYER met2 ;
        RECT 57.530 32.520 70.960 32.720 ;
        RECT 57.530 -13.020 57.680 32.520 ;
        RECT 57.470 -13.340 57.730 -13.020 ;
        RECT 57.530 -49.095 57.680 -13.340 ;
        RECT 57.530 -49.245 61.040 -49.095 ;
        RECT 60.875 -50.550 61.040 -49.245 ;
        RECT 60.870 -50.930 61.165 -50.550 ;
        RECT 65.430 -50.970 65.795 -50.530 ;
        RECT 74.050 -50.950 74.455 -50.545 ;
        RECT 82.705 -50.945 83.090 -50.550 ;
        RECT 91.320 -50.955 91.725 -50.560 ;
      LAYER via2 ;
        RECT 60.880 -50.885 61.160 -50.595 ;
        RECT 65.460 -50.925 65.750 -50.575 ;
        RECT 74.095 -50.905 74.410 -50.590 ;
        RECT 82.750 -50.900 83.045 -50.595 ;
        RECT 91.370 -50.910 91.675 -50.610 ;
      LAYER met3 ;
        RECT 60.850 -50.595 61.185 -50.550 ;
        RECT 65.430 -50.585 65.795 -50.530 ;
        RECT 74.050 -50.585 74.455 -50.545 ;
        RECT 82.705 -50.585 83.090 -50.550 ;
        RECT 91.320 -50.585 91.725 -50.560 ;
        RECT 65.215 -50.595 91.725 -50.585 ;
        RECT 60.850 -50.920 91.725 -50.595 ;
        RECT 60.850 -50.930 61.185 -50.920 ;
        RECT 65.430 -50.970 65.795 -50.920 ;
        RECT 74.050 -50.950 74.455 -50.920 ;
        RECT 82.705 -50.945 83.090 -50.920 ;
        RECT 91.320 -50.955 91.725 -50.920 ;
    END
  END phi1b
  PIN phi2b
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 17.060 -14.030 17.230 -12.700 ;
        RECT 25.760 -14.030 25.930 -12.700 ;
        RECT 31.710 -14.030 31.880 -12.700 ;
        RECT 82.630 -14.030 82.800 -12.700 ;
        RECT 88.580 -14.030 88.750 -12.700 ;
        RECT 97.280 -14.030 97.450 -12.700 ;
        RECT 16.980 -14.200 17.310 -14.030 ;
        RECT 25.680 -14.200 26.010 -14.030 ;
        RECT 31.630 -14.200 31.960 -14.030 ;
        RECT 82.550 -14.200 82.880 -14.030 ;
        RECT 88.500 -14.200 88.830 -14.030 ;
        RECT 97.200 -14.200 97.530 -14.030 ;
      LAYER mcon ;
        RECT 17.060 -12.870 17.230 -12.700 ;
        RECT 25.760 -12.870 25.930 -12.700 ;
        RECT 31.710 -12.870 31.880 -12.700 ;
        RECT 82.630 -12.870 82.800 -12.700 ;
        RECT 88.580 -12.870 88.750 -12.700 ;
        RECT 97.280 -12.870 97.450 -12.700 ;
      LAYER met1 ;
        RECT 17.000 -12.730 17.290 -12.640 ;
        RECT 25.700 -12.730 25.990 -12.640 ;
        RECT 31.650 -12.730 31.940 -12.670 ;
        RECT 57.830 -12.730 58.090 -12.560 ;
        RECT 82.570 -12.730 82.860 -12.670 ;
        RECT 88.520 -12.730 88.810 -12.640 ;
        RECT 97.220 -12.730 97.510 -12.640 ;
        RECT 17.000 -12.870 97.510 -12.730 ;
        RECT 17.000 -12.900 17.290 -12.870 ;
        RECT 25.700 -12.900 25.990 -12.870 ;
        RECT 31.650 -12.900 31.940 -12.870 ;
        RECT 57.830 -12.880 58.090 -12.870 ;
        RECT 82.570 -12.900 82.860 -12.870 ;
        RECT 88.520 -12.900 88.810 -12.870 ;
        RECT 97.220 -12.900 97.510 -12.870 ;
      LAYER via ;
        RECT 57.830 -12.850 58.090 -12.590 ;
      LAYER met2 ;
        RECT 57.880 31.380 78.840 31.580 ;
        RECT 57.880 -12.560 58.030 31.380 ;
        RECT 57.830 -12.880 58.090 -12.560 ;
    END
  END phi2b
  PIN vbotm
    PORT
      LAYER met1 ;
        RECT 58.170 -15.850 58.430 -15.780 ;
        RECT 59.260 -15.850 59.530 -15.760 ;
        RECT 58.170 -15.990 59.530 -15.850 ;
        RECT 58.170 -16.100 58.430 -15.990 ;
        RECT 59.260 -16.080 59.530 -15.990 ;
      LAYER via ;
        RECT 58.170 -16.070 58.430 -15.810 ;
        RECT 59.260 -16.050 59.530 -15.790 ;
      LAYER met2 ;
        RECT 58.230 30.440 85.010 30.640 ;
        RECT 58.230 -15.780 58.380 30.440 ;
        RECT 58.170 -16.100 58.430 -15.780 ;
        RECT 59.230 -16.140 59.570 -15.700 ;
      LAYER via2 ;
        RECT 59.230 -16.090 59.570 -15.750 ;
      LAYER met3 ;
        RECT 58.570 -17.970 60.210 -15.020 ;
        RECT 58.450 -48.250 83.740 -17.970 ;
      LAYER via3 ;
        RECT 59.230 -16.090 59.570 -15.750 ;
      LAYER met4 ;
        RECT 58.770 -16.460 59.950 -15.280 ;
      LAYER met5 ;
        RECT 58.570 -18.050 60.210 -15.020 ;
        RECT 58.580 -19.780 60.210 -18.050 ;
    END
  END vbotm
  PIN vbotp
    PORT
      LAYER met1 ;
        RECT 54.980 -15.850 55.250 -15.760 ;
        RECT 57.130 -15.850 57.390 -15.780 ;
        RECT 54.980 -15.990 57.390 -15.850 ;
        RECT 54.980 -16.080 55.250 -15.990 ;
        RECT 57.130 -16.100 57.390 -15.990 ;
      LAYER via ;
        RECT 54.980 -16.050 55.250 -15.790 ;
        RECT 57.130 -16.070 57.390 -15.810 ;
      LAYER met2 ;
        RECT 54.940 -16.140 55.280 -15.700 ;
        RECT 57.180 -15.780 57.330 37.200 ;
        RECT 57.130 -16.100 57.390 -15.780 ;
      LAYER via2 ;
        RECT 54.940 -16.090 55.280 -15.750 ;
      LAYER met3 ;
        RECT 54.300 -17.970 55.940 -15.020 ;
        RECT 30.770 -48.250 56.060 -17.970 ;
      LAYER via3 ;
        RECT 54.940 -16.090 55.280 -15.750 ;
      LAYER met4 ;
        RECT 54.560 -16.460 55.740 -15.280 ;
      LAYER met5 ;
        RECT 54.300 -18.050 55.940 -15.020 ;
        RECT 54.300 -19.780 55.930 -18.050 ;
    END
  END vbotp
  PIN vdda1
    ANTENNADIFFAREA 11.214825 ;
    PORT
      LAYER nwell ;
        RECT 8.430 -15.050 32.650 -14.210 ;
        RECT 81.860 -15.050 106.080 -14.210 ;
        RECT 65.095 -49.370 107.235 -48.575 ;
        RECT 56.790 -50.220 107.235 -49.370 ;
        RECT 65.095 -50.440 107.235 -50.220 ;
      LAYER li1 ;
        RECT 18.390 -13.500 18.560 -13.470 ;
        RECT 27.090 -13.500 27.260 -13.470 ;
        RECT 32.280 -13.500 32.450 -13.470 ;
        RECT 82.060 -13.500 82.230 -13.470 ;
        RECT 87.250 -13.500 87.420 -13.470 ;
        RECT 95.950 -13.500 96.120 -13.470 ;
        RECT 9.460 -13.670 9.740 -13.500 ;
        RECT 18.360 -13.670 18.590 -13.500 ;
        RECT 27.060 -13.670 27.290 -13.500 ;
        RECT 32.250 -13.670 32.480 -13.500 ;
        RECT 82.030 -13.670 82.260 -13.500 ;
        RECT 87.220 -13.670 87.450 -13.500 ;
        RECT 95.920 -13.670 96.150 -13.500 ;
        RECT 104.770 -13.670 105.050 -13.500 ;
        RECT 9.520 -14.810 9.690 -13.670 ;
        RECT 18.390 -14.810 18.560 -13.670 ;
        RECT 27.090 -14.810 27.260 -13.670 ;
        RECT 32.280 -14.810 32.450 -13.670 ;
        RECT 82.060 -14.810 82.230 -13.670 ;
        RECT 87.250 -14.810 87.420 -13.670 ;
        RECT 95.950 -14.810 96.120 -13.670 ;
        RECT 104.820 -14.810 104.990 -13.670 ;
        RECT 56.490 -48.850 107.045 -48.680 ;
        RECT 57.470 -49.630 57.640 -48.850 ;
        RECT 57.430 -49.960 57.680 -49.630 ;
        RECT 59.960 -49.960 60.230 -49.630 ;
        RECT 61.260 -49.980 61.430 -48.850 ;
        RECT 62.200 -49.680 62.370 -48.850 ;
        RECT 62.170 -50.010 62.420 -49.680 ;
        RECT 63.260 -49.890 63.430 -48.850 ;
        RECT 64.070 -49.680 64.240 -48.850 ;
        RECT 65.380 -49.435 65.710 -48.850 ;
        RECT 64.040 -50.010 64.290 -49.680 ;
        RECT 66.875 -49.810 67.205 -48.850 ;
        RECT 69.260 -49.470 69.590 -48.850 ;
        RECT 71.435 -50.120 71.815 -48.850 ;
        RECT 72.620 -50.280 72.900 -48.850 ;
        RECT 73.505 -50.280 73.740 -48.850 ;
        RECT 74.020 -49.435 74.350 -48.850 ;
        RECT 75.515 -49.810 75.845 -48.850 ;
        RECT 77.900 -49.470 78.230 -48.850 ;
        RECT 80.075 -50.120 80.455 -48.850 ;
        RECT 81.260 -50.280 81.540 -48.850 ;
        RECT 82.145 -50.280 82.380 -48.850 ;
        RECT 82.660 -49.435 82.990 -48.850 ;
        RECT 84.155 -49.810 84.485 -48.850 ;
        RECT 86.540 -49.470 86.870 -48.850 ;
        RECT 88.715 -50.120 89.095 -48.850 ;
        RECT 89.900 -50.280 90.180 -48.850 ;
        RECT 90.785 -50.280 91.020 -48.850 ;
        RECT 91.300 -49.435 91.630 -48.850 ;
        RECT 92.795 -49.810 93.125 -48.850 ;
        RECT 95.180 -49.470 95.510 -48.850 ;
        RECT 97.355 -50.120 97.735 -48.850 ;
        RECT 98.540 -50.280 98.820 -48.850 ;
        RECT 99.425 -50.280 99.660 -48.850 ;
        RECT 100.835 -49.690 101.115 -48.850 ;
        RECT 101.810 -49.180 102.140 -48.850 ;
        RECT 103.625 -50.140 103.955 -48.850 ;
        RECT 104.750 -49.835 105.080 -48.850 ;
        RECT 106.190 -50.150 106.520 -48.850 ;
      LAYER mcon ;
        RECT 9.520 -13.670 9.690 -13.500 ;
        RECT 18.390 -13.670 18.560 -13.500 ;
        RECT 27.090 -13.670 27.260 -13.500 ;
        RECT 32.280 -13.670 32.450 -13.500 ;
        RECT 82.060 -13.670 82.230 -13.500 ;
        RECT 87.250 -13.670 87.420 -13.500 ;
        RECT 95.950 -13.670 96.120 -13.500 ;
        RECT 104.820 -13.670 104.990 -13.500 ;
        RECT 56.800 -48.850 56.970 -48.680 ;
        RECT 57.280 -48.850 57.450 -48.680 ;
        RECT 57.760 -48.850 57.930 -48.680 ;
        RECT 58.240 -48.850 58.410 -48.680 ;
        RECT 58.720 -48.850 58.890 -48.680 ;
        RECT 59.200 -48.850 59.370 -48.680 ;
        RECT 59.680 -48.850 59.850 -48.680 ;
        RECT 60.160 -48.850 60.330 -48.680 ;
        RECT 60.640 -48.850 60.810 -48.680 ;
        RECT 61.120 -48.850 61.290 -48.680 ;
        RECT 61.600 -48.850 61.770 -48.680 ;
        RECT 62.080 -48.850 62.250 -48.680 ;
        RECT 62.560 -48.850 62.730 -48.680 ;
        RECT 63.040 -48.850 63.210 -48.680 ;
        RECT 63.520 -48.850 63.690 -48.680 ;
        RECT 64.000 -48.850 64.170 -48.680 ;
        RECT 64.480 -48.850 64.650 -48.680 ;
        RECT 64.960 -48.850 65.130 -48.680 ;
        RECT 65.440 -48.850 65.610 -48.680 ;
        RECT 65.920 -48.850 66.090 -48.680 ;
        RECT 66.400 -48.850 66.570 -48.680 ;
        RECT 66.880 -48.850 67.050 -48.680 ;
        RECT 67.360 -48.850 67.530 -48.680 ;
        RECT 67.840 -48.850 68.010 -48.680 ;
        RECT 68.320 -48.850 68.490 -48.680 ;
        RECT 68.800 -48.850 68.970 -48.680 ;
        RECT 69.280 -48.850 69.450 -48.680 ;
        RECT 69.760 -48.850 69.930 -48.680 ;
        RECT 70.240 -48.850 70.410 -48.680 ;
        RECT 70.720 -48.850 70.890 -48.680 ;
        RECT 71.200 -48.850 71.370 -48.680 ;
        RECT 71.680 -48.850 71.850 -48.680 ;
        RECT 72.160 -48.850 72.330 -48.680 ;
        RECT 72.640 -48.850 72.810 -48.680 ;
        RECT 73.120 -48.850 73.290 -48.680 ;
        RECT 73.600 -48.850 73.770 -48.680 ;
        RECT 74.080 -48.850 74.250 -48.680 ;
        RECT 74.560 -48.850 74.730 -48.680 ;
        RECT 75.040 -48.850 75.210 -48.680 ;
        RECT 75.520 -48.850 75.690 -48.680 ;
        RECT 76.000 -48.850 76.170 -48.680 ;
        RECT 76.480 -48.850 76.650 -48.680 ;
        RECT 76.960 -48.850 77.130 -48.680 ;
        RECT 77.440 -48.850 77.610 -48.680 ;
        RECT 77.920 -48.850 78.090 -48.680 ;
        RECT 78.400 -48.850 78.570 -48.680 ;
        RECT 78.880 -48.850 79.050 -48.680 ;
        RECT 79.360 -48.850 79.530 -48.680 ;
        RECT 79.840 -48.850 80.010 -48.680 ;
        RECT 80.320 -48.850 80.490 -48.680 ;
        RECT 80.800 -48.850 80.970 -48.680 ;
        RECT 81.280 -48.850 81.450 -48.680 ;
        RECT 81.760 -48.850 81.930 -48.680 ;
        RECT 82.240 -48.850 82.410 -48.680 ;
        RECT 82.720 -48.850 82.890 -48.680 ;
        RECT 83.200 -48.850 83.370 -48.680 ;
        RECT 83.680 -48.850 83.850 -48.680 ;
        RECT 84.160 -48.850 84.330 -48.680 ;
        RECT 84.640 -48.850 84.810 -48.680 ;
        RECT 85.120 -48.850 85.290 -48.680 ;
        RECT 85.600 -48.850 85.770 -48.680 ;
        RECT 86.080 -48.850 86.250 -48.680 ;
        RECT 86.560 -48.850 86.730 -48.680 ;
        RECT 87.040 -48.850 87.210 -48.680 ;
        RECT 87.520 -48.850 87.690 -48.680 ;
        RECT 88.000 -48.850 88.170 -48.680 ;
        RECT 88.480 -48.850 88.650 -48.680 ;
        RECT 88.960 -48.850 89.130 -48.680 ;
        RECT 89.440 -48.850 89.610 -48.680 ;
        RECT 89.920 -48.850 90.090 -48.680 ;
        RECT 90.400 -48.850 90.570 -48.680 ;
        RECT 90.880 -48.850 91.050 -48.680 ;
        RECT 91.360 -48.850 91.530 -48.680 ;
        RECT 91.840 -48.850 92.010 -48.680 ;
        RECT 92.320 -48.850 92.490 -48.680 ;
        RECT 92.800 -48.850 92.970 -48.680 ;
        RECT 93.280 -48.850 93.450 -48.680 ;
        RECT 93.760 -48.850 93.930 -48.680 ;
        RECT 94.240 -48.850 94.410 -48.680 ;
        RECT 94.720 -48.850 94.890 -48.680 ;
        RECT 95.200 -48.850 95.370 -48.680 ;
        RECT 95.680 -48.850 95.850 -48.680 ;
        RECT 96.160 -48.850 96.330 -48.680 ;
        RECT 96.640 -48.850 96.810 -48.680 ;
        RECT 97.120 -48.850 97.290 -48.680 ;
        RECT 97.600 -48.850 97.770 -48.680 ;
        RECT 98.080 -48.850 98.250 -48.680 ;
        RECT 98.560 -48.850 98.730 -48.680 ;
        RECT 99.040 -48.850 99.210 -48.680 ;
        RECT 99.520 -48.850 99.690 -48.680 ;
        RECT 100.000 -48.850 100.170 -48.680 ;
        RECT 100.480 -48.850 100.650 -48.680 ;
        RECT 100.960 -48.850 101.130 -48.680 ;
        RECT 101.440 -48.850 101.610 -48.680 ;
        RECT 101.920 -48.850 102.090 -48.680 ;
        RECT 102.400 -48.850 102.570 -48.680 ;
        RECT 102.880 -48.850 103.050 -48.680 ;
        RECT 103.360 -48.850 103.530 -48.680 ;
        RECT 103.840 -48.850 104.010 -48.680 ;
        RECT 104.320 -48.850 104.490 -48.680 ;
        RECT 104.800 -48.850 104.970 -48.680 ;
        RECT 105.280 -48.850 105.450 -48.680 ;
        RECT 105.760 -48.850 105.930 -48.680 ;
        RECT 106.240 -48.850 106.410 -48.680 ;
        RECT 106.720 -48.850 106.890 -48.680 ;
        RECT 60.000 -49.880 60.170 -49.710 ;
      LAYER met1 ;
        RECT 9.490 -13.500 9.720 -13.470 ;
        RECT 18.360 -13.500 18.590 -13.470 ;
        RECT 27.060 -13.500 27.290 -13.470 ;
        RECT 32.250 -13.500 32.480 -13.470 ;
        RECT 56.000 -13.500 56.260 -13.440 ;
        RECT 82.030 -13.500 82.260 -13.470 ;
        RECT 87.220 -13.500 87.450 -13.470 ;
        RECT 95.920 -13.500 96.150 -13.470 ;
        RECT 104.790 -13.500 105.020 -13.470 ;
        RECT 9.460 -13.670 105.050 -13.500 ;
        RECT 9.490 -13.700 9.720 -13.670 ;
        RECT 18.360 -13.700 18.590 -13.670 ;
        RECT 27.060 -13.700 27.290 -13.670 ;
        RECT 32.250 -13.700 32.480 -13.670 ;
        RECT 56.000 -13.760 56.260 -13.670 ;
        RECT 82.030 -13.700 82.260 -13.670 ;
        RECT 87.220 -13.700 87.450 -13.670 ;
        RECT 95.920 -13.700 96.150 -13.670 ;
        RECT 104.790 -13.700 105.020 -13.670 ;
        RECT 56.040 -49.010 107.045 -48.520 ;
        RECT 60.000 -49.680 60.170 -49.010 ;
        RECT 59.970 -49.940 60.200 -49.680 ;
      LAYER via ;
        RECT 56.000 -13.730 56.260 -13.470 ;
        RECT 56.075 -48.860 56.335 -48.600 ;
      LAYER met2 ;
        RECT 28.130 30.440 56.280 30.640 ;
        RECT 56.130 -13.440 56.280 30.440 ;
        RECT 56.000 -13.760 56.280 -13.440 ;
        RECT 56.130 -48.520 56.280 -13.760 ;
        RECT 56.040 -49.010 56.340 -48.520 ;
    END
  END vdda1
  PIN phi1
    ANTENNAGATEAREA 0.567000 ;
    PORT
      LAYER li1 ;
        RECT 8.950 -16.240 9.120 -16.210 ;
        RECT 105.390 -16.240 105.560 -16.210 ;
        RECT 8.870 -16.410 9.200 -16.240 ;
        RECT 17.740 -16.410 18.070 -16.240 ;
        RECT 26.440 -16.410 26.770 -16.240 ;
        RECT 87.740 -16.410 88.070 -16.240 ;
        RECT 96.440 -16.410 96.770 -16.240 ;
        RECT 105.310 -16.410 105.640 -16.240 ;
        RECT 8.950 -16.440 9.120 -16.410 ;
        RECT 17.820 -17.480 17.990 -16.410 ;
        RECT 26.520 -17.480 26.690 -16.410 ;
        RECT 87.820 -17.480 87.990 -16.410 ;
        RECT 96.520 -17.480 96.690 -16.410 ;
        RECT 105.390 -16.440 105.560 -16.410 ;
        RECT 58.510 -50.710 58.840 -50.540 ;
      LAYER mcon ;
        RECT 8.950 -16.410 9.120 -16.240 ;
        RECT 105.390 -16.410 105.560 -16.240 ;
        RECT 17.820 -17.390 17.990 -17.220 ;
        RECT 96.520 -17.390 96.690 -17.220 ;
        RECT 58.590 -50.710 58.760 -50.540 ;
      LAYER met1 ;
        RECT 8.920 -16.440 9.150 -16.180 ;
        RECT 105.360 -16.440 105.590 -16.180 ;
        RECT 8.950 -17.340 9.120 -16.440 ;
        RECT 17.730 -17.340 18.050 -17.140 ;
        RECT 26.460 -17.340 26.750 -17.240 ;
        RECT 56.425 -17.340 56.685 -17.150 ;
        RECT 87.760 -17.340 88.050 -17.240 ;
        RECT 96.460 -17.340 96.780 -17.140 ;
        RECT 105.390 -17.340 105.560 -16.440 ;
        RECT 8.950 -17.480 105.560 -17.340 ;
        RECT 26.460 -17.520 26.750 -17.480 ;
        RECT 87.760 -17.520 88.050 -17.480 ;
        RECT 58.475 -50.765 58.870 -50.480 ;
      LAYER via ;
        RECT 56.425 -17.440 56.685 -17.180 ;
        RECT 58.510 -50.765 58.815 -50.480 ;
      LAYER met2 ;
        RECT 36.680 31.390 56.630 31.590 ;
        RECT 56.480 -17.150 56.630 31.390 ;
        RECT 56.425 -17.470 56.685 -17.150 ;
        RECT 56.475 -17.480 56.685 -17.470 ;
        RECT 56.480 -17.485 56.685 -17.480 ;
        RECT 56.480 -50.040 56.630 -17.485 ;
        RECT 56.480 -50.185 58.855 -50.040 ;
        RECT 58.620 -50.480 58.855 -50.185 ;
        RECT 58.475 -50.765 58.870 -50.480 ;
    END
  END phi1
  PIN phi2
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 16.980 -16.410 17.310 -16.240 ;
        RECT 25.680 -16.410 26.010 -16.240 ;
        RECT 31.630 -16.410 31.960 -16.240 ;
        RECT 82.550 -16.410 82.880 -16.240 ;
        RECT 88.500 -16.410 88.830 -16.240 ;
        RECT 97.200 -16.410 97.530 -16.240 ;
        RECT 17.060 -17.820 17.230 -16.410 ;
        RECT 25.760 -17.820 25.930 -16.410 ;
        RECT 31.710 -17.820 31.880 -16.410 ;
        RECT 82.630 -17.820 82.800 -16.410 ;
        RECT 88.580 -17.820 88.750 -16.410 ;
        RECT 97.280 -17.820 97.450 -16.410 ;
      LAYER met1 ;
        RECT 17.000 -17.660 17.290 -17.620 ;
        RECT 25.700 -17.660 26.000 -17.620 ;
        RECT 31.650 -17.660 31.940 -17.620 ;
        RECT 56.830 -17.660 57.090 -17.620 ;
        RECT 82.570 -17.660 82.860 -17.620 ;
        RECT 88.510 -17.660 88.810 -17.620 ;
        RECT 97.220 -17.660 97.510 -17.620 ;
        RECT 17.000 -17.800 97.510 -17.660 ;
        RECT 17.000 -17.880 17.290 -17.800 ;
        RECT 25.700 -17.910 26.000 -17.800 ;
        RECT 31.650 -17.880 31.940 -17.800 ;
        RECT 56.830 -17.940 57.090 -17.800 ;
        RECT 82.570 -17.880 82.860 -17.800 ;
        RECT 88.510 -17.910 88.810 -17.800 ;
        RECT 97.220 -17.880 97.510 -17.800 ;
      LAYER via ;
        RECT 56.830 -17.910 57.090 -17.650 ;
      LAYER met2 ;
        RECT 44.650 32.510 56.980 32.710 ;
        RECT 56.830 -17.620 56.980 32.510 ;
        RECT 56.830 -17.940 57.090 -17.620 ;
    END
  END phi2
  PIN events
    ANTENNADIFFAREA 0.556500 ;
    PORT
      LAYER li1 ;
        RECT 106.690 -50.230 106.960 -49.020 ;
        RECT 106.785 -51.065 106.960 -50.230 ;
        RECT 106.690 -51.840 106.960 -51.065 ;
      LAYER mcon ;
        RECT 106.700 -51.320 106.880 -51.130 ;
      LAYER met1 ;
        RECT 106.640 -51.140 106.940 -51.070 ;
        RECT 107.470 -51.140 135.830 -51.110 ;
        RECT 106.640 -51.310 135.830 -51.140 ;
        RECT 106.640 -51.385 106.940 -51.310 ;
    END
  END events
  PIN polxevent
    ANTENNADIFFAREA 0.581700 ;
    PORT
      LAYER li1 ;
        RECT 105.250 -51.115 105.520 -49.020 ;
        RECT 104.955 -51.840 105.520 -51.115 ;
      LAYER mcon ;
        RECT 105.260 -49.735 105.430 -49.565 ;
      LAYER met1 ;
        RECT 105.195 -49.565 105.510 -49.505 ;
        RECT 107.435 -49.565 135.820 -49.535 ;
        RECT 105.195 -49.735 135.820 -49.565 ;
        RECT 105.195 -49.795 105.510 -49.735 ;
    END
  END polxevent
  OBS
      LAYER li1 ;
        RECT 8.710 -15.990 8.880 -14.480 ;
        RECT 9.180 -15.200 9.350 -14.480 ;
        RECT 9.180 -15.370 9.430 -15.200 ;
        RECT 9.180 -15.990 9.350 -15.370 ;
        RECT 16.820 -15.990 16.990 -14.480 ;
        RECT 17.290 -15.990 17.750 -14.480 ;
        RECT 18.050 -15.200 18.220 -14.480 ;
        RECT 18.050 -15.370 18.300 -15.200 ;
        RECT 18.050 -15.990 18.220 -15.370 ;
        RECT 25.520 -15.990 25.690 -14.480 ;
        RECT 25.990 -15.990 26.450 -14.480 ;
        RECT 26.750 -15.200 26.920 -14.480 ;
        RECT 31.470 -15.190 31.640 -14.480 ;
        RECT 26.750 -15.370 27.000 -15.200 ;
        RECT 31.380 -15.360 31.640 -15.190 ;
        RECT 26.750 -15.990 26.920 -15.370 ;
        RECT 31.470 -15.990 31.640 -15.360 ;
        RECT 31.940 -15.200 32.110 -14.480 ;
        RECT 82.400 -15.200 82.570 -14.480 ;
        RECT 31.940 -15.370 32.190 -15.200 ;
        RECT 82.320 -15.370 82.570 -15.200 ;
        RECT 31.940 -15.990 32.110 -15.370 ;
        RECT 82.400 -15.990 82.570 -15.370 ;
        RECT 82.870 -15.190 83.040 -14.480 ;
        RECT 82.870 -15.360 83.130 -15.190 ;
        RECT 87.590 -15.200 87.760 -14.480 ;
        RECT 82.870 -15.990 83.040 -15.360 ;
        RECT 87.510 -15.370 87.760 -15.200 ;
        RECT 87.590 -15.990 87.760 -15.370 ;
        RECT 88.060 -15.990 88.520 -14.480 ;
        RECT 88.820 -15.990 88.990 -14.480 ;
        RECT 96.290 -15.200 96.460 -14.480 ;
        RECT 96.210 -15.370 96.460 -15.200 ;
        RECT 96.290 -15.990 96.460 -15.370 ;
        RECT 96.760 -15.990 97.220 -14.480 ;
        RECT 97.520 -15.990 97.690 -14.480 ;
        RECT 105.160 -15.200 105.330 -14.480 ;
        RECT 105.080 -15.370 105.330 -15.200 ;
        RECT 105.160 -15.990 105.330 -15.370 ;
        RECT 105.630 -15.990 105.800 -14.480 ;
        RECT 57.950 -49.190 60.430 -49.020 ;
        RECT 57.950 -49.630 58.120 -49.190 ;
        RECT 60.100 -49.290 60.430 -49.190 ;
        RECT 56.830 -49.960 57.240 -49.630 ;
        RECT 57.870 -49.640 58.120 -49.630 ;
        RECT 57.870 -49.960 58.260 -49.640 ;
        RECT 56.830 -51.130 57.000 -49.960 ;
        RECT 57.190 -50.890 57.360 -50.550 ;
        RECT 57.720 -50.890 57.890 -50.550 ;
        RECT 58.090 -51.130 58.260 -49.960 ;
        RECT 58.600 -50.020 58.830 -49.690 ;
        RECT 59.080 -49.960 59.330 -49.630 ;
        RECT 59.520 -49.960 59.770 -49.630 ;
        RECT 60.400 -49.960 60.650 -49.630 ;
        RECT 60.840 -49.960 61.090 -49.630 ;
        RECT 59.080 -50.260 59.250 -49.960 ;
        RECT 60.240 -50.260 60.410 -50.180 ;
        RECT 60.880 -50.210 61.050 -49.960 ;
        RECT 61.760 -50.010 61.970 -49.680 ;
        RECT 63.630 -50.010 63.840 -49.680 ;
        RECT 64.480 -50.010 64.900 -49.680 ;
        RECT 59.080 -50.430 60.410 -50.260 ;
        RECT 59.420 -51.130 59.590 -50.430 ;
        RECT 60.240 -50.510 60.410 -50.430 ;
        RECT 60.580 -50.380 61.050 -50.210 ;
        RECT 59.760 -50.690 59.930 -50.610 ;
        RECT 60.580 -50.690 60.750 -50.380 ;
        RECT 61.460 -50.620 61.630 -50.290 ;
        RECT 61.800 -50.560 61.970 -50.010 ;
        RECT 62.430 -50.560 62.600 -50.480 ;
        RECT 59.760 -50.860 60.750 -50.690 ;
        RECT 59.760 -50.940 59.930 -50.860 ;
        RECT 60.450 -50.930 60.750 -50.860 ;
        RECT 61.800 -50.730 62.600 -50.560 ;
        RECT 63.330 -50.620 63.500 -50.290 ;
        RECT 63.670 -50.560 63.840 -50.010 ;
        RECT 64.300 -50.560 64.470 -50.480 ;
        RECT 60.450 -51.130 60.620 -50.930 ;
        RECT 61.800 -51.130 61.970 -50.730 ;
        RECT 62.430 -50.810 62.600 -50.730 ;
        RECT 63.670 -50.730 64.470 -50.560 ;
        RECT 63.670 -51.130 63.840 -50.730 ;
        RECT 64.300 -50.810 64.470 -50.730 ;
        RECT 64.730 -51.130 64.900 -50.010 ;
        RECT 56.830 -51.460 57.080 -51.130 ;
        RECT 57.420 -51.460 57.670 -51.130 ;
        RECT 58.000 -51.300 58.260 -51.130 ;
        RECT 58.000 -51.460 58.250 -51.300 ;
        RECT 58.570 -51.460 58.810 -51.130 ;
        RECT 59.420 -51.300 59.770 -51.130 ;
        RECT 59.520 -51.460 59.770 -51.300 ;
        RECT 60.400 -51.460 60.650 -51.130 ;
        RECT 61.760 -51.460 61.970 -51.130 ;
        RECT 63.630 -51.460 63.840 -51.130 ;
        RECT 64.480 -51.460 64.900 -51.130 ;
        RECT 57.450 -51.640 57.620 -51.460 ;
        RECT 58.570 -51.640 58.740 -51.460 ;
        RECT 57.450 -51.810 58.740 -51.640 ;
        RECT 65.880 -51.765 66.325 -49.045 ;
        RECT 66.495 -49.990 66.705 -49.230 ;
        RECT 67.375 -49.335 68.975 -49.155 ;
        RECT 67.375 -49.990 67.555 -49.335 ;
        RECT 66.495 -50.160 67.555 -49.990 ;
        RECT 66.495 -51.455 66.870 -50.160 ;
        RECT 67.725 -50.875 67.915 -49.505 ;
        RECT 68.085 -50.710 68.255 -49.335 ;
        RECT 68.425 -50.870 68.635 -49.505 ;
        RECT 68.805 -49.640 68.975 -49.335 ;
        RECT 68.805 -49.810 70.450 -49.640 ;
        RECT 68.890 -50.180 70.100 -49.980 ;
        RECT 68.890 -50.690 69.220 -50.180 ;
        RECT 69.460 -50.870 69.710 -50.420 ;
        RECT 67.725 -51.125 67.905 -50.875 ;
        RECT 68.425 -51.040 69.710 -50.870 ;
        RECT 68.425 -51.060 68.625 -51.040 ;
        RECT 67.510 -51.455 67.905 -51.125 ;
        RECT 68.075 -51.230 68.625 -51.060 ;
        RECT 68.075 -51.455 68.345 -51.230 ;
        RECT 69.880 -51.510 70.090 -50.180 ;
        RECT 70.270 -50.540 70.450 -49.810 ;
        RECT 70.620 -50.220 70.940 -49.340 ;
        RECT 70.270 -50.620 70.590 -50.540 ;
        RECT 70.260 -50.800 70.590 -50.620 ;
        RECT 70.770 -50.800 70.940 -50.220 ;
        RECT 72.035 -50.290 72.450 -49.340 ;
        RECT 71.310 -50.450 72.450 -50.290 ;
        RECT 71.310 -50.460 72.720 -50.450 ;
        RECT 71.310 -50.630 71.640 -50.460 ;
        RECT 71.850 -50.800 72.110 -50.640 ;
        RECT 70.770 -50.970 72.110 -50.800 ;
        RECT 72.280 -50.670 72.720 -50.460 ;
        RECT 70.430 -51.450 70.940 -50.970 ;
        RECT 72.280 -51.150 72.450 -50.670 ;
        RECT 71.975 -51.680 72.450 -51.150 ;
        RECT 73.070 -51.720 73.335 -49.020 ;
        RECT 74.520 -51.765 74.965 -49.045 ;
        RECT 75.135 -49.990 75.345 -49.230 ;
        RECT 76.015 -49.335 77.615 -49.155 ;
        RECT 76.015 -49.990 76.195 -49.335 ;
        RECT 75.135 -50.160 76.195 -49.990 ;
        RECT 75.135 -51.455 75.510 -50.160 ;
        RECT 75.865 -50.955 76.195 -50.330 ;
        RECT 76.365 -50.875 76.555 -49.505 ;
        RECT 76.725 -50.710 76.895 -49.335 ;
        RECT 77.065 -50.870 77.275 -49.505 ;
        RECT 77.445 -49.640 77.615 -49.335 ;
        RECT 77.445 -49.810 79.090 -49.640 ;
        RECT 77.530 -50.180 78.740 -49.980 ;
        RECT 77.530 -50.690 77.860 -50.180 ;
        RECT 78.100 -50.870 78.350 -50.420 ;
        RECT 76.365 -51.125 76.545 -50.875 ;
        RECT 77.065 -51.040 78.350 -50.870 ;
        RECT 77.065 -51.060 77.265 -51.040 ;
        RECT 76.150 -51.455 76.545 -51.125 ;
        RECT 76.715 -51.230 77.265 -51.060 ;
        RECT 76.715 -51.455 76.985 -51.230 ;
        RECT 78.520 -51.510 78.730 -50.180 ;
        RECT 78.910 -50.540 79.090 -49.810 ;
        RECT 79.260 -50.220 79.580 -49.340 ;
        RECT 78.910 -50.620 79.230 -50.540 ;
        RECT 78.900 -50.800 79.230 -50.620 ;
        RECT 79.410 -50.800 79.580 -50.220 ;
        RECT 80.675 -50.290 81.090 -49.340 ;
        RECT 79.950 -50.450 81.090 -50.290 ;
        RECT 79.950 -50.460 81.360 -50.450 ;
        RECT 79.950 -50.630 80.280 -50.460 ;
        RECT 80.490 -50.800 80.750 -50.640 ;
        RECT 79.410 -50.970 80.750 -50.800 ;
        RECT 80.920 -50.670 81.360 -50.460 ;
        RECT 79.070 -51.450 79.580 -50.970 ;
        RECT 80.920 -51.150 81.090 -50.670 ;
        RECT 80.615 -51.680 81.090 -51.150 ;
        RECT 81.710 -51.720 81.975 -49.020 ;
        RECT 83.160 -51.765 83.605 -49.045 ;
        RECT 83.775 -49.990 83.985 -49.230 ;
        RECT 84.655 -49.335 86.255 -49.155 ;
        RECT 84.655 -49.990 84.835 -49.335 ;
        RECT 83.775 -50.160 84.835 -49.990 ;
        RECT 83.775 -51.455 84.150 -50.160 ;
        RECT 84.505 -50.955 84.835 -50.330 ;
        RECT 85.005 -50.875 85.195 -49.505 ;
        RECT 85.365 -50.710 85.535 -49.335 ;
        RECT 85.705 -50.870 85.915 -49.505 ;
        RECT 86.085 -49.640 86.255 -49.335 ;
        RECT 86.085 -49.810 87.730 -49.640 ;
        RECT 86.170 -50.180 87.380 -49.980 ;
        RECT 86.170 -50.690 86.500 -50.180 ;
        RECT 86.740 -50.870 86.990 -50.420 ;
        RECT 85.005 -51.125 85.185 -50.875 ;
        RECT 85.705 -51.040 86.990 -50.870 ;
        RECT 85.705 -51.060 85.905 -51.040 ;
        RECT 84.790 -51.455 85.185 -51.125 ;
        RECT 85.355 -51.230 85.905 -51.060 ;
        RECT 85.355 -51.455 85.625 -51.230 ;
        RECT 87.160 -51.510 87.370 -50.180 ;
        RECT 87.550 -50.540 87.730 -49.810 ;
        RECT 87.900 -50.220 88.220 -49.340 ;
        RECT 87.550 -50.620 87.870 -50.540 ;
        RECT 87.540 -50.800 87.870 -50.620 ;
        RECT 88.050 -50.800 88.220 -50.220 ;
        RECT 89.315 -50.290 89.730 -49.340 ;
        RECT 88.590 -50.450 89.730 -50.290 ;
        RECT 88.590 -50.460 90.000 -50.450 ;
        RECT 88.590 -50.630 88.920 -50.460 ;
        RECT 89.130 -50.800 89.390 -50.640 ;
        RECT 88.050 -50.970 89.390 -50.800 ;
        RECT 89.560 -50.670 90.000 -50.460 ;
        RECT 87.710 -51.450 88.220 -50.970 ;
        RECT 89.560 -51.150 89.730 -50.670 ;
        RECT 89.255 -51.680 89.730 -51.150 ;
        RECT 90.350 -51.720 90.615 -49.020 ;
        RECT 91.800 -51.765 92.245 -49.045 ;
        RECT 92.415 -49.990 92.625 -49.230 ;
        RECT 93.295 -49.335 94.895 -49.155 ;
        RECT 93.295 -49.990 93.475 -49.335 ;
        RECT 92.415 -50.160 93.475 -49.990 ;
        RECT 92.415 -51.455 92.790 -50.160 ;
        RECT 93.145 -50.955 93.475 -50.330 ;
        RECT 93.645 -50.875 93.835 -49.505 ;
        RECT 94.005 -50.710 94.175 -49.335 ;
        RECT 94.345 -50.870 94.555 -49.505 ;
        RECT 94.725 -49.640 94.895 -49.335 ;
        RECT 94.725 -49.810 96.370 -49.640 ;
        RECT 94.810 -50.180 96.020 -49.980 ;
        RECT 94.810 -50.690 95.140 -50.180 ;
        RECT 95.380 -50.870 95.630 -50.420 ;
        RECT 93.645 -51.125 93.825 -50.875 ;
        RECT 94.345 -51.040 95.630 -50.870 ;
        RECT 94.345 -51.060 94.545 -51.040 ;
        RECT 93.430 -51.455 93.825 -51.125 ;
        RECT 93.995 -51.230 94.545 -51.060 ;
        RECT 93.995 -51.455 94.265 -51.230 ;
        RECT 95.800 -51.510 96.010 -50.180 ;
        RECT 96.190 -50.540 96.370 -49.810 ;
        RECT 96.540 -50.220 96.860 -49.340 ;
        RECT 96.190 -50.620 96.510 -50.540 ;
        RECT 96.180 -50.800 96.510 -50.620 ;
        RECT 96.690 -50.800 96.860 -50.220 ;
        RECT 97.955 -50.290 98.370 -49.340 ;
        RECT 97.230 -50.450 98.370 -50.290 ;
        RECT 97.230 -50.460 98.640 -50.450 ;
        RECT 97.230 -50.630 97.560 -50.460 ;
        RECT 97.770 -50.800 98.030 -50.640 ;
        RECT 96.690 -50.970 98.030 -50.800 ;
        RECT 98.200 -50.670 98.640 -50.460 ;
        RECT 96.350 -51.450 96.860 -50.970 ;
        RECT 98.200 -51.150 98.370 -50.670 ;
        RECT 97.895 -51.680 98.370 -51.150 ;
        RECT 98.990 -51.720 99.255 -49.020 ;
        RECT 100.015 -49.860 100.345 -49.020 ;
        RECT 101.285 -49.350 101.615 -49.020 ;
        RECT 102.780 -49.350 103.110 -49.170 ;
        RECT 101.285 -49.520 103.110 -49.350 ;
        RECT 101.285 -49.690 101.615 -49.520 ;
        RECT 101.785 -49.860 103.080 -49.690 ;
        RECT 100.015 -50.030 101.955 -49.860 ;
        RECT 99.930 -50.370 101.960 -50.200 ;
        RECT 102.350 -50.300 102.680 -50.030 ;
        RECT 102.350 -50.345 102.580 -50.300 ;
        RECT 99.930 -50.885 100.300 -50.370 ;
        RECT 100.470 -50.885 101.610 -50.540 ;
        RECT 101.780 -50.750 101.960 -50.370 ;
        RECT 102.130 -50.525 102.580 -50.345 ;
        RECT 102.910 -50.470 103.080 -49.860 ;
        RECT 104.125 -50.005 104.455 -49.810 ;
        RECT 104.125 -50.175 105.080 -50.005 ;
        RECT 102.130 -50.930 102.300 -50.525 ;
        RECT 102.750 -50.695 103.080 -50.470 ;
        RECT 103.290 -50.605 104.070 -50.345 ;
        RECT 104.240 -50.605 104.640 -50.345 ;
        RECT 100.445 -51.225 101.715 -51.055 ;
        RECT 100.445 -51.760 100.705 -51.225 ;
        RECT 101.545 -51.670 101.715 -51.225 ;
        RECT 101.885 -51.500 102.300 -50.930 ;
        RECT 102.470 -50.865 103.080 -50.695 ;
        RECT 104.830 -50.775 105.080 -50.175 ;
        RECT 105.700 -50.320 106.020 -49.610 ;
        RECT 105.700 -50.390 106.540 -50.320 ;
        RECT 105.700 -50.490 106.615 -50.390 ;
        RECT 102.470 -51.670 102.640 -50.865 ;
        RECT 103.625 -50.945 105.080 -50.775 ;
        RECT 105.690 -50.905 106.040 -50.660 ;
        RECT 106.350 -50.910 106.615 -50.490 ;
        RECT 103.625 -51.395 103.955 -50.945 ;
        RECT 106.350 -51.075 106.520 -50.910 ;
        RECT 105.700 -51.245 106.520 -51.075 ;
        RECT 105.700 -51.405 106.020 -51.245 ;
        RECT 101.545 -51.840 102.640 -51.670 ;
      LAYER mcon ;
        RECT 8.710 -15.340 8.880 -15.170 ;
        RECT 9.260 -15.370 9.430 -15.200 ;
        RECT 16.820 -15.340 16.990 -15.170 ;
        RECT 17.290 -15.380 17.460 -15.210 ;
        RECT 18.130 -15.370 18.300 -15.200 ;
        RECT 25.520 -15.340 25.690 -15.170 ;
        RECT 25.990 -15.380 26.160 -15.210 ;
        RECT 26.830 -15.370 27.000 -15.200 ;
        RECT 32.020 -15.370 32.190 -15.200 ;
        RECT 82.960 -15.360 83.130 -15.190 ;
        RECT 88.350 -15.380 88.520 -15.210 ;
        RECT 88.820 -15.340 88.990 -15.170 ;
        RECT 97.050 -15.380 97.220 -15.210 ;
        RECT 97.520 -15.340 97.690 -15.170 ;
        RECT 105.630 -15.340 105.800 -15.170 ;
        RECT 57.030 -49.880 57.200 -49.710 ;
        RECT 57.190 -50.810 57.360 -50.640 ;
        RECT 57.720 -50.810 57.890 -50.640 ;
        RECT 58.630 -49.940 58.800 -49.770 ;
        RECT 60.240 -50.430 60.410 -50.260 ;
        RECT 61.460 -50.540 61.630 -50.370 ;
        RECT 63.330 -50.540 63.500 -50.370 ;
        RECT 73.120 -50.165 73.290 -49.995 ;
        RECT 75.945 -50.545 76.115 -50.375 ;
        RECT 81.760 -49.760 81.930 -49.590 ;
        RECT 84.585 -50.545 84.755 -50.375 ;
        RECT 90.410 -50.275 90.580 -50.105 ;
        RECT 93.225 -50.545 93.395 -50.375 ;
        RECT 99.030 -50.850 99.220 -50.665 ;
        RECT 102.430 -50.220 102.600 -50.050 ;
        RECT 100.025 -50.810 100.225 -50.640 ;
        RECT 100.900 -50.745 101.070 -50.575 ;
        RECT 103.480 -50.595 103.660 -50.415 ;
        RECT 104.355 -50.565 104.545 -50.395 ;
        RECT 101.965 -51.120 102.135 -50.950 ;
        RECT 105.815 -50.895 105.995 -50.705 ;
      LAYER met1 ;
        RECT 8.640 -15.120 8.940 -15.110 ;
        RECT 8.610 -15.490 9.040 -15.120 ;
        RECT 9.800 -15.160 10.100 -15.150 ;
        RECT 9.180 -15.400 10.130 -15.160 ;
        RECT 9.700 -15.530 10.130 -15.400 ;
        RECT 16.350 -15.460 17.020 -15.090 ;
        RECT 17.240 -15.160 17.580 -15.130 ;
        RECT 18.670 -15.160 18.970 -15.150 ;
        RECT 17.230 -15.460 17.580 -15.160 ;
        RECT 18.050 -15.400 19.000 -15.160 ;
        RECT 16.380 -15.470 16.680 -15.460 ;
        RECT 17.240 -15.490 17.580 -15.460 ;
        RECT 18.570 -15.530 19.000 -15.400 ;
        RECT 25.050 -15.460 25.720 -15.090 ;
        RECT 25.940 -15.160 26.280 -15.130 ;
        RECT 27.370 -15.160 27.670 -15.150 ;
        RECT 25.930 -15.460 26.280 -15.160 ;
        RECT 26.750 -15.400 27.700 -15.160 ;
        RECT 25.080 -15.470 25.380 -15.460 ;
        RECT 25.940 -15.490 26.280 -15.460 ;
        RECT 27.270 -15.530 27.700 -15.400 ;
        RECT 31.220 -15.460 31.650 -15.090 ;
        RECT 32.560 -15.160 32.860 -15.150 ;
        RECT 81.650 -15.160 81.950 -15.150 ;
        RECT 31.940 -15.400 32.890 -15.160 ;
        RECT 31.250 -15.470 31.550 -15.460 ;
        RECT 32.460 -15.530 32.890 -15.400 ;
        RECT 81.620 -15.400 82.570 -15.160 ;
        RECT 81.620 -15.530 82.050 -15.400 ;
        RECT 82.860 -15.460 83.290 -15.090 ;
        RECT 86.840 -15.160 87.140 -15.150 ;
        RECT 88.230 -15.160 88.570 -15.130 ;
        RECT 86.810 -15.400 87.760 -15.160 ;
        RECT 82.960 -15.470 83.260 -15.460 ;
        RECT 86.810 -15.530 87.240 -15.400 ;
        RECT 88.230 -15.460 88.580 -15.160 ;
        RECT 88.790 -15.460 89.460 -15.090 ;
        RECT 95.540 -15.160 95.840 -15.150 ;
        RECT 96.930 -15.160 97.270 -15.130 ;
        RECT 95.510 -15.400 96.460 -15.160 ;
        RECT 88.230 -15.490 88.570 -15.460 ;
        RECT 89.130 -15.470 89.430 -15.460 ;
        RECT 95.510 -15.530 95.940 -15.400 ;
        RECT 96.930 -15.460 97.280 -15.160 ;
        RECT 97.490 -15.460 98.160 -15.090 ;
        RECT 105.570 -15.120 105.870 -15.110 ;
        RECT 104.410 -15.160 104.710 -15.150 ;
        RECT 104.380 -15.400 105.330 -15.160 ;
        RECT 96.930 -15.490 97.270 -15.460 ;
        RECT 97.830 -15.470 98.130 -15.460 ;
        RECT 104.380 -15.530 104.810 -15.400 ;
        RECT 105.470 -15.490 105.900 -15.120 ;
        RECT 81.700 -49.605 81.990 -49.530 ;
        RECT 84.525 -49.605 100.960 -49.595 ;
        RECT 56.970 -49.700 57.240 -49.670 ;
        RECT 56.970 -49.890 58.830 -49.700 ;
        RECT 81.700 -49.765 100.960 -49.605 ;
        RECT 81.700 -49.820 81.990 -49.765 ;
        RECT 56.970 -49.920 57.240 -49.890 ;
        RECT 58.600 -50.010 58.830 -49.890 ;
        RECT 73.060 -49.995 73.355 -49.960 ;
        RECT 73.060 -50.165 76.195 -49.995 ;
        RECT 60.190 -50.260 60.460 -50.180 ;
        RECT 73.060 -50.205 73.355 -50.165 ;
        RECT 60.190 -50.430 61.680 -50.260 ;
        RECT 60.190 -50.510 60.460 -50.430 ;
        RECT 57.100 -50.550 57.360 -50.535 ;
        RECT 57.725 -50.545 58.105 -50.515 ;
        RECT 57.100 -50.890 57.440 -50.550 ;
        RECT 57.650 -50.890 58.105 -50.545 ;
        RECT 57.100 -50.905 57.360 -50.890 ;
        RECT 57.725 -50.925 58.105 -50.890 ;
        RECT 59.710 -50.940 59.980 -50.600 ;
        RECT 61.410 -50.620 61.680 -50.430 ;
        RECT 63.300 -50.620 63.550 -50.260 ;
        RECT 75.870 -50.575 76.195 -50.165 ;
        RECT 84.580 -50.325 84.795 -49.765 ;
        RECT 90.345 -50.105 90.650 -50.045 ;
        RECT 90.345 -50.275 93.425 -50.105 ;
        RECT 84.525 -50.580 84.825 -50.325 ;
        RECT 90.345 -50.335 90.650 -50.275 ;
        RECT 59.760 -51.210 59.930 -50.940 ;
        RECT 63.330 -51.210 63.500 -50.620 ;
        RECT 93.165 -50.675 93.425 -50.275 ;
        RECT 100.775 -50.490 100.960 -49.765 ;
        RECT 102.365 -50.195 104.620 -50.005 ;
        RECT 102.365 -50.250 102.680 -50.195 ;
        RECT 100.625 -50.500 101.565 -50.490 ;
        RECT 103.290 -50.500 104.015 -50.350 ;
        RECT 99.000 -50.920 100.295 -50.595 ;
        RECT 100.625 -50.745 104.015 -50.500 ;
        RECT 104.245 -50.605 104.620 -50.195 ;
        RECT 100.625 -50.825 101.565 -50.745 ;
        RECT 101.895 -50.940 102.205 -50.895 ;
        RECT 105.755 -50.940 106.055 -50.620 ;
        RECT 101.895 -51.120 106.055 -50.940 ;
        RECT 101.895 -51.190 102.205 -51.120 ;
        RECT 59.760 -51.380 63.500 -51.210 ;
      LAYER via ;
        RECT 8.660 -15.400 8.920 -15.140 ;
        RECT 9.820 -15.440 10.080 -15.180 ;
        RECT 16.400 -15.440 16.660 -15.180 ;
        RECT 17.260 -15.440 17.520 -15.180 ;
        RECT 18.690 -15.440 18.950 -15.180 ;
        RECT 25.100 -15.440 25.360 -15.180 ;
        RECT 25.960 -15.440 26.220 -15.180 ;
        RECT 27.390 -15.440 27.650 -15.180 ;
        RECT 31.270 -15.440 31.530 -15.180 ;
        RECT 32.580 -15.440 32.840 -15.180 ;
        RECT 81.670 -15.440 81.930 -15.180 ;
        RECT 82.980 -15.440 83.240 -15.180 ;
        RECT 86.860 -15.440 87.120 -15.180 ;
        RECT 88.290 -15.440 88.550 -15.180 ;
        RECT 89.150 -15.440 89.410 -15.180 ;
        RECT 95.560 -15.440 95.820 -15.180 ;
        RECT 96.990 -15.440 97.250 -15.180 ;
        RECT 97.850 -15.440 98.110 -15.180 ;
        RECT 104.430 -15.440 104.690 -15.180 ;
        RECT 105.590 -15.400 105.850 -15.140 ;
        RECT 57.100 -50.840 57.360 -50.580 ;
        RECT 57.720 -50.845 57.980 -50.585 ;
      LAYER met2 ;
        RECT 8.610 -15.460 8.970 -15.080 ;
        RECT 9.770 -15.500 10.130 -15.120 ;
        RECT 16.350 -15.500 16.710 -15.120 ;
        RECT 17.200 -15.490 17.580 -15.130 ;
        RECT 18.640 -15.500 19.000 -15.120 ;
        RECT 25.050 -15.500 25.410 -15.120 ;
        RECT 25.900 -15.490 26.280 -15.130 ;
        RECT 27.340 -15.500 27.700 -15.120 ;
        RECT 31.220 -15.500 31.580 -15.120 ;
        RECT 32.530 -15.500 32.890 -15.120 ;
        RECT 81.620 -15.500 81.980 -15.120 ;
        RECT 82.930 -15.500 83.290 -15.120 ;
        RECT 86.810 -15.500 87.170 -15.120 ;
        RECT 88.230 -15.490 88.610 -15.130 ;
        RECT 89.100 -15.500 89.460 -15.120 ;
        RECT 95.510 -15.500 95.870 -15.120 ;
        RECT 96.930 -15.490 97.310 -15.130 ;
        RECT 97.800 -15.500 98.160 -15.120 ;
        RECT 104.380 -15.500 104.740 -15.120 ;
        RECT 105.540 -15.460 105.900 -15.080 ;
        RECT 57.030 -50.925 57.360 -50.525 ;
        RECT 57.725 -50.555 58.105 -50.515 ;
        RECT 57.720 -50.875 58.105 -50.555 ;
        RECT 57.725 -50.925 58.105 -50.875 ;
      LAYER via2 ;
        RECT 8.650 -15.410 8.930 -15.130 ;
        RECT 9.810 -15.450 10.090 -15.170 ;
        RECT 16.390 -15.450 16.670 -15.170 ;
        RECT 17.250 -15.450 17.530 -15.170 ;
        RECT 18.680 -15.450 18.960 -15.170 ;
        RECT 25.090 -15.450 25.370 -15.170 ;
        RECT 25.950 -15.450 26.230 -15.170 ;
        RECT 27.380 -15.450 27.660 -15.170 ;
        RECT 31.260 -15.450 31.540 -15.170 ;
        RECT 32.570 -15.450 32.850 -15.170 ;
        RECT 81.660 -15.450 81.940 -15.170 ;
        RECT 82.970 -15.450 83.250 -15.170 ;
        RECT 86.850 -15.450 87.130 -15.170 ;
        RECT 88.280 -15.450 88.560 -15.170 ;
        RECT 89.140 -15.450 89.420 -15.170 ;
        RECT 95.550 -15.450 95.830 -15.170 ;
        RECT 96.980 -15.450 97.260 -15.170 ;
        RECT 97.840 -15.450 98.120 -15.170 ;
        RECT 104.420 -15.450 104.700 -15.170 ;
        RECT 105.580 -15.410 105.860 -15.130 ;
        RECT 57.030 -50.880 57.315 -50.570 ;
        RECT 57.775 -50.880 58.055 -50.560 ;
      LAYER met3 ;
        RECT 8.550 -15.490 9.040 -15.010 ;
        RECT 8.600 -15.530 9.040 -15.490 ;
        RECT 9.700 -15.570 10.190 -15.050 ;
        RECT 16.290 -15.570 16.780 -15.050 ;
        RECT 17.130 -15.560 17.650 -15.070 ;
        RECT 18.570 -15.570 19.060 -15.050 ;
        RECT 24.990 -15.570 25.480 -15.050 ;
        RECT 25.830 -15.560 26.350 -15.070 ;
        RECT 27.270 -15.570 27.760 -15.050 ;
        RECT 31.160 -15.570 31.650 -15.050 ;
        RECT 32.460 -15.510 32.950 -15.050 ;
        RECT 81.560 -15.510 82.050 -15.050 ;
        RECT 32.460 -15.570 32.880 -15.510 ;
        RECT 81.630 -15.570 82.050 -15.510 ;
        RECT 82.860 -15.570 83.350 -15.050 ;
        RECT 86.750 -15.570 87.240 -15.050 ;
        RECT 88.160 -15.560 88.680 -15.070 ;
        RECT 89.030 -15.570 89.520 -15.050 ;
        RECT 95.450 -15.570 95.940 -15.050 ;
        RECT 96.860 -15.560 97.380 -15.070 ;
        RECT 97.730 -15.570 98.220 -15.050 ;
        RECT 104.320 -15.570 104.810 -15.050 ;
        RECT 105.470 -15.490 105.960 -15.010 ;
        RECT 105.470 -15.530 105.910 -15.490 ;
        RECT 56.575 -50.910 57.360 -50.535 ;
        RECT 57.720 -50.910 58.505 -50.535 ;
      LAYER via3 ;
        RECT 8.630 -15.430 8.950 -15.110 ;
        RECT 9.790 -15.470 10.110 -15.150 ;
        RECT 16.370 -15.470 16.690 -15.150 ;
        RECT 17.230 -15.470 17.550 -15.150 ;
        RECT 18.660 -15.470 18.980 -15.150 ;
        RECT 25.070 -15.470 25.390 -15.150 ;
        RECT 25.930 -15.470 26.250 -15.150 ;
        RECT 27.360 -15.470 27.680 -15.150 ;
        RECT 31.240 -15.470 31.560 -15.150 ;
        RECT 32.550 -15.470 32.870 -15.150 ;
        RECT 81.640 -15.470 81.960 -15.150 ;
        RECT 82.950 -15.470 83.270 -15.150 ;
        RECT 86.830 -15.470 87.150 -15.150 ;
        RECT 88.260 -15.470 88.580 -15.150 ;
        RECT 89.120 -15.470 89.440 -15.150 ;
        RECT 95.530 -15.470 95.850 -15.150 ;
        RECT 96.960 -15.470 97.280 -15.150 ;
        RECT 97.820 -15.470 98.140 -15.150 ;
        RECT 104.400 -15.470 104.720 -15.150 ;
        RECT 105.560 -15.430 105.880 -15.110 ;
        RECT 56.990 -50.890 57.315 -50.555 ;
        RECT 57.775 -50.885 58.095 -50.550 ;
      LAYER met4 ;
        RECT -24.120 -15.110 -23.820 31.030 ;
        RECT -20.900 -12.500 56.060 28.620 ;
        RECT 58.450 -12.500 135.410 28.620 ;
        RECT 8.530 -15.110 8.960 -15.080 ;
        RECT -24.120 -15.410 8.960 -15.110 ;
        RECT 8.530 -15.440 8.960 -15.410 ;
        RECT 9.780 -15.480 11.300 -15.120 ;
        RECT 10.920 -15.500 11.300 -15.480 ;
        RECT 15.200 -15.140 15.580 -15.130 ;
        RECT 15.200 -15.500 16.700 -15.140 ;
        RECT 17.200 -15.480 17.560 -12.500 ;
        RECT 18.650 -15.480 20.120 -15.120 ;
        RECT 24.060 -15.500 25.400 -15.140 ;
        RECT 25.900 -15.480 26.260 -15.130 ;
        RECT 27.350 -15.480 28.780 -15.120 ;
        RECT 15.200 -15.510 15.580 -15.500 ;
        RECT 25.930 -17.970 26.250 -15.480 ;
        RECT 30.260 -15.500 31.570 -15.140 ;
        RECT 32.500 -17.970 33.000 -15.090 ;
        RECT 81.510 -17.970 82.010 -15.090 ;
        RECT 82.940 -15.500 84.250 -15.140 ;
        RECT 85.730 -15.480 87.160 -15.120 ;
        RECT 88.250 -15.480 88.610 -15.130 ;
        RECT 88.260 -17.970 88.580 -15.480 ;
        RECT 89.110 -15.500 90.450 -15.140 ;
        RECT 94.390 -15.480 95.860 -15.120 ;
        RECT 96.950 -15.480 97.310 -12.500 ;
        RECT 105.550 -15.110 105.980 -15.080 ;
        RECT 138.330 -15.110 138.630 31.030 ;
        RECT 98.930 -15.140 99.310 -15.130 ;
        RECT 97.810 -15.500 99.310 -15.140 ;
        RECT 103.210 -15.480 104.730 -15.120 ;
        RECT 105.550 -15.410 138.630 -15.110 ;
        RECT 105.550 -15.440 105.980 -15.410 ;
        RECT 103.210 -15.500 103.590 -15.480 ;
        RECT 98.930 -15.510 99.310 -15.500 ;
        RECT -20.910 -48.250 30.210 -17.970 ;
        RECT 30.770 -48.250 56.060 -17.970 ;
        RECT 58.450 -47.760 83.740 -17.970 ;
        RECT 58.070 -48.250 83.740 -47.760 ;
        RECT 84.300 -48.250 135.420 -17.970 ;
        RECT 55.630 -50.560 55.930 -48.250 ;
        RECT 58.070 -50.240 58.370 -48.250 ;
        RECT 57.980 -50.535 58.370 -50.240 ;
        RECT 56.970 -50.560 57.330 -50.545 ;
        RECT 55.630 -50.860 57.330 -50.560 ;
        RECT 56.970 -50.900 57.330 -50.860 ;
        RECT 57.760 -50.895 58.370 -50.535 ;
  END
END filter_p_m_fin
END LIBRARY

