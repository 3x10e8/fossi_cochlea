magic
tech sky130A
magscale 1 2
timestamp 1654658877
<< error_p >>
rect -963 27652 -862 28197
rect -643 28015 -542 28304
rect 51063 28015 51164 28304
rect -643 27652 -481 28015
rect -619 27610 -481 27652
rect -862 27374 -481 27610
rect -619 27342 -481 27374
rect 51002 27652 51164 28015
rect 51383 27652 51484 28197
rect 51002 27610 51140 27652
rect 51002 27374 51383 27610
rect 51002 27342 51140 27374
rect -963 27012 -862 27332
rect -643 27012 -542 27332
rect 7217 27015 7344 27050
rect -862 26734 -481 26970
rect 7157 26955 7404 26990
rect -619 26692 -481 26734
rect 14147 26725 14556 27045
rect 35965 26725 36374 27045
rect 43177 27015 43304 27050
rect 51063 27012 51164 27332
rect 51383 27012 51484 27332
rect 43117 26955 43364 26990
rect 51002 26734 51383 26970
rect -963 26372 -862 26692
rect -643 26372 -481 26692
rect -619 26330 -481 26372
rect -862 26094 -481 26330
rect 51002 26692 51140 26734
rect 51002 26372 51164 26692
rect 51383 26372 51484 26692
rect 51002 26330 51140 26372
rect -619 26052 -481 26094
rect -963 25732 -862 26052
rect -643 25732 -481 26052
rect 14156 25875 14565 26195
rect 35956 25875 36365 26195
rect 51002 26094 51383 26330
rect 51002 26052 51140 26094
rect -619 25690 -481 25732
rect -862 25454 -481 25690
rect -619 25436 -481 25454
rect 51002 25732 51164 26052
rect 51383 25732 51484 26052
rect 51002 25690 51140 25732
rect 51002 25454 51383 25690
rect 51002 25436 51140 25454
rect -963 25092 -862 25412
rect -643 25250 -542 25412
rect -963 24930 -542 25092
rect 14148 25023 14557 25343
rect 35964 25023 36373 25343
rect 51063 25250 51164 25412
rect 51383 25092 51484 25412
rect 51063 24930 51484 25092
rect 14143 23322 14552 23642
rect 35969 23322 36378 23642
rect 14153 22427 14562 22747
rect 35959 22427 36368 22747
rect 14144 21544 14553 21864
rect 35968 21544 36377 21864
rect 14163 19840 14572 20160
rect 35949 19840 36358 20160
rect 14158 18958 14567 19278
rect 35954 18958 36363 19278
rect 14169 18061 14578 18381
rect 35943 18061 36352 18381
rect 14158 16368 14567 16688
rect 35954 16368 36363 16688
rect 14164 15470 14573 15790
rect 35948 15470 36357 15790
rect 14167 14577 14576 14897
rect 35945 14577 36354 14897
rect 14172 12881 14581 13201
rect 35940 12881 36349 13201
rect 14167 11988 14576 12308
rect 35945 11988 36354 12308
rect 14173 11093 14582 11413
rect 35939 11093 36348 11413
rect 14171 9395 14580 9715
rect 35941 9395 36350 9715
rect 14168 8502 14577 8822
rect 35944 8502 36353 8822
rect 14164 7610 14566 7930
rect 35955 7610 36357 7930
rect 14166 5914 14568 6234
rect 35953 5914 36355 6234
rect 14170 5020 14572 5340
rect 35949 5020 36351 5340
rect 14162 4126 14564 4446
rect 35957 4126 36359 4446
rect 14170 2430 14572 2750
rect 35949 2430 36351 2750
rect 14161 1541 14570 1861
rect 35951 1541 36360 1861
rect 14152 676 14561 996
rect 35960 676 36369 996
<< error_s >>
rect 25000 -342 25201 -318
rect 24722 -578 25201 -342
rect 25320 -342 25521 -318
rect 25320 -578 25799 -342
rect 25042 -1218 25479 -898
rect 24722 -1774 25201 -1538
rect 25000 -1798 25201 -1774
rect 25320 -1774 25799 -1538
rect 25320 -1798 25521 -1774
use comparator  comparator_0 ~/Documents/fossi_cochlea/mag/final_designs/comparator
timestamp 1654474334
transform 1 0 25121 0 1 28763
box -690 -1057 969 1108
use filter  filter_0
timestamp 1654658877
transform 1 0 358 0 1 0
box -1800 -1798 25922 29716
use filter  filter_1
timestamp 1654658877
transform -1 0 50163 0 1 0
box -1800 -1798 25922 29716
<< end >>
