magic
tech sky130B
magscale 1 2
timestamp 1662790266
<< obsli1 >>
rect 1104 2159 190808 17425
<< obsm1 >>
rect 1104 1572 190968 17672
<< metal2 >>
rect 4986 19200 5042 20000
rect 12898 19200 12954 20000
rect 20810 19200 20866 20000
rect 28722 19200 28778 20000
rect 36634 19200 36690 20000
rect 44546 19200 44602 20000
rect 52458 19200 52514 20000
rect 60370 19200 60426 20000
rect 68282 19200 68338 20000
rect 76194 19200 76250 20000
rect 84106 19200 84162 20000
rect 92018 19200 92074 20000
rect 99930 19200 99986 20000
rect 107842 19200 107898 20000
rect 115754 19200 115810 20000
rect 123666 19200 123722 20000
rect 131578 19200 131634 20000
rect 139490 19200 139546 20000
rect 147402 19200 147458 20000
rect 155314 19200 155370 20000
rect 163226 19200 163282 20000
rect 171138 19200 171194 20000
rect 179050 19200 179106 20000
rect 186962 19200 187018 20000
rect 4986 0 5042 800
rect 12898 0 12954 800
rect 20810 0 20866 800
rect 28722 0 28778 800
rect 36634 0 36690 800
rect 44546 0 44602 800
rect 52458 0 52514 800
rect 60370 0 60426 800
rect 68282 0 68338 800
rect 76194 0 76250 800
rect 84106 0 84162 800
rect 92018 0 92074 800
rect 99930 0 99986 800
rect 107842 0 107898 800
rect 115754 0 115810 800
rect 123666 0 123722 800
rect 131578 0 131634 800
rect 139490 0 139546 800
rect 147402 0 147458 800
rect 155314 0 155370 800
rect 163226 0 163282 800
rect 171138 0 171194 800
rect 179050 0 179106 800
rect 186962 0 187018 800
<< obsm2 >>
rect 1582 19144 4930 19258
rect 5098 19144 12842 19258
rect 13010 19144 20754 19258
rect 20922 19144 28666 19258
rect 28834 19144 36578 19258
rect 36746 19144 44490 19258
rect 44658 19144 52402 19258
rect 52570 19144 60314 19258
rect 60482 19144 68226 19258
rect 68394 19144 76138 19258
rect 76306 19144 84050 19258
rect 84218 19144 91962 19258
rect 92130 19144 99874 19258
rect 100042 19144 107786 19258
rect 107954 19144 115698 19258
rect 115866 19144 123610 19258
rect 123778 19144 131522 19258
rect 131690 19144 139434 19258
rect 139602 19144 147346 19258
rect 147514 19144 155258 19258
rect 155426 19144 163170 19258
rect 163338 19144 171082 19258
rect 171250 19144 178994 19258
rect 179162 19144 186906 19258
rect 187074 19144 190962 19258
rect 1582 856 190962 19144
rect 1582 800 4930 856
rect 5098 800 12842 856
rect 13010 800 20754 856
rect 20922 800 28666 856
rect 28834 800 36578 856
rect 36746 800 44490 856
rect 44658 800 52402 856
rect 52570 800 60314 856
rect 60482 800 68226 856
rect 68394 800 76138 856
rect 76306 800 84050 856
rect 84218 800 91962 856
rect 92130 800 99874 856
rect 100042 800 107786 856
rect 107954 800 115698 856
rect 115866 800 123610 856
rect 123778 800 131522 856
rect 131690 800 139434 856
rect 139602 800 147346 856
rect 147514 800 155258 856
rect 155426 800 163170 856
rect 163338 800 171082 856
rect 171250 800 178994 856
rect 179162 800 186906 856
rect 187074 800 190962 856
<< metal3 >>
rect 191200 17280 192000 17400
rect 0 16600 800 16720
rect 191200 12384 192000 12504
rect 0 9936 800 10056
rect 191200 7488 192000 7608
rect 0 3272 800 3392
rect 191200 2592 192000 2712
<< obsm3 >>
rect 800 17200 191120 17441
rect 800 16800 191200 17200
rect 880 16520 191200 16800
rect 800 12584 191200 16520
rect 800 12304 191120 12584
rect 800 10136 191200 12304
rect 880 9856 191200 10136
rect 800 7688 191200 9856
rect 800 7408 191120 7688
rect 800 3472 191200 7408
rect 880 3192 191200 3472
rect 800 2792 191200 3192
rect 800 2512 191120 2792
rect 800 1939 191200 2512
<< metal4 >>
rect 24657 2128 24977 17456
rect 48370 2128 48690 17456
rect 72083 2128 72403 17456
rect 95796 2128 96116 17456
rect 119509 2128 119829 17456
rect 143222 2128 143542 17456
rect 166935 2128 167255 17456
rect 190648 2128 190968 17456
<< obsm4 >>
rect 51579 2211 72003 13293
rect 72483 2211 82741 13293
<< labels >>
rlabel metal2 s 28722 19200 28778 20000 6 cclk_I[0]
port 1 nsew signal output
rlabel metal2 s 76194 19200 76250 20000 6 cclk_I[1]
port 2 nsew signal output
rlabel metal2 s 123666 19200 123722 20000 6 cclk_I[2]
port 3 nsew signal output
rlabel metal2 s 171138 19200 171194 20000 6 cclk_I[3]
port 4 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 cclk_Q[0]
port 5 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 cclk_Q[1]
port 6 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 cclk_Q[2]
port 7 nsew signal output
rlabel metal2 s 171138 0 171194 800 6 cclk_Q[3]
port 8 nsew signal output
rlabel metal3 s 0 3272 800 3392 6 clk_master
port 9 nsew signal input
rlabel metal2 s 20810 19200 20866 20000 6 clkdiv2_I[0]
port 10 nsew signal output
rlabel metal2 s 68282 19200 68338 20000 6 clkdiv2_I[1]
port 11 nsew signal output
rlabel metal2 s 115754 19200 115810 20000 6 clkdiv2_I[2]
port 12 nsew signal output
rlabel metal2 s 163226 19200 163282 20000 6 clkdiv2_I[3]
port 13 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 clkdiv2_Q[0]
port 14 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 clkdiv2_Q[1]
port 15 nsew signal output
rlabel metal2 s 115754 0 115810 800 6 clkdiv2_Q[2]
port 16 nsew signal output
rlabel metal2 s 163226 0 163282 800 6 clkdiv2_Q[3]
port 17 nsew signal output
rlabel metal2 s 44546 19200 44602 20000 6 comp_high_I[0]
port 18 nsew signal input
rlabel metal2 s 92018 19200 92074 20000 6 comp_high_I[1]
port 19 nsew signal input
rlabel metal2 s 139490 19200 139546 20000 6 comp_high_I[2]
port 20 nsew signal input
rlabel metal2 s 186962 19200 187018 20000 6 comp_high_I[3]
port 21 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 comp_high_Q[0]
port 22 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 comp_high_Q[1]
port 23 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 comp_high_Q[2]
port 24 nsew signal input
rlabel metal2 s 186962 0 187018 800 6 comp_high_Q[3]
port 25 nsew signal input
rlabel metal2 s 4986 19200 5042 20000 6 cos_out[0]
port 26 nsew signal output
rlabel metal2 s 52458 19200 52514 20000 6 cos_out[1]
port 27 nsew signal output
rlabel metal2 s 99930 19200 99986 20000 6 cos_out[2]
port 28 nsew signal output
rlabel metal2 s 147402 19200 147458 20000 6 cos_out[3]
port 29 nsew signal output
rlabel metal2 s 12898 19200 12954 20000 6 fb1_I[0]
port 30 nsew signal output
rlabel metal2 s 60370 19200 60426 20000 6 fb1_I[1]
port 31 nsew signal output
rlabel metal2 s 107842 19200 107898 20000 6 fb1_I[2]
port 32 nsew signal output
rlabel metal2 s 155314 19200 155370 20000 6 fb1_I[3]
port 33 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 fb1_Q[0]
port 34 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 fb1_Q[1]
port 35 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 fb1_Q[2]
port 36 nsew signal output
rlabel metal2 s 155314 0 155370 800 6 fb1_Q[3]
port 37 nsew signal output
rlabel metal2 s 36634 19200 36690 20000 6 phi1b_dig_I[0]
port 38 nsew signal input
rlabel metal2 s 84106 19200 84162 20000 6 phi1b_dig_I[1]
port 39 nsew signal input
rlabel metal2 s 131578 19200 131634 20000 6 phi1b_dig_I[2]
port 40 nsew signal input
rlabel metal2 s 179050 19200 179106 20000 6 phi1b_dig_I[3]
port 41 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 phi1b_dig_Q[0]
port 42 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 phi1b_dig_Q[1]
port 43 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 phi1b_dig_Q[2]
port 44 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 phi1b_dig_Q[3]
port 45 nsew signal input
rlabel metal3 s 191200 17280 192000 17400 6 read_out_I[0]
port 46 nsew signal output
rlabel metal3 s 191200 12384 192000 12504 6 read_out_I[1]
port 47 nsew signal output
rlabel metal3 s 191200 7488 192000 7608 6 read_out_Q[0]
port 48 nsew signal output
rlabel metal3 s 191200 2592 192000 2712 6 read_out_Q[1]
port 49 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 rstb
port 50 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 sin_out[0]
port 51 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 sin_out[1]
port 52 nsew signal output
rlabel metal2 s 99930 0 99986 800 6 sin_out[2]
port 53 nsew signal output
rlabel metal2 s 147402 0 147458 800 6 sin_out[3]
port 54 nsew signal output
rlabel metal3 s 0 9936 800 10056 6 ud_en
port 55 nsew signal input
rlabel metal4 s 24657 2128 24977 17456 6 vccd1
port 56 nsew power bidirectional
rlabel metal4 s 72083 2128 72403 17456 6 vccd1
port 56 nsew power bidirectional
rlabel metal4 s 119509 2128 119829 17456 6 vccd1
port 56 nsew power bidirectional
rlabel metal4 s 166935 2128 167255 17456 6 vccd1
port 56 nsew power bidirectional
rlabel metal4 s 48370 2128 48690 17456 6 vssd1
port 57 nsew ground bidirectional
rlabel metal4 s 95796 2128 96116 17456 6 vssd1
port 57 nsew ground bidirectional
rlabel metal4 s 143222 2128 143542 17456 6 vssd1
port 57 nsew ground bidirectional
rlabel metal4 s 190648 2128 190968 17456 6 vssd1
port 57 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 192000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7416256
string GDS_FILE /local_disk/fossi_cochlea/openlane/digital_unison/runs/22_09_09_23_08/results/signoff/digital_unison.magic.gds
string GDS_START 579666
<< end >>

