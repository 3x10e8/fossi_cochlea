magic
tech sky130A
magscale 1 2
timestamp 1654658877
<< error_p >>
rect 25000 71517 25201 71541
rect 24722 71281 25201 71517
rect 25320 71517 25521 71541
rect 25320 71281 25799 71517
rect 25042 70641 25479 70961
rect 24722 70085 25201 70321
rect 25000 70061 25201 70085
rect 25320 70085 25799 70321
rect 25320 70061 25521 70085
rect 14152 68747 14561 69067
rect 35960 68747 36369 69067
rect 14161 67882 14570 68202
rect 35951 67882 36360 68202
rect 14170 66993 14572 67313
rect 35949 66993 36351 67313
rect 14162 65297 14564 65617
rect 35957 65297 36359 65617
rect 14170 64403 14572 64723
rect 35949 64403 36351 64723
rect 14166 63509 14568 63829
rect 35953 63509 36355 63829
rect 14164 61813 14566 62133
rect 35955 61813 36357 62133
rect 14168 60921 14577 61241
rect 35944 60921 36353 61241
rect 14171 60028 14580 60348
rect 35941 60028 36350 60348
rect 14173 58330 14582 58650
rect 35939 58330 36348 58650
rect 14167 57435 14576 57755
rect 35945 57435 36354 57755
rect 14172 56542 14581 56862
rect 35940 56542 36349 56862
rect 14167 54846 14576 55166
rect 35945 54846 36354 55166
rect 14164 53953 14573 54273
rect 35948 53953 36357 54273
rect 14158 53055 14567 53375
rect 35954 53055 36363 53375
rect 14169 51362 14578 51682
rect 35943 51362 36352 51682
rect 14158 50465 14567 50785
rect 35954 50465 36363 50785
rect 14163 49583 14572 49903
rect 35949 49583 36358 49903
rect 14144 47879 14553 48199
rect 35968 47879 36377 48199
rect 14153 46996 14562 47316
rect 35959 46996 36368 47316
rect 14143 46101 14552 46421
rect 35969 46101 36378 46421
rect -963 44651 -542 44813
rect -963 44331 -862 44651
rect -643 44331 -542 44493
rect -222 44331 -200 44507
rect 14148 44400 14557 44720
rect 35964 44400 36373 44720
rect 51063 44651 51484 44813
rect -619 44289 -347 44307
rect -862 44053 -347 44289
rect -297 44187 -200 44331
rect -619 44011 -347 44053
rect -222 44011 -200 44187
rect 50721 44331 50743 44507
rect 51063 44331 51164 44493
rect 51383 44331 51484 44651
rect 50721 44187 50818 44331
rect 50868 44289 51140 44307
rect 50721 44011 50743 44187
rect 50868 44053 51383 44289
rect 50868 44011 51140 44053
rect -963 43691 -862 44011
rect -643 43691 -347 44011
rect -619 43649 -347 43691
rect -862 43413 -347 43649
rect -619 43371 -347 43413
rect -321 43371 -222 43691
rect 14156 43548 14565 43868
rect 35956 43548 36365 43868
rect 50868 43691 51164 44011
rect 51383 43691 51484 44011
rect 50743 43371 50842 43691
rect 50868 43649 51140 43691
rect 50868 43413 51383 43649
rect 50868 43371 51140 43413
rect -963 43051 -862 43371
rect -643 43051 -347 43371
rect 50868 43051 51164 43371
rect 51383 43051 51484 43371
rect -619 43009 -347 43051
rect -862 42974 -347 43009
rect -222 42974 -200 43051
rect -862 42773 -383 42974
rect -321 42731 -222 42974
rect 7157 42753 7404 42788
rect -963 42411 -862 42731
rect -643 42411 -542 42731
rect -222 42411 -200 42731
rect 7217 42693 7344 42728
rect 14147 42698 14556 43018
rect 35965 42698 36374 43018
rect 50721 42974 50743 43051
rect 50868 43009 51140 43051
rect 50868 42974 51383 43009
rect 43117 42753 43364 42788
rect 50743 42731 50842 42974
rect 50904 42773 51383 42974
rect 43177 42693 43304 42728
rect 50721 42411 50743 42731
rect 51063 42411 51164 42731
rect 51383 42411 51484 42731
rect -321 42401 -222 42411
rect 50743 42401 50842 42411
rect -619 42369 -347 42401
rect -862 42133 -347 42369
rect -619 42091 -347 42133
rect -222 42091 -200 42401
rect 50721 42091 50743 42401
rect 50868 42369 51140 42401
rect 50868 42133 51383 42369
rect 50868 42091 51140 42133
rect -963 41546 -862 42091
rect -643 41735 -347 42091
rect -241 41771 -200 42081
rect 50721 41771 50762 42081
rect -241 41759 -222 41771
rect 50743 41759 50762 41771
rect -222 41735 -200 41759
rect -643 41728 -354 41735
rect -306 41729 -200 41735
rect -643 41439 -542 41728
rect -222 41582 -200 41729
rect 50721 41735 50743 41759
rect 50868 41735 51164 42091
rect 50721 41729 50827 41735
rect 50721 41582 50743 41729
rect 50875 41728 51164 41735
rect -222 41451 -163 41582
rect 50684 41451 50743 41582
rect 51063 41439 51164 41728
rect 51383 41546 51484 42091
rect -963 27520 -862 28065
rect -643 27883 -542 28172
rect -222 28029 -163 28160
rect 50684 28029 50743 28160
rect -643 27876 -354 27883
rect -222 27882 -200 28029
rect -306 27876 -200 27882
rect -643 27520 -347 27876
rect -222 27852 -200 27876
rect 50721 27882 50743 28029
rect 51063 27883 51164 28172
rect 50721 27876 50827 27882
rect 50875 27876 51164 27883
rect 50721 27852 50743 27876
rect -241 27840 -222 27852
rect 50743 27840 50762 27852
rect -241 27530 -200 27840
rect 50721 27530 50762 27840
rect 50868 27520 51164 27876
rect 51383 27520 51484 28065
rect -619 27478 -347 27520
rect -862 27242 -347 27478
rect -619 27210 -347 27242
rect -222 27210 -200 27520
rect 50721 27210 50743 27520
rect 50868 27478 51140 27520
rect 50868 27242 51383 27478
rect 50868 27210 51140 27242
rect -321 27200 -222 27210
rect 50743 27200 50842 27210
rect -963 26880 -862 27200
rect -643 26880 -542 27200
rect -222 26880 -200 27200
rect 7217 26883 7344 26918
rect -862 26637 -383 26838
rect -321 26637 -222 26880
rect 7157 26823 7404 26858
rect -862 26602 -347 26637
rect -619 26560 -347 26602
rect -222 26560 -200 26637
rect 14147 26593 14556 26913
rect 35965 26593 36374 26913
rect 43177 26883 43304 26918
rect 50721 26880 50743 27200
rect 51063 26880 51164 27200
rect 51383 26880 51484 27200
rect 43117 26823 43364 26858
rect 50743 26637 50842 26880
rect 50904 26637 51383 26838
rect 50721 26560 50743 26637
rect 50868 26602 51383 26637
rect 50868 26560 51140 26602
rect -963 26240 -862 26560
rect -643 26240 -347 26560
rect 50868 26240 51164 26560
rect 51383 26240 51484 26560
rect -619 26198 -347 26240
rect -862 25962 -347 26198
rect -619 25920 -347 25962
rect -321 25920 -222 26240
rect -963 25600 -862 25920
rect -643 25600 -347 25920
rect 14156 25743 14565 26063
rect 35956 25743 36365 26063
rect 50743 25920 50842 26240
rect 50868 26198 51140 26240
rect 50868 25962 51383 26198
rect 50868 25920 51140 25962
rect 50868 25600 51164 25920
rect 51383 25600 51484 25920
rect -619 25558 -347 25600
rect -862 25322 -347 25558
rect -222 25424 -200 25600
rect -619 25304 -347 25322
rect -297 25280 -200 25424
rect -963 24960 -862 25280
rect -643 25118 -542 25280
rect -222 25104 -200 25280
rect 50721 25424 50743 25600
rect 50868 25558 51140 25600
rect 50721 25280 50818 25424
rect 50868 25322 51383 25558
rect 50868 25304 51140 25322
rect -963 24798 -542 24960
rect 14148 24891 14557 25211
rect 35964 24891 36373 25211
rect 50721 25104 50743 25280
rect 51063 25118 51164 25280
rect 51383 24960 51484 25280
rect 51063 24798 51484 24960
rect 14143 23190 14552 23510
rect 35969 23190 36378 23510
rect 14153 22295 14562 22615
rect 35959 22295 36368 22615
rect 14144 21412 14553 21732
rect 35968 21412 36377 21732
rect 14163 19708 14572 20028
rect 35949 19708 36358 20028
rect 14158 18826 14567 19146
rect 35954 18826 36363 19146
rect 14169 17929 14578 18249
rect 35943 17929 36352 18249
rect 14158 16236 14567 16556
rect 35954 16236 36363 16556
rect 14164 15338 14573 15658
rect 35948 15338 36357 15658
rect 14167 14445 14576 14765
rect 35945 14445 36354 14765
rect 14172 12749 14581 13069
rect 35940 12749 36349 13069
rect 14167 11856 14576 12176
rect 35945 11856 36354 12176
rect 14173 10961 14582 11281
rect 35939 10961 36348 11281
rect 14171 9263 14580 9583
rect 35941 9263 36350 9583
rect 14168 8370 14577 8690
rect 35944 8370 36353 8690
rect 14164 7478 14566 7798
rect 35955 7478 36357 7798
rect 14166 5782 14568 6102
rect 35953 5782 36355 6102
rect 14170 4888 14572 5208
rect 35949 4888 36351 5208
rect 14162 3994 14564 4314
rect 35957 3994 36359 4314
rect 14170 2298 14572 2618
rect 35949 2298 36351 2618
rect 14161 1409 14570 1729
rect 35951 1409 36360 1729
rect 14152 544 14561 864
rect 35960 544 36369 864
rect 25000 -474 25201 -450
rect 24722 -710 25201 -474
rect 25320 -474 25521 -450
rect 25320 -710 25799 -474
rect 25042 -1350 25479 -1030
rect 24722 -1906 25201 -1670
rect 25000 -1930 25201 -1906
rect 25320 -1906 25799 -1670
rect 25320 -1930 25521 -1906
use filter_p_m  filter_p_m_0
timestamp 1654658877
transform 1 0 0 0 -1 69743
box -1442 -1798 51963 29871
use filter_p_m  filter_p_m_1
timestamp 1654658877
transform 1 0 0 0 1 -132
box -1442 -1798 51963 29871
<< end >>
