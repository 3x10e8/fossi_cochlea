magic
tech TECHNAME
magscale 1 2
timestamp 1650466559
<< nwell >>
rect -10 -900 390 0
rect -10 -2485 390 -2125
<< nmos >>
rect 120 -2665 320 -2635
<< pmos >>
rect 120 -2365 320 -2335
<< mvnmos >>
rect 120 -1160 320 -1060
rect 120 -1350 320 -1250
rect 120 -1540 320 -1440
rect 120 -1730 320 -1630
<< mvpmos >>
rect 120 -400 320 -300
rect 120 -740 320 -640
<< ndiff >>
rect 120 -2575 320 -2555
rect 120 -2615 150 -2575
rect 290 -2615 320 -2575
rect 120 -2635 320 -2615
rect 120 -2690 320 -2665
rect 120 -2730 150 -2690
rect 290 -2730 320 -2690
rect 120 -2745 320 -2730
<< pdiff >>
rect 120 -2275 320 -2255
rect 120 -2315 150 -2275
rect 290 -2315 320 -2275
rect 120 -2335 320 -2315
rect 120 -2385 320 -2365
rect 120 -2425 150 -2385
rect 290 -2425 320 -2385
rect 120 -2445 320 -2425
<< mvndiff >>
rect 120 -990 320 -970
rect 120 -1040 150 -990
rect 290 -1040 320 -990
rect 120 -1060 320 -1040
rect 120 -1180 320 -1160
rect 120 -1230 150 -1180
rect 290 -1230 320 -1180
rect 120 -1250 320 -1230
rect 120 -1370 320 -1350
rect 120 -1420 150 -1370
rect 290 -1420 320 -1370
rect 120 -1440 320 -1420
rect 120 -1560 320 -1540
rect 120 -1610 150 -1560
rect 290 -1610 320 -1560
rect 120 -1630 320 -1610
rect 120 -1750 320 -1730
rect 120 -1800 150 -1750
rect 290 -1800 320 -1750
rect 120 -1820 320 -1800
<< mvpdiff >>
rect 120 -230 320 -210
rect 120 -280 150 -230
rect 290 -280 320 -230
rect 120 -300 320 -280
rect 120 -420 320 -400
rect 120 -470 150 -420
rect 290 -470 320 -420
rect 120 -490 320 -470
rect 120 -570 320 -550
rect 120 -620 150 -570
rect 290 -620 320 -570
rect 120 -640 320 -620
rect 120 -760 320 -740
rect 120 -810 150 -760
rect 290 -810 320 -760
rect 120 -830 320 -810
<< ndiffc >>
rect 150 -2615 290 -2575
rect 150 -2730 290 -2690
<< pdiffc >>
rect 150 -2315 290 -2275
rect 150 -2425 290 -2385
<< mvndiffc >>
rect 150 -1040 290 -990
rect 150 -1230 290 -1180
rect 150 -1420 290 -1370
rect 150 -1610 290 -1560
rect 150 -1800 290 -1750
<< mvpdiffc >>
rect 150 -280 290 -230
rect 150 -470 290 -420
rect 150 -620 290 -570
rect 150 -810 290 -760
<< psubdiff >>
rect 120 -2765 320 -2745
rect 120 -2805 150 -2765
rect 290 -2805 320 -2765
rect 120 -2835 320 -2805
<< nsubdiff >>
rect 120 -2195 320 -2165
rect 120 -2235 150 -2195
rect 290 -2235 320 -2195
rect 120 -2255 320 -2235
<< mvpsubdiff >>
rect 120 -1840 320 -1820
rect 120 -1930 150 -1840
rect 290 -1930 320 -1840
rect 120 -1960 320 -1930
<< mvnsubdiff >>
rect 120 -110 320 -70
rect 120 -180 150 -110
rect 290 -180 320 -110
rect 120 -210 320 -180
<< psubdiffcont >>
rect 150 -2805 290 -2765
<< nsubdiffcont >>
rect 150 -2235 290 -2195
<< mvpsubdiffcont >>
rect 150 -1930 290 -1840
<< mvnsubdiffcont >>
rect 150 -180 290 -110
<< poly >>
rect 0 -320 120 -300
rect 0 -380 10 -320
rect 70 -380 120 -320
rect 0 -400 120 -380
rect 320 -400 350 -300
rect 0 -660 120 -640
rect 0 -720 10 -660
rect 70 -720 120 -660
rect 0 -740 120 -720
rect 320 -740 350 -640
rect 0 -1080 120 -1060
rect 0 -1140 10 -1080
rect 70 -1140 120 -1080
rect 0 -1160 120 -1140
rect 320 -1160 350 -1060
rect 0 -1270 120 -1250
rect 0 -1330 10 -1270
rect 70 -1330 120 -1270
rect 0 -1350 120 -1330
rect 320 -1350 350 -1250
rect 0 -1460 120 -1440
rect 0 -1520 10 -1460
rect 70 -1520 120 -1460
rect 0 -1540 120 -1520
rect 320 -1540 350 -1440
rect 0 -1650 120 -1630
rect 0 -1710 10 -1650
rect 70 -1710 120 -1650
rect 0 -1730 120 -1710
rect 320 -1730 350 -1630
rect 0 -2325 70 -2305
rect 0 -2375 10 -2325
rect 60 -2335 70 -2325
rect 60 -2365 120 -2335
rect 320 -2365 350 -2335
rect 60 -2375 70 -2365
rect 0 -2395 70 -2375
rect 0 -2625 70 -2605
rect 0 -2675 10 -2625
rect 60 -2635 70 -2625
rect 60 -2665 120 -2635
rect 320 -2665 350 -2635
rect 60 -2675 70 -2665
rect 0 -2695 70 -2675
<< polycont >>
rect 10 -380 70 -320
rect 10 -720 70 -660
rect 10 -1140 70 -1080
rect 10 -1330 70 -1270
rect 10 -1520 70 -1460
rect 10 -1710 70 -1650
rect 10 -2375 60 -2325
rect 10 -2675 60 -2625
<< locali >>
rect 130 -110 310 -80
rect 130 -180 150 -110
rect 290 -180 310 -110
rect 130 -230 310 -180
rect 130 -280 150 -230
rect 290 -280 310 -230
rect 130 -290 310 -280
rect -10 -320 90 -310
rect -10 -380 10 -320
rect 70 -380 90 -320
rect -10 -390 90 -380
rect 20 -570 60 -390
rect 130 -420 310 -410
rect 130 -470 150 -420
rect 290 -470 310 -420
rect 130 -480 310 -470
rect 130 -570 310 -560
rect 20 -610 150 -570
rect 130 -620 150 -610
rect 290 -620 310 -570
rect 130 -630 310 -620
rect -10 -660 90 -650
rect -10 -720 10 -660
rect 70 -720 90 -660
rect -10 -730 90 -720
rect 130 -760 310 -750
rect 130 -810 150 -760
rect 290 -810 310 -760
rect 130 -820 310 -810
rect 130 -990 310 -980
rect 130 -1040 150 -990
rect 290 -1040 310 -990
rect 130 -1050 310 -1040
rect -10 -1080 90 -1070
rect -10 -1140 10 -1080
rect 70 -1140 90 -1080
rect -10 -1150 90 -1140
rect 130 -1180 310 -1170
rect 130 -1230 150 -1180
rect 290 -1230 310 -1180
rect 130 -1240 310 -1230
rect -10 -1270 95 -1260
rect -10 -1330 10 -1270
rect 70 -1330 95 -1270
rect -10 -1340 95 -1330
rect 130 -1370 310 -1360
rect 130 -1420 150 -1370
rect 290 -1420 310 -1370
rect 130 -1430 310 -1420
rect -10 -1460 90 -1450
rect -10 -1520 10 -1460
rect 70 -1520 90 -1460
rect -10 -1530 90 -1520
rect 130 -1560 310 -1550
rect 130 -1610 150 -1560
rect 290 -1610 310 -1560
rect 130 -1620 310 -1610
rect -10 -1650 95 -1640
rect -10 -1710 10 -1650
rect 70 -1710 95 -1650
rect -10 -1720 95 -1710
rect 130 -1750 310 -1740
rect 130 -1800 150 -1750
rect 290 -1800 310 -1750
rect 130 -1840 310 -1800
rect 130 -1930 150 -1840
rect 290 -1930 310 -1840
rect 130 -1950 310 -1930
rect 130 -2195 310 -2175
rect 130 -2235 150 -2195
rect 290 -2235 310 -2195
rect 130 -2275 310 -2235
rect -10 -2325 70 -2305
rect 130 -2315 150 -2275
rect 290 -2315 310 -2275
rect 130 -2325 310 -2315
rect -10 -2375 10 -2325
rect 60 -2375 70 -2325
rect -10 -2395 70 -2375
rect 130 -2385 310 -2375
rect 10 -2435 50 -2395
rect 130 -2425 150 -2385
rect 290 -2425 310 -2385
rect 130 -2435 310 -2425
rect 0 -2455 80 -2435
rect 0 -2545 10 -2455
rect 70 -2545 80 -2455
rect 0 -2565 80 -2545
rect 180 -2455 260 -2435
rect 180 -2545 190 -2455
rect 250 -2545 260 -2455
rect 180 -2565 260 -2545
rect 10 -2605 50 -2565
rect 130 -2575 310 -2565
rect -10 -2625 70 -2605
rect 130 -2615 150 -2575
rect 290 -2615 310 -2575
rect 130 -2625 310 -2615
rect -10 -2675 10 -2625
rect 60 -2675 70 -2625
rect -10 -2695 70 -2675
rect 130 -2690 310 -2675
rect 130 -2730 150 -2690
rect 290 -2730 310 -2690
rect 130 -2765 310 -2730
rect 130 -2805 150 -2765
rect 290 -2805 310 -2765
rect 130 -2825 310 -2805
<< viali >>
rect 150 -180 290 -110
rect 150 -470 290 -420
rect 150 -620 290 -570
rect 10 -720 70 -660
rect 150 -810 290 -760
rect 150 -1040 290 -990
rect 10 -1140 70 -1080
rect 150 -1230 290 -1180
rect 10 -1330 70 -1270
rect 150 -1420 290 -1370
rect 10 -1520 70 -1460
rect 150 -1610 290 -1560
rect 10 -1710 70 -1650
rect 150 -1930 290 -1840
rect 150 -2235 290 -2195
rect 10 -2545 70 -2455
rect 190 -2545 250 -2455
rect 150 -2805 290 -2765
<< metal1 >>
rect 120 -110 320 -100
rect 120 -115 150 -110
rect -10 -175 150 -115
rect 120 -180 150 -175
rect 290 -115 320 -110
rect 290 -175 390 -115
rect 290 -180 310 -175
rect 120 -190 310 -180
rect 130 -420 310 -410
rect 130 -425 150 -420
rect 18 -465 150 -425
rect 18 -650 62 -465
rect 130 -470 150 -465
rect 290 -470 310 -420
rect 130 -480 310 -470
rect 265 -560 335 -550
rect 130 -570 270 -560
rect 130 -620 150 -570
rect 130 -630 270 -620
rect 330 -630 335 -560
rect 265 -640 335 -630
rect -10 -660 90 -650
rect -10 -720 10 -660
rect 70 -720 90 -660
rect -10 -730 90 -720
rect 130 -760 310 -750
rect -10 -810 150 -760
rect 290 -810 390 -760
rect 130 -820 310 -810
rect 130 -990 310 -980
rect -10 -1040 150 -990
rect 290 -1040 390 -990
rect 130 -1050 310 -1040
rect -10 -1080 90 -1070
rect -10 -1140 10 -1080
rect 70 -1140 90 -1080
rect -10 -1150 90 -1140
rect 130 -1180 180 -1170
rect 240 -1180 310 -1170
rect 130 -1230 150 -1180
rect 290 -1230 310 -1180
rect 130 -1240 310 -1230
rect -10 -1270 95 -1260
rect -10 -1330 10 -1270
rect 70 -1325 95 -1270
rect 156 -1325 166 -1272
rect 70 -1326 166 -1325
rect 70 -1330 95 -1326
rect -10 -1340 95 -1330
rect 130 -1370 310 -1360
rect -10 -1420 150 -1370
rect 290 -1420 390 -1370
rect 130 -1430 310 -1420
rect -10 -1460 90 -1450
rect -10 -1520 10 -1460
rect 70 -1520 170 -1460
rect 230 -1520 240 -1460
rect -10 -1530 90 -1520
rect 270 -1550 340 -1540
rect 130 -1560 270 -1550
rect 130 -1610 150 -1560
rect 130 -1620 270 -1610
rect 330 -1620 340 -1550
rect 270 -1630 340 -1620
rect -10 -1650 95 -1640
rect -10 -1710 5 -1650
rect 75 -1710 95 -1650
rect -10 -1720 95 -1710
rect 130 -1840 310 -1820
rect 130 -1850 150 -1840
rect -10 -1920 150 -1850
rect 130 -1930 150 -1920
rect 290 -1850 310 -1840
rect 290 -1920 390 -1850
rect 290 -1930 310 -1920
rect 130 -1950 310 -1930
rect 130 -2185 310 -2175
rect -10 -2195 390 -2185
rect -10 -2235 150 -2195
rect 290 -2235 390 -2195
rect -10 -2245 390 -2235
rect 130 -2255 310 -2245
rect 0 -2455 80 -2435
rect 0 -2545 10 -2455
rect 70 -2545 80 -2455
rect 0 -2565 80 -2545
rect 180 -2455 260 -2425
rect 180 -2545 190 -2455
rect 250 -2545 260 -2455
rect 180 -2575 260 -2545
rect 130 -2755 310 -2745
rect -10 -2765 390 -2755
rect -10 -2805 150 -2765
rect 290 -2805 390 -2765
rect -10 -2815 390 -2805
rect 130 -2825 310 -2815
<< via1 >>
rect 270 -570 330 -560
rect 270 -620 290 -570
rect 290 -620 330 -570
rect 270 -630 330 -620
rect 10 -720 70 -660
rect 10 -1140 70 -1080
rect 180 -1180 240 -1170
rect 180 -1230 240 -1180
rect 95 -1325 156 -1272
rect 10 -1520 70 -1460
rect 170 -1520 230 -1460
rect 270 -1560 330 -1550
rect 270 -1610 290 -1560
rect 290 -1610 330 -1560
rect 270 -1620 330 -1610
rect 5 -1710 10 -1650
rect 10 -1710 70 -1650
rect 70 -1710 75 -1650
rect 10 -2545 70 -2455
rect 190 -2545 250 -2455
<< metal2 >>
rect 265 -560 335 -550
rect 265 -630 270 -560
rect 330 -630 335 -560
rect 265 -640 335 -630
rect -10 -660 90 -650
rect -10 -720 10 -660
rect 70 -670 90 -660
rect 70 -710 230 -670
rect 70 -720 90 -710
rect -10 -730 90 -720
rect 10 -1080 70 -1070
rect 10 -1150 70 -1140
rect 20 -1450 60 -1150
rect 190 -1170 230 -710
rect 170 -1230 180 -1170
rect 240 -1230 250 -1170
rect 90 -1272 170 -1260
rect 90 -1325 95 -1272
rect 156 -1325 170 -1272
rect 90 -1340 170 -1325
rect 10 -1460 70 -1450
rect 10 -1530 70 -1520
rect 100 -1650 140 -1340
rect 170 -1460 230 -1450
rect 170 -1530 230 -1520
rect -5 -1710 5 -1650
rect 75 -1710 140 -1650
rect 20 -2435 60 -1710
rect 180 -2435 220 -1530
rect 280 -1540 320 -640
rect 260 -1550 340 -1540
rect 260 -1620 270 -1550
rect 330 -1620 340 -1550
rect 260 -1630 340 -1620
rect 0 -2455 80 -2435
rect 0 -2545 10 -2455
rect 70 -2545 80 -2455
rect 0 -2565 80 -2545
rect 180 -2455 260 -2435
rect 180 -2545 190 -2455
rect 250 -2545 260 -2455
rect 180 -2565 260 -2545
rect 20 -2835 60 -2565
<< labels >>
rlabel metal1 -10 -150 -10 -150 7 vdda1
port 4 w
rlabel metal1 -10 -1020 -10 -1020 7 vssd1
port 3 w
rlabel metal1 -10 -786 -10 -786 7 vdda1
rlabel metal1 -10 -1396 -10 -1396 7 vdda1
rlabel metal1 -10 -1886 -10 -1886 7 vssd1
rlabel polycont 40 -350 40 -350 1 outb
port 5 n
rlabel viali 220 -444 220 -444 1 out
port 6 n
rlabel metal1 390 -2791 390 -2791 7 vssd1
rlabel metal1 390 -2215 390 -2215 7 vccd1
port 2 w
rlabel metal1 -10 -2791 -10 -2791 7 vssd1
rlabel metal2 40 -2835 40 -2835 5 in
port 1 s
rlabel metal1 -10 -2215 -10 -2215 7 vccd1
port 2 w
<< end >>
