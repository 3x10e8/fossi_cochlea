magic
tech sky130A
magscale 1 2
timestamp 1654714494
<< obsli1 >>
rect 1104 2159 78844 57681
<< obsm1 >>
rect 1104 2128 78844 59152
<< metal2 >>
rect 1674 59200 1730 60000
rect 5078 59200 5134 60000
rect 8574 59200 8630 60000
rect 12070 59200 12126 60000
rect 15566 59200 15622 60000
rect 19062 59200 19118 60000
rect 22466 59200 22522 60000
rect 25962 59200 26018 60000
rect 29458 59200 29514 60000
rect 32954 59200 33010 60000
rect 36450 59200 36506 60000
rect 39946 59200 40002 60000
rect 43350 59200 43406 60000
rect 46846 59200 46902 60000
rect 50342 59200 50398 60000
rect 53838 59200 53894 60000
rect 57334 59200 57390 60000
rect 60830 59200 60886 60000
rect 64234 59200 64290 60000
rect 67730 59200 67786 60000
rect 71226 59200 71282 60000
rect 74722 59200 74778 60000
rect 78218 59200 78274 60000
rect 2226 0 2282 800
rect 6642 0 6698 800
rect 11058 0 11114 800
rect 15566 0 15622 800
rect 19982 0 20038 800
rect 24398 0 24454 800
rect 28906 0 28962 800
rect 33322 0 33378 800
rect 37738 0 37794 800
rect 42246 0 42302 800
rect 46662 0 46718 800
rect 51078 0 51134 800
rect 55586 0 55642 800
rect 60002 0 60058 800
rect 64418 0 64474 800
rect 68926 0 68982 800
rect 73342 0 73398 800
rect 77758 0 77814 800
<< obsm2 >>
rect 1398 59144 1618 59945
rect 1786 59144 5022 59945
rect 5190 59144 8518 59945
rect 8686 59144 12014 59945
rect 12182 59144 15510 59945
rect 15678 59144 19006 59945
rect 19174 59144 22410 59945
rect 22578 59144 25906 59945
rect 26074 59144 29402 59945
rect 29570 59144 32898 59945
rect 33066 59144 36394 59945
rect 36562 59144 39890 59945
rect 40058 59144 43294 59945
rect 43462 59144 46790 59945
rect 46958 59144 50286 59945
rect 50454 59144 53782 59945
rect 53950 59144 57278 59945
rect 57446 59144 60774 59945
rect 60942 59144 64178 59945
rect 64346 59144 67674 59945
rect 67842 59144 71170 59945
rect 71338 59144 74666 59945
rect 74834 59144 78162 59945
rect 78330 59144 78550 59945
rect 1398 856 78550 59144
rect 1398 800 2170 856
rect 2338 800 6586 856
rect 6754 800 11002 856
rect 11170 800 15510 856
rect 15678 800 19926 856
rect 20094 800 24342 856
rect 24510 800 28850 856
rect 29018 800 33266 856
rect 33434 800 37682 856
rect 37850 800 42190 856
rect 42358 800 46606 856
rect 46774 800 51022 856
rect 51190 800 55530 856
rect 55698 800 59946 856
rect 60114 800 64362 856
rect 64530 800 68870 856
rect 69038 800 73286 856
rect 73454 800 77702 856
rect 77870 800 78550 856
<< metal3 >>
rect 0 57400 800 57520
rect 79200 55632 80000 55752
rect 0 52368 800 52488
rect 0 47336 800 47456
rect 79200 47064 80000 47184
rect 0 42440 800 42560
rect 79200 38496 80000 38616
rect 0 37408 800 37528
rect 0 32376 800 32496
rect 79200 29928 80000 30048
rect 0 27344 800 27464
rect 0 22448 800 22568
rect 79200 21360 80000 21480
rect 0 17416 800 17536
rect 79200 12792 80000 12912
rect 0 12384 800 12504
rect 0 7352 800 7472
rect 79200 4224 80000 4344
rect 0 2456 800 2576
<< obsm3 >>
rect 800 57600 79200 59941
rect 880 57320 79200 57600
rect 800 55832 79200 57320
rect 800 55552 79120 55832
rect 800 52568 79200 55552
rect 880 52288 79200 52568
rect 800 47536 79200 52288
rect 880 47264 79200 47536
rect 880 47256 79120 47264
rect 800 46984 79120 47256
rect 800 42640 79200 46984
rect 880 42360 79200 42640
rect 800 38696 79200 42360
rect 800 38416 79120 38696
rect 800 37608 79200 38416
rect 880 37328 79200 37608
rect 800 32576 79200 37328
rect 880 32296 79200 32576
rect 800 30128 79200 32296
rect 800 29848 79120 30128
rect 800 27544 79200 29848
rect 880 27264 79200 27544
rect 800 22648 79200 27264
rect 880 22368 79200 22648
rect 800 21560 79200 22368
rect 800 21280 79120 21560
rect 800 17616 79200 21280
rect 880 17336 79200 17616
rect 800 12992 79200 17336
rect 800 12712 79120 12992
rect 800 12584 79200 12712
rect 880 12304 79200 12584
rect 800 7552 79200 12304
rect 880 7272 79200 7552
rect 800 4424 79200 7272
rect 800 4144 79120 4424
rect 800 2656 79200 4144
rect 880 2376 79200 2656
rect 800 2143 79200 2376
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
rect 65648 2128 65968 57712
<< obsm4 >>
rect 5395 57792 75933 59941
rect 5395 2891 19488 57792
rect 19968 2891 34848 57792
rect 35328 2891 50208 57792
rect 50688 2891 65568 57792
rect 66048 2891 75933 57792
<< labels >>
rlabel metal2 s 33322 0 33378 800 6 cclk_I[0]
port 1 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 cclk_I[1]
port 2 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 cclk_Q[0]
port 3 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 cclk_Q[1]
port 4 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 clk_master
port 5 nsew signal input
rlabel metal2 s 25962 59200 26018 60000 6 clk_master_out
port 6 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 clkdiv2_I[0]
port 7 nsew signal output
rlabel metal2 s 64234 59200 64290 60000 6 clkdiv2_I[1]
port 8 nsew signal output
rlabel metal2 s 53838 59200 53894 60000 6 clkdiv2_Q[0]
port 9 nsew signal output
rlabel metal3 s 0 47336 800 47456 6 clkdiv2_Q[1]
port 10 nsew signal output
rlabel metal3 s 0 27344 800 27464 6 comp_high_I[0]
port 11 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 comp_high_I[1]
port 12 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 comp_high_Q[0]
port 13 nsew signal input
rlabel metal2 s 67730 59200 67786 60000 6 comp_high_Q[1]
port 14 nsew signal input
rlabel metal2 s 57334 59200 57390 60000 6 cos_out[0]
port 15 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 cos_out[1]
port 16 nsew signal output
rlabel metal2 s 42246 0 42302 800 6 cos_outb[0]
port 17 nsew signal output
rlabel metal2 s 71226 59200 71282 60000 6 cos_outb[1]
port 18 nsew signal output
rlabel metal2 s 22466 59200 22522 60000 6 div2out
port 19 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 fb1_I[0]
port 20 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 fb1_I[1]
port 21 nsew signal output
rlabel metal3 s 79200 29928 80000 30048 6 fb1_Q[0]
port 22 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 fb1_Q[1]
port 23 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 fb2_I[0]
port 24 nsew signal output
rlabel metal3 s 79200 55632 80000 55752 6 fb2_I[1]
port 25 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 fb2_Q[0]
port 26 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 fb2_Q[1]
port 27 nsew signal output
rlabel metal3 s 79200 21360 80000 21480 6 gray_clk_out[10]
port 28 nsew signal output
rlabel metal2 s 29458 59200 29514 60000 6 gray_clk_out[1]
port 29 nsew signal output
rlabel metal2 s 32954 59200 33010 60000 6 gray_clk_out[2]
port 30 nsew signal output
rlabel metal2 s 36450 59200 36506 60000 6 gray_clk_out[3]
port 31 nsew signal output
rlabel metal2 s 39946 59200 40002 60000 6 gray_clk_out[4]
port 32 nsew signal output
rlabel metal2 s 43350 59200 43406 60000 6 gray_clk_out[5]
port 33 nsew signal output
rlabel metal2 s 46846 59200 46902 60000 6 gray_clk_out[6]
port 34 nsew signal output
rlabel metal2 s 50342 59200 50398 60000 6 gray_clk_out[7]
port 35 nsew signal output
rlabel metal3 s 79200 4224 80000 4344 6 gray_clk_out[8]
port 36 nsew signal output
rlabel metal3 s 79200 12792 80000 12912 6 gray_clk_out[9]
port 37 nsew signal output
rlabel metal3 s 0 2456 800 2576 6 no_ones_below_out[0]
port 38 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 no_ones_below_out[1]
port 39 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 no_ones_below_out[2]
port 40 nsew signal output
rlabel metal3 s 79200 38496 80000 38616 6 phi1b_dig_I[0]
port 41 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 phi1b_dig_I[1]
port 42 nsew signal input
rlabel metal3 s 79200 47064 80000 47184 6 phi1b_dig_Q[0]
port 43 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 phi1b_dig_Q[1]
port 44 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 read_out_I[0]
port 45 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 read_out_I[1]
port 46 nsew signal output
rlabel metal2 s 1674 59200 1730 60000 6 read_out_I_top[0]
port 47 nsew signal output
rlabel metal2 s 5078 59200 5134 60000 6 read_out_I_top[1]
port 48 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 read_out_Q[0]
port 49 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 read_out_Q[1]
port 50 nsew signal output
rlabel metal2 s 8574 59200 8630 60000 6 read_out_Q_top[0]
port 51 nsew signal output
rlabel metal2 s 12070 59200 12126 60000 6 read_out_Q_top[1]
port 52 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 rstb
port 53 nsew signal input
rlabel metal2 s 15566 59200 15622 60000 6 rstb_out
port 54 nsew signal output
rlabel metal2 s 60830 59200 60886 60000 6 sin_out[0]
port 55 nsew signal output
rlabel metal2 s 74722 59200 74778 60000 6 sin_out[1]
port 56 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 sin_outb[0]
port 57 nsew signal output
rlabel metal2 s 78218 59200 78274 60000 6 sin_outb[1]
port 58 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 ud_en
port 59 nsew signal input
rlabel metal2 s 19062 59200 19118 60000 6 ud_en_out
port 60 nsew signal output
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 61 nsew power input
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 61 nsew power input
rlabel metal4 s 65648 2128 65968 57712 6 vccd1
port 61 nsew power input
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 62 nsew ground input
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 62 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 80000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7900218
string GDS_FILE /Volumes/export/isn/abhinav/fossi_cochlea/openlane/first_dual_core/runs/first_dual_core/results/finishing/first_dual_core.magic.gds
string GDS_START 464388
<< end >>

