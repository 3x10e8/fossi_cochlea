magic
tech sky130A
timestamp 1647479110
<< nwell >>
rect 2694 -1643 3074 -1555
<< nmos >>
rect 2739 -1803 2754 -1761
rect 2783 -1803 2798 -1761
rect 2827 -1803 2842 -1761
rect 2871 -1803 2886 -1761
rect 2915 -1803 2930 -1761
rect 2959 -1803 2974 -1761
<< pmos >>
rect 2739 -1625 2754 -1583
rect 2783 -1625 2798 -1583
rect 2827 -1625 2842 -1583
rect 2871 -1625 2886 -1583
rect 2915 -1625 2930 -1583
rect 2959 -1625 2974 -1583
<< ndiff >>
rect 2712 -1773 2739 -1761
rect 2712 -1790 2716 -1773
rect 2733 -1790 2739 -1773
rect 2712 -1803 2739 -1790
rect 2754 -1773 2783 -1761
rect 2754 -1790 2760 -1773
rect 2777 -1790 2783 -1773
rect 2754 -1803 2783 -1790
rect 2798 -1773 2827 -1761
rect 2798 -1790 2804 -1773
rect 2821 -1790 2827 -1773
rect 2798 -1803 2827 -1790
rect 2842 -1773 2871 -1761
rect 2842 -1790 2848 -1773
rect 2865 -1790 2871 -1773
rect 2842 -1803 2871 -1790
rect 2886 -1773 2915 -1761
rect 2886 -1790 2892 -1773
rect 2909 -1790 2915 -1773
rect 2886 -1803 2915 -1790
rect 2930 -1773 2959 -1761
rect 2930 -1790 2936 -1773
rect 2953 -1790 2959 -1773
rect 2930 -1803 2959 -1790
rect 2974 -1773 3001 -1761
rect 2974 -1790 2980 -1773
rect 2997 -1790 3001 -1773
rect 2974 -1803 3001 -1790
<< pdiff >>
rect 2712 -1595 2739 -1583
rect 2712 -1612 2716 -1595
rect 2733 -1612 2739 -1595
rect 2712 -1625 2739 -1612
rect 2754 -1595 2783 -1583
rect 2754 -1612 2760 -1595
rect 2777 -1612 2783 -1595
rect 2754 -1625 2783 -1612
rect 2798 -1595 2827 -1583
rect 2798 -1612 2804 -1595
rect 2821 -1612 2827 -1595
rect 2798 -1625 2827 -1612
rect 2842 -1595 2871 -1583
rect 2842 -1612 2848 -1595
rect 2865 -1612 2871 -1595
rect 2842 -1625 2871 -1612
rect 2886 -1595 2915 -1583
rect 2886 -1612 2892 -1595
rect 2909 -1612 2915 -1595
rect 2886 -1625 2915 -1612
rect 2930 -1595 2959 -1583
rect 2930 -1612 2936 -1595
rect 2953 -1612 2959 -1595
rect 2930 -1625 2959 -1612
rect 2974 -1595 3001 -1583
rect 2974 -1612 2980 -1595
rect 2997 -1612 3001 -1595
rect 2974 -1625 3001 -1612
<< ndiffc >>
rect 2716 -1790 2733 -1773
rect 2760 -1790 2777 -1773
rect 2804 -1790 2821 -1773
rect 2848 -1790 2865 -1773
rect 2892 -1790 2909 -1773
rect 2936 -1790 2953 -1773
rect 2980 -1790 2997 -1773
<< pdiffc >>
rect 2716 -1612 2733 -1595
rect 2760 -1612 2777 -1595
rect 2804 -1612 2821 -1595
rect 2848 -1612 2865 -1595
rect 2892 -1612 2909 -1595
rect 2936 -1612 2953 -1595
rect 2980 -1612 2997 -1595
<< psubdiff >>
rect 2716 -1879 2743 -1866
rect 2716 -1896 2721 -1879
rect 2738 -1896 2743 -1879
rect 2716 -1908 2743 -1896
<< nsubdiff >>
rect 3029 -1596 3056 -1583
rect 3029 -1613 3034 -1596
rect 3051 -1613 3056 -1596
rect 3029 -1625 3056 -1613
<< psubdiffcont >>
rect 2721 -1896 2738 -1879
<< nsubdiffcont >>
rect 3034 -1613 3051 -1596
<< poly >>
rect 2735 -1531 2762 -1523
rect 2735 -1548 2740 -1531
rect 2757 -1534 2762 -1531
rect 2757 -1548 2930 -1534
rect 2735 -1549 2930 -1548
rect 2735 -1557 2762 -1549
rect 2739 -1583 2754 -1557
rect 2783 -1583 2798 -1570
rect 2827 -1583 2842 -1549
rect 2871 -1583 2886 -1570
rect 2915 -1583 2930 -1549
rect 2959 -1583 2974 -1570
rect 2739 -1638 2754 -1625
rect 2675 -1653 2702 -1645
rect 2675 -1670 2680 -1653
rect 2697 -1659 2702 -1653
rect 2783 -1659 2798 -1625
rect 2827 -1638 2842 -1625
rect 2871 -1659 2886 -1625
rect 2915 -1638 2930 -1625
rect 2959 -1659 2974 -1625
rect 2697 -1670 2974 -1659
rect 2675 -1674 2974 -1670
rect 2675 -1679 2702 -1674
rect 2675 -1709 2702 -1701
rect 2675 -1726 2680 -1709
rect 2697 -1712 2702 -1709
rect 2697 -1726 2930 -1712
rect 2675 -1727 2930 -1726
rect 2675 -1735 2702 -1727
rect 2739 -1761 2754 -1727
rect 2783 -1761 2798 -1748
rect 2827 -1761 2842 -1727
rect 2871 -1761 2886 -1748
rect 2915 -1761 2930 -1727
rect 2959 -1761 2974 -1748
rect 2739 -1816 2754 -1803
rect 2783 -1823 2798 -1803
rect 2827 -1816 2842 -1803
rect 2779 -1831 2806 -1823
rect 2779 -1848 2784 -1831
rect 2801 -1837 2806 -1831
rect 2871 -1837 2886 -1803
rect 2915 -1816 2930 -1803
rect 2959 -1837 2974 -1803
rect 2801 -1848 2974 -1837
rect 2779 -1852 2974 -1848
rect 2779 -1857 2806 -1852
<< polycont >>
rect 2740 -1548 2757 -1531
rect 2680 -1670 2697 -1653
rect 2680 -1726 2697 -1709
rect 2784 -1848 2801 -1831
<< locali >>
rect 2798 -1326 2828 -1319
rect 2798 -1344 2804 -1326
rect 2822 -1344 2828 -1326
rect 2798 -1351 2828 -1344
rect 2695 -1483 2718 -1477
rect 2695 -1500 2698 -1483
rect 2715 -1500 2718 -1483
rect 2695 -1506 2718 -1500
rect 2698 -1569 2715 -1506
rect 2736 -1531 2761 -1523
rect 2736 -1548 2740 -1531
rect 2757 -1548 2761 -1531
rect 2736 -1557 2761 -1548
rect 2698 -1574 2718 -1569
rect 2698 -1586 2731 -1574
rect 2701 -1587 2731 -1586
rect 2804 -1587 2821 -1351
rect 3035 -1426 3052 -1423
rect 2977 -1486 3000 -1480
rect 2977 -1503 2980 -1486
rect 2997 -1503 3000 -1486
rect 2977 -1509 3000 -1503
rect 2980 -1587 2997 -1509
rect 3035 -1583 3052 -1443
rect 2701 -1591 2735 -1587
rect 2714 -1595 2735 -1591
rect 2714 -1612 2716 -1595
rect 2733 -1612 2735 -1595
rect 2714 -1620 2735 -1612
rect 2758 -1595 2779 -1587
rect 2758 -1612 2760 -1595
rect 2777 -1612 2779 -1595
rect 2758 -1620 2779 -1612
rect 2802 -1595 2823 -1587
rect 2802 -1612 2804 -1595
rect 2821 -1612 2823 -1595
rect 2802 -1620 2823 -1612
rect 2846 -1595 2867 -1587
rect 2846 -1612 2848 -1595
rect 2865 -1612 2867 -1595
rect 2846 -1620 2867 -1612
rect 2890 -1595 2911 -1587
rect 2890 -1612 2892 -1595
rect 2909 -1612 2911 -1595
rect 2890 -1620 2911 -1612
rect 2934 -1595 2955 -1587
rect 2934 -1612 2936 -1595
rect 2953 -1612 2955 -1595
rect 2934 -1620 2955 -1612
rect 2978 -1595 2999 -1587
rect 2978 -1612 2980 -1595
rect 2997 -1612 2999 -1595
rect 2978 -1620 2999 -1612
rect 3029 -1596 3056 -1583
rect 3029 -1613 3034 -1596
rect 3051 -1613 3056 -1596
rect 2676 -1653 2701 -1645
rect 2676 -1670 2680 -1653
rect 2697 -1670 2701 -1653
rect 2676 -1679 2701 -1670
rect 2676 -1709 2701 -1701
rect 2676 -1726 2680 -1709
rect 2697 -1726 2701 -1709
rect 2676 -1735 2701 -1726
rect 2718 -1765 2735 -1620
rect 2760 -1765 2777 -1620
rect 2804 -1765 2821 -1620
rect 2848 -1765 2865 -1620
rect 2892 -1765 2909 -1620
rect 2936 -1765 2953 -1620
rect 2980 -1765 2997 -1620
rect 3029 -1625 3056 -1613
rect 2714 -1773 2735 -1765
rect 2714 -1790 2716 -1773
rect 2733 -1790 2735 -1773
rect 2714 -1798 2735 -1790
rect 2758 -1773 2779 -1765
rect 2758 -1790 2760 -1773
rect 2777 -1790 2779 -1773
rect 2758 -1798 2779 -1790
rect 2802 -1773 2823 -1765
rect 2802 -1790 2804 -1773
rect 2821 -1790 2823 -1773
rect 2802 -1798 2823 -1790
rect 2846 -1773 2867 -1765
rect 2846 -1790 2848 -1773
rect 2865 -1790 2867 -1773
rect 2846 -1798 2867 -1790
rect 2890 -1773 2911 -1765
rect 2890 -1790 2892 -1773
rect 2909 -1790 2911 -1773
rect 2890 -1798 2911 -1790
rect 2934 -1772 2955 -1765
rect 2934 -1790 2936 -1772
rect 2954 -1790 2955 -1772
rect 2934 -1798 2955 -1790
rect 2978 -1773 2999 -1765
rect 2978 -1790 2980 -1773
rect 2997 -1778 2999 -1773
rect 2997 -1790 3137 -1778
rect 2978 -1795 3137 -1790
rect 2978 -1798 2999 -1795
rect 2780 -1831 2805 -1823
rect 2780 -1848 2784 -1831
rect 2801 -1848 2805 -1831
rect 2780 -1857 2805 -1848
rect 2716 -1879 2743 -1866
rect 2716 -1896 2721 -1879
rect 2738 -1896 2743 -1879
rect 2716 -1908 2743 -1896
rect 2892 -1976 2909 -1798
rect 3120 -1976 3137 -1795
rect 2885 -1983 2915 -1976
rect 2885 -2001 2891 -1983
rect 2909 -2001 2915 -1983
rect 2885 -2008 2915 -2001
rect 3113 -1983 3143 -1976
rect 3113 -2001 3119 -1983
rect 3137 -2001 3143 -1983
rect 3113 -2008 3143 -2001
<< viali >>
rect 2804 -1344 2822 -1326
rect 2698 -1500 2715 -1483
rect 2740 -1548 2757 -1531
rect 3035 -1443 3052 -1426
rect 2980 -1503 2997 -1486
rect 2760 -1612 2777 -1595
rect 2680 -1670 2697 -1653
rect 2680 -1726 2697 -1709
rect 2848 -1790 2865 -1773
rect 2936 -1773 2954 -1772
rect 2936 -1790 2953 -1773
rect 2953 -1790 2954 -1773
rect 2784 -1848 2801 -1831
rect 2721 -1896 2738 -1879
rect 2891 -2001 2909 -1983
rect 3119 -2001 3137 -1983
<< metal1 >>
rect 2798 -1322 2828 -1319
rect 2798 -1348 2800 -1322
rect 2826 -1348 2828 -1322
rect 2798 -1351 2828 -1348
rect 3032 -1426 3056 -1423
rect -2201 -1443 3035 -1426
rect 3052 -1443 5603 -1426
rect -2201 -1446 5603 -1443
rect 2695 -1483 2718 -1477
rect 2695 -1486 2698 -1483
rect -2201 -1500 2698 -1486
rect 2715 -1500 2718 -1483
rect 2695 -1506 2718 -1500
rect 2977 -1486 3000 -1480
rect 2977 -1503 2980 -1486
rect 2997 -1500 5603 -1486
rect 2997 -1503 3000 -1500
rect 2977 -1509 3000 -1503
rect 2734 -1531 2763 -1526
rect 2734 -1532 2740 -1531
rect -2201 -1546 2740 -1532
rect 2734 -1548 2740 -1546
rect 2757 -1532 2763 -1531
rect 2757 -1546 5603 -1532
rect 2757 -1548 2763 -1546
rect 2734 -1552 2763 -1548
rect 2636 -1587 2679 -1578
rect 2636 -1613 2641 -1587
rect 2667 -1591 2679 -1587
rect 2757 -1591 2783 -1590
rect 2667 -1595 2783 -1591
rect 2667 -1612 2760 -1595
rect 2777 -1612 2783 -1595
rect 2667 -1613 2783 -1612
rect 2636 -1615 2783 -1613
rect 2639 -1616 2669 -1615
rect 2757 -1616 2783 -1615
rect 2674 -1653 2703 -1649
rect 2674 -1654 2680 -1653
rect -2201 -1668 2680 -1654
rect 2674 -1670 2680 -1668
rect 2697 -1654 2703 -1653
rect 2697 -1668 5603 -1654
rect 2697 -1670 2703 -1668
rect 2674 -1675 2703 -1670
rect 2674 -1709 2703 -1706
rect 2674 -1710 2680 -1709
rect -2201 -1724 2680 -1710
rect 2674 -1726 2680 -1724
rect 2697 -1710 2703 -1709
rect 2697 -1724 5603 -1710
rect 2697 -1726 2703 -1724
rect 2674 -1732 2703 -1726
rect 3172 -1766 3202 -1763
rect 2845 -1771 2871 -1769
rect 2636 -1773 2871 -1771
rect 2636 -1780 2848 -1773
rect 2636 -1806 2641 -1780
rect 2667 -1790 2848 -1780
rect 2865 -1790 2871 -1773
rect 2667 -1792 2871 -1790
rect 2667 -1806 2672 -1792
rect 2845 -1794 2871 -1792
rect 2930 -1771 2959 -1769
rect 3172 -1771 3174 -1766
rect 2930 -1772 3174 -1771
rect 2930 -1790 2936 -1772
rect 2954 -1790 3174 -1772
rect 2930 -1792 3174 -1790
rect 3200 -1771 3202 -1766
rect 3200 -1792 3205 -1771
rect 2930 -1793 2959 -1792
rect 3172 -1795 3202 -1792
rect 2639 -1809 2669 -1806
rect 2778 -1831 2807 -1826
rect 2778 -1832 2784 -1831
rect -2201 -1846 2784 -1832
rect 2778 -1848 2784 -1846
rect 2801 -1832 2807 -1831
rect 2801 -1846 5603 -1832
rect 2801 -1848 2807 -1846
rect 2778 -1852 2807 -1848
rect -2059 -1878 -1892 -1877
rect 2718 -1878 2741 -1876
rect -2201 -1879 5603 -1878
rect -2201 -1895 2721 -1879
rect -2201 -1898 -2005 -1895
rect -2059 -1954 -2005 -1898
rect -1940 -1896 2721 -1895
rect 2738 -1896 5603 -1879
rect -1940 -1898 5603 -1896
rect -1940 -1954 -1892 -1898
rect 2718 -1899 2741 -1898
rect -2059 -1984 -1892 -1954
rect 2885 -1979 2915 -1976
rect 2885 -2005 2887 -1979
rect 2913 -2005 2915 -1979
rect 2885 -2008 2915 -2005
rect 3113 -1979 3143 -1976
rect 3113 -2005 3115 -1979
rect 3141 -2005 3143 -1979
rect 3113 -2008 3143 -2005
<< via1 >>
rect 2800 -1326 2826 -1322
rect 2800 -1344 2804 -1326
rect 2804 -1344 2822 -1326
rect 2822 -1344 2826 -1326
rect 2800 -1348 2826 -1344
rect 2641 -1613 2667 -1587
rect 2641 -1806 2667 -1780
rect 3174 -1792 3200 -1766
rect -2005 -1954 -1940 -1895
rect 2887 -1983 2913 -1979
rect 2887 -2001 2891 -1983
rect 2891 -2001 2909 -1983
rect 2909 -2001 2913 -1983
rect 2887 -2005 2913 -2001
rect 3115 -1983 3141 -1979
rect 3115 -2001 3119 -1983
rect 3119 -2001 3137 -1983
rect 3137 -2001 3141 -1983
rect 3115 -2005 3141 -2001
<< metal2 >>
rect 2795 -1321 2831 -1316
rect 2795 -1349 2799 -1321
rect 2827 -1349 2831 -1321
rect 2795 -1354 2831 -1349
rect 2636 -1586 2672 -1581
rect 2636 -1614 2640 -1586
rect 2668 -1614 2672 -1586
rect 2636 -1619 2672 -1614
rect 3169 -1765 3205 -1760
rect 2636 -1779 2672 -1774
rect 2636 -1807 2640 -1779
rect 2668 -1807 2672 -1779
rect 3169 -1793 3173 -1765
rect 3201 -1793 3205 -1765
rect 3169 -1798 3205 -1793
rect 2636 -1812 2672 -1807
rect -2011 -1895 -1934 -1888
rect -2011 -1954 -2005 -1895
rect -1940 -1954 -1934 -1895
rect -2011 -1961 -1934 -1954
rect 2882 -1978 2918 -1973
rect 2882 -2006 2886 -1978
rect 2914 -2006 2918 -1978
rect 2882 -2011 2918 -2006
rect 3110 -1978 3146 -1973
rect 3110 -2006 3114 -1978
rect 3142 -2006 3146 -1978
rect 3110 -2011 3146 -2006
<< via2 >>
rect 2799 -1322 2827 -1321
rect 2799 -1348 2800 -1322
rect 2800 -1348 2826 -1322
rect 2826 -1348 2827 -1322
rect 2799 -1349 2827 -1348
rect 2640 -1587 2668 -1586
rect 2640 -1613 2641 -1587
rect 2641 -1613 2667 -1587
rect 2667 -1613 2668 -1587
rect 2640 -1614 2668 -1613
rect 2640 -1780 2668 -1779
rect 2640 -1806 2641 -1780
rect 2641 -1806 2667 -1780
rect 2667 -1806 2668 -1780
rect 2640 -1807 2668 -1806
rect 3173 -1766 3201 -1765
rect 3173 -1792 3174 -1766
rect 3174 -1792 3200 -1766
rect 3200 -1792 3201 -1766
rect 3173 -1793 3201 -1792
rect -2005 -1954 -1940 -1895
rect 2886 -1979 2914 -1978
rect 2886 -2005 2887 -1979
rect 2887 -2005 2913 -1979
rect 2913 -2005 2914 -1979
rect 2886 -2006 2914 -2005
rect 3114 -1979 3142 -1978
rect 3114 -2005 3115 -1979
rect 3115 -2005 3141 -1979
rect 3141 -2005 3142 -1979
rect 3114 -2006 3142 -2005
<< metal3 >>
rect -2092 -1250 5604 2862
rect -2059 -1895 -1892 -1250
rect 2057 -1306 2090 -1250
rect 2057 -1734 2585 -1306
rect 2788 -1319 2837 -1309
rect 2788 -1351 2797 -1319
rect 2829 -1351 2837 -1319
rect 2788 -1361 2837 -1351
rect 2630 -1584 2679 -1574
rect 2630 -1616 2638 -1584
rect 2670 -1616 2679 -1584
rect 2630 -1626 2679 -1616
rect 3163 -1763 3212 -1753
rect 2630 -1777 2679 -1767
rect -2059 -1954 -2005 -1895
rect -1940 -1954 -1892 -1895
rect -2059 -2077 -1892 -1954
rect 2057 -2021 2585 -1793
rect 2630 -1809 2638 -1777
rect 2670 -1809 2679 -1777
rect 3163 -1795 3171 -1763
rect 3203 -1795 3212 -1763
rect 3163 -1805 3212 -1795
rect 2630 -1819 2679 -1809
rect 2876 -1976 2925 -1966
rect 2876 -2008 2884 -1976
rect 2916 -2008 2925 -1976
rect 2876 -2018 2925 -2008
rect 3104 -1976 3153 -1966
rect 3104 -2008 3112 -1976
rect 3144 -2008 3153 -1976
rect 3104 -2018 3153 -2008
rect 3243 -2021 3521 -1793
rect 2057 -2077 2090 -2021
rect 3243 -2077 3276 -2021
rect -2093 -2675 3019 -2077
rect 3075 -2675 5604 -2077
rect -2093 -3034 5604 -2675
rect -2093 -5105 3019 -3034
rect 3075 -5105 5604 -3034
<< via3 >>
rect 2797 -1321 2829 -1319
rect 2797 -1349 2799 -1321
rect 2799 -1349 2827 -1321
rect 2827 -1349 2829 -1321
rect 2797 -1351 2829 -1349
rect 2638 -1586 2670 -1584
rect 2638 -1614 2640 -1586
rect 2640 -1614 2668 -1586
rect 2668 -1614 2670 -1586
rect 2638 -1616 2670 -1614
rect -2005 -1954 -1940 -1895
rect 2638 -1779 2670 -1777
rect 2638 -1807 2640 -1779
rect 2640 -1807 2668 -1779
rect 2668 -1807 2670 -1779
rect 2638 -1809 2670 -1807
rect 3171 -1765 3203 -1763
rect 3171 -1793 3173 -1765
rect 3173 -1793 3201 -1765
rect 3201 -1793 3203 -1765
rect 3171 -1795 3203 -1793
rect 2884 -1978 2916 -1976
rect 2884 -2006 2886 -1978
rect 2886 -2006 2914 -1978
rect 2914 -2006 2916 -1978
rect 2884 -2008 2916 -2006
rect 3112 -1978 3144 -1976
rect 3112 -2006 3114 -1978
rect 3114 -2006 3142 -1978
rect 3142 -2006 3144 -1978
rect 3112 -2008 3144 -2006
<< mimcap >>
rect -2078 1187 922 2848
rect -2078 1069 757 1187
rect 875 1069 922 1187
rect -2078 848 922 1069
rect 1006 1184 4006 2848
rect 1006 1066 1059 1184
rect 1177 1161 4006 1184
rect 1177 1066 3847 1161
rect 1006 1043 3847 1066
rect 3965 1043 4006 1161
rect 1006 848 4006 1043
rect 4090 1194 5590 2848
rect 4090 1076 4143 1194
rect 4261 1076 5590 1194
rect 4090 848 5590 1076
rect -2078 540 922 764
rect -2078 422 767 540
rect 885 422 922 540
rect -2078 -1071 922 422
rect -2078 -1189 -1858 -1071
rect -1740 -1189 922 -1071
rect -2078 -1236 922 -1189
rect 1006 547 4006 764
rect 1006 429 1040 547
rect 1158 505 4006 547
rect 1158 429 3825 505
rect 1006 387 3825 429
rect 3943 387 4006 505
rect 1006 -1236 4006 387
rect 4090 488 5590 764
rect 4090 370 4133 488
rect 4251 370 5590 488
rect 4090 -1236 5590 370
rect 2071 -1584 2571 -1320
rect 2071 -1618 2529 -1584
rect 2563 -1618 2571 -1584
rect 2071 -1720 2571 -1618
rect 2071 -1841 2571 -1807
rect 2071 -1875 2527 -1841
rect 2561 -1875 2571 -1841
rect 2071 -2007 2571 -1875
rect 3257 -1828 3507 -1807
rect 3257 -1860 3265 -1828
rect 3297 -1860 3507 -1828
rect 3257 -2007 3507 -1860
rect -2079 -2144 421 -2091
rect -2079 -2262 -1843 -2144
rect -1725 -2262 421 -2144
rect -2079 -5091 421 -2262
rect 505 -2127 3005 -2091
rect 505 -2245 725 -2127
rect 843 -2245 3005 -2127
rect 505 -5091 3005 -2245
rect 3089 -2144 5590 -2091
rect 3089 -2262 3327 -2144
rect 3445 -2262 5590 -2144
rect 3089 -5091 5590 -2262
<< mimcapcontact >>
rect 757 1069 875 1187
rect 1059 1066 1177 1184
rect 3847 1043 3965 1161
rect 4143 1076 4261 1194
rect 767 422 885 540
rect -1858 -1189 -1740 -1071
rect 1040 429 1158 547
rect 3825 387 3943 505
rect 4133 370 4251 488
rect 2529 -1618 2563 -1584
rect 2527 -1875 2561 -1841
rect 3265 -1860 3297 -1828
rect -1843 -2262 -1725 -2144
rect 725 -2245 843 -2127
rect 3327 -2262 3445 -2144
<< metal4 >>
rect -2092 1194 5604 2862
rect -2092 1187 4143 1194
rect -2092 1069 757 1187
rect 875 1184 4143 1187
rect 875 1069 1059 1184
rect -2092 1066 1059 1069
rect 1177 1161 4143 1184
rect 1177 1066 3847 1161
rect -2092 1043 3847 1066
rect 3965 1076 4143 1161
rect 4261 1076 5604 1194
rect 3965 1043 5604 1076
rect -2092 547 5604 1043
rect -2092 540 1040 547
rect -2092 422 767 540
rect 885 429 1040 540
rect 1158 505 5604 547
rect 1158 429 3825 505
rect 885 422 3825 429
rect -2092 387 3825 422
rect 3943 488 5604 505
rect 3943 387 4133 488
rect -2092 370 4133 387
rect 4251 370 5604 488
rect -2092 -1071 5604 370
rect -2092 -1189 -1858 -1071
rect -1740 -1189 5604 -1071
rect -2092 -1250 5604 -1189
rect 2798 -1315 2828 -1250
rect 2796 -1319 2830 -1315
rect 2796 -1351 2797 -1319
rect 2829 -1351 2830 -1319
rect 2796 -1352 2830 -1351
rect 2528 -1584 2671 -1583
rect 2528 -1618 2529 -1584
rect 2563 -1616 2638 -1584
rect 2670 -1616 2671 -1584
rect 2563 -1618 2671 -1616
rect 2528 -1619 2671 -1618
rect 3170 -1763 3204 -1762
rect 2637 -1777 2671 -1776
rect 2637 -1809 2638 -1777
rect 2670 -1809 2671 -1777
rect 3170 -1795 3171 -1763
rect 3203 -1795 3204 -1763
rect 3170 -1799 3204 -1795
rect 2637 -1813 2671 -1809
rect 2526 -1841 2562 -1840
rect 2526 -1875 2527 -1841
rect 2561 -1843 2562 -1841
rect 2639 -1843 2669 -1813
rect 2561 -1873 2669 -1843
rect 3172 -1829 3202 -1799
rect 3262 -1828 3298 -1827
rect 3262 -1829 3265 -1828
rect 3172 -1859 3265 -1829
rect 3262 -1860 3265 -1859
rect 3297 -1860 3298 -1828
rect 3262 -1861 3298 -1860
rect 2561 -1875 2562 -1873
rect 2526 -1876 2562 -1875
rect 2883 -1976 2917 -1975
rect 2883 -2008 2884 -1976
rect 2916 -2008 2917 -1976
rect 2883 -2012 2917 -2008
rect 3111 -1976 3145 -1975
rect 3111 -2008 3112 -1976
rect 3144 -2008 3145 -1976
rect 3111 -2012 3145 -2008
rect 2885 -2077 2915 -2012
rect 3113 -2077 3143 -2012
rect -2093 -2127 3019 -2077
rect -2093 -2144 725 -2127
rect -2093 -2262 -1843 -2144
rect -1725 -2245 725 -2144
rect 843 -2245 3019 -2127
rect -1725 -2262 3019 -2245
rect -2093 -5105 3019 -2262
rect 3075 -2144 5604 -2077
rect 3075 -2262 3327 -2144
rect 3445 -2262 5604 -2144
rect 3075 -5105 5604 -2262
<< via4 >>
rect -2030 -1895 -1908 -1853
rect -2030 -1954 -2005 -1895
rect -2005 -1954 -1940 -1895
rect -1940 -1954 -1908 -1895
rect -2030 -1976 -1908 -1954
<< mimcap2 >>
rect -2078 1003 922 2848
rect -2078 885 763 1003
rect 881 885 922 1003
rect -2078 848 922 885
rect 1006 1005 4006 2848
rect 1006 887 1047 1005
rect 1165 987 4006 1005
rect 1165 887 3833 987
rect 1006 869 3833 887
rect 3951 869 4006 987
rect 1006 848 4006 869
rect 4090 992 5590 2848
rect 4090 874 4124 992
rect 4242 874 5590 992
rect 4090 848 5590 874
rect -2078 726 922 764
rect -2078 608 762 726
rect 880 608 922 726
rect -2078 -1070 922 608
rect -2078 -1188 -2022 -1070
rect -1904 -1188 922 -1070
rect -2078 -1236 922 -1188
rect 1006 729 4006 764
rect 1006 611 1044 729
rect 1162 708 4006 729
rect 1162 611 3830 708
rect 1006 590 3830 611
rect 3948 590 4006 708
rect 1006 -1236 4006 590
rect 4090 706 5590 764
rect 4090 588 4122 706
rect 4240 588 5590 706
rect 4090 -1236 5590 588
rect -2079 -2122 421 -2091
rect -2079 -2240 -2037 -2122
rect -1919 -2145 421 -2122
rect -1919 -2240 241 -2145
rect -2079 -2263 241 -2240
rect 359 -2263 421 -2145
rect -2079 -5091 421 -2263
rect 505 -2133 3005 -2091
rect 505 -2145 2841 -2133
rect 505 -2263 554 -2145
rect 672 -2251 2841 -2145
rect 2959 -2251 3005 -2133
rect 672 -2263 3005 -2251
rect 505 -5091 3005 -2263
rect 3089 -2132 5590 -2091
rect 3089 -2250 3134 -2132
rect 3252 -2250 5590 -2132
rect 3089 -5091 5590 -2250
<< mimcap2contact >>
rect 763 885 881 1003
rect 1047 887 1165 1005
rect 3833 869 3951 987
rect 4124 874 4242 992
rect 762 608 880 726
rect -2022 -1188 -1904 -1070
rect 1044 611 1162 729
rect 3830 590 3948 708
rect 4122 588 4240 706
rect -2037 -2240 -1919 -2122
rect 241 -2263 359 -2145
rect 554 -2263 672 -2145
rect 2841 -2251 2959 -2133
rect 3134 -2250 3252 -2132
<< metal5 >>
rect 730 1005 1188 1029
rect 730 1003 1047 1005
rect 730 885 763 1003
rect 881 887 1047 1003
rect 1165 887 1188 1005
rect 881 885 1188 887
rect 730 729 1188 885
rect 730 726 1044 729
rect 730 608 762 726
rect 880 611 1044 726
rect 1162 611 1188 729
rect 880 608 1188 611
rect 730 592 1188 608
rect 3809 992 4266 1013
rect 3809 987 4124 992
rect 3809 869 3833 987
rect 3951 874 4124 987
rect 4242 874 4266 992
rect 3951 869 4266 874
rect 3809 708 4266 869
rect 3809 590 3830 708
rect 3948 706 4266 708
rect 3948 590 4122 706
rect 3809 588 4122 590
rect 4240 588 4266 706
rect 3809 569 4266 588
rect -2059 -1070 -1892 -1058
rect -2059 -1188 -2022 -1070
rect -1904 -1188 -1892 -1070
rect -2059 -1853 -1892 -1188
rect -2059 -1976 -2030 -1853
rect -1908 -1976 -1892 -1853
rect -2059 -2122 -1892 -1976
rect -2059 -2240 -2037 -2122
rect -1919 -2240 -1892 -2122
rect -2059 -2263 -1892 -2240
rect 218 -2145 700 -2119
rect 218 -2263 241 -2145
rect 359 -2263 554 -2145
rect 672 -2263 700 -2145
rect 218 -2280 700 -2263
rect 2819 -2132 3275 -2104
rect 2819 -2133 3134 -2132
rect 2819 -2251 2841 -2133
rect 2959 -2250 3134 -2133
rect 3252 -2250 3275 -2132
rect 2959 -2251 3275 -2250
rect 2819 -2279 3275 -2251
<< labels >>
rlabel metal1 -2201 -1890 -2201 -1890 7 GND
rlabel metal1 -2201 -1839 -2201 -1839 7 PHI2
rlabel metal1 -2201 -1717 -2201 -1717 7 PHI1
rlabel metal1 -2201 -1662 -2201 -1662 7 PHI2b
rlabel metal1 -2201 -1540 -2201 -1540 7 PHI1b
rlabel metal1 -2201 -1436 -2201 -1436 7 VDD
rlabel metal4 2614 -1619 2614 -1619 5 cs1
rlabel metal4 2639 -1825 2639 -1825 7 cs2
rlabel metal4 3214 -1859 3214 -1859 5 cs3
rlabel locali 2821 -1388 2821 -1388 3 c1
rlabel locali 2909 -1946 2909 -1946 3 c2
rlabel locali 3120 -1946 3120 -1946 7 c3
rlabel metal1 -2201 -1493 -2201 -1493 7 in
rlabel metal1 5603 -1493 5603 -1493 3 out
<< end >>
