magic
tech sky130A
timestamp 1654307754
<< metal3 >>
rect -22 1024 138 1368
rect -34 1023 138 1024
rect 412 1023 572 1368
rect 846 1024 1006 1368
rect 846 1023 1019 1024
rect -34 1011 1019 1023
rect -34 851 1363 1011
rect -34 577 1018 851
rect -34 417 1363 577
rect -34 143 1018 417
rect -34 -17 1363 143
rect -34 -29 1019 -17
rect -34 -30 138 -29
rect -22 -374 138 -30
rect 412 -374 572 -29
rect 846 -30 1019 -29
rect 846 -374 1006 -30
<< mimcap >>
rect -8 893 992 997
rect -8 101 96 893
rect 168 533 456 821
rect 528 533 816 821
rect 168 173 456 461
rect 528 173 816 461
rect 888 101 992 893
rect -8 -3 992 101
<< mimcapcontact >>
rect 96 821 888 893
rect 96 533 168 821
rect 456 533 528 821
rect 816 533 888 821
rect 96 461 888 533
rect 96 173 168 461
rect 456 173 528 461
rect 816 173 888 461
rect 96 101 888 173
<< metal4 >>
rect 18 1011 98 1368
rect 452 1011 532 1368
rect 886 1011 966 1368
rect -22 971 1006 1011
rect -34 893 1363 971
rect -34 891 96 893
rect -22 537 96 891
rect 888 891 1363 893
rect -34 457 96 537
rect 168 533 456 821
rect 528 533 816 821
rect 888 537 1006 891
rect -22 103 96 457
rect 168 173 456 461
rect 528 173 816 461
rect 888 457 1363 537
rect -34 101 96 103
rect 888 103 1006 457
rect 888 101 1363 103
rect -34 23 1363 101
rect -22 -17 1006 23
rect 18 -374 98 -17
rect 452 -374 532 -17
rect 886 -374 966 -17
<< mimcap2 >>
rect -8 906 992 997
rect -8 788 83 906
rect 201 788 258 906
rect 376 788 433 906
rect 551 788 608 906
rect 726 788 783 906
rect 901 788 992 906
rect -8 731 992 788
rect -8 613 83 731
rect 201 613 433 731
rect 551 613 783 731
rect 901 613 992 731
rect -8 556 992 613
rect -8 438 83 556
rect 201 438 258 556
rect 376 438 433 556
rect 551 438 608 556
rect 726 438 783 556
rect 901 438 992 556
rect -8 381 992 438
rect -8 263 83 381
rect 201 263 433 381
rect 551 263 783 381
rect 901 263 992 381
rect -8 206 992 263
rect -8 88 83 206
rect 201 88 258 206
rect 376 88 433 206
rect 551 88 608 206
rect 726 88 783 206
rect 901 88 992 206
rect -8 -3 992 88
<< mimcap2contact >>
rect 83 788 201 906
rect 258 788 376 906
rect 433 788 551 906
rect 608 788 726 906
rect 783 788 901 906
rect 83 613 201 731
rect 433 613 551 731
rect 783 613 901 731
rect 83 438 201 556
rect 258 438 376 556
rect 433 438 551 556
rect 608 438 726 556
rect 783 438 901 556
rect 83 263 201 381
rect 433 263 551 381
rect 783 263 901 381
rect 83 88 201 206
rect 258 88 376 206
rect 433 88 551 206
rect 608 88 726 206
rect 783 88 901 206
<< metal5 >>
rect -22 1024 138 1368
rect -34 1023 138 1024
rect 412 1023 572 1368
rect 846 1024 1006 1368
rect 846 1023 1019 1024
rect -34 1011 1019 1023
rect -34 906 1363 1011
rect -34 788 83 906
rect 201 788 258 906
rect 376 788 433 906
rect 551 788 608 906
rect 726 788 783 906
rect 901 851 1363 906
rect 901 788 1018 851
rect -34 731 1018 788
rect -34 613 83 731
rect 201 613 433 731
rect 551 613 783 731
rect 901 613 1018 731
rect -34 577 1018 613
rect -34 556 1363 577
rect -34 438 83 556
rect 201 438 258 556
rect 376 438 433 556
rect 551 438 608 556
rect 726 438 783 556
rect 901 438 1363 556
rect -34 417 1363 438
rect -34 381 1018 417
rect -34 263 83 381
rect 201 263 433 381
rect 551 263 783 381
rect 901 263 1018 381
rect -34 206 1018 263
rect -34 88 83 206
rect 201 88 258 206
rect 376 88 433 206
rect 551 88 608 206
rect 726 88 783 206
rect 901 143 1018 206
rect 901 88 1363 143
rect -34 -17 1363 88
rect -34 -29 1019 -17
rect -34 -30 138 -29
rect -22 -374 138 -30
rect 412 -374 572 -29
rect 846 -30 1019 -29
rect 846 -374 1006 -30
<< end >>
