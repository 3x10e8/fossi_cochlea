magic
tech TECHNAME
magscale 1 2
timestamp 1650467753
<< nwell >>
rect 272 5540 332 5592
rect 12 5320 72 5388
<< metal1 >>
rect 12 5382 72 5388
rect 12 5326 14 5382
rect 70 5326 72 5382
rect 12 5320 72 5326
rect 20 5100 64 5320
rect 206 2200 208 2262
<< via1 >>
rect 14 5326 70 5382
rect 146 2200 206 2262
<< metal2 >>
rect 264 5602 342 5614
rect 112 5600 342 5602
rect 12 5382 72 5592
rect 112 5542 274 5600
rect 332 5542 342 5600
rect 264 5530 342 5542
rect 12 5326 14 5382
rect 70 5326 72 5382
rect 12 5320 72 5326
rect 2 5042 82 5054
rect 2 4982 12 5042
rect 72 4982 336 5042
rect 2 4970 82 4982
rect 2 2790 82 2804
rect 2 2726 12 2790
rect 72 2726 82 2790
rect 2 2716 82 2726
rect 138 2262 212 2272
rect 138 2200 146 2262
rect 206 2200 212 2262
rect 138 2190 212 2200
rect 22 -161 62 -63
<< via2 >>
rect 274 5542 332 5600
rect 12 4982 72 5042
rect 12 2726 72 2790
rect 146 2200 206 2262
rect 272 2044 332 2114
<< metal3 >>
rect 12 5054 72 5740
rect 2 5042 82 5054
rect 2 4982 12 5042
rect 72 4982 82 5042
rect 2 4970 82 4982
rect 2 2790 82 2804
rect 2 2726 12 2790
rect 72 2726 82 2790
rect 2 2716 82 2726
rect 12 -161 72 2716
rect 142 2272 202 5612
rect 264 5600 342 5614
rect 264 5542 274 5600
rect 332 5542 342 5600
rect 264 5530 342 5542
rect 138 2262 212 2272
rect 138 2200 146 2262
rect 206 2200 212 2262
rect 138 2190 212 2200
rect 272 2124 332 5530
rect 262 2114 342 2124
rect 262 2044 272 2114
rect 332 2044 342 2114
rect 262 2034 342 2044
use level_up_shifter  level_up_shifter_0
timestamp 1650466559
transform 1 0 2 0 1 2674
box -10 -2835 390 0
use level_up_shifter  level_up_shifter_1
timestamp 1650466559
transform 1 0 2 0 1 5592
box -10 -2835 390 0
<< labels >>
rlabel metal3 174 5592 174 5592 1 Bup
rlabel metal2 136 5592 136 5592 1 Bupb
rlabel metal3 54 5592 54 5592 1 Aupb
rlabel metal2 40 5592 40 5592 1 Aup
rlabel metal3 20 -156 20 -156 7 A
rlabel metal2 42 -156 42 -156 7 B
<< end >>
