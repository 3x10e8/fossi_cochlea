magic
tech sky130A
magscale 1 2
timestamp 1647622803
<< error_s >>
rect 1134 364 1150 368
rect 1168 330 1184 334
<< nwell >>
rect 984 416 1056 588
use sky130_fd_sc_lp__buf_0  sky130_fd_sc_lp__buf_0_0 ~/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1626515395
transform 1 0 1082 0 1 43
box -38 -49 326 715
use comp_42_15_single_tail  comp_42_15_single_tail_0
timestamp 1647622143
transform 1 0 546 0 1 424
box -572 -430 536 334
<< end >>
