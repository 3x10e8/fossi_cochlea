magic
tech sky130A
magscale 1 2
timestamp 1654751242
<< obsli1 >>
rect 1104 2159 78844 95761
<< obsm1 >>
rect 1104 2128 78844 95872
<< metal2 >>
rect 1950 97200 2006 98000
rect 5906 97200 5962 98000
rect 9954 97200 10010 98000
rect 13910 97200 13966 98000
rect 17958 97200 18014 98000
rect 21914 97200 21970 98000
rect 25962 97200 26018 98000
rect 29918 97200 29974 98000
rect 33966 97200 34022 98000
rect 37922 97200 37978 98000
rect 41970 97200 42026 98000
rect 45926 97200 45982 98000
rect 49974 97200 50030 98000
rect 53930 97200 53986 98000
rect 57978 97200 58034 98000
rect 61934 97200 61990 98000
rect 65982 97200 66038 98000
rect 69938 97200 69994 98000
rect 73986 97200 74042 98000
rect 77942 97200 77998 98000
rect 4986 0 5042 800
rect 14922 0 14978 800
rect 24950 0 25006 800
rect 34978 0 35034 800
rect 45006 0 45062 800
rect 54942 0 54998 800
rect 64970 0 65026 800
rect 74998 0 75054 800
<< obsm2 >>
rect 1398 97144 1894 97322
rect 2062 97144 5850 97322
rect 6018 97144 9898 97322
rect 10066 97144 13854 97322
rect 14022 97144 17902 97322
rect 18070 97144 21858 97322
rect 22026 97144 25906 97322
rect 26074 97144 29862 97322
rect 30030 97144 33910 97322
rect 34078 97144 37866 97322
rect 38034 97144 41914 97322
rect 42082 97144 45870 97322
rect 46038 97144 49918 97322
rect 50086 97144 53874 97322
rect 54042 97144 57922 97322
rect 58090 97144 61878 97322
rect 62046 97144 65926 97322
rect 66094 97144 69882 97322
rect 70050 97144 73930 97322
rect 74098 97144 77886 97322
rect 78054 97144 78826 97322
rect 1398 856 78826 97144
rect 1398 734 4930 856
rect 5098 734 14866 856
rect 15034 734 24894 856
rect 25062 734 34922 856
rect 35090 734 44950 856
rect 45118 734 54886 856
rect 55054 734 64914 856
rect 65082 734 74942 856
rect 75110 734 78826 856
<< metal3 >>
rect 0 94800 800 94920
rect 79200 94800 80000 94920
rect 0 88680 800 88800
rect 79200 88680 80000 88800
rect 0 82560 800 82680
rect 79200 82560 80000 82680
rect 0 76440 800 76560
rect 79200 76440 80000 76560
rect 0 70320 800 70440
rect 79200 70320 80000 70440
rect 0 64200 800 64320
rect 79200 64200 80000 64320
rect 0 58080 800 58200
rect 79200 58080 80000 58200
rect 0 51960 800 52080
rect 79200 51960 80000 52080
rect 0 45840 800 45960
rect 79200 45840 80000 45960
rect 0 39720 800 39840
rect 79200 39720 80000 39840
rect 0 33600 800 33720
rect 79200 33600 80000 33720
rect 0 27480 800 27600
rect 79200 27480 80000 27600
rect 0 21360 800 21480
rect 79200 21360 80000 21480
rect 0 15240 800 15360
rect 79200 15240 80000 15360
rect 0 9120 800 9240
rect 79200 9120 80000 9240
rect 0 3000 800 3120
rect 79200 3000 80000 3120
<< obsm3 >>
rect 800 95000 79200 96525
rect 880 94720 79120 95000
rect 800 88880 79200 94720
rect 880 88600 79120 88880
rect 800 82760 79200 88600
rect 880 82480 79120 82760
rect 800 76640 79200 82480
rect 880 76360 79120 76640
rect 800 70520 79200 76360
rect 880 70240 79120 70520
rect 800 64400 79200 70240
rect 880 64120 79120 64400
rect 800 58280 79200 64120
rect 880 58000 79120 58280
rect 800 52160 79200 58000
rect 880 51880 79120 52160
rect 800 46040 79200 51880
rect 880 45760 79120 46040
rect 800 39920 79200 45760
rect 880 39640 79120 39920
rect 800 33800 79200 39640
rect 880 33520 79120 33800
rect 800 27680 79200 33520
rect 880 27400 79120 27680
rect 800 21560 79200 27400
rect 880 21280 79120 21560
rect 800 15440 79200 21280
rect 880 15160 79120 15440
rect 800 9320 79200 15160
rect 880 9040 79120 9320
rect 800 3200 79200 9040
rect 880 2920 79120 3200
rect 800 2143 79200 2920
<< metal4 >>
rect 4208 2128 4528 95792
rect 19568 2128 19888 95792
rect 34928 2128 35248 95792
rect 50288 2128 50608 95792
rect 65648 2128 65968 95792
<< obsm4 >>
rect 9443 95872 76117 96525
rect 9443 35531 19488 95872
rect 19968 35531 34848 95872
rect 35328 35531 50208 95872
rect 50688 35531 65568 95872
rect 66048 35531 76117 95872
<< labels >>
rlabel metal3 s 0 33600 800 33720 6 cclk_I[0]
port 1 nsew signal output
rlabel metal3 s 0 76440 800 76560 6 cclk_I[1]
port 2 nsew signal output
rlabel metal3 s 79200 9120 80000 9240 6 cclk_Q[0]
port 3 nsew signal output
rlabel metal3 s 79200 51960 80000 52080 6 cclk_Q[1]
port 4 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 clk_master
port 5 nsew signal input
rlabel metal2 s 5906 97200 5962 98000 6 clk_master_out
port 6 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 clkdiv2_I[0]
port 7 nsew signal output
rlabel metal3 s 0 70320 800 70440 6 clkdiv2_I[1]
port 8 nsew signal output
rlabel metal3 s 79200 15240 80000 15360 6 clkdiv2_Q[0]
port 9 nsew signal output
rlabel metal3 s 79200 58080 80000 58200 6 clkdiv2_Q[1]
port 10 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 comp_high_I[0]
port 11 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 comp_high_I[1]
port 12 nsew signal input
rlabel metal3 s 79200 21360 80000 21480 6 comp_high_Q[0]
port 13 nsew signal input
rlabel metal3 s 79200 64200 80000 64320 6 comp_high_Q[1]
port 14 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 cos_out[0]
port 15 nsew signal output
rlabel metal3 s 0 82560 800 82680 6 cos_out[1]
port 16 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 cos_outb[0]
port 17 nsew signal output
rlabel metal3 s 0 45840 800 45960 6 cos_outb[1]
port 18 nsew signal output
rlabel metal2 s 13910 97200 13966 98000 6 div2out
port 19 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 fb1_I[0]
port 20 nsew signal output
rlabel metal3 s 0 51960 800 52080 6 fb1_I[1]
port 21 nsew signal output
rlabel metal3 s 79200 33600 80000 33720 6 fb1_Q[0]
port 22 nsew signal output
rlabel metal3 s 79200 76440 80000 76560 6 fb1_Q[1]
port 23 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 fb2_I[0]
port 24 nsew signal output
rlabel metal2 s 73986 97200 74042 98000 6 fb2_I[1]
port 25 nsew signal output
rlabel metal2 s 69938 97200 69994 98000 6 fb2_Q[0]
port 26 nsew signal output
rlabel metal2 s 77942 97200 77998 98000 6 fb2_Q[1]
port 27 nsew signal output
rlabel metal2 s 53930 97200 53986 98000 6 gray_clk_out[10]
port 28 nsew signal output
rlabel metal2 s 17958 97200 18014 98000 6 gray_clk_out[1]
port 29 nsew signal output
rlabel metal2 s 21914 97200 21970 98000 6 gray_clk_out[2]
port 30 nsew signal output
rlabel metal2 s 25962 97200 26018 98000 6 gray_clk_out[3]
port 31 nsew signal output
rlabel metal2 s 29918 97200 29974 98000 6 gray_clk_out[4]
port 32 nsew signal output
rlabel metal2 s 33966 97200 34022 98000 6 gray_clk_out[5]
port 33 nsew signal output
rlabel metal2 s 37922 97200 37978 98000 6 gray_clk_out[6]
port 34 nsew signal output
rlabel metal2 s 41970 97200 42026 98000 6 gray_clk_out[7]
port 35 nsew signal output
rlabel metal2 s 45926 97200 45982 98000 6 gray_clk_out[8]
port 36 nsew signal output
rlabel metal2 s 49974 97200 50030 98000 6 gray_clk_out[9]
port 37 nsew signal output
rlabel metal2 s 57978 97200 58034 98000 6 no_ones_below_out[0]
port 38 nsew signal output
rlabel metal2 s 61934 97200 61990 98000 6 no_ones_below_out[1]
port 39 nsew signal output
rlabel metal2 s 65982 97200 66038 98000 6 no_ones_below_out[2]
port 40 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 phi1b_dig_I[0]
port 41 nsew signal input
rlabel metal3 s 0 58080 800 58200 6 phi1b_dig_I[1]
port 42 nsew signal input
rlabel metal3 s 79200 27480 80000 27600 6 phi1b_dig_Q[0]
port 43 nsew signal input
rlabel metal3 s 79200 70320 80000 70440 6 phi1b_dig_Q[1]
port 44 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 read_out_I[0]
port 45 nsew signal output
rlabel metal2 s 14922 0 14978 800 6 read_out_I[1]
port 46 nsew signal output
rlabel metal3 s 0 88680 800 88800 6 read_out_I_top[0]
port 47 nsew signal output
rlabel metal3 s 0 94800 800 94920 6 read_out_I_top[1]
port 48 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 read_out_Q[0]
port 49 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 read_out_Q[1]
port 50 nsew signal output
rlabel metal3 s 79200 88680 80000 88800 6 read_out_Q_top[0]
port 51 nsew signal output
rlabel metal3 s 79200 94800 80000 94920 6 read_out_Q_top[1]
port 52 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 rstb
port 53 nsew signal input
rlabel metal2 s 1950 97200 2006 98000 6 rstb_out
port 54 nsew signal output
rlabel metal3 s 79200 3000 80000 3120 6 sin_out[0]
port 55 nsew signal output
rlabel metal3 s 79200 45840 80000 45960 6 sin_out[1]
port 56 nsew signal output
rlabel metal3 s 79200 39720 80000 39840 6 sin_outb[0]
port 57 nsew signal output
rlabel metal3 s 79200 82560 80000 82680 6 sin_outb[1]
port 58 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 ud_en
port 59 nsew signal input
rlabel metal2 s 9954 97200 10010 98000 6 ud_en_out
port 60 nsew signal output
rlabel metal4 s 4208 2128 4528 95792 6 vccd1
port 61 nsew power input
rlabel metal4 s 34928 2128 35248 95792 6 vccd1
port 61 nsew power input
rlabel metal4 s 65648 2128 65968 95792 6 vccd1
port 61 nsew power input
rlabel metal4 s 19568 2128 19888 95792 6 vssd1
port 62 nsew ground input
rlabel metal4 s 50288 2128 50608 95792 6 vssd1
port 62 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 80000 98000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8568854
string GDS_FILE /Volumes/export/isn/abhinav/fossi_cochlea/openlane/first_dual_core/runs/first_dual_core/results/finishing/first_dual_core.magic.gds
string GDS_START 446370
<< end >>

