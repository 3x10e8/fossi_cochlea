* NGSPICE file created from cap_12pF.ext - technology: sky130B

.subckt cap_10_10_edge_x2 m3_n712_n702# c1_n16_n6#
X0 m3_n712_n702# c1_n16_n6# sky130_fd_pr__cap_mim_m3_2 l=1e+07u w=1e+07u
X1 c1_n16_n6# m3_n712_n702# sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
.ends

.subckt cap_10_10_x2 c2_n16_n6# m3_n376_n34# c1_n16_n6#
X0 c2_n16_n6# c1_n16_n6# sky130_fd_pr__cap_mim_m3_2 l=1e+07u w=1e+07u
X1 c1_n16_n6# m3_n376_n34# sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
.ends

.subckt cap_10_10__side_x2 m3_n712_n366# c1_n16_n6#
X0 m3_n712_n366# c1_n16_n6# sky130_fd_pr__cap_mim_m3_2 l=1e+07u w=1e+07u
X1 c1_n16_n6# m3_n712_n366# sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
.ends

.subckt cap_12pF sig vss
Xcap_10_10_edge_x2_1 vss sig cap_10_10_edge_x2
Xcap_10_10_edge_x2_0 vss sig cap_10_10_edge_x2
Xcap_10_10_edge_x2_2 vss sig cap_10_10_edge_x2
Xcap_10_10_x2_0[0|0] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[1|0] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[0|1] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[1|1] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[0|2] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[1|2] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[0|3] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[1|3] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[0|4] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[1|4] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[0|5] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[1|5] vss vss sig cap_10_10_x2
Xcap_10_10_edge_x2_3 vss sig cap_10_10_edge_x2
Xcap_10_10__side_x2_0[0] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_0[1] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_0[2] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_0[3] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_0[4] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_0[5] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[0] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[1] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[2] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[3] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[4] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[5] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_2 vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_3 vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_5 vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_4 vss sig cap_10_10__side_x2
.ends

