magic
tech sky130A
magscale 1 2
timestamp 1647845704
<< nwell >>
rect -512 -6 518 164
<< pmos >>
rect -418 34 -388 118
rect -330 34 -300 118
rect 0 34 30 118
rect 88 34 118 118
rect 176 34 206 118
rect 264 34 294 118
<< nmoslvt >>
rect -430 -266 -400 -182
rect -324 -266 -294 -182
rect -104 -266 -74 -182
rect 0 -266 30 -182
rect 88 -266 118 -182
rect 176 -266 206 -182
rect 264 -266 294 -182
<< ndiff >>
rect -504 -204 -430 -182
rect -504 -238 -496 -204
rect -462 -238 -430 -204
rect -504 -266 -430 -238
rect -400 -204 -324 -182
rect -400 -238 -378 -204
rect -344 -238 -324 -204
rect -400 -266 -324 -238
rect -294 -204 -220 -182
rect -294 -238 -262 -204
rect -228 -238 -220 -204
rect -294 -266 -220 -238
rect -158 -204 -104 -182
rect -158 -238 -150 -204
rect -116 -238 -104 -204
rect -158 -266 -104 -238
rect -74 -216 0 -182
rect -74 -250 -60 -216
rect -26 -250 0 -216
rect -74 -266 0 -250
rect 30 -204 88 -182
rect 30 -238 42 -204
rect 76 -238 88 -204
rect 30 -266 88 -238
rect 118 -204 176 -182
rect 118 -238 130 -204
rect 164 -238 176 -204
rect 118 -266 176 -238
rect 206 -204 264 -182
rect 206 -238 218 -204
rect 252 -238 264 -204
rect 206 -266 264 -238
rect 294 -204 354 -182
rect 294 -238 306 -204
rect 340 -238 354 -204
rect 294 -266 354 -238
<< pdiff >>
rect -476 96 -418 118
rect -476 62 -464 96
rect -430 62 -418 96
rect -476 34 -418 62
rect -388 96 -330 118
rect -388 62 -376 96
rect -342 62 -330 96
rect -388 34 -330 62
rect -300 96 -246 118
rect -300 62 -288 96
rect -254 62 -246 96
rect -300 34 -246 62
rect -54 96 0 118
rect -54 62 -46 96
rect -12 62 0 96
rect -54 34 0 62
rect 30 96 88 118
rect 30 62 42 96
rect 76 62 88 96
rect 30 34 88 62
rect 118 96 176 118
rect 118 62 130 96
rect 164 62 176 96
rect 118 34 176 62
rect 206 96 264 118
rect 206 62 218 96
rect 252 62 264 96
rect 206 34 264 62
rect 294 96 354 118
rect 294 62 306 96
rect 340 62 354 96
rect 294 34 354 62
<< ndiffc >>
rect -496 -238 -462 -204
rect -378 -238 -344 -204
rect -262 -238 -228 -204
rect -150 -238 -116 -204
rect -60 -250 -26 -216
rect 42 -238 76 -204
rect 130 -238 164 -204
rect 218 -238 252 -204
rect 306 -238 340 -204
<< pdiffc >>
rect -464 62 -430 96
rect -376 62 -342 96
rect -288 62 -254 96
rect -46 62 -12 96
rect 42 62 76 96
rect 130 62 164 96
rect 218 62 252 96
rect 306 62 340 96
<< psubdiff >>
rect 354 -206 416 -182
rect 354 -240 382 -206
rect 354 -266 416 -240
<< nsubdiff >>
rect 354 92 416 118
rect 354 58 382 92
rect 354 34 416 58
<< psubdiffcont >>
rect 382 -240 416 -206
<< nsubdiffcont >>
rect 382 58 416 92
<< poly >>
rect 150 230 216 246
rect 150 196 166 230
rect 200 226 216 230
rect 200 196 294 226
rect 150 186 216 196
rect -418 118 -388 144
rect -330 118 -300 144
rect 0 118 30 144
rect 88 118 118 144
rect 176 118 206 144
rect 264 118 294 196
rect -154 84 -70 100
rect -154 50 -144 84
rect -110 50 -70 84
rect -154 34 -70 50
rect -418 14 -388 34
rect -330 14 -300 34
rect -418 -16 -204 14
rect -100 12 -70 34
rect 0 12 30 34
rect -246 -26 -172 -16
rect -100 -18 30 12
rect -246 -30 -170 -26
rect -236 -46 -170 -30
rect -204 -60 -170 -46
rect -204 -70 -100 -60
rect -446 -90 -382 -72
rect -446 -124 -432 -90
rect -398 -124 -382 -90
rect -446 -140 -382 -124
rect -340 -90 -278 -72
rect -340 -124 -326 -90
rect -292 -124 -278 -90
rect -340 -140 -278 -124
rect -204 -104 -152 -70
rect -118 -104 -100 -70
rect 88 -78 118 34
rect 176 2 206 34
rect 264 8 294 34
rect 168 -14 222 2
rect 168 -48 178 -14
rect 212 -48 222 -14
rect 168 -64 222 -48
rect -204 -114 -100 -104
rect 72 -84 118 -78
rect 72 -100 126 -84
rect -430 -182 -400 -140
rect -324 -182 -294 -140
rect -430 -292 -400 -266
rect -324 -292 -294 -266
rect -204 -282 -174 -114
rect 72 -134 82 -100
rect 116 -134 126 -100
rect 72 -150 126 -134
rect -104 -182 -74 -156
rect 0 -182 30 -156
rect 88 -182 118 -150
rect 176 -182 206 -64
rect 304 -94 358 -78
rect 304 -114 314 -94
rect 264 -128 314 -114
rect 348 -128 358 -94
rect 264 -144 358 -128
rect 264 -182 294 -144
rect -104 -282 -74 -266
rect -204 -312 -74 -282
rect 0 -334 30 -266
rect 88 -292 118 -266
rect 176 -292 206 -266
rect 264 -334 294 -266
rect 0 -364 294 -334
<< polycont >>
rect 166 196 200 230
rect -144 50 -110 84
rect -432 -124 -398 -90
rect -326 -124 -292 -90
rect -152 -104 -118 -70
rect 178 -48 212 -14
rect 82 -134 116 -100
rect 314 -128 348 -94
<< locali >>
rect -572 268 -510 302
rect -476 268 -414 302
rect -380 268 -318 302
rect -284 268 -222 302
rect -188 268 -126 302
rect -92 268 -30 302
rect 4 268 66 302
rect 100 268 162 302
rect 196 268 258 302
rect 292 268 354 302
rect 388 268 450 302
rect 484 268 546 302
rect -376 112 -342 268
rect -280 230 216 234
rect -280 200 166 230
rect -280 112 -246 200
rect 150 196 166 200
rect 200 196 216 230
rect 150 180 216 196
rect -504 96 -422 112
rect -504 62 -464 96
rect -430 62 -422 96
rect -504 46 -422 62
rect -384 96 -334 112
rect -384 62 -376 96
rect -342 62 -334 96
rect -384 46 -334 62
rect -296 110 -246 112
rect -296 96 -218 110
rect -296 62 -288 96
rect -254 62 -218 96
rect -296 46 -218 62
rect -504 -188 -470 46
rect -432 -90 -398 -72
rect -432 -140 -398 -124
rect -326 -90 -292 -72
rect -326 -140 -292 -124
rect -252 -188 -218 46
rect -150 84 -104 100
rect -150 50 -144 84
rect -110 50 -104 84
rect -150 34 -104 50
rect -54 96 -4 112
rect -54 62 -46 96
rect -12 62 -4 96
rect -54 46 -4 62
rect 34 96 84 112
rect 34 62 42 96
rect 76 62 84 96
rect 34 46 84 62
rect 122 96 176 112
rect 122 62 130 96
rect 164 62 176 96
rect 122 46 176 62
rect 210 96 260 112
rect 210 62 218 96
rect 252 62 260 96
rect 210 46 260 62
rect 298 96 348 112
rect 298 62 306 96
rect 340 62 348 96
rect 298 46 348 62
rect 382 92 416 268
rect -54 -14 -20 46
rect 178 -14 212 2
rect 306 -4 340 46
rect 382 42 416 58
rect -54 -48 178 -14
rect -168 -104 -152 -70
rect -118 -104 -102 -70
rect 14 -188 48 -48
rect 178 -64 212 -48
rect 246 -38 340 -4
rect 82 -100 116 -84
rect 246 -100 280 -38
rect 116 -134 280 -100
rect 82 -150 116 -134
rect 220 -148 280 -134
rect 314 -94 348 -78
rect 314 -144 348 -128
rect 220 -188 254 -148
rect -504 -204 -454 -188
rect -504 -238 -496 -204
rect -462 -238 -454 -204
rect -504 -254 -454 -238
rect -386 -204 -336 -188
rect -386 -238 -378 -204
rect -344 -238 -336 -204
rect -386 -254 -336 -238
rect -270 -204 -218 -188
rect -270 -238 -262 -204
rect -228 -222 -218 -204
rect -156 -204 -108 -188
rect -228 -238 -220 -222
rect -270 -254 -220 -238
rect -156 -238 -150 -204
rect -116 -238 -108 -204
rect -156 -254 -108 -238
rect -66 -216 -20 -200
rect -66 -250 -60 -216
rect -26 -250 -20 -216
rect 14 -204 84 -188
rect 14 -222 42 -204
rect -380 -290 -346 -254
rect -156 -290 -122 -254
rect -66 -266 -20 -250
rect 34 -238 42 -222
rect 76 -238 84 -204
rect 34 -254 84 -238
rect 122 -204 172 -188
rect 122 -238 130 -204
rect 164 -238 172 -204
rect 122 -254 172 -238
rect 210 -204 260 -188
rect 210 -238 218 -204
rect 252 -238 260 -204
rect 210 -254 260 -238
rect 298 -204 348 -188
rect 298 -238 306 -204
rect 340 -238 348 -204
rect 298 -254 348 -238
rect 382 -206 416 -188
rect -380 -324 -122 -290
rect -54 -364 -20 -266
rect 132 -364 166 -254
rect 308 -364 342 -254
rect 382 -364 416 -240
rect -572 -398 -510 -364
rect -476 -398 -414 -364
rect -380 -398 -318 -364
rect -284 -398 -222 -364
rect -188 -398 -126 -364
rect -92 -398 -30 -364
rect 4 -398 66 -364
rect 100 -398 162 -364
rect 196 -398 258 -364
rect 292 -398 354 -364
rect 388 -398 450 -364
rect 484 -398 546 -364
<< viali >>
rect -510 268 -476 302
rect -414 268 -380 302
rect -318 268 -284 302
rect -222 268 -188 302
rect -126 268 -92 302
rect -30 268 4 302
rect 66 268 100 302
rect 162 268 196 302
rect 258 268 292 302
rect 354 268 388 302
rect 450 268 484 302
rect -464 62 -430 96
rect -144 50 -110 84
rect 130 62 164 96
rect -510 -398 -476 -364
rect -414 -398 -380 -364
rect -318 -398 -284 -364
rect -222 -398 -188 -364
rect -126 -398 -92 -364
rect -30 -398 4 -364
rect 66 -398 100 -364
rect 162 -398 196 -364
rect 258 -398 292 -364
rect 354 -398 388 -364
rect 450 -398 484 -364
<< metal1 >>
rect -572 302 546 334
rect -572 268 -510 302
rect -476 268 -414 302
rect -380 268 -318 302
rect -284 268 -222 302
rect -188 268 -126 302
rect -92 268 -30 302
rect 4 268 66 302
rect 100 268 162 302
rect 196 268 258 302
rect 292 268 354 302
rect 388 268 450 302
rect 484 268 546 302
rect -572 236 546 268
rect -476 98 -422 104
rect 130 102 164 236
rect -476 96 -104 98
rect -476 62 -464 96
rect -430 84 -104 96
rect -430 62 -144 84
rect -476 60 -144 62
rect -476 54 -422 60
rect -150 50 -144 60
rect -110 50 -104 84
rect 124 96 170 102
rect 124 62 130 96
rect 164 62 170 96
rect 124 50 170 62
rect -150 36 -104 50
rect -572 -364 546 -332
rect -572 -398 -510 -364
rect -476 -398 -414 -364
rect -380 -398 -318 -364
rect -284 -398 -222 -364
rect -188 -398 -126 -364
rect -92 -398 -30 -364
rect 4 -398 66 -364
rect 100 -398 162 -364
rect 196 -398 258 -364
rect 292 -398 354 -364
rect 388 -398 450 -364
rect 484 -398 546 -364
rect -572 -430 546 -398
use sky130_fd_sc_lp__dfxtp_lp  sky130_fd_sc_lp__dfxtp_lp_0 ~/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1626515395
transform 1 0 546 0 1 -381
box -38 -49 2246 715
<< labels >>
flabel polycont 178 -48 212 -14 0 FreeSans 112 0 0 0 high
flabel polycont 82 -134 116 -100 0 FreeSans 112 0 0 0 low
flabel polycont 314 -128 348 -94 0 FreeSans 112 0 0 0 phi1b
flabel polycont -152 -104 -118 -70 0 FreeSans 112 0 0 0 phi1
rlabel locali -102 -88 -102 -88 3 phi1
rlabel locali 236 112 236 112 1 pfete
rlabel locali 60 112 60 112 1 pfetw
rlabel locali 236 -188 236 -188 1 low
rlabel locali 60 -188 60 -188 1 high
rlabel locali 330 -78 330 -78 1 phi1b
rlabel locali -208 -290 -208 -290 1 tail
rlabel locali -310 -74 -310 -74 1 inm
flabel polycont -326 -124 -292 -90 0 FreeSans 112 0 0 0 inm
flabel polycont -432 -124 -398 -90 0 FreeSans 112 0 0 0 inp
rlabel locali -414 -72 -414 -72 1 inp
rlabel locali -470 -40 -470 -40 3 FP
rlabel locali -252 -46 -252 -46 7 FN
rlabel locali 546 288 546 288 3 VDD
rlabel locali 546 -382 546 -382 3 GND
<< end >>
