VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital_unison
  CLASS BLOCK ;
  FOREIGN digital_unison ;
  ORIGIN 0.000 0.000 ;
  SIZE 1920.000 BY 120.000 ;
  PIN cclk_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 116.000 148.950 120.000 ;
    END
  END cclk_I[0]
  PIN cclk_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 116.000 386.310 120.000 ;
    END
  END cclk_I[1]
  PIN cclk_I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 116.000 623.670 120.000 ;
    END
  END cclk_I[2]
  PIN cclk_I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.750 116.000 861.030 120.000 ;
    END
  END cclk_I[3]
  PIN cclk_I[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 116.000 1098.390 120.000 ;
    END
  END cclk_I[4]
  PIN cclk_I[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.470 116.000 1335.750 120.000 ;
    END
  END cclk_I[5]
  PIN cclk_I[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.830 116.000 1573.110 120.000 ;
    END
  END cclk_I[6]
  PIN cclk_I[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.190 116.000 1810.470 120.000 ;
    END
  END cclk_I[7]
  PIN cclk_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END cclk_Q[0]
  PIN cclk_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END cclk_Q[1]
  PIN cclk_Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 0.000 623.670 4.000 ;
    END
  END cclk_Q[2]
  PIN cclk_Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.750 0.000 861.030 4.000 ;
    END
  END cclk_Q[3]
  PIN cclk_Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END cclk_Q[4]
  PIN cclk_Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.470 0.000 1335.750 4.000 ;
    END
  END cclk_Q[5]
  PIN cclk_Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.830 0.000 1573.110 4.000 ;
    END
  END cclk_Q[6]
  PIN cclk_Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.190 0.000 1810.470 4.000 ;
    END
  END cclk_Q[7]
  PIN clk_master
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END clk_master
  PIN clkdiv2_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 116.000 109.390 120.000 ;
    END
  END clkdiv2_I[0]
  PIN clkdiv2_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 116.000 346.750 120.000 ;
    END
  END clkdiv2_I[1]
  PIN clkdiv2_I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 116.000 584.110 120.000 ;
    END
  END clkdiv2_I[2]
  PIN clkdiv2_I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 116.000 821.470 120.000 ;
    END
  END clkdiv2_I[3]
  PIN clkdiv2_I[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.550 116.000 1058.830 120.000 ;
    END
  END clkdiv2_I[4]
  PIN clkdiv2_I[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1295.910 116.000 1296.190 120.000 ;
    END
  END clkdiv2_I[5]
  PIN clkdiv2_I[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.270 116.000 1533.550 120.000 ;
    END
  END clkdiv2_I[6]
  PIN clkdiv2_I[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.630 116.000 1770.910 120.000 ;
    END
  END clkdiv2_I[7]
  PIN clkdiv2_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END clkdiv2_Q[0]
  PIN clkdiv2_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END clkdiv2_Q[1]
  PIN clkdiv2_Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 0.000 584.110 4.000 ;
    END
  END clkdiv2_Q[2]
  PIN clkdiv2_Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 0.000 821.470 4.000 ;
    END
  END clkdiv2_Q[3]
  PIN clkdiv2_Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.550 0.000 1058.830 4.000 ;
    END
  END clkdiv2_Q[4]
  PIN clkdiv2_Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1295.910 0.000 1296.190 4.000 ;
    END
  END clkdiv2_Q[5]
  PIN clkdiv2_Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.270 0.000 1533.550 4.000 ;
    END
  END clkdiv2_Q[6]
  PIN clkdiv2_Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.630 0.000 1770.910 4.000 ;
    END
  END clkdiv2_Q[7]
  PIN comp_high_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 116.000 228.070 120.000 ;
    END
  END comp_high_I[0]
  PIN comp_high_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 116.000 465.430 120.000 ;
    END
  END comp_high_I[1]
  PIN comp_high_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 116.000 702.790 120.000 ;
    END
  END comp_high_I[2]
  PIN comp_high_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.870 116.000 940.150 120.000 ;
    END
  END comp_high_I[3]
  PIN comp_high_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.230 116.000 1177.510 120.000 ;
    END
  END comp_high_I[4]
  PIN comp_high_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.590 116.000 1414.870 120.000 ;
    END
  END comp_high_I[5]
  PIN comp_high_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.950 116.000 1652.230 120.000 ;
    END
  END comp_high_I[6]
  PIN comp_high_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1889.310 116.000 1889.590 120.000 ;
    END
  END comp_high_I[7]
  PIN comp_high_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END comp_high_Q[0]
  PIN comp_high_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 0.000 465.430 4.000 ;
    END
  END comp_high_Q[1]
  PIN comp_high_Q[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END comp_high_Q[2]
  PIN comp_high_Q[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.870 0.000 940.150 4.000 ;
    END
  END comp_high_Q[3]
  PIN comp_high_Q[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.230 0.000 1177.510 4.000 ;
    END
  END comp_high_Q[4]
  PIN comp_high_Q[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.590 0.000 1414.870 4.000 ;
    END
  END comp_high_Q[5]
  PIN comp_high_Q[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.950 0.000 1652.230 4.000 ;
    END
  END comp_high_Q[6]
  PIN comp_high_Q[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1889.310 0.000 1889.590 4.000 ;
    END
  END comp_high_Q[7]
  PIN cos_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 116.000 30.270 120.000 ;
    END
  END cos_out[0]
  PIN cos_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 116.000 267.630 120.000 ;
    END
  END cos_out[1]
  PIN cos_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 116.000 504.990 120.000 ;
    END
  END cos_out[2]
  PIN cos_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 116.000 742.350 120.000 ;
    END
  END cos_out[3]
  PIN cos_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.430 116.000 979.710 120.000 ;
    END
  END cos_out[4]
  PIN cos_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.790 116.000 1217.070 120.000 ;
    END
  END cos_out[5]
  PIN cos_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.150 116.000 1454.430 120.000 ;
    END
  END cos_out[6]
  PIN cos_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.510 116.000 1691.790 120.000 ;
    END
  END cos_out[7]
  PIN fb1_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 116.000 69.830 120.000 ;
    END
  END fb1_I[0]
  PIN fb1_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 116.000 307.190 120.000 ;
    END
  END fb1_I[1]
  PIN fb1_I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 116.000 544.550 120.000 ;
    END
  END fb1_I[2]
  PIN fb1_I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.630 116.000 781.910 120.000 ;
    END
  END fb1_I[3]
  PIN fb1_I[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.990 116.000 1019.270 120.000 ;
    END
  END fb1_I[4]
  PIN fb1_I[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.350 116.000 1256.630 120.000 ;
    END
  END fb1_I[5]
  PIN fb1_I[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1493.710 116.000 1493.990 120.000 ;
    END
  END fb1_I[6]
  PIN fb1_I[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1731.070 116.000 1731.350 120.000 ;
    END
  END fb1_I[7]
  PIN fb1_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END fb1_Q[0]
  PIN fb1_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END fb1_Q[1]
  PIN fb1_Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END fb1_Q[2]
  PIN fb1_Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.630 0.000 781.910 4.000 ;
    END
  END fb1_Q[3]
  PIN fb1_Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.990 0.000 1019.270 4.000 ;
    END
  END fb1_Q[4]
  PIN fb1_Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.350 0.000 1256.630 4.000 ;
    END
  END fb1_Q[5]
  PIN fb1_Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1493.710 0.000 1493.990 4.000 ;
    END
  END fb1_Q[6]
  PIN fb1_Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1731.070 0.000 1731.350 4.000 ;
    END
  END fb1_Q[7]
  PIN phi1b_dig_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 116.000 188.510 120.000 ;
    END
  END phi1b_dig_I[0]
  PIN phi1b_dig_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 116.000 425.870 120.000 ;
    END
  END phi1b_dig_I[1]
  PIN phi1b_dig_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.950 116.000 663.230 120.000 ;
    END
  END phi1b_dig_I[2]
  PIN phi1b_dig_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.310 116.000 900.590 120.000 ;
    END
  END phi1b_dig_I[3]
  PIN phi1b_dig_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.670 116.000 1137.950 120.000 ;
    END
  END phi1b_dig_I[4]
  PIN phi1b_dig_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 116.000 1375.310 120.000 ;
    END
  END phi1b_dig_I[5]
  PIN phi1b_dig_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.390 116.000 1612.670 120.000 ;
    END
  END phi1b_dig_I[6]
  PIN phi1b_dig_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1849.750 116.000 1850.030 120.000 ;
    END
  END phi1b_dig_I[7]
  PIN phi1b_dig_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END phi1b_dig_Q[0]
  PIN phi1b_dig_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END phi1b_dig_Q[1]
  PIN phi1b_dig_Q[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.950 0.000 663.230 4.000 ;
    END
  END phi1b_dig_Q[2]
  PIN phi1b_dig_Q[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.310 0.000 900.590 4.000 ;
    END
  END phi1b_dig_Q[3]
  PIN phi1b_dig_Q[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.670 0.000 1137.950 4.000 ;
    END
  END phi1b_dig_Q[4]
  PIN phi1b_dig_Q[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 0.000 1375.310 4.000 ;
    END
  END phi1b_dig_Q[5]
  PIN phi1b_dig_Q[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.390 0.000 1612.670 4.000 ;
    END
  END phi1b_dig_Q[6]
  PIN phi1b_dig_Q[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1849.750 0.000 1850.030 4.000 ;
    END
  END phi1b_dig_Q[7]
  PIN read_out_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1916.000 104.080 1920.000 104.680 ;
    END
  END read_out_I[0]
  PIN read_out_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1916.000 74.160 1920.000 74.760 ;
    END
  END read_out_I[1]
  PIN read_out_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1916.000 44.240 1920.000 44.840 ;
    END
  END read_out_Q[0]
  PIN read_out_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1916.000 14.320 1920.000 14.920 ;
    END
  END read_out_Q[1]
  PIN rstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END rstb
  PIN sin_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END sin_out[0]
  PIN sin_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END sin_out[1]
  PIN sin_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 0.000 504.990 4.000 ;
    END
  END sin_out[2]
  PIN sin_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 0.000 742.350 4.000 ;
    END
  END sin_out[3]
  PIN sin_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.430 0.000 979.710 4.000 ;
    END
  END sin_out[4]
  PIN sin_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.790 0.000 1217.070 4.000 ;
    END
  END sin_out[5]
  PIN sin_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.150 0.000 1454.430 4.000 ;
    END
  END sin_out[6]
  PIN sin_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.510 0.000 1691.790 4.000 ;
    END
  END sin_out[7]
  PIN ud_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END ud_en
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 243.285 10.640 244.885 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 720.420 10.640 722.020 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.555 10.640 1199.155 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1674.690 10.640 1676.290 109.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 481.850 10.640 483.450 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 958.985 10.640 960.585 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1436.120 10.640 1437.720 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1913.255 10.640 1914.855 109.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1914.060 108.885 ;
      LAYER met1 ;
        RECT 5.520 4.460 1914.855 109.780 ;
      LAYER met2 ;
        RECT 7.910 115.720 29.710 116.690 ;
        RECT 30.550 115.720 69.270 116.690 ;
        RECT 70.110 115.720 108.830 116.690 ;
        RECT 109.670 115.720 148.390 116.690 ;
        RECT 149.230 115.720 187.950 116.690 ;
        RECT 188.790 115.720 227.510 116.690 ;
        RECT 228.350 115.720 267.070 116.690 ;
        RECT 267.910 115.720 306.630 116.690 ;
        RECT 307.470 115.720 346.190 116.690 ;
        RECT 347.030 115.720 385.750 116.690 ;
        RECT 386.590 115.720 425.310 116.690 ;
        RECT 426.150 115.720 464.870 116.690 ;
        RECT 465.710 115.720 504.430 116.690 ;
        RECT 505.270 115.720 543.990 116.690 ;
        RECT 544.830 115.720 583.550 116.690 ;
        RECT 584.390 115.720 623.110 116.690 ;
        RECT 623.950 115.720 662.670 116.690 ;
        RECT 663.510 115.720 702.230 116.690 ;
        RECT 703.070 115.720 741.790 116.690 ;
        RECT 742.630 115.720 781.350 116.690 ;
        RECT 782.190 115.720 820.910 116.690 ;
        RECT 821.750 115.720 860.470 116.690 ;
        RECT 861.310 115.720 900.030 116.690 ;
        RECT 900.870 115.720 939.590 116.690 ;
        RECT 940.430 115.720 979.150 116.690 ;
        RECT 979.990 115.720 1018.710 116.690 ;
        RECT 1019.550 115.720 1058.270 116.690 ;
        RECT 1059.110 115.720 1097.830 116.690 ;
        RECT 1098.670 115.720 1137.390 116.690 ;
        RECT 1138.230 115.720 1176.950 116.690 ;
        RECT 1177.790 115.720 1216.510 116.690 ;
        RECT 1217.350 115.720 1256.070 116.690 ;
        RECT 1256.910 115.720 1295.630 116.690 ;
        RECT 1296.470 115.720 1335.190 116.690 ;
        RECT 1336.030 115.720 1374.750 116.690 ;
        RECT 1375.590 115.720 1414.310 116.690 ;
        RECT 1415.150 115.720 1453.870 116.690 ;
        RECT 1454.710 115.720 1493.430 116.690 ;
        RECT 1494.270 115.720 1532.990 116.690 ;
        RECT 1533.830 115.720 1572.550 116.690 ;
        RECT 1573.390 115.720 1612.110 116.690 ;
        RECT 1612.950 115.720 1651.670 116.690 ;
        RECT 1652.510 115.720 1691.230 116.690 ;
        RECT 1692.070 115.720 1730.790 116.690 ;
        RECT 1731.630 115.720 1770.350 116.690 ;
        RECT 1771.190 115.720 1809.910 116.690 ;
        RECT 1810.750 115.720 1849.470 116.690 ;
        RECT 1850.310 115.720 1889.030 116.690 ;
        RECT 1889.870 115.720 1914.825 116.690 ;
        RECT 7.910 4.280 1914.825 115.720 ;
        RECT 7.910 3.670 29.710 4.280 ;
        RECT 30.550 3.670 69.270 4.280 ;
        RECT 70.110 3.670 108.830 4.280 ;
        RECT 109.670 3.670 148.390 4.280 ;
        RECT 149.230 3.670 187.950 4.280 ;
        RECT 188.790 3.670 227.510 4.280 ;
        RECT 228.350 3.670 267.070 4.280 ;
        RECT 267.910 3.670 306.630 4.280 ;
        RECT 307.470 3.670 346.190 4.280 ;
        RECT 347.030 3.670 385.750 4.280 ;
        RECT 386.590 3.670 425.310 4.280 ;
        RECT 426.150 3.670 464.870 4.280 ;
        RECT 465.710 3.670 504.430 4.280 ;
        RECT 505.270 3.670 543.990 4.280 ;
        RECT 544.830 3.670 583.550 4.280 ;
        RECT 584.390 3.670 623.110 4.280 ;
        RECT 623.950 3.670 662.670 4.280 ;
        RECT 663.510 3.670 702.230 4.280 ;
        RECT 703.070 3.670 741.790 4.280 ;
        RECT 742.630 3.670 781.350 4.280 ;
        RECT 782.190 3.670 820.910 4.280 ;
        RECT 821.750 3.670 860.470 4.280 ;
        RECT 861.310 3.670 900.030 4.280 ;
        RECT 900.870 3.670 939.590 4.280 ;
        RECT 940.430 3.670 979.150 4.280 ;
        RECT 979.990 3.670 1018.710 4.280 ;
        RECT 1019.550 3.670 1058.270 4.280 ;
        RECT 1059.110 3.670 1097.830 4.280 ;
        RECT 1098.670 3.670 1137.390 4.280 ;
        RECT 1138.230 3.670 1176.950 4.280 ;
        RECT 1177.790 3.670 1216.510 4.280 ;
        RECT 1217.350 3.670 1256.070 4.280 ;
        RECT 1256.910 3.670 1295.630 4.280 ;
        RECT 1296.470 3.670 1335.190 4.280 ;
        RECT 1336.030 3.670 1374.750 4.280 ;
        RECT 1375.590 3.670 1414.310 4.280 ;
        RECT 1415.150 3.670 1453.870 4.280 ;
        RECT 1454.710 3.670 1493.430 4.280 ;
        RECT 1494.270 3.670 1532.990 4.280 ;
        RECT 1533.830 3.670 1572.550 4.280 ;
        RECT 1573.390 3.670 1612.110 4.280 ;
        RECT 1612.950 3.670 1651.670 4.280 ;
        RECT 1652.510 3.670 1691.230 4.280 ;
        RECT 1692.070 3.670 1730.790 4.280 ;
        RECT 1731.630 3.670 1770.350 4.280 ;
        RECT 1771.190 3.670 1809.910 4.280 ;
        RECT 1810.750 3.670 1849.470 4.280 ;
        RECT 1850.310 3.670 1889.030 4.280 ;
        RECT 1889.870 3.670 1914.825 4.280 ;
      LAYER met3 ;
        RECT 4.000 105.080 1916.000 108.965 ;
        RECT 4.000 103.680 1915.600 105.080 ;
        RECT 4.000 99.640 1916.000 103.680 ;
        RECT 4.400 98.240 1916.000 99.640 ;
        RECT 4.000 75.160 1916.000 98.240 ;
        RECT 4.000 73.760 1915.600 75.160 ;
        RECT 4.000 60.200 1916.000 73.760 ;
        RECT 4.400 58.800 1916.000 60.200 ;
        RECT 4.000 45.240 1916.000 58.800 ;
        RECT 4.000 43.840 1915.600 45.240 ;
        RECT 4.000 20.760 1916.000 43.840 ;
        RECT 4.400 19.360 1916.000 20.760 ;
        RECT 4.000 15.320 1916.000 19.360 ;
        RECT 4.000 13.920 1915.600 15.320 ;
        RECT 4.000 9.015 1916.000 13.920 ;
      LAYER met4 ;
        RECT 510.895 10.240 720.020 106.585 ;
        RECT 722.420 10.240 958.585 106.585 ;
        RECT 960.985 10.240 1197.155 106.585 ;
        RECT 1199.555 10.240 1401.785 106.585 ;
        RECT 510.895 9.695 1401.785 10.240 ;
  END
END digital_unison
END LIBRARY

