magic
tech sky130B
magscale 1 2
timestamp 1662952954
<< nwell >>
rect 25556 33458 25620 33522
<< psubdiff >>
rect 25260 32921 25311 32971
<< locali >>
rect 25260 32921 25311 32971
rect 22218 28813 22252 29386
rect 25824 28777 25858 29363
<< viali >>
rect 22218 29386 22252 29420
<< metal1 >>
rect 24646 34322 24698 34328
rect 23265 34272 24646 34316
rect 24646 34264 24698 34270
rect 24403 33834 24455 33840
rect 23252 33785 24403 33829
rect 24403 33776 24455 33782
rect 11806 33392 12084 33488
rect 13174 33484 14830 33488
rect 13174 33396 14592 33484
rect 14824 33396 14830 33484
rect 23531 33465 24319 33544
rect 25556 33515 25620 33522
rect 25556 33463 25562 33515
rect 25614 33463 25620 33515
rect 25556 33458 25620 33463
rect 13174 33392 14830 33396
rect 11806 32400 11906 33392
rect 19238 33336 19270 33344
rect 19130 33254 19270 33336
rect 11958 32944 12128 32950
rect 19238 32918 19270 33254
rect 24210 33213 24262 33219
rect 23256 33165 24210 33209
rect 24210 33155 24262 33161
rect 23547 32923 24335 33002
rect 25260 32921 25311 32971
rect 11958 32842 12128 32848
rect 23757 32741 23810 32747
rect 23250 32697 23757 32741
rect 23810 32689 24300 32735
rect 23757 32683 24300 32689
rect 23789 32681 24300 32683
rect 11806 32304 12114 32400
rect 23538 32371 24326 32450
rect 23593 32116 23646 32122
rect 23229 32059 23593 32116
rect 23645 32059 23646 32116
rect 23593 32053 23646 32059
rect 23225 31714 23277 31720
rect 23225 31547 23277 31553
rect 13786 30310 22323 30350
rect 25813 30311 25866 30350
rect 25881 30311 34418 30350
rect 25884 30310 34418 30311
rect 13796 30190 22333 30230
rect 22335 30190 22387 30230
rect 25686 30190 25738 30230
rect 25744 30190 34281 30230
rect 24402 30120 24456 30126
rect 24402 30068 24403 30120
rect 24455 30068 24456 30120
rect 24402 30062 24456 30068
rect 24645 29997 24697 30003
rect 24645 29939 24697 29945
rect 23758 29880 23810 29886
rect 23758 29822 23810 29828
rect 24209 29756 24261 29762
rect 24209 29698 24261 29704
rect 23593 28713 23645 28719
rect 22201 28666 23593 28711
rect 23645 28666 25876 28711
rect 23593 28654 23645 28661
rect 23224 28544 23276 28550
rect 22279 28496 23224 28541
rect 23276 28496 25793 28541
rect 23224 28486 23276 28492
rect 24645 28453 24697 28459
rect 23390 28447 23442 28453
rect 22206 28406 23390 28440
rect 23442 28406 24645 28440
rect 24697 28406 25871 28440
rect 24645 28395 24697 28401
rect 23390 28389 23442 28395
<< via1 >>
rect 24646 34270 24698 34322
rect 24403 33782 24455 33834
rect 14592 33396 14824 33484
rect 25562 33463 25614 33515
rect 11958 32848 12128 32944
rect 24210 33161 24262 33213
rect 26207 33158 26259 33210
rect 23757 32689 23810 32741
rect 26208 32684 26260 32736
rect 12278 32312 12510 32390
rect 13992 32312 14224 32390
rect 25478 32362 25690 32450
rect 23593 32059 23645 32116
rect 23225 31553 23277 31714
rect 24403 30068 24455 30120
rect 24645 29945 24697 29997
rect 23758 29828 23810 29880
rect 24209 29704 24261 29756
rect 23593 28661 23645 28713
rect 23224 28492 23276 28544
rect 23390 28395 23442 28447
rect 24645 28401 24697 28453
rect 24018 26706 24070 26758
<< metal2 >>
rect 24646 34322 24698 34328
rect 24646 34264 24698 34270
rect 24403 33834 24455 33840
rect 24403 33776 24455 33782
rect 14592 33484 14824 33490
rect 11958 32944 12128 32950
rect 11958 29658 12128 32848
rect 12205 32670 12239 33030
rect 12278 32390 12510 32400
rect 12278 30998 12510 32312
rect 13285 31160 13319 32880
rect 13804 31320 13838 32868
rect 13992 32390 14224 32400
rect 13776 31312 13866 31320
rect 13776 31242 13786 31312
rect 13856 31242 13866 31312
rect 13776 31234 13866 31242
rect 13256 31152 13346 31160
rect 13256 31082 13266 31152
rect 13336 31082 13346 31152
rect 13256 31074 13346 31082
rect 12268 30990 12520 30998
rect 12268 30886 12278 30990
rect 12510 30886 12520 30990
rect 12268 30876 12520 30886
rect 11916 29648 12168 29658
rect 13992 29656 14224 32312
rect 11916 29550 11926 29648
rect 12158 29550 12168 29648
rect 11916 29540 12168 29550
rect 13982 29648 14234 29656
rect 13982 29550 13992 29648
rect 14224 29550 14234 29648
rect 13982 29540 14234 29550
rect 14592 29472 14824 33396
rect 24210 33213 24262 33219
rect 24210 33155 24262 33161
rect 23757 32741 23810 32747
rect 23757 32683 23810 32689
rect 23593 32116 23646 32122
rect 23645 32059 23646 32116
rect 23593 32053 23646 32059
rect 23225 31714 23277 31720
rect 23225 31547 23277 31553
rect 21701 30758 21757 30767
rect 21701 30693 21757 30702
rect 21714 30481 21748 30693
rect 22096 30579 22130 30580
rect 22085 30570 22141 30579
rect 22085 30505 22141 30514
rect 14582 29456 14834 29472
rect 14582 29358 14592 29456
rect 14824 29358 14834 29456
rect 14582 29348 14834 29358
rect 21713 28443 21749 30481
rect 21713 28405 21922 28443
rect 22095 28442 22131 30505
rect 22202 28666 22240 28717
rect 23227 28551 23275 31547
rect 23594 28719 23644 32053
rect 23758 29880 23810 32683
rect 23758 29809 23810 29828
rect 24009 30958 24080 30970
rect 24009 30902 24017 30958
rect 24073 30902 24080 30958
rect 23593 28713 23645 28719
rect 23593 28654 23645 28661
rect 23224 28544 23276 28551
rect 23224 28486 23276 28492
rect 23390 28447 23442 28453
rect 23390 28389 23442 28395
rect 23400 26902 23434 28389
rect 24009 26758 24080 30902
rect 24211 29762 24260 33155
rect 24404 30126 24454 33776
rect 24402 30120 24456 30126
rect 24402 30068 24403 30120
rect 24455 30068 24456 30120
rect 24402 30062 24456 30068
rect 24404 30060 24454 30062
rect 24647 30003 24696 34264
rect 25560 33519 25618 33528
rect 25560 33452 25618 33461
rect 26195 33218 26275 33227
rect 26195 33155 26204 33218
rect 26266 33155 26275 33218
rect 26195 33146 26275 33155
rect 26206 32738 26262 32747
rect 26206 32673 26262 32682
rect 25468 32450 25700 32458
rect 25468 32362 25478 32450
rect 25690 32362 25700 32450
rect 25468 30986 25700 32362
rect 25468 30886 25474 30986
rect 25694 30886 25700 30986
rect 25468 30876 25700 30886
rect 25935 30765 25991 30774
rect 25935 30700 25991 30709
rect 24645 29997 24697 30003
rect 24645 29939 24697 29945
rect 24647 29925 24696 29939
rect 24209 29756 24261 29762
rect 24209 29698 24261 29704
rect 25820 28683 25861 28717
rect 24645 28453 24697 28459
rect 25946 28432 25980 30700
rect 26315 30568 26371 30578
rect 26315 30503 26371 30512
rect 26328 28440 26362 30503
rect 26152 28403 26362 28440
rect 24645 28395 24697 28401
rect 24656 26902 24690 28395
rect 24009 26706 24018 26758
rect 24070 26706 24080 26758
rect 24009 26700 24080 26706
rect 46310 26270 47033 26314
rect 24015 26077 24071 26081
rect 46310 26064 46355 26270
rect 1063 26007 1751 26051
<< via2 >>
rect 13786 31242 13856 31312
rect 13266 31082 13336 31152
rect 12278 30886 12510 30990
rect 11926 29550 12158 29648
rect 13992 29550 14224 29648
rect 21701 30702 21757 30758
rect 22085 30514 22141 30570
rect 14592 29358 14824 29456
rect 24017 30902 24073 30958
rect 25560 33515 25618 33519
rect 25560 33463 25562 33515
rect 25562 33463 25614 33515
rect 25614 33463 25618 33515
rect 25560 33461 25618 33463
rect 26204 33210 26266 33218
rect 26204 33158 26207 33210
rect 26207 33158 26259 33210
rect 26259 33158 26266 33210
rect 26204 33155 26266 33158
rect 26206 32736 26262 32738
rect 26206 32684 26208 32736
rect 26208 32684 26260 32736
rect 26260 32684 26262 32736
rect 26206 32682 26262 32684
rect 25478 32362 25690 32450
rect 25474 30886 25694 30986
rect 25935 30709 25991 30765
rect 26315 30512 26371 30568
<< metal3 >>
rect 25540 33522 25640 33539
rect 25540 33458 25556 33522
rect 25620 33458 25640 33522
rect 25540 33440 25640 33458
rect 26179 33227 26288 33244
rect 26179 33146 26195 33227
rect 26275 33146 26288 33227
rect 26179 33136 26288 33146
rect 26181 32744 26283 32760
rect 26181 32680 26201 32744
rect 26267 32680 26283 32744
rect 26181 32658 26283 32680
rect 25468 32450 25700 32458
rect 25468 32362 25478 32450
rect 25690 32362 25700 32450
rect 25468 32354 25700 32362
rect 13776 31312 13866 31320
rect 5834 31308 5920 31310
rect 5834 31244 5840 31308
rect 5914 31306 5920 31308
rect 13776 31306 13786 31312
rect 5914 31246 13786 31306
rect 5914 31244 5920 31246
rect 5834 31242 5920 31244
rect 13776 31242 13786 31246
rect 13856 31242 13866 31312
rect 13776 31234 13866 31242
rect 13256 31152 13346 31160
rect 13256 31082 13266 31152
rect 13336 31146 13346 31152
rect 42156 31148 42242 31150
rect 42156 31146 42162 31148
rect 13336 31086 42162 31146
rect 13336 31082 13346 31086
rect 42156 31084 42162 31086
rect 42236 31084 42242 31148
rect 42156 31082 42242 31084
rect 13256 31074 13346 31082
rect 12268 30990 12520 30998
rect 12268 30986 12278 30990
rect 17 30886 12278 30986
rect 12510 30986 12520 30990
rect 25468 30986 25700 30996
rect 12510 30971 25474 30986
rect 12510 30895 18624 30971
rect 18710 30958 25474 30971
rect 18710 30902 24017 30958
rect 24073 30902 25474 30958
rect 18710 30895 25474 30902
rect 12510 30886 25474 30895
rect 25694 30886 48059 30986
rect 12268 30876 12520 30886
rect 25468 30876 25700 30886
rect 21701 30758 21757 30767
rect 21701 30693 21757 30702
rect 25935 30765 25991 30774
rect 25935 30700 25991 30709
rect 17 30570 48059 30586
rect 17 30514 22085 30570
rect 22141 30568 48059 30570
rect 22141 30514 26315 30568
rect 17 30512 26315 30514
rect 26371 30512 48059 30568
rect 17 30486 48059 30512
rect 11916 29649 12168 29658
rect 13982 29649 14234 29656
rect 1242 29648 23388 29649
rect 1242 29550 11926 29648
rect 12158 29550 13992 29648
rect 14224 29636 23388 29648
rect 14224 29565 22940 29636
rect 23014 29565 23388 29636
rect 14224 29550 23388 29565
rect 1242 29549 23388 29550
rect 11916 29540 12168 29549
rect 13982 29540 14234 29549
rect 14582 29456 14834 29472
rect 14582 29358 14592 29456
rect 14824 29358 14834 29456
rect 28122 29358 33044 29458
rect 14582 29348 14834 29358
rect 23278 26637 23355 26642
rect 23278 26571 23284 26637
rect 23349 26571 23355 26637
rect 23278 26566 23355 26571
rect 24730 26636 24807 26642
rect 24730 26572 24737 26636
rect 24801 26572 24807 26636
rect 24730 26566 24807 26572
rect 24004 26083 24081 26092
rect 24004 26019 24010 26083
rect 24074 26019 24081 26083
rect 24004 26013 24081 26019
<< via3 >>
rect 25556 33519 25620 33522
rect 25556 33461 25560 33519
rect 25560 33461 25618 33519
rect 25618 33461 25620 33519
rect 25556 33458 25620 33461
rect 26195 33218 26275 33227
rect 26195 33155 26204 33218
rect 26204 33155 26266 33218
rect 26266 33155 26275 33218
rect 26195 33146 26275 33155
rect 26201 32738 26267 32744
rect 26201 32682 26206 32738
rect 26206 32682 26262 32738
rect 26262 32682 26267 32738
rect 26201 32680 26267 32682
rect 25478 32362 25690 32450
rect 5840 31244 5914 31308
rect 42162 31084 42236 31148
rect 18624 30895 18710 30971
rect 22940 29565 23014 29636
rect 22483 29373 22555 29445
rect 23284 26571 23349 26637
rect 24737 26572 24801 26636
rect 24010 26019 24074 26083
<< metal4 >>
rect 25550 33522 25625 33523
rect 25550 33458 25556 33522
rect 25620 33458 25625 33522
rect 25550 32458 25625 33458
rect 26179 33227 26288 33244
rect 26179 33221 26195 33227
rect 26043 33148 26195 33221
rect 25468 32450 25700 32458
rect 25468 32362 25478 32450
rect 25690 32362 25700 32450
rect 25468 32354 25700 32362
rect 26044 31948 26111 33148
rect 26179 33146 26195 33148
rect 26275 33146 26288 33227
rect 26179 33136 26288 33146
rect 26181 32744 26510 32754
rect 26181 32680 26201 32744
rect 26267 32680 26510 32744
rect 26181 32653 26510 32680
rect 24241 31876 26111 31948
rect 5834 31308 5920 31310
rect 5834 31244 5840 31308
rect 5914 31244 5920 31308
rect 5834 31242 5920 31244
rect 5840 25993 5914 31242
rect 18618 30971 18716 31705
rect 18618 30895 18624 30971
rect 18710 30895 18716 30971
rect 18618 30886 18716 30895
rect 22481 29445 22558 31376
rect 22933 29636 23019 31287
rect 22933 29565 22940 29636
rect 23014 29565 23019 29636
rect 22933 29532 23019 29565
rect 22481 29373 22483 29445
rect 22555 29373 22558 29445
rect 22481 29341 22558 29373
rect 24241 27210 24316 31876
rect 26444 31586 26508 32653
rect 23824 27124 24316 27210
rect 24737 31522 26508 31586
rect 23284 26642 23349 26769
rect 23278 26637 23355 26642
rect 23278 26571 23284 26637
rect 23349 26571 23355 26637
rect 23278 26566 23355 26571
rect 24010 26089 24076 27124
rect 24737 26642 24801 31522
rect 26444 31521 26508 31522
rect 42156 31148 42242 31150
rect 42156 31084 42162 31148
rect 42236 31084 42242 31148
rect 42156 31082 42242 31084
rect 24730 26636 24807 26642
rect 24730 26572 24737 26636
rect 24801 26572 24807 26636
rect 24730 26566 24807 26572
rect 24004 26083 24081 26089
rect 24004 26019 24010 26083
rect 24074 26019 24081 26083
rect 24004 26013 24081 26019
rect 42162 25993 42236 31082
use comparator  comparator_0
timestamp 1662929294
transform 1 0 23898 0 1 26079
box -1669 -1057 1961 897
use filter  filter_0
timestamp 1662946268
transform 1 0 1272 0 1 -2522
box -1298 2522 22766 33508
use filter  filter_1
timestamp 1662946268
transform -1 0 46804 0 1 -2522
box -1298 2522 22766 33508
use filter_clkgen  filter_clkgen_0
timestamp 1662952756
transform 1 0 20194 0 1 33421
box -1661 -2136 3360 1229
use level_shifter_low  level_shifter_low_0
timestamp 1662946268
transform 1 0 24311 0 1 32944
box -71 -46 2139 722
use level_shifter_low  level_shifter_low_1
timestamp 1662946268
transform 1 0 24311 0 -1 32948
box -71 -46 2139 722
use level_up_shifter_d_a  level_up_shifter_d_a_0
timestamp 1662952756
transform 1 0 11668 0 1 31806
box 402 498 2794 1683
<< labels >>
flabel metal2 13804 32480 13838 32868 1 FreeSans 1600 0 0 0 fb_inv
flabel metal2 13285 32481 13319 32868 1 FreeSans 1600 0 0 0 fb
flabel metal2 12205 32670 12239 33030 1 FreeSans 1600 0 0 0 fb1
port 1 n default input
flabel metal3 17 30886 48059 30986 1 FreeSans 3200 0 0 0 vccd
port 3 n default bidirectional
flabel metal3 28122 29358 33044 29458 1 FreeSans 3200 0 0 0 vdda
port 4 n default bidirectional
flabel metal3 1242 29549 23388 29649 1 FreeSans 3200 0 0 0 vssd
port 2 n default bidirectional
<< end >>
