magic
tech sky130B
magscale 1 2
timestamp 1654748254
<< error_p >>
rect 239 1920 291 1960
rect 385 1800 437 1840
rect 273 1024 307 1030
rect 273 1002 279 1024
rect 301 1002 307 1024
rect 273 996 307 1002
<< nwell >>
rect -125 328 357 497
<< nmos >>
rect 0 -10 30 74
rect 96 -10 126 74
<< pmos >>
rect 0 365 30 449
rect 96 365 126 449
<< ndiff >>
rect -66 48 0 74
rect -66 14 -57 48
rect -23 14 0 48
rect -66 -10 0 14
rect 30 49 96 74
rect 30 15 49 49
rect 83 15 96 49
rect 30 -10 96 15
rect 126 52 192 74
rect 126 18 150 52
rect 184 18 192 52
rect 126 -10 192 18
<< pdiff >>
rect -66 425 0 449
rect -66 391 -57 425
rect -23 391 0 425
rect -66 365 0 391
rect 30 424 96 449
rect 30 390 49 424
rect 83 390 96 424
rect 30 365 96 390
rect 126 421 192 449
rect 126 387 150 421
rect 184 387 192 421
rect 126 365 192 387
<< ndiffc >>
rect -57 14 -23 48
rect 49 15 83 49
rect 150 18 184 52
<< pdiffc >>
rect -57 391 -23 425
rect 49 390 83 424
rect 150 387 184 421
<< psubdiff >>
rect 256 50 305 74
rect 256 16 264 50
rect 298 16 305 50
rect 256 -8 305 16
<< nsubdiff >>
rect 260 424 317 449
rect 260 390 273 424
rect 307 390 317 424
rect 260 366 317 390
<< psubdiffcont >>
rect 264 16 298 50
<< nsubdiffcont >>
rect 273 390 307 424
<< poly >>
rect 0 449 30 475
rect 96 449 126 475
rect 0 328 30 365
rect -24 318 30 328
rect 96 328 126 365
rect 96 318 150 328
rect -30 284 -14 318
rect 20 284 36 318
rect 90 284 106 318
rect 140 284 156 318
rect -24 274 32 284
rect 96 274 150 284
rect 2 232 32 274
rect 2 202 126 232
rect 96 156 126 202
rect -24 146 30 156
rect 96 146 150 156
rect -30 112 -14 146
rect 20 112 36 146
rect 90 112 106 146
rect 140 112 156 146
rect -24 102 30 112
rect 0 74 30 102
rect 96 102 150 112
rect 96 74 126 102
rect 0 -36 30 -10
rect 96 -36 126 -10
<< polycont >>
rect -14 284 20 318
rect 106 284 140 318
rect -14 112 20 146
rect 106 112 140 146
<< locali >>
rect 273 1030 307 1057
rect -66 425 -11 449
rect -66 391 -57 425
rect -23 391 -11 425
rect -66 373 -11 391
rect 40 424 86 449
rect 40 390 49 424
rect 83 390 86 424
rect 40 373 86 390
rect 132 421 192 449
rect 132 387 150 421
rect 184 387 192 421
rect 132 365 192 387
rect 273 424 307 996
rect 273 374 307 390
rect -30 284 -14 318
rect 20 284 36 318
rect 90 284 106 318
rect 140 284 265 318
rect 299 284 302 318
rect 94 234 128 284
rect -14 200 128 234
rect -14 146 20 200
rect -30 112 -14 146
rect 20 112 36 146
rect 90 112 106 146
rect 140 112 395 146
rect 429 112 435 146
rect -66 48 -11 66
rect -66 14 -57 48
rect -23 14 -11 48
rect -66 -10 -11 14
rect 40 49 86 66
rect 40 15 49 49
rect 83 15 86 49
rect 40 -10 86 15
rect 132 52 192 74
rect 132 18 150 52
rect 184 18 192 52
rect 132 -10 192 18
rect 264 50 298 66
rect 264 0 298 16
<< viali >>
rect 273 996 307 1030
rect -57 391 -23 425
rect 49 390 83 424
rect 150 387 184 421
rect 265 284 299 318
rect 395 112 429 146
rect -57 14 -23 48
rect 49 15 83 49
rect 150 18 184 52
<< metal1 >>
rect 239 1920 291 1960
rect 385 1800 437 1840
rect -65 437 -13 441
rect -69 435 -11 437
rect -69 383 -65 435
rect -13 383 -11 435
rect 35 424 94 440
rect 139 433 191 438
rect 35 390 49 424
rect 83 390 94 424
rect -65 377 -13 383
rect 35 378 94 390
rect 138 432 196 433
rect 138 380 139 432
rect 191 380 196 432
rect -57 60 -23 377
rect 49 61 83 378
rect 138 375 196 380
rect 139 374 191 375
rect 150 64 184 374
rect 254 327 314 331
rect 252 275 258 327
rect 310 275 316 327
rect 254 270 314 275
rect 384 155 444 158
rect 382 103 388 155
rect 440 103 446 155
rect 384 98 444 103
rect -69 48 -11 60
rect -69 14 -57 48
rect -23 14 -11 48
rect -69 2 -11 14
rect 37 49 95 61
rect 37 15 49 49
rect 83 15 95 49
rect 37 3 95 15
rect 138 52 196 64
rect 138 18 150 52
rect 184 18 196 52
rect 138 6 196 18
<< via1 >>
rect -65 425 -13 435
rect -65 391 -57 425
rect -57 391 -23 425
rect -23 391 -13 425
rect -65 383 -13 391
rect 139 421 191 432
rect 139 387 150 421
rect 150 387 184 421
rect 184 387 191 421
rect 139 380 191 387
rect 258 318 310 327
rect 258 284 265 318
rect 265 284 299 318
rect 299 284 310 318
rect 258 275 310 284
rect 388 146 440 155
rect 388 112 395 146
rect 395 112 429 146
rect 429 112 440 146
rect 388 103 440 112
<< metal2 >>
rect -231 425 -197 2013
rect -65 435 -13 441
rect 151 438 185 2107
rect -231 391 -65 425
rect -65 377 -13 383
rect 139 432 191 438
rect 139 374 191 380
rect 252 275 258 327
rect 310 275 316 327
rect 382 103 388 155
rect 440 103 446 155
<< labels >>
flabel metal1 150 18 184 52 0 FreeSans 160 0 0 0 vref2
flabel metal1 -57 14 -23 48 0 FreeSans 160 0 0 0 vref1
flabel metal2 382 103 446 155 0 FreeSans 160 0 0 0 cclkb
flabel metal2 252 275 316 327 0 FreeSans 160 0 0 0 cclk
<< end >>
