magic
tech sky130A
magscale 1 2
timestamp 1647910269
<< error_s >>
rect 6881 6852 6887 6858
rect 9673 6852 9679 6858
rect 1870 6843 1890 6849
rect 4262 6843 4282 6849
rect 6913 6828 6917 6848
rect 9643 6828 9647 6848
rect 2415 6817 2424 6827
rect 4807 6817 4816 6827
rect 5627 6825 5640 6827
rect 5674 6825 5693 6827
rect 5674 6817 5675 6825
rect 1848 6795 1849 6807
rect 4240 6795 4241 6807
rect 2381 6783 2390 6793
rect 4773 6783 4782 6793
rect 5593 6791 5606 6793
rect 5708 6791 5727 6793
rect 5708 6783 5709 6791
rect 1819 6765 1831 6777
rect 4211 6765 4223 6777
rect 2087 6744 2099 6753
rect 4479 6744 4491 6753
rect 6955 6740 6959 6760
rect 9601 6740 9605 6760
rect 6911 6718 6917 6724
rect 9643 6718 9649 6724
rect 2125 6706 2137 6715
rect 4517 6706 4529 6715
rect 1263 6691 1280 6697
rect 3655 6691 3672 6697
rect 625 6362 631 6368
rect 1519 6362 1536 6363
rect 657 6338 661 6358
rect 1553 6328 1570 6329
rect 699 6250 703 6270
rect 6537 6263 6553 6265
rect 8169 6263 8182 6265
rect 8284 6263 8303 6265
rect 655 6228 661 6234
rect 6503 6229 6519 6231
rect 8203 6229 8216 6231
rect 8250 6229 8269 6231
rect 1487 5737 1500 5739
rect 1534 5737 1553 5739
rect 4523 5737 4536 5739
rect 4570 5737 4589 5739
rect 5899 5737 5918 5739
rect 5952 5737 5965 5739
rect 7463 5737 7482 5739
rect 7516 5737 7529 5739
rect 9447 5737 9463 5739
rect 1534 5729 1535 5737
rect 1453 5703 1466 5705
rect 1568 5703 1587 5705
rect 4489 5703 4502 5705
rect 4604 5703 4623 5705
rect 5865 5703 5884 5705
rect 5986 5703 5999 5705
rect 7429 5703 7448 5705
rect 7550 5703 7563 5705
rect 9481 5703 9497 5705
rect 1568 5695 1569 5703
rect 9857 5274 9863 5280
rect 1166 5253 1167 5259
rect 9827 5250 9831 5270
rect 1200 5219 1201 5225
rect 5791 5177 5792 5185
rect 1085 5175 1098 5177
rect 1200 5175 1219 5177
rect 2581 5175 2597 5177
rect 4029 5175 4042 5177
rect 4144 5175 4163 5177
rect 5773 5175 5792 5177
rect 5894 5175 5907 5177
rect 6419 5175 6435 5177
rect 8445 5175 8458 5177
rect 8560 5175 8579 5177
rect 9087 5175 9103 5177
rect 9785 5162 9789 5182
rect 5825 5143 5826 5151
rect 1119 5141 1132 5143
rect 1166 5141 1185 5143
rect 2547 5141 2563 5143
rect 4063 5141 4076 5143
rect 4110 5141 4129 5143
rect 5807 5141 5826 5143
rect 5860 5141 5873 5143
rect 6453 5141 6469 5143
rect 8479 5141 8492 5143
rect 8526 5141 8545 5143
rect 9121 5141 9137 5143
rect 9827 5140 9833 5146
rect 1839 4848 1848 4854
rect 1811 4820 1820 4826
rect 625 4676 631 4682
rect 657 4652 661 4672
rect 3603 4649 3616 4651
rect 3650 4649 3669 4651
rect 3569 4615 3582 4617
rect 3684 4615 3703 4617
rect 699 4564 703 4584
rect 655 4542 661 4548
rect 9262 4221 9279 4227
rect 8443 4165 8455 4174
rect 8791 4145 8803 4157
rect 8481 4127 8493 4136
rect 8761 4103 8762 4115
rect 1201 4087 1217 4089
rect 3199 4087 3215 4089
rect 4485 4087 4504 4089
rect 4606 4087 4619 4089
rect 8190 4087 8199 4097
rect 8732 4073 8752 4079
rect 1167 4053 1183 4055
rect 3233 4053 3249 4055
rect 4519 4053 4538 4055
rect 4572 4053 4585 4055
rect 8156 4053 8165 4063
rect 9008 3760 9016 3766
rect 9036 3732 9044 3738
rect 1238 3579 1258 3585
rect 704 3553 713 3563
rect 5307 3561 5323 3563
rect 5951 3561 5967 3563
rect 7007 3561 7020 3563
rect 7054 3561 7073 3563
rect 8567 3561 8586 3563
rect 8620 3561 8633 3563
rect 1279 3531 1280 3543
rect 738 3519 747 3529
rect 5341 3527 5357 3529
rect 5985 3527 6001 3529
rect 6973 3527 6986 3529
rect 7088 3527 7107 3529
rect 8533 3527 8552 3529
rect 8654 3527 8667 3529
rect 1297 3501 1309 3513
rect 1029 3480 1041 3489
rect 991 3442 1003 3451
rect 1848 3427 1865 3433
rect 1945 3133 1962 3139
rect 7514 3133 7531 3139
rect 625 3098 631 3104
rect 4245 3098 4251 3104
rect 8753 3098 8759 3104
rect 9733 3098 9739 3104
rect 657 3074 661 3094
rect 2769 3077 2781 3086
rect 4215 3074 4219 3094
rect 6695 3077 6707 3086
rect 8723 3074 8727 3094
rect 9765 3074 9769 3094
rect 2421 3057 2433 3069
rect 7043 3057 7055 3069
rect 2731 3039 2743 3048
rect 6733 3039 6745 3048
rect 2462 3015 2463 3027
rect 7013 3015 7014 3027
rect 699 2986 703 3006
rect 3025 2999 3034 3009
rect 2472 2985 2492 2991
rect 4173 2986 4177 3006
rect 6442 2999 6451 3009
rect 6984 2985 7004 2991
rect 8681 2986 8685 3006
rect 9807 2986 9811 3006
rect 655 2964 661 2970
rect 3059 2965 3068 2975
rect 4215 2964 4221 2970
rect 6408 2965 6417 2975
rect 8723 2964 8729 2970
rect 9763 2964 9769 2970
rect 4354 2491 4374 2497
rect 9322 2491 9342 2497
rect 4899 2465 4908 2475
rect 6913 2473 6929 2475
rect 9867 2465 9876 2475
rect 4332 2443 4333 2455
rect 9300 2443 9301 2455
rect 4865 2431 4874 2441
rect 6879 2439 6895 2441
rect 9833 2431 9842 2441
rect 4303 2413 4315 2425
rect 9271 2413 9283 2425
rect 4571 2392 4583 2401
rect 9539 2392 9551 2401
rect 1650 2375 1667 2376
rect 4609 2354 4621 2363
rect 9577 2354 9589 2363
rect 1684 2341 1701 2342
rect 3747 2339 3764 2345
rect 8715 2339 8732 2345
<< viali >>
rect 9505 6953 9539 6987
rect 7021 6885 7055 6919
rect 673 6817 707 6851
rect 949 6817 983 6851
rect 5641 6817 5675 6851
rect 3065 6749 3099 6783
rect 5549 6749 5583 6783
rect 5733 6749 5767 6783
rect 6837 6749 6871 6783
rect 8125 6749 8159 6783
rect 8309 6749 8343 6783
rect 9689 6749 9723 6783
rect 3341 6681 3375 6715
rect 2421 6613 2455 6647
rect 4813 6613 4847 6647
rect 8217 6613 8251 6647
rect 765 6409 799 6443
rect 1501 6409 1535 6443
rect 8217 6409 8251 6443
rect 9781 6341 9815 6375
rect 581 6273 615 6307
rect 1685 6273 1719 6307
rect 2145 6273 2179 6307
rect 2329 6273 2363 6307
rect 4077 6273 4111 6307
rect 5549 6273 5583 6307
rect 5641 6273 5675 6307
rect 5825 6273 5859 6307
rect 6469 6273 6503 6307
rect 6561 6273 6595 6307
rect 7021 6273 7055 6307
rect 7205 6273 7239 6307
rect 8125 6273 8159 6307
rect 8309 6273 8343 6307
rect 8769 6273 8803 6307
rect 8953 6273 8987 6307
rect 9045 6295 9079 6329
rect 9505 6273 9539 6307
rect 9597 6273 9631 6307
rect 4353 6205 4387 6239
rect 5733 6137 5767 6171
rect 8769 6137 8803 6171
rect 9505 6137 9539 6171
rect 2329 6069 2363 6103
rect 7021 6069 7055 6103
rect 2973 5865 3007 5899
rect 4537 5865 4571 5899
rect 5917 5865 5951 5899
rect 8585 5865 8619 5899
rect 9413 5865 9447 5899
rect 2053 5797 2087 5831
rect 5273 5797 5307 5831
rect 1501 5729 1535 5763
rect 765 5661 799 5695
rect 949 5661 983 5695
rect 1409 5661 1443 5695
rect 1593 5661 1627 5695
rect 2053 5661 2087 5695
rect 2145 5661 2179 5695
rect 2973 5661 3007 5695
rect 3157 5661 3191 5695
rect 4445 5661 4479 5695
rect 4629 5661 4663 5695
rect 5089 5661 5123 5695
rect 5825 5661 5859 5695
rect 6009 5661 6043 5695
rect 7389 5661 7423 5695
rect 7573 5661 7607 5695
rect 8125 5661 8159 5695
rect 8401 5661 8435 5695
rect 9505 5661 9539 5695
rect 2329 5593 2363 5627
rect 5181 5593 5215 5627
rect 5365 5593 5399 5627
rect 857 5525 891 5559
rect 7481 5525 7515 5559
rect 8217 5525 8251 5559
rect 2513 5321 2547 5355
rect 3157 5321 3191 5355
rect 4077 5321 4111 5355
rect 8493 5321 8527 5355
rect 1133 5253 1167 5287
rect 7757 5253 7791 5287
rect 7941 5253 7975 5287
rect 1041 5185 1075 5219
rect 1225 5185 1259 5219
rect 1685 5185 1719 5219
rect 1869 5185 1903 5219
rect 1961 5185 1995 5219
rect 2605 5185 2639 5219
rect 3065 5185 3099 5219
rect 3249 5185 3283 5219
rect 3985 5185 4019 5219
rect 4169 5185 4203 5219
rect 4813 5185 4847 5219
rect 4997 5185 5031 5219
rect 5733 5185 5767 5219
rect 5917 5185 5951 5219
rect 6377 5185 6411 5219
rect 7021 5185 7055 5219
rect 7205 5185 7239 5219
rect 7665 5185 7699 5219
rect 8401 5185 8435 5219
rect 8585 5185 8619 5219
rect 9045 5185 9079 5219
rect 9873 5185 9907 5219
rect 5825 5117 5859 5151
rect 7113 5117 7147 5151
rect 9137 5117 9171 5151
rect 1961 5049 1995 5083
rect 7665 5049 7699 5083
rect 9689 5049 9723 5083
rect 4813 4981 4847 5015
rect 6469 4981 6503 5015
rect 1961 4777 1995 4811
rect 3617 4777 3651 4811
rect 4353 4777 4387 4811
rect 4997 4777 5031 4811
rect 9597 4777 9631 4811
rect 7389 4709 7423 4743
rect 8401 4709 8435 4743
rect 581 4573 615 4607
rect 1593 4573 1627 4607
rect 1685 4573 1719 4607
rect 1777 4573 1811 4607
rect 3525 4573 3559 4607
rect 3709 4573 3743 4607
rect 4169 4573 4203 4607
rect 4353 4573 4387 4607
rect 4997 4573 5031 4607
rect 5273 4573 5307 4607
rect 6101 4573 6135 4607
rect 6285 4573 6319 4607
rect 6745 4573 6779 4607
rect 6929 4573 6963 4607
rect 7389 4573 7423 4607
rect 7573 4573 7607 4607
rect 8309 4573 8343 4607
rect 8401 4573 8435 4607
rect 8861 4573 8895 4607
rect 9137 4573 9171 4607
rect 9597 4573 9631 4607
rect 9689 4573 9723 4607
rect 5089 4505 5123 4539
rect 8125 4505 8159 4539
rect 8953 4505 8987 4539
rect 9873 4505 9907 4539
rect 765 4437 799 4471
rect 6193 4437 6227 4471
rect 6837 4437 6871 4471
rect 9045 4437 9079 4471
rect 1777 4233 1811 4267
rect 4537 4233 4571 4267
rect 5549 4233 5583 4267
rect 1869 4165 1903 4199
rect 5641 4165 5675 4199
rect 6837 4165 6871 4199
rect 7021 4165 7055 4199
rect 1225 4097 1259 4131
rect 1685 4097 1719 4131
rect 1961 4097 1995 4131
rect 2410 4097 2444 4131
rect 3157 4097 3191 4131
rect 4445 4097 4479 4131
rect 4629 4097 4663 4131
rect 5549 4097 5583 4131
rect 5825 4097 5859 4131
rect 6745 4097 6779 4131
rect 2697 4029 2731 4063
rect 8125 4029 8159 4063
rect 9597 4029 9631 4063
rect 9873 4029 9907 4063
rect 1133 3961 1167 3995
rect 2513 3961 2547 3995
rect 6745 3961 6779 3995
rect 2605 3893 2639 3927
rect 3249 3893 3283 3927
rect 4353 3689 4387 3723
rect 5273 3689 5307 3723
rect 5917 3689 5951 3723
rect 7021 3689 7055 3723
rect 8585 3689 8619 3723
rect 9137 3689 9171 3723
rect 673 3553 707 3587
rect 3617 3553 3651 3587
rect 2421 3485 2455 3519
rect 3065 3485 3099 3519
rect 4169 3485 4203 3519
rect 4353 3485 4387 3519
rect 5365 3485 5399 3519
rect 6009 3485 6043 3519
rect 6929 3485 6963 3519
rect 7113 3485 7147 3519
rect 8493 3485 8527 3519
rect 8677 3485 8711 3519
rect 9137 3485 9171 3519
rect 9321 3485 9355 3519
rect 2145 3417 2179 3451
rect 4077 3145 4111 3179
rect 6377 3145 6411 3179
rect 9873 3145 9907 3179
rect 1593 3077 1627 3111
rect 7849 3077 7883 3111
rect 581 3009 615 3043
rect 4261 3009 4295 3043
rect 8769 3009 8803 3043
rect 9689 3009 9723 3043
rect 1317 2941 1351 2975
rect 8125 2941 8159 2975
rect 765 2873 799 2907
rect 3065 2873 3099 2907
rect 8585 2873 8619 2907
rect 4905 2601 4939 2635
rect 6929 2601 6963 2635
rect 9873 2601 9907 2635
rect 3157 2465 3191 2499
rect 3433 2465 3467 2499
rect 8401 2465 8435 2499
rect 581 2397 615 2431
rect 1501 2397 1535 2431
rect 5641 2397 5675 2431
rect 6193 2397 6227 2431
rect 6837 2397 6871 2431
rect 8125 2397 8159 2431
rect 857 2329 891 2363
rect 1685 2261 1719 2295
<< metal1 >>
rect 276 7098 10580 7120
rect 276 7046 1839 7098
rect 1891 7046 1903 7098
rect 1955 7046 1967 7098
rect 2019 7046 2031 7098
rect 2083 7046 2095 7098
rect 2147 7046 5274 7098
rect 5326 7046 5338 7098
rect 5390 7046 5402 7098
rect 5454 7046 5466 7098
rect 5518 7046 5530 7098
rect 5582 7046 8708 7098
rect 8760 7046 8772 7098
rect 8824 7046 8836 7098
rect 8888 7046 8900 7098
rect 8952 7046 8964 7098
rect 9016 7046 10580 7098
rect 276 7024 10580 7046
rect 2866 6984 2872 6996
rect 676 6956 2872 6984
rect 676 6860 704 6956
rect 2866 6944 2872 6956
rect 2924 6944 2930 6996
rect 9493 6987 9551 6993
rect 9493 6984 9505 6987
rect 3160 6956 9505 6984
rect 658 6848 664 6860
rect 571 6820 664 6848
rect 658 6808 664 6820
rect 716 6808 722 6860
rect 937 6851 995 6857
rect 937 6817 949 6851
rect 983 6848 995 6851
rect 3160 6848 3188 6956
rect 9493 6953 9505 6956
rect 9539 6953 9551 6987
rect 9493 6947 9551 6953
rect 7009 6919 7067 6925
rect 7009 6885 7021 6919
rect 7055 6916 7067 6919
rect 7834 6916 7840 6928
rect 7055 6888 7840 6916
rect 7055 6885 7067 6888
rect 7009 6879 7067 6885
rect 7834 6876 7840 6888
rect 7892 6876 7898 6928
rect 983 6820 3188 6848
rect 983 6817 995 6820
rect 937 6811 995 6817
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 5629 6851 5687 6857
rect 5629 6848 5641 6851
rect 3476 6820 5641 6848
rect 3476 6808 3482 6820
rect 5629 6817 5641 6820
rect 5675 6817 5687 6851
rect 5629 6811 5687 6817
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 3053 6783 3111 6789
rect 3053 6780 3065 6783
rect 2832 6752 3065 6780
rect 2832 6740 2838 6752
rect 3053 6749 3065 6752
rect 3099 6749 3111 6783
rect 3053 6743 3111 6749
rect 5166 6740 5172 6792
rect 5224 6780 5230 6792
rect 5537 6783 5595 6789
rect 5537 6780 5549 6783
rect 5224 6752 5549 6780
rect 5224 6740 5230 6752
rect 5537 6749 5549 6752
rect 5583 6749 5595 6783
rect 5718 6780 5724 6792
rect 5679 6752 5724 6780
rect 5537 6743 5595 6749
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 6730 6740 6736 6792
rect 6788 6780 6794 6792
rect 6825 6783 6883 6789
rect 6825 6780 6837 6783
rect 6788 6752 6837 6780
rect 6788 6740 6794 6752
rect 6825 6749 6837 6752
rect 6871 6749 6883 6783
rect 6825 6743 6883 6749
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6780 8171 6783
rect 8202 6780 8208 6792
rect 8159 6752 8208 6780
rect 8159 6749 8171 6752
rect 8113 6743 8171 6749
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 8297 6783 8355 6789
rect 8297 6749 8309 6783
rect 8343 6780 8355 6783
rect 8754 6780 8760 6792
rect 8343 6752 8760 6780
rect 8343 6749 8355 6752
rect 8297 6743 8355 6749
rect 8754 6740 8760 6752
rect 8812 6740 8818 6792
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9456 6752 9689 6780
rect 9456 6740 9462 6752
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 2314 6712 2320 6724
rect 2162 6684 2320 6712
rect 2314 6672 2320 6684
rect 2372 6712 2378 6724
rect 2372 6684 2774 6712
rect 2372 6672 2378 6684
rect 2222 6604 2228 6656
rect 2280 6644 2286 6656
rect 2409 6647 2467 6653
rect 2409 6644 2421 6647
rect 2280 6616 2421 6644
rect 2280 6604 2286 6616
rect 2409 6613 2421 6616
rect 2455 6613 2467 6647
rect 2746 6644 2774 6684
rect 2866 6672 2872 6724
rect 2924 6712 2930 6724
rect 3329 6715 3387 6721
rect 3329 6712 3341 6715
rect 2924 6684 3341 6712
rect 2924 6672 2930 6684
rect 3329 6681 3341 6684
rect 3375 6681 3387 6715
rect 3329 6675 3387 6681
rect 3436 6684 3818 6712
rect 3436 6644 3464 6684
rect 2746 6616 3464 6644
rect 4801 6647 4859 6653
rect 2409 6607 2467 6613
rect 4801 6613 4813 6647
rect 4847 6644 4859 6647
rect 5902 6644 5908 6656
rect 4847 6616 5908 6644
rect 4847 6613 4859 6616
rect 4801 6607 4859 6613
rect 5902 6604 5908 6616
rect 5960 6644 5966 6656
rect 6546 6644 6552 6656
rect 5960 6616 6552 6644
rect 5960 6604 5966 6616
rect 6546 6604 6552 6616
rect 6604 6604 6610 6656
rect 7374 6604 7380 6656
rect 7432 6644 7438 6656
rect 8205 6647 8263 6653
rect 8205 6644 8217 6647
rect 7432 6616 8217 6644
rect 7432 6604 7438 6616
rect 8205 6613 8217 6616
rect 8251 6613 8263 6647
rect 8205 6607 8263 6613
rect 276 6554 10580 6576
rect 276 6502 3556 6554
rect 3608 6502 3620 6554
rect 3672 6502 3684 6554
rect 3736 6502 3748 6554
rect 3800 6502 3812 6554
rect 3864 6502 6991 6554
rect 7043 6502 7055 6554
rect 7107 6502 7119 6554
rect 7171 6502 7183 6554
rect 7235 6502 7247 6554
rect 7299 6502 10580 6554
rect 276 6480 10580 6502
rect 658 6400 664 6452
rect 716 6440 722 6452
rect 753 6443 811 6449
rect 753 6440 765 6443
rect 716 6412 765 6440
rect 716 6400 722 6412
rect 753 6409 765 6412
rect 799 6409 811 6443
rect 753 6403 811 6409
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 1489 6443 1547 6449
rect 1489 6440 1501 6443
rect 1452 6412 1501 6440
rect 1452 6400 1458 6412
rect 1489 6409 1501 6412
rect 1535 6409 1547 6443
rect 7374 6440 7380 6452
rect 1489 6403 1547 6409
rect 2746 6412 7380 6440
rect 2746 6372 2774 6412
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 8202 6440 8208 6452
rect 8163 6412 8208 6440
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 9582 6440 9588 6452
rect 8312 6412 9588 6440
rect 8312 6372 8340 6412
rect 9582 6400 9588 6412
rect 9640 6400 9646 6452
rect 1688 6344 2774 6372
rect 6472 6344 7052 6372
rect 566 6304 572 6316
rect 527 6276 572 6304
rect 566 6264 572 6276
rect 624 6264 630 6316
rect 1688 6313 1716 6344
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 2133 6307 2191 6313
rect 2133 6273 2145 6307
rect 2179 6304 2191 6307
rect 2222 6304 2228 6316
rect 2179 6276 2228 6304
rect 2179 6273 2191 6276
rect 2133 6267 2191 6273
rect 2222 6264 2228 6276
rect 2280 6264 2286 6316
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6304 2375 6307
rect 2958 6304 2964 6316
rect 2363 6276 2964 6304
rect 2363 6273 2375 6276
rect 2317 6267 2375 6273
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 3970 6264 3976 6316
rect 4028 6304 4034 6316
rect 4065 6307 4123 6313
rect 4065 6304 4077 6307
rect 4028 6276 4077 6304
rect 4028 6264 4034 6276
rect 4065 6273 4077 6276
rect 4111 6273 4123 6307
rect 4065 6267 4123 6273
rect 4522 6264 4528 6316
rect 4580 6304 4586 6316
rect 5537 6307 5595 6313
rect 5537 6304 5549 6307
rect 4580 6276 5549 6304
rect 4580 6264 4586 6276
rect 5537 6273 5549 6276
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 5626 6264 5632 6316
rect 5684 6304 5690 6316
rect 6472 6313 6500 6344
rect 5813 6307 5871 6313
rect 5684 6276 5729 6304
rect 5684 6264 5690 6276
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 6457 6307 6515 6313
rect 6457 6304 6469 6307
rect 5859 6276 6469 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 6457 6273 6469 6276
rect 6503 6273 6515 6307
rect 6457 6267 6515 6273
rect 6546 6264 6552 6316
rect 6604 6304 6610 6316
rect 7024 6313 7052 6344
rect 7116 6344 8340 6372
rect 7009 6307 7067 6313
rect 6604 6276 6649 6304
rect 6604 6264 6610 6276
rect 7009 6273 7021 6307
rect 7055 6273 7067 6307
rect 7009 6267 7067 6273
rect 4154 6196 4160 6248
rect 4212 6236 4218 6248
rect 4341 6239 4399 6245
rect 4341 6236 4353 6239
rect 4212 6208 4353 6236
rect 4212 6196 4218 6208
rect 4341 6205 4353 6208
rect 4387 6236 4399 6239
rect 7116 6236 7144 6344
rect 9030 6332 9036 6384
rect 9088 6332 9094 6384
rect 9122 6332 9128 6384
rect 9180 6372 9186 6384
rect 9398 6372 9404 6384
rect 9180 6344 9404 6372
rect 9180 6332 9186 6344
rect 9398 6332 9404 6344
rect 9456 6372 9462 6384
rect 9769 6375 9827 6381
rect 9769 6372 9781 6375
rect 9456 6344 9781 6372
rect 9456 6332 9462 6344
rect 9769 6341 9781 6344
rect 9815 6341 9827 6375
rect 9769 6335 9827 6341
rect 9033 6329 9091 6332
rect 7193 6307 7251 6313
rect 7193 6273 7205 6307
rect 7239 6304 7251 6307
rect 7374 6304 7380 6316
rect 7239 6276 7380 6304
rect 7239 6273 7251 6276
rect 7193 6267 7251 6273
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 8018 6264 8024 6316
rect 8076 6304 8082 6316
rect 8113 6307 8171 6313
rect 8113 6304 8125 6307
rect 8076 6276 8125 6304
rect 8076 6264 8082 6276
rect 8113 6273 8125 6276
rect 8159 6273 8171 6307
rect 8294 6304 8300 6316
rect 8255 6276 8300 6304
rect 8113 6267 8171 6273
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 8757 6307 8815 6313
rect 8757 6273 8769 6307
rect 8803 6304 8815 6307
rect 8846 6304 8852 6316
rect 8803 6276 8852 6304
rect 8803 6273 8815 6276
rect 8757 6267 8815 6273
rect 8846 6264 8852 6276
rect 8904 6264 8910 6316
rect 8941 6307 8999 6313
rect 8941 6273 8953 6307
rect 8987 6273 8999 6307
rect 9033 6295 9045 6329
rect 9079 6295 9091 6329
rect 9033 6289 9091 6295
rect 8941 6267 8999 6273
rect 4387 6208 7144 6236
rect 4387 6205 4399 6208
rect 4341 6199 4399 6205
rect 5718 6168 5724 6180
rect 5679 6140 5724 6168
rect 5718 6128 5724 6140
rect 5776 6128 5782 6180
rect 8754 6168 8760 6180
rect 8715 6140 8760 6168
rect 8754 6128 8760 6140
rect 8812 6128 8818 6180
rect 8846 6128 8852 6180
rect 8904 6128 8910 6180
rect 8956 6168 8984 6267
rect 9306 6264 9312 6316
rect 9364 6304 9370 6316
rect 9493 6307 9551 6313
rect 9493 6304 9505 6307
rect 9364 6276 9505 6304
rect 9364 6264 9370 6276
rect 9493 6273 9505 6276
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 9585 6307 9643 6313
rect 9585 6273 9597 6307
rect 9631 6273 9643 6307
rect 9585 6267 9643 6273
rect 9600 6236 9628 6267
rect 9766 6236 9772 6248
rect 9600 6208 9772 6236
rect 9214 6168 9220 6180
rect 8956 6140 9220 6168
rect 9214 6128 9220 6140
rect 9272 6128 9278 6180
rect 9490 6168 9496 6180
rect 9451 6140 9496 6168
rect 9490 6128 9496 6140
rect 9548 6128 9554 6180
rect 842 6060 848 6112
rect 900 6100 906 6112
rect 2317 6103 2375 6109
rect 2317 6100 2329 6103
rect 900 6072 2329 6100
rect 900 6060 906 6072
rect 2317 6069 2329 6072
rect 2363 6069 2375 6103
rect 2317 6063 2375 6069
rect 7009 6103 7067 6109
rect 7009 6069 7021 6103
rect 7055 6100 7067 6103
rect 7558 6100 7564 6112
rect 7055 6072 7564 6100
rect 7055 6069 7067 6072
rect 7009 6063 7067 6069
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 8864 6100 8892 6128
rect 9600 6100 9628 6208
rect 9766 6196 9772 6208
rect 9824 6196 9830 6248
rect 8864 6072 9628 6100
rect 276 6010 10580 6032
rect 276 5958 1839 6010
rect 1891 5958 1903 6010
rect 1955 5958 1967 6010
rect 2019 5958 2031 6010
rect 2083 5958 2095 6010
rect 2147 5958 5274 6010
rect 5326 5958 5338 6010
rect 5390 5958 5402 6010
rect 5454 5958 5466 6010
rect 5518 5958 5530 6010
rect 5582 5958 8708 6010
rect 8760 5958 8772 6010
rect 8824 5958 8836 6010
rect 8888 5958 8900 6010
rect 8952 5958 8964 6010
rect 9016 5958 10580 6010
rect 276 5936 10580 5958
rect 2958 5896 2964 5908
rect 2919 5868 2964 5896
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 4522 5896 4528 5908
rect 4483 5868 4528 5896
rect 4522 5856 4528 5868
rect 4580 5856 4586 5908
rect 5905 5899 5963 5905
rect 5905 5896 5917 5899
rect 5092 5868 5917 5896
rect 2041 5831 2099 5837
rect 2041 5797 2053 5831
rect 2087 5797 2099 5831
rect 2041 5791 2099 5797
rect 1489 5763 1547 5769
rect 1489 5760 1501 5763
rect 952 5732 1501 5760
rect 753 5695 811 5701
rect 753 5661 765 5695
rect 799 5692 811 5695
rect 842 5692 848 5704
rect 799 5664 848 5692
rect 799 5661 811 5664
rect 753 5655 811 5661
rect 842 5652 848 5664
rect 900 5652 906 5704
rect 952 5701 980 5732
rect 1489 5729 1501 5732
rect 1535 5729 1547 5763
rect 2056 5760 2084 5791
rect 5092 5760 5120 5868
rect 5905 5865 5917 5868
rect 5951 5865 5963 5899
rect 5905 5859 5963 5865
rect 8573 5899 8631 5905
rect 8573 5865 8585 5899
rect 8619 5896 8631 5899
rect 9214 5896 9220 5908
rect 8619 5868 9220 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 9398 5896 9404 5908
rect 9359 5868 9404 5896
rect 9398 5856 9404 5868
rect 9456 5856 9462 5908
rect 5166 5788 5172 5840
rect 5224 5828 5230 5840
rect 5261 5831 5319 5837
rect 5261 5828 5273 5831
rect 5224 5800 5273 5828
rect 5224 5788 5230 5800
rect 5261 5797 5273 5800
rect 5307 5797 5319 5831
rect 8478 5828 8484 5840
rect 5261 5791 5319 5797
rect 5920 5800 8484 5828
rect 5920 5760 5948 5800
rect 8478 5788 8484 5800
rect 8536 5788 8542 5840
rect 8570 5760 8576 5772
rect 1489 5723 1547 5729
rect 1596 5732 2084 5760
rect 4632 5732 5120 5760
rect 5184 5732 5672 5760
rect 1596 5701 1624 5732
rect 937 5695 995 5701
rect 937 5661 949 5695
rect 983 5661 995 5695
rect 937 5655 995 5661
rect 1397 5695 1455 5701
rect 1397 5661 1409 5695
rect 1443 5661 1455 5695
rect 1397 5655 1455 5661
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5661 1639 5695
rect 2038 5692 2044 5704
rect 1999 5664 2044 5692
rect 1581 5655 1639 5661
rect 1412 5624 1440 5655
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5692 2191 5695
rect 2222 5692 2228 5704
rect 2179 5664 2228 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 2222 5652 2228 5664
rect 2280 5652 2286 5704
rect 2958 5692 2964 5704
rect 2919 5664 2964 5692
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5692 3203 5695
rect 3418 5692 3424 5704
rect 3191 5664 3424 5692
rect 3191 5661 3203 5664
rect 3145 5655 3203 5661
rect 3418 5652 3424 5664
rect 3476 5652 3482 5704
rect 4430 5692 4436 5704
rect 4391 5664 4436 5692
rect 4430 5652 4436 5664
rect 4488 5652 4494 5704
rect 4632 5701 4660 5732
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5661 5135 5695
rect 5077 5655 5135 5661
rect 2317 5627 2375 5633
rect 1412 5596 2268 5624
rect 2240 5568 2268 5596
rect 2317 5593 2329 5627
rect 2363 5624 2375 5627
rect 2682 5624 2688 5636
rect 2363 5596 2688 5624
rect 2363 5593 2375 5596
rect 2317 5587 2375 5593
rect 2682 5584 2688 5596
rect 2740 5584 2746 5636
rect 5092 5568 5120 5655
rect 5184 5633 5212 5732
rect 5644 5692 5672 5732
rect 5828 5732 5948 5760
rect 6012 5732 8576 5760
rect 5828 5701 5856 5732
rect 6012 5704 6040 5732
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 5813 5695 5871 5701
rect 5813 5692 5825 5695
rect 5276 5664 5580 5692
rect 5644 5664 5825 5692
rect 5169 5627 5227 5633
rect 5169 5593 5181 5627
rect 5215 5593 5227 5627
rect 5169 5587 5227 5593
rect 845 5559 903 5565
rect 845 5525 857 5559
rect 891 5556 903 5559
rect 1486 5556 1492 5568
rect 891 5528 1492 5556
rect 891 5525 903 5528
rect 845 5519 903 5525
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 2222 5516 2228 5568
rect 2280 5516 2286 5568
rect 5074 5556 5080 5568
rect 4987 5528 5080 5556
rect 5074 5516 5080 5528
rect 5132 5556 5138 5568
rect 5276 5556 5304 5664
rect 5353 5627 5411 5633
rect 5353 5593 5365 5627
rect 5399 5593 5411 5627
rect 5552 5624 5580 5664
rect 5813 5661 5825 5664
rect 5859 5661 5871 5695
rect 5994 5692 6000 5704
rect 5955 5664 6000 5692
rect 5813 5655 5871 5661
rect 5994 5652 6000 5664
rect 6052 5652 6058 5704
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5661 7435 5695
rect 7558 5692 7564 5704
rect 7519 5664 7564 5692
rect 7377 5655 7435 5661
rect 7392 5624 7420 5655
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 8110 5692 8116 5704
rect 8071 5664 8116 5692
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5692 8447 5695
rect 9030 5692 9036 5704
rect 8435 5664 9036 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 9490 5692 9496 5704
rect 9451 5664 9496 5692
rect 9490 5652 9496 5664
rect 9548 5652 9554 5704
rect 5552 5596 7420 5624
rect 5353 5587 5411 5593
rect 5132 5528 5304 5556
rect 5368 5556 5396 5587
rect 6454 5556 6460 5568
rect 5368 5528 6460 5556
rect 5132 5516 5138 5528
rect 6454 5516 6460 5528
rect 6512 5516 6518 5568
rect 7469 5559 7527 5565
rect 7469 5525 7481 5559
rect 7515 5556 7527 5559
rect 8205 5559 8263 5565
rect 8205 5556 8217 5559
rect 7515 5528 8217 5556
rect 7515 5525 7527 5528
rect 7469 5519 7527 5525
rect 8205 5525 8217 5528
rect 8251 5525 8263 5559
rect 8205 5519 8263 5525
rect 276 5466 10580 5488
rect 276 5414 3556 5466
rect 3608 5414 3620 5466
rect 3672 5414 3684 5466
rect 3736 5414 3748 5466
rect 3800 5414 3812 5466
rect 3864 5414 6991 5466
rect 7043 5414 7055 5466
rect 7107 5414 7119 5466
rect 7171 5414 7183 5466
rect 7235 5414 7247 5466
rect 7299 5414 10580 5466
rect 276 5392 10580 5414
rect 2038 5312 2044 5364
rect 2096 5352 2102 5364
rect 2501 5355 2559 5361
rect 2501 5352 2513 5355
rect 2096 5324 2513 5352
rect 2096 5312 2102 5324
rect 2501 5321 2513 5324
rect 2547 5321 2559 5355
rect 2501 5315 2559 5321
rect 2682 5312 2688 5364
rect 2740 5352 2746 5364
rect 3145 5355 3203 5361
rect 3145 5352 3157 5355
rect 2740 5324 3157 5352
rect 2740 5312 2746 5324
rect 3145 5321 3157 5324
rect 3191 5321 3203 5355
rect 3145 5315 3203 5321
rect 4065 5355 4123 5361
rect 4065 5321 4077 5355
rect 4111 5352 4123 5355
rect 5074 5352 5080 5364
rect 4111 5324 5080 5352
rect 4111 5321 4123 5324
rect 4065 5315 4123 5321
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 5718 5312 5724 5364
rect 5776 5352 5782 5364
rect 7374 5352 7380 5364
rect 5776 5324 7380 5352
rect 5776 5312 5782 5324
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 8481 5355 8539 5361
rect 8481 5352 8493 5355
rect 8168 5324 8493 5352
rect 8168 5312 8174 5324
rect 8481 5321 8493 5324
rect 8527 5321 8539 5355
rect 8481 5315 8539 5321
rect 1121 5287 1179 5293
rect 1121 5253 1133 5287
rect 1167 5284 1179 5287
rect 1167 5256 3280 5284
rect 1167 5253 1179 5256
rect 1121 5247 1179 5253
rect 1029 5219 1087 5225
rect 1029 5185 1041 5219
rect 1075 5185 1087 5219
rect 1029 5179 1087 5185
rect 1213 5219 1271 5225
rect 1213 5185 1225 5219
rect 1259 5216 1271 5219
rect 1578 5216 1584 5228
rect 1259 5188 1584 5216
rect 1259 5185 1271 5188
rect 1213 5179 1271 5185
rect 1044 5148 1072 5179
rect 1578 5176 1584 5188
rect 1636 5176 1642 5228
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5185 1731 5219
rect 1854 5216 1860 5228
rect 1815 5188 1860 5216
rect 1673 5179 1731 5185
rect 1688 5148 1716 5179
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 2593 5219 2651 5225
rect 2593 5185 2605 5219
rect 2639 5185 2651 5219
rect 2593 5179 2651 5185
rect 1044 5120 1716 5148
rect 1688 5012 1716 5120
rect 1762 5108 1768 5160
rect 1820 5148 1826 5160
rect 1964 5148 1992 5179
rect 1820 5120 1992 5148
rect 2608 5148 2636 5179
rect 2866 5176 2872 5228
rect 2924 5216 2930 5228
rect 3252 5225 3280 5256
rect 4338 5244 4344 5296
rect 4396 5284 4402 5296
rect 7742 5284 7748 5296
rect 4396 5256 7748 5284
rect 4396 5244 4402 5256
rect 7742 5244 7748 5256
rect 7800 5244 7806 5296
rect 7929 5287 7987 5293
rect 7929 5253 7941 5287
rect 7975 5284 7987 5287
rect 9122 5284 9128 5296
rect 7975 5256 9128 5284
rect 7975 5253 7987 5256
rect 7929 5247 7987 5253
rect 9122 5244 9128 5256
rect 9180 5244 9186 5296
rect 3053 5219 3111 5225
rect 3053 5216 3065 5219
rect 2924 5188 3065 5216
rect 2924 5176 2930 5188
rect 3053 5185 3065 5188
rect 3099 5185 3111 5219
rect 3053 5179 3111 5185
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5185 3295 5219
rect 3237 5179 3295 5185
rect 3602 5176 3608 5228
rect 3660 5216 3666 5228
rect 3973 5219 4031 5225
rect 3973 5216 3985 5219
rect 3660 5188 3985 5216
rect 3660 5176 3666 5188
rect 3973 5185 3985 5188
rect 4019 5185 4031 5219
rect 3973 5179 4031 5185
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5216 4215 5219
rect 4706 5216 4712 5228
rect 4203 5188 4712 5216
rect 4203 5185 4215 5188
rect 4157 5179 4215 5185
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 4801 5219 4859 5225
rect 4801 5185 4813 5219
rect 4847 5185 4859 5219
rect 4801 5179 4859 5185
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5216 5043 5219
rect 5626 5216 5632 5228
rect 5031 5188 5632 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 3418 5148 3424 5160
rect 2608 5120 3424 5148
rect 1820 5108 1826 5120
rect 3418 5108 3424 5120
rect 3476 5108 3482 5160
rect 4816 5148 4844 5179
rect 5626 5176 5632 5188
rect 5684 5176 5690 5228
rect 5718 5176 5724 5228
rect 5776 5216 5782 5228
rect 5776 5188 5821 5216
rect 5776 5176 5782 5188
rect 5902 5176 5908 5228
rect 5960 5216 5966 5228
rect 6365 5219 6423 5225
rect 5960 5188 6005 5216
rect 5960 5176 5966 5188
rect 6365 5185 6377 5219
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 5813 5151 5871 5157
rect 5813 5148 5825 5151
rect 4816 5120 5825 5148
rect 5813 5117 5825 5120
rect 5859 5148 5871 5151
rect 6380 5148 6408 5179
rect 6546 5176 6552 5228
rect 6604 5216 6610 5228
rect 7009 5219 7067 5225
rect 7009 5216 7021 5219
rect 6604 5188 7021 5216
rect 6604 5176 6610 5188
rect 7009 5185 7021 5188
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 7193 5219 7251 5225
rect 7193 5185 7205 5219
rect 7239 5216 7251 5219
rect 7374 5216 7380 5228
rect 7239 5188 7380 5216
rect 7239 5185 7251 5188
rect 7193 5179 7251 5185
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 7558 5176 7564 5228
rect 7616 5216 7622 5228
rect 7653 5219 7711 5225
rect 7653 5216 7665 5219
rect 7616 5188 7665 5216
rect 7616 5176 7622 5188
rect 7653 5185 7665 5188
rect 7699 5185 7711 5219
rect 7653 5179 7711 5185
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5185 8447 5219
rect 8570 5216 8576 5228
rect 8531 5188 8576 5216
rect 8389 5179 8447 5185
rect 5859 5120 6408 5148
rect 7101 5151 7159 5157
rect 5859 5117 5871 5120
rect 5813 5111 5871 5117
rect 7101 5117 7113 5151
rect 7147 5148 7159 5151
rect 8294 5148 8300 5160
rect 7147 5120 8300 5148
rect 7147 5117 7159 5120
rect 7101 5111 7159 5117
rect 8294 5108 8300 5120
rect 8352 5148 8358 5160
rect 8404 5148 8432 5179
rect 8570 5176 8576 5188
rect 8628 5176 8634 5228
rect 9030 5216 9036 5228
rect 8991 5188 9036 5216
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 9398 5176 9404 5228
rect 9456 5216 9462 5228
rect 9861 5219 9919 5225
rect 9861 5216 9873 5219
rect 9456 5188 9873 5216
rect 9456 5176 9462 5188
rect 9861 5185 9873 5188
rect 9907 5185 9919 5219
rect 9861 5179 9919 5185
rect 8352 5120 8432 5148
rect 8352 5108 8358 5120
rect 8478 5108 8484 5160
rect 8536 5148 8542 5160
rect 9125 5151 9183 5157
rect 9125 5148 9137 5151
rect 8536 5120 9137 5148
rect 8536 5108 8542 5120
rect 9125 5117 9137 5120
rect 9171 5117 9183 5151
rect 9125 5111 9183 5117
rect 1949 5083 2007 5089
rect 1949 5049 1961 5083
rect 1995 5080 2007 5083
rect 2958 5080 2964 5092
rect 1995 5052 2964 5080
rect 1995 5049 2007 5052
rect 1949 5043 2007 5049
rect 2958 5040 2964 5052
rect 3016 5040 3022 5092
rect 7653 5083 7711 5089
rect 7653 5080 7665 5083
rect 3988 5052 7665 5080
rect 3988 5012 4016 5052
rect 7653 5049 7665 5052
rect 7699 5049 7711 5083
rect 7653 5043 7711 5049
rect 8386 5040 8392 5092
rect 8444 5080 8450 5092
rect 9677 5083 9735 5089
rect 9677 5080 9689 5083
rect 8444 5052 9689 5080
rect 8444 5040 8450 5052
rect 9677 5049 9689 5052
rect 9723 5049 9735 5083
rect 9677 5043 9735 5049
rect 4798 5012 4804 5024
rect 1688 4984 4016 5012
rect 4759 4984 4804 5012
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 4890 4972 4896 5024
rect 4948 5012 4954 5024
rect 5994 5012 6000 5024
rect 4948 4984 6000 5012
rect 4948 4972 4954 4984
rect 5994 4972 6000 4984
rect 6052 5012 6058 5024
rect 6270 5012 6276 5024
rect 6052 4984 6276 5012
rect 6052 4972 6058 4984
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6454 5012 6460 5024
rect 6367 4984 6460 5012
rect 6454 4972 6460 4984
rect 6512 5012 6518 5024
rect 8570 5012 8576 5024
rect 6512 4984 8576 5012
rect 6512 4972 6518 4984
rect 8570 4972 8576 4984
rect 8628 4972 8634 5024
rect 276 4922 10580 4944
rect 276 4870 1839 4922
rect 1891 4870 1903 4922
rect 1955 4870 1967 4922
rect 2019 4870 2031 4922
rect 2083 4870 2095 4922
rect 2147 4870 5274 4922
rect 5326 4870 5338 4922
rect 5390 4870 5402 4922
rect 5454 4870 5466 4922
rect 5518 4870 5530 4922
rect 5582 4870 8708 4922
rect 8760 4870 8772 4922
rect 8824 4870 8836 4922
rect 8888 4870 8900 4922
rect 8952 4870 8964 4922
rect 9016 4870 10580 4922
rect 276 4848 10580 4870
rect 1762 4768 1768 4820
rect 1820 4808 1826 4820
rect 1949 4811 2007 4817
rect 1949 4808 1961 4811
rect 1820 4780 1961 4808
rect 1820 4768 1826 4780
rect 1949 4777 1961 4780
rect 1995 4777 2007 4811
rect 3602 4808 3608 4820
rect 3563 4780 3608 4808
rect 1949 4771 2007 4777
rect 3602 4768 3608 4780
rect 3660 4768 3666 4820
rect 4338 4808 4344 4820
rect 4299 4780 4344 4808
rect 4338 4768 4344 4780
rect 4396 4768 4402 4820
rect 4430 4768 4436 4820
rect 4488 4808 4494 4820
rect 4985 4811 5043 4817
rect 4985 4808 4997 4811
rect 4488 4780 4997 4808
rect 4488 4768 4494 4780
rect 4985 4777 4997 4780
rect 5031 4777 5043 4811
rect 4985 4771 5043 4777
rect 9490 4768 9496 4820
rect 9548 4808 9554 4820
rect 9585 4811 9643 4817
rect 9585 4808 9597 4811
rect 9548 4780 9597 4808
rect 9548 4768 9554 4780
rect 9585 4777 9597 4780
rect 9631 4777 9643 4811
rect 9585 4771 9643 4777
rect 7377 4743 7435 4749
rect 5000 4712 6408 4740
rect 2314 4672 2320 4684
rect 1596 4644 2320 4672
rect 566 4604 572 4616
rect 527 4576 572 4604
rect 566 4564 572 4576
rect 624 4564 630 4616
rect 1596 4613 1624 4644
rect 2314 4632 2320 4644
rect 2372 4632 2378 4684
rect 4062 4672 4068 4684
rect 3528 4644 4068 4672
rect 1581 4607 1639 4613
rect 1581 4573 1593 4607
rect 1627 4573 1639 4607
rect 1581 4567 1639 4573
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4573 1731 4607
rect 1673 4567 1731 4573
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4604 1823 4607
rect 1854 4604 1860 4616
rect 1811 4576 1860 4604
rect 1811 4573 1823 4576
rect 1765 4567 1823 4573
rect 753 4471 811 4477
rect 753 4437 765 4471
rect 799 4468 811 4471
rect 1394 4468 1400 4480
rect 799 4440 1400 4468
rect 799 4437 811 4440
rect 753 4431 811 4437
rect 1394 4428 1400 4440
rect 1452 4428 1458 4480
rect 1688 4468 1716 4567
rect 1854 4564 1860 4576
rect 1912 4604 1918 4616
rect 3528 4613 3556 4644
rect 4062 4632 4068 4644
rect 4120 4672 4126 4684
rect 4120 4644 4384 4672
rect 4120 4632 4126 4644
rect 4356 4613 4384 4644
rect 3513 4607 3571 4613
rect 3513 4604 3525 4607
rect 1912 4576 3525 4604
rect 1912 4564 1918 4576
rect 3513 4573 3525 4576
rect 3559 4573 3571 4607
rect 3513 4567 3571 4573
rect 3697 4607 3755 4613
rect 3697 4573 3709 4607
rect 3743 4604 3755 4607
rect 4157 4607 4215 4613
rect 4157 4604 4169 4607
rect 3743 4576 4169 4604
rect 3743 4573 3755 4576
rect 3697 4567 3755 4573
rect 4157 4573 4169 4576
rect 4203 4573 4215 4607
rect 4157 4567 4215 4573
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 4172 4536 4200 4567
rect 4522 4564 4528 4616
rect 4580 4604 4586 4616
rect 5000 4613 5028 4712
rect 5644 4644 6316 4672
rect 5644 4616 5672 4644
rect 4985 4607 5043 4613
rect 4985 4604 4997 4607
rect 4580 4576 4997 4604
rect 4580 4564 4586 4576
rect 4985 4573 4997 4576
rect 5031 4573 5043 4607
rect 4985 4567 5043 4573
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4604 5319 4607
rect 5626 4604 5632 4616
rect 5307 4576 5632 4604
rect 5307 4573 5319 4576
rect 5261 4567 5319 4573
rect 5626 4564 5632 4576
rect 5684 4564 5690 4616
rect 6288 4613 6316 4644
rect 6089 4607 6147 4613
rect 6089 4604 6101 4607
rect 5736 4576 6101 4604
rect 5074 4536 5080 4548
rect 4172 4508 5080 4536
rect 5074 4496 5080 4508
rect 5132 4496 5138 4548
rect 1762 4468 1768 4480
rect 1688 4440 1768 4468
rect 1762 4428 1768 4440
rect 1820 4428 1826 4480
rect 5092 4468 5120 4496
rect 5736 4468 5764 4576
rect 6089 4573 6101 4576
rect 6135 4573 6147 4607
rect 6089 4567 6147 4573
rect 6273 4607 6331 4613
rect 6273 4573 6285 4607
rect 6319 4573 6331 4607
rect 6273 4567 6331 4573
rect 6380 4536 6408 4712
rect 7377 4709 7389 4743
rect 7423 4740 7435 4743
rect 8389 4743 8447 4749
rect 7423 4712 8340 4740
rect 7423 4709 7435 4712
rect 7377 4703 7435 4709
rect 6546 4632 6552 4684
rect 6604 4672 6610 4684
rect 8312 4672 8340 4712
rect 8389 4709 8401 4743
rect 8435 4740 8447 4743
rect 8435 4712 9628 4740
rect 8435 4709 8447 4712
rect 8389 4703 8447 4709
rect 9600 4672 9628 4712
rect 6604 4644 7512 4672
rect 8312 4644 8432 4672
rect 6604 4632 6610 4644
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 6733 4607 6791 4613
rect 6733 4604 6745 4607
rect 6696 4576 6745 4604
rect 6696 4564 6702 4576
rect 6733 4573 6745 4576
rect 6779 4573 6791 4607
rect 6914 4604 6920 4616
rect 6875 4576 6920 4604
rect 6733 4567 6791 4573
rect 6914 4564 6920 4576
rect 6972 4564 6978 4616
rect 7374 4604 7380 4616
rect 7335 4576 7380 4604
rect 7374 4564 7380 4576
rect 7432 4564 7438 4616
rect 7484 4604 7512 4644
rect 7561 4607 7619 4613
rect 7561 4604 7573 4607
rect 7484 4576 7573 4604
rect 7561 4573 7573 4576
rect 7607 4573 7619 4607
rect 8294 4604 8300 4616
rect 8255 4576 8300 4604
rect 7561 4567 7619 4573
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 8404 4613 8432 4644
rect 8496 4644 9260 4672
rect 9600 4644 9720 4672
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 8113 4539 8171 4545
rect 8113 4536 8125 4539
rect 6380 4508 8125 4536
rect 8113 4505 8125 4508
rect 8159 4505 8171 4539
rect 8113 4499 8171 4505
rect 8202 4496 8208 4548
rect 8260 4536 8266 4548
rect 8496 4536 8524 4644
rect 8570 4564 8576 4616
rect 8628 4604 8634 4616
rect 8849 4607 8907 4613
rect 8849 4604 8861 4607
rect 8628 4576 8861 4604
rect 8628 4564 8634 4576
rect 8849 4573 8861 4576
rect 8895 4573 8907 4607
rect 9122 4604 9128 4616
rect 9083 4576 9128 4604
rect 8849 4567 8907 4573
rect 9122 4564 9128 4576
rect 9180 4564 9186 4616
rect 9232 4604 9260 4644
rect 9692 4613 9720 4644
rect 9585 4607 9643 4613
rect 9585 4604 9597 4607
rect 9232 4576 9597 4604
rect 9585 4573 9597 4576
rect 9631 4573 9643 4607
rect 9585 4567 9643 4573
rect 9677 4607 9735 4613
rect 9677 4573 9689 4607
rect 9723 4573 9735 4607
rect 9677 4567 9735 4573
rect 8260 4508 8524 4536
rect 8941 4539 8999 4545
rect 8260 4496 8266 4508
rect 8941 4505 8953 4539
rect 8987 4505 8999 4539
rect 8941 4499 8999 4505
rect 9861 4539 9919 4545
rect 9861 4505 9873 4539
rect 9907 4505 9919 4539
rect 9861 4499 9919 4505
rect 6178 4468 6184 4480
rect 5092 4440 5764 4468
rect 6139 4440 6184 4468
rect 6178 4428 6184 4440
rect 6236 4428 6242 4480
rect 6822 4468 6828 4480
rect 6783 4440 6828 4468
rect 6822 4428 6828 4440
rect 6880 4428 6886 4480
rect 7742 4428 7748 4480
rect 7800 4468 7806 4480
rect 8956 4468 8984 4499
rect 7800 4440 8984 4468
rect 9033 4471 9091 4477
rect 7800 4428 7806 4440
rect 9033 4437 9045 4471
rect 9079 4468 9091 4471
rect 9876 4468 9904 4499
rect 9079 4440 9904 4468
rect 9079 4437 9091 4440
rect 9033 4431 9091 4437
rect 276 4378 10580 4400
rect 276 4326 3556 4378
rect 3608 4326 3620 4378
rect 3672 4326 3684 4378
rect 3736 4326 3748 4378
rect 3800 4326 3812 4378
rect 3864 4326 6991 4378
rect 7043 4326 7055 4378
rect 7107 4326 7119 4378
rect 7171 4326 7183 4378
rect 7235 4326 7247 4378
rect 7299 4326 10580 4378
rect 276 4304 10580 4326
rect 1670 4224 1676 4276
rect 1728 4264 1734 4276
rect 1765 4267 1823 4273
rect 1765 4264 1777 4267
rect 1728 4236 1777 4264
rect 1728 4224 1734 4236
rect 1765 4233 1777 4236
rect 1811 4233 1823 4267
rect 2314 4264 2320 4276
rect 2227 4236 2320 4264
rect 1765 4227 1823 4233
rect 2314 4224 2320 4236
rect 2372 4264 2378 4276
rect 4522 4264 4528 4276
rect 2372 4236 3372 4264
rect 4483 4236 4528 4264
rect 2372 4224 2378 4236
rect 1854 4196 1860 4208
rect 1815 4168 1860 4196
rect 1854 4156 1860 4168
rect 1912 4156 1918 4208
rect 1213 4131 1271 4137
rect 1213 4097 1225 4131
rect 1259 4128 1271 4131
rect 1670 4128 1676 4140
rect 1259 4100 1676 4128
rect 1259 4097 1271 4100
rect 1213 4091 1271 4097
rect 1670 4088 1676 4100
rect 1728 4088 1734 4140
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4097 2007 4131
rect 2332 4128 2360 4224
rect 3344 4196 3372 4236
rect 4522 4224 4528 4236
rect 4580 4224 4586 4276
rect 5537 4267 5595 4273
rect 5537 4233 5549 4267
rect 5583 4233 5595 4267
rect 9490 4264 9496 4276
rect 5537 4227 5595 4233
rect 5920 4236 6960 4264
rect 5552 4196 5580 4227
rect 5920 4208 5948 4236
rect 2976 4168 3280 4196
rect 3344 4168 5580 4196
rect 5629 4199 5687 4205
rect 2398 4131 2456 4137
rect 2398 4128 2410 4131
rect 2332 4100 2410 4128
rect 1949 4091 2007 4097
rect 2398 4097 2410 4100
rect 2444 4097 2456 4131
rect 2976 4128 3004 4168
rect 2398 4091 2456 4097
rect 2516 4100 3004 4128
rect 1964 4060 1992 4091
rect 2516 4060 2544 4100
rect 3050 4088 3056 4140
rect 3108 4128 3114 4140
rect 3145 4131 3203 4137
rect 3145 4128 3157 4131
rect 3108 4100 3157 4128
rect 3108 4088 3114 4100
rect 3145 4097 3157 4100
rect 3191 4097 3203 4131
rect 3252 4128 3280 4168
rect 5629 4165 5641 4199
rect 5675 4196 5687 4199
rect 5902 4196 5908 4208
rect 5675 4168 5908 4196
rect 5675 4165 5687 4168
rect 5629 4159 5687 4165
rect 5902 4156 5908 4168
rect 5960 4156 5966 4208
rect 6546 4196 6552 4208
rect 6012 4168 6552 4196
rect 6012 4140 6040 4168
rect 6546 4156 6552 4168
rect 6604 4156 6610 4208
rect 6822 4196 6828 4208
rect 6783 4168 6828 4196
rect 6822 4156 6828 4168
rect 6880 4156 6886 4208
rect 6932 4196 6960 4236
rect 8312 4236 9496 4264
rect 7009 4199 7067 4205
rect 7009 4196 7021 4199
rect 6932 4168 7021 4196
rect 7009 4165 7021 4168
rect 7055 4165 7067 4199
rect 7009 4159 7067 4165
rect 8018 4156 8024 4208
rect 8076 4196 8082 4208
rect 8312 4196 8340 4236
rect 9490 4224 9496 4236
rect 9548 4224 9554 4276
rect 8076 4168 8418 4196
rect 8076 4156 8082 4168
rect 3252 4100 3832 4128
rect 3145 4091 3203 4097
rect 1964 4032 2544 4060
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4060 2743 4063
rect 3234 4060 3240 4072
rect 2731 4032 3240 4060
rect 2731 4029 2743 4032
rect 2685 4023 2743 4029
rect 3234 4020 3240 4032
rect 3292 4020 3298 4072
rect 3804 4060 3832 4100
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 4433 4131 4491 4137
rect 4433 4128 4445 4131
rect 4120 4100 4445 4128
rect 4120 4088 4126 4100
rect 4433 4097 4445 4100
rect 4479 4097 4491 4131
rect 4614 4128 4620 4140
rect 4575 4100 4620 4128
rect 4433 4091 4491 4097
rect 4614 4088 4620 4100
rect 4672 4128 4678 4140
rect 4672 4100 5120 4128
rect 4672 4088 4678 4100
rect 4798 4060 4804 4072
rect 3804 4032 4804 4060
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 5092 4060 5120 4100
rect 5166 4088 5172 4140
rect 5224 4128 5230 4140
rect 5537 4131 5595 4137
rect 5537 4128 5549 4131
rect 5224 4100 5549 4128
rect 5224 4088 5230 4100
rect 5537 4097 5549 4100
rect 5583 4097 5595 4131
rect 5537 4091 5595 4097
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 5994 4128 6000 4140
rect 5859 4100 6000 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 5994 4088 6000 4100
rect 6052 4088 6058 4140
rect 6178 4088 6184 4140
rect 6236 4128 6242 4140
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 6236 4100 6745 4128
rect 6236 4088 6242 4100
rect 6733 4097 6745 4100
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 6638 4060 6644 4072
rect 5092 4032 6644 4060
rect 6638 4020 6644 4032
rect 6696 4060 6702 4072
rect 8113 4063 8171 4069
rect 8113 4060 8125 4063
rect 6696 4032 8125 4060
rect 6696 4020 6702 4032
rect 8113 4029 8125 4032
rect 8159 4060 8171 4063
rect 8570 4060 8576 4072
rect 8159 4032 8576 4060
rect 8159 4029 8171 4032
rect 8113 4023 8171 4029
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 9582 4060 9588 4072
rect 9543 4032 9588 4060
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 9858 4060 9864 4072
rect 9819 4032 9864 4060
rect 9858 4020 9864 4032
rect 9916 4020 9922 4072
rect 1121 3995 1179 4001
rect 1121 3961 1133 3995
rect 1167 3992 1179 3995
rect 2501 3995 2559 4001
rect 2501 3992 2513 3995
rect 1167 3964 2513 3992
rect 1167 3961 1179 3964
rect 1121 3955 1179 3961
rect 2501 3961 2513 3964
rect 2547 3961 2559 3995
rect 2501 3955 2559 3961
rect 6733 3995 6791 4001
rect 6733 3961 6745 3995
rect 6779 3992 6791 3995
rect 8202 3992 8208 4004
rect 6779 3964 8208 3992
rect 6779 3961 6791 3964
rect 6733 3955 6791 3961
rect 8202 3952 8208 3964
rect 8260 3952 8266 4004
rect 2593 3927 2651 3933
rect 2593 3893 2605 3927
rect 2639 3924 2651 3927
rect 2866 3924 2872 3936
rect 2639 3896 2872 3924
rect 2639 3893 2651 3896
rect 2593 3887 2651 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 3234 3924 3240 3936
rect 3147 3896 3240 3924
rect 3234 3884 3240 3896
rect 3292 3924 3298 3936
rect 6914 3924 6920 3936
rect 3292 3896 6920 3924
rect 3292 3884 3298 3896
rect 6914 3884 6920 3896
rect 6972 3884 6978 3936
rect 276 3834 10580 3856
rect 276 3782 1839 3834
rect 1891 3782 1903 3834
rect 1955 3782 1967 3834
rect 2019 3782 2031 3834
rect 2083 3782 2095 3834
rect 2147 3782 5274 3834
rect 5326 3782 5338 3834
rect 5390 3782 5402 3834
rect 5454 3782 5466 3834
rect 5518 3782 5530 3834
rect 5582 3782 8708 3834
rect 8760 3782 8772 3834
rect 8824 3782 8836 3834
rect 8888 3782 8900 3834
rect 8952 3782 8964 3834
rect 9016 3782 10580 3834
rect 276 3760 10580 3782
rect 1670 3680 1676 3732
rect 1728 3720 1734 3732
rect 4341 3723 4399 3729
rect 4341 3720 4353 3723
rect 1728 3692 4353 3720
rect 1728 3680 1734 3692
rect 4341 3689 4353 3692
rect 4387 3689 4399 3723
rect 4341 3683 4399 3689
rect 5166 3680 5172 3732
rect 5224 3720 5230 3732
rect 5261 3723 5319 3729
rect 5261 3720 5273 3723
rect 5224 3692 5273 3720
rect 5224 3680 5230 3692
rect 5261 3689 5273 3692
rect 5307 3689 5319 3723
rect 5261 3683 5319 3689
rect 5626 3680 5632 3732
rect 5684 3720 5690 3732
rect 5905 3723 5963 3729
rect 5905 3720 5917 3723
rect 5684 3692 5917 3720
rect 5684 3680 5690 3692
rect 5905 3689 5917 3692
rect 5951 3689 5963 3723
rect 5905 3683 5963 3689
rect 6270 3680 6276 3732
rect 6328 3720 6334 3732
rect 7009 3723 7067 3729
rect 7009 3720 7021 3723
rect 6328 3692 7021 3720
rect 6328 3680 6334 3692
rect 7009 3689 7021 3692
rect 7055 3689 7067 3723
rect 7009 3683 7067 3689
rect 8573 3723 8631 3729
rect 8573 3689 8585 3723
rect 8619 3720 8631 3723
rect 9030 3720 9036 3732
rect 8619 3692 9036 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 9030 3680 9036 3692
rect 9088 3680 9094 3732
rect 9122 3680 9128 3732
rect 9180 3720 9186 3732
rect 9180 3692 9225 3720
rect 9180 3680 9186 3692
rect 661 3587 719 3593
rect 661 3553 673 3587
rect 707 3584 719 3587
rect 3605 3587 3663 3593
rect 707 3556 3096 3584
rect 707 3553 719 3556
rect 661 3547 719 3553
rect 3068 3528 3096 3556
rect 3605 3553 3617 3587
rect 3651 3584 3663 3587
rect 4062 3584 4068 3596
rect 3651 3556 4068 3584
rect 3651 3553 3663 3556
rect 3605 3547 3663 3553
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 6012 3556 9352 3584
rect 6012 3528 6040 3556
rect 2409 3519 2467 3525
rect 2409 3485 2421 3519
rect 2455 3516 2467 3519
rect 3050 3516 3056 3528
rect 2455 3488 2912 3516
rect 3011 3488 3056 3516
rect 2455 3485 2467 3488
rect 2409 3479 2467 3485
rect 2133 3451 2191 3457
rect 1702 3420 2084 3448
rect 2056 3380 2084 3420
rect 2133 3417 2145 3451
rect 2179 3448 2191 3451
rect 2774 3448 2780 3460
rect 2179 3420 2780 3448
rect 2179 3417 2191 3420
rect 2133 3411 2191 3417
rect 2774 3408 2780 3420
rect 2832 3408 2838 3460
rect 2884 3448 2912 3488
rect 3050 3476 3056 3488
rect 3108 3476 3114 3528
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3485 4215 3519
rect 4157 3479 4215 3485
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3516 4399 3519
rect 4614 3516 4620 3528
rect 4387 3488 4620 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 4062 3448 4068 3460
rect 2884 3420 4068 3448
rect 4062 3408 4068 3420
rect 4120 3408 4126 3460
rect 4172 3448 4200 3479
rect 4614 3476 4620 3488
rect 4672 3476 4678 3528
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3516 5411 3519
rect 5718 3516 5724 3528
rect 5399 3488 5724 3516
rect 5399 3485 5411 3488
rect 5353 3479 5411 3485
rect 5718 3476 5724 3488
rect 5776 3476 5782 3528
rect 5994 3516 6000 3528
rect 5955 3488 6000 3516
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 6914 3516 6920 3528
rect 6875 3488 6920 3516
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7101 3519 7159 3525
rect 7101 3485 7113 3519
rect 7147 3516 7159 3519
rect 7374 3516 7380 3528
rect 7147 3488 7380 3516
rect 7147 3485 7159 3488
rect 7101 3479 7159 3485
rect 7374 3476 7380 3488
rect 7432 3476 7438 3528
rect 8496 3525 8524 3556
rect 8481 3519 8539 3525
rect 8481 3485 8493 3519
rect 8527 3485 8539 3519
rect 8481 3479 8539 3485
rect 8570 3476 8576 3528
rect 8628 3516 8634 3528
rect 9324 3525 9352 3556
rect 8665 3519 8723 3525
rect 8665 3516 8677 3519
rect 8628 3488 8677 3516
rect 8628 3476 8634 3488
rect 8665 3485 8677 3488
rect 8711 3516 8723 3519
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 8711 3488 9137 3516
rect 8711 3485 8723 3488
rect 8665 3479 8723 3485
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 5074 3448 5080 3460
rect 4172 3420 5080 3448
rect 5074 3408 5080 3420
rect 5132 3408 5138 3460
rect 2222 3380 2228 3392
rect 2056 3352 2228 3380
rect 2222 3340 2228 3352
rect 2280 3380 2286 3392
rect 2682 3380 2688 3392
rect 2280 3352 2688 3380
rect 2280 3340 2286 3352
rect 2682 3340 2688 3352
rect 2740 3340 2746 3392
rect 276 3290 10580 3312
rect 276 3238 3556 3290
rect 3608 3238 3620 3290
rect 3672 3238 3684 3290
rect 3736 3238 3748 3290
rect 3800 3238 3812 3290
rect 3864 3238 6991 3290
rect 7043 3238 7055 3290
rect 7107 3238 7119 3290
rect 7171 3238 7183 3290
rect 7235 3238 7247 3290
rect 7299 3238 10580 3290
rect 276 3216 10580 3238
rect 1394 3136 1400 3188
rect 1452 3136 1458 3188
rect 2866 3136 2872 3188
rect 2924 3176 2930 3188
rect 4065 3179 4123 3185
rect 4065 3176 4077 3179
rect 2924 3148 4077 3176
rect 2924 3136 2930 3148
rect 4065 3145 4077 3148
rect 4111 3145 4123 3179
rect 4065 3139 4123 3145
rect 5718 3136 5724 3188
rect 5776 3176 5782 3188
rect 6365 3179 6423 3185
rect 6365 3176 6377 3179
rect 5776 3148 6377 3176
rect 5776 3136 5782 3148
rect 6365 3145 6377 3148
rect 6411 3145 6423 3179
rect 9858 3176 9864 3188
rect 9819 3148 9864 3176
rect 6365 3139 6423 3145
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 1412 3108 1440 3136
rect 1581 3111 1639 3117
rect 1581 3108 1593 3111
rect 1412 3080 1593 3108
rect 1581 3077 1593 3080
rect 1627 3077 1639 3111
rect 1581 3071 1639 3077
rect 6822 3068 6828 3120
rect 6880 3068 6886 3120
rect 7834 3108 7840 3120
rect 7795 3080 7840 3108
rect 7834 3068 7840 3080
rect 7892 3068 7898 3120
rect 566 3040 572 3052
rect 527 3012 572 3040
rect 566 3000 572 3012
rect 624 3000 630 3052
rect 2682 3000 2688 3052
rect 2740 3000 2746 3052
rect 3970 3000 3976 3052
rect 4028 3040 4034 3052
rect 4249 3043 4307 3049
rect 4249 3040 4261 3043
rect 4028 3012 4261 3040
rect 4028 3000 4034 3012
rect 4249 3009 4261 3012
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 8757 3043 8815 3049
rect 8757 3009 8769 3043
rect 8803 3009 8815 3043
rect 9674 3040 9680 3052
rect 9635 3012 9680 3040
rect 8757 3003 8815 3009
rect 1305 2975 1363 2981
rect 1305 2941 1317 2975
rect 1351 2941 1363 2975
rect 1305 2935 1363 2941
rect 753 2907 811 2913
rect 753 2873 765 2907
rect 799 2904 811 2907
rect 1320 2904 1348 2935
rect 3418 2932 3424 2984
rect 3476 2972 3482 2984
rect 8113 2975 8171 2981
rect 8113 2972 8125 2975
rect 3476 2944 8125 2972
rect 3476 2932 3482 2944
rect 8113 2941 8125 2944
rect 8159 2972 8171 2975
rect 8159 2944 8616 2972
rect 8159 2941 8171 2944
rect 8113 2935 8171 2941
rect 799 2876 1348 2904
rect 3053 2907 3111 2913
rect 799 2873 811 2876
rect 753 2867 811 2873
rect 3053 2873 3065 2907
rect 3099 2904 3111 2907
rect 6178 2904 6184 2916
rect 3099 2876 6184 2904
rect 3099 2873 3111 2876
rect 3053 2867 3111 2873
rect 6178 2864 6184 2876
rect 6236 2864 6242 2916
rect 8588 2913 8616 2944
rect 8573 2907 8631 2913
rect 8573 2873 8585 2907
rect 8619 2873 8631 2907
rect 8573 2867 8631 2873
rect 6730 2796 6736 2848
rect 6788 2836 6794 2848
rect 8772 2836 8800 3003
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 6788 2808 8800 2836
rect 6788 2796 6794 2808
rect 276 2746 10580 2768
rect 276 2694 1839 2746
rect 1891 2694 1903 2746
rect 1955 2694 1967 2746
rect 2019 2694 2031 2746
rect 2083 2694 2095 2746
rect 2147 2694 5274 2746
rect 5326 2694 5338 2746
rect 5390 2694 5402 2746
rect 5454 2694 5466 2746
rect 5518 2694 5530 2746
rect 5582 2694 8708 2746
rect 8760 2694 8772 2746
rect 8824 2694 8836 2746
rect 8888 2694 8900 2746
rect 8952 2694 8964 2746
rect 9016 2694 10580 2746
rect 276 2672 10580 2694
rect 4893 2635 4951 2641
rect 4893 2601 4905 2635
rect 4939 2632 4951 2635
rect 5994 2632 6000 2644
rect 4939 2604 6000 2632
rect 4939 2601 4951 2604
rect 4893 2595 4951 2601
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 6917 2635 6975 2641
rect 6917 2601 6929 2635
rect 6963 2632 6975 2635
rect 7374 2632 7380 2644
rect 6963 2604 7380 2632
rect 6963 2601 6975 2604
rect 6917 2595 6975 2601
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 9490 2632 9496 2644
rect 8036 2604 9496 2632
rect 6822 2524 6828 2576
rect 6880 2564 6886 2576
rect 8036 2564 8064 2604
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 9766 2592 9772 2644
rect 9824 2632 9830 2644
rect 9861 2635 9919 2641
rect 9861 2632 9873 2635
rect 9824 2604 9873 2632
rect 9824 2592 9830 2604
rect 9861 2601 9873 2604
rect 9907 2601 9919 2635
rect 9861 2595 9919 2601
rect 6880 2536 8064 2564
rect 6880 2524 6886 2536
rect 1394 2456 1400 2508
rect 1452 2496 1458 2508
rect 3145 2499 3203 2505
rect 3145 2496 3157 2499
rect 1452 2468 3157 2496
rect 1452 2456 1458 2468
rect 3145 2465 3157 2468
rect 3191 2465 3203 2499
rect 3418 2496 3424 2508
rect 3379 2468 3424 2496
rect 3145 2459 3203 2465
rect 3418 2456 3424 2468
rect 3476 2456 3482 2508
rect 8386 2496 8392 2508
rect 8347 2468 8392 2496
rect 8386 2456 8392 2468
rect 8444 2456 8450 2508
rect 566 2428 572 2440
rect 527 2400 572 2428
rect 566 2388 572 2400
rect 624 2388 630 2440
rect 1486 2428 1492 2440
rect 1447 2400 1492 2428
rect 1486 2388 1492 2400
rect 1544 2388 1550 2440
rect 5074 2388 5080 2440
rect 5132 2428 5138 2440
rect 5629 2431 5687 2437
rect 5629 2428 5641 2431
rect 5132 2400 5641 2428
rect 5132 2388 5138 2400
rect 5629 2397 5641 2400
rect 5675 2397 5687 2431
rect 6178 2428 6184 2440
rect 6139 2400 6184 2428
rect 5629 2391 5687 2397
rect 6178 2388 6184 2400
rect 6236 2428 6242 2440
rect 6825 2431 6883 2437
rect 6825 2428 6837 2431
rect 6236 2400 6837 2428
rect 6236 2388 6242 2400
rect 6825 2397 6837 2400
rect 6871 2397 6883 2431
rect 6825 2391 6883 2397
rect 7834 2388 7840 2440
rect 7892 2428 7898 2440
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 7892 2400 8125 2428
rect 7892 2388 7898 2400
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 9490 2388 9496 2440
rect 9548 2388 9554 2440
rect 845 2363 903 2369
rect 845 2329 857 2363
rect 891 2360 903 2363
rect 891 2332 2728 2360
rect 4646 2332 6868 2360
rect 891 2329 903 2332
rect 845 2323 903 2329
rect 2700 2304 2728 2332
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 1360 2264 1685 2292
rect 1360 2252 1366 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 2682 2252 2688 2304
rect 2740 2292 2746 2304
rect 4724 2292 4752 2332
rect 6840 2304 6868 2332
rect 2740 2264 4752 2292
rect 2740 2252 2746 2264
rect 6822 2252 6828 2304
rect 6880 2252 6886 2304
rect 276 2202 10580 2224
rect 276 2150 3556 2202
rect 3608 2150 3620 2202
rect 3672 2150 3684 2202
rect 3736 2150 3748 2202
rect 3800 2150 3812 2202
rect 3864 2150 6991 2202
rect 7043 2150 7055 2202
rect 7107 2150 7119 2202
rect 7171 2150 7183 2202
rect 7235 2150 7247 2202
rect 7299 2150 10580 2202
rect 276 2128 10580 2150
<< via1 >>
rect 1839 7046 1891 7098
rect 1903 7046 1955 7098
rect 1967 7046 2019 7098
rect 2031 7046 2083 7098
rect 2095 7046 2147 7098
rect 5274 7046 5326 7098
rect 5338 7046 5390 7098
rect 5402 7046 5454 7098
rect 5466 7046 5518 7098
rect 5530 7046 5582 7098
rect 8708 7046 8760 7098
rect 8772 7046 8824 7098
rect 8836 7046 8888 7098
rect 8900 7046 8952 7098
rect 8964 7046 9016 7098
rect 2872 6944 2924 6996
rect 664 6851 716 6860
rect 664 6817 673 6851
rect 673 6817 707 6851
rect 707 6817 716 6851
rect 664 6808 716 6817
rect 7840 6876 7892 6928
rect 3424 6808 3476 6860
rect 2780 6740 2832 6792
rect 5172 6740 5224 6792
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 6736 6740 6788 6792
rect 8208 6740 8260 6792
rect 8760 6740 8812 6792
rect 9404 6740 9456 6792
rect 2320 6672 2372 6724
rect 2228 6604 2280 6656
rect 2872 6672 2924 6724
rect 5908 6604 5960 6656
rect 6552 6604 6604 6656
rect 7380 6604 7432 6656
rect 3556 6502 3608 6554
rect 3620 6502 3672 6554
rect 3684 6502 3736 6554
rect 3748 6502 3800 6554
rect 3812 6502 3864 6554
rect 6991 6502 7043 6554
rect 7055 6502 7107 6554
rect 7119 6502 7171 6554
rect 7183 6502 7235 6554
rect 7247 6502 7299 6554
rect 664 6400 716 6452
rect 1400 6400 1452 6452
rect 7380 6400 7432 6452
rect 8208 6443 8260 6452
rect 8208 6409 8217 6443
rect 8217 6409 8251 6443
rect 8251 6409 8260 6443
rect 8208 6400 8260 6409
rect 9588 6400 9640 6452
rect 572 6307 624 6316
rect 572 6273 581 6307
rect 581 6273 615 6307
rect 615 6273 624 6307
rect 572 6264 624 6273
rect 2228 6264 2280 6316
rect 2964 6264 3016 6316
rect 3976 6264 4028 6316
rect 4528 6264 4580 6316
rect 5632 6307 5684 6316
rect 5632 6273 5641 6307
rect 5641 6273 5675 6307
rect 5675 6273 5684 6307
rect 5632 6264 5684 6273
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 4160 6196 4212 6248
rect 9036 6332 9088 6384
rect 9128 6332 9180 6384
rect 9404 6332 9456 6384
rect 7380 6264 7432 6316
rect 8024 6264 8076 6316
rect 8300 6307 8352 6316
rect 8300 6273 8309 6307
rect 8309 6273 8343 6307
rect 8343 6273 8352 6307
rect 8300 6264 8352 6273
rect 8852 6264 8904 6316
rect 5724 6171 5776 6180
rect 5724 6137 5733 6171
rect 5733 6137 5767 6171
rect 5767 6137 5776 6171
rect 5724 6128 5776 6137
rect 8760 6171 8812 6180
rect 8760 6137 8769 6171
rect 8769 6137 8803 6171
rect 8803 6137 8812 6171
rect 8760 6128 8812 6137
rect 8852 6128 8904 6180
rect 9312 6264 9364 6316
rect 9220 6128 9272 6180
rect 9496 6171 9548 6180
rect 9496 6137 9505 6171
rect 9505 6137 9539 6171
rect 9539 6137 9548 6171
rect 9496 6128 9548 6137
rect 848 6060 900 6112
rect 7564 6060 7616 6112
rect 9772 6196 9824 6248
rect 1839 5958 1891 6010
rect 1903 5958 1955 6010
rect 1967 5958 2019 6010
rect 2031 5958 2083 6010
rect 2095 5958 2147 6010
rect 5274 5958 5326 6010
rect 5338 5958 5390 6010
rect 5402 5958 5454 6010
rect 5466 5958 5518 6010
rect 5530 5958 5582 6010
rect 8708 5958 8760 6010
rect 8772 5958 8824 6010
rect 8836 5958 8888 6010
rect 8900 5958 8952 6010
rect 8964 5958 9016 6010
rect 2964 5899 3016 5908
rect 2964 5865 2973 5899
rect 2973 5865 3007 5899
rect 3007 5865 3016 5899
rect 2964 5856 3016 5865
rect 4528 5899 4580 5908
rect 4528 5865 4537 5899
rect 4537 5865 4571 5899
rect 4571 5865 4580 5899
rect 4528 5856 4580 5865
rect 848 5652 900 5704
rect 9220 5856 9272 5908
rect 9404 5899 9456 5908
rect 9404 5865 9413 5899
rect 9413 5865 9447 5899
rect 9447 5865 9456 5899
rect 9404 5856 9456 5865
rect 5172 5788 5224 5840
rect 8484 5788 8536 5840
rect 2044 5695 2096 5704
rect 2044 5661 2053 5695
rect 2053 5661 2087 5695
rect 2087 5661 2096 5695
rect 2044 5652 2096 5661
rect 2228 5652 2280 5704
rect 2964 5695 3016 5704
rect 2964 5661 2973 5695
rect 2973 5661 3007 5695
rect 3007 5661 3016 5695
rect 2964 5652 3016 5661
rect 3424 5652 3476 5704
rect 4436 5695 4488 5704
rect 4436 5661 4445 5695
rect 4445 5661 4479 5695
rect 4479 5661 4488 5695
rect 4436 5652 4488 5661
rect 2688 5584 2740 5636
rect 8576 5720 8628 5772
rect 1492 5516 1544 5568
rect 2228 5516 2280 5568
rect 5080 5516 5132 5568
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 7564 5695 7616 5704
rect 7564 5661 7573 5695
rect 7573 5661 7607 5695
rect 7607 5661 7616 5695
rect 7564 5652 7616 5661
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 9036 5652 9088 5704
rect 9496 5695 9548 5704
rect 9496 5661 9505 5695
rect 9505 5661 9539 5695
rect 9539 5661 9548 5695
rect 9496 5652 9548 5661
rect 6460 5516 6512 5568
rect 3556 5414 3608 5466
rect 3620 5414 3672 5466
rect 3684 5414 3736 5466
rect 3748 5414 3800 5466
rect 3812 5414 3864 5466
rect 6991 5414 7043 5466
rect 7055 5414 7107 5466
rect 7119 5414 7171 5466
rect 7183 5414 7235 5466
rect 7247 5414 7299 5466
rect 2044 5312 2096 5364
rect 2688 5312 2740 5364
rect 5080 5312 5132 5364
rect 5724 5312 5776 5364
rect 7380 5312 7432 5364
rect 8116 5312 8168 5364
rect 1584 5176 1636 5228
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 1768 5108 1820 5160
rect 2872 5176 2924 5228
rect 4344 5244 4396 5296
rect 7748 5287 7800 5296
rect 7748 5253 7757 5287
rect 7757 5253 7791 5287
rect 7791 5253 7800 5287
rect 7748 5244 7800 5253
rect 9128 5244 9180 5296
rect 3608 5176 3660 5228
rect 4712 5176 4764 5228
rect 3424 5108 3476 5160
rect 5632 5176 5684 5228
rect 5724 5219 5776 5228
rect 5724 5185 5733 5219
rect 5733 5185 5767 5219
rect 5767 5185 5776 5219
rect 5724 5176 5776 5185
rect 5908 5219 5960 5228
rect 5908 5185 5917 5219
rect 5917 5185 5951 5219
rect 5951 5185 5960 5219
rect 5908 5176 5960 5185
rect 6552 5176 6604 5228
rect 7380 5176 7432 5228
rect 7564 5176 7616 5228
rect 8576 5219 8628 5228
rect 8300 5108 8352 5160
rect 8576 5185 8585 5219
rect 8585 5185 8619 5219
rect 8619 5185 8628 5219
rect 8576 5176 8628 5185
rect 9036 5219 9088 5228
rect 9036 5185 9045 5219
rect 9045 5185 9079 5219
rect 9079 5185 9088 5219
rect 9036 5176 9088 5185
rect 9404 5176 9456 5228
rect 8484 5108 8536 5160
rect 2964 5040 3016 5092
rect 8392 5040 8444 5092
rect 4804 5015 4856 5024
rect 4804 4981 4813 5015
rect 4813 4981 4847 5015
rect 4847 4981 4856 5015
rect 4804 4972 4856 4981
rect 4896 4972 4948 5024
rect 6000 4972 6052 5024
rect 6276 4972 6328 5024
rect 6460 5015 6512 5024
rect 6460 4981 6469 5015
rect 6469 4981 6503 5015
rect 6503 4981 6512 5015
rect 6460 4972 6512 4981
rect 8576 4972 8628 5024
rect 1839 4870 1891 4922
rect 1903 4870 1955 4922
rect 1967 4870 2019 4922
rect 2031 4870 2083 4922
rect 2095 4870 2147 4922
rect 5274 4870 5326 4922
rect 5338 4870 5390 4922
rect 5402 4870 5454 4922
rect 5466 4870 5518 4922
rect 5530 4870 5582 4922
rect 8708 4870 8760 4922
rect 8772 4870 8824 4922
rect 8836 4870 8888 4922
rect 8900 4870 8952 4922
rect 8964 4870 9016 4922
rect 1768 4768 1820 4820
rect 3608 4811 3660 4820
rect 3608 4777 3617 4811
rect 3617 4777 3651 4811
rect 3651 4777 3660 4811
rect 3608 4768 3660 4777
rect 4344 4811 4396 4820
rect 4344 4777 4353 4811
rect 4353 4777 4387 4811
rect 4387 4777 4396 4811
rect 4344 4768 4396 4777
rect 4436 4768 4488 4820
rect 9496 4768 9548 4820
rect 572 4607 624 4616
rect 572 4573 581 4607
rect 581 4573 615 4607
rect 615 4573 624 4607
rect 572 4564 624 4573
rect 2320 4632 2372 4684
rect 1400 4428 1452 4480
rect 1860 4564 1912 4616
rect 4068 4632 4120 4684
rect 4528 4564 4580 4616
rect 5632 4564 5684 4616
rect 5080 4539 5132 4548
rect 5080 4505 5089 4539
rect 5089 4505 5123 4539
rect 5123 4505 5132 4539
rect 5080 4496 5132 4505
rect 1768 4428 1820 4480
rect 6552 4632 6604 4684
rect 6644 4564 6696 4616
rect 6920 4607 6972 4616
rect 6920 4573 6929 4607
rect 6929 4573 6963 4607
rect 6963 4573 6972 4607
rect 6920 4564 6972 4573
rect 7380 4607 7432 4616
rect 7380 4573 7389 4607
rect 7389 4573 7423 4607
rect 7423 4573 7432 4607
rect 7380 4564 7432 4573
rect 8300 4607 8352 4616
rect 8300 4573 8309 4607
rect 8309 4573 8343 4607
rect 8343 4573 8352 4607
rect 8300 4564 8352 4573
rect 8208 4496 8260 4548
rect 8576 4564 8628 4616
rect 9128 4607 9180 4616
rect 9128 4573 9137 4607
rect 9137 4573 9171 4607
rect 9171 4573 9180 4607
rect 9128 4564 9180 4573
rect 6184 4471 6236 4480
rect 6184 4437 6193 4471
rect 6193 4437 6227 4471
rect 6227 4437 6236 4471
rect 6184 4428 6236 4437
rect 6828 4471 6880 4480
rect 6828 4437 6837 4471
rect 6837 4437 6871 4471
rect 6871 4437 6880 4471
rect 6828 4428 6880 4437
rect 7748 4428 7800 4480
rect 3556 4326 3608 4378
rect 3620 4326 3672 4378
rect 3684 4326 3736 4378
rect 3748 4326 3800 4378
rect 3812 4326 3864 4378
rect 6991 4326 7043 4378
rect 7055 4326 7107 4378
rect 7119 4326 7171 4378
rect 7183 4326 7235 4378
rect 7247 4326 7299 4378
rect 1676 4224 1728 4276
rect 2320 4224 2372 4276
rect 4528 4267 4580 4276
rect 1860 4199 1912 4208
rect 1860 4165 1869 4199
rect 1869 4165 1903 4199
rect 1903 4165 1912 4199
rect 1860 4156 1912 4165
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 4528 4233 4537 4267
rect 4537 4233 4571 4267
rect 4571 4233 4580 4267
rect 4528 4224 4580 4233
rect 3056 4088 3108 4140
rect 5908 4156 5960 4208
rect 6552 4156 6604 4208
rect 6828 4199 6880 4208
rect 6828 4165 6837 4199
rect 6837 4165 6871 4199
rect 6871 4165 6880 4199
rect 6828 4156 6880 4165
rect 8024 4156 8076 4208
rect 9496 4224 9548 4276
rect 3240 4020 3292 4072
rect 4068 4088 4120 4140
rect 4620 4131 4672 4140
rect 4620 4097 4629 4131
rect 4629 4097 4663 4131
rect 4663 4097 4672 4131
rect 4620 4088 4672 4097
rect 4804 4020 4856 4072
rect 5172 4088 5224 4140
rect 6000 4088 6052 4140
rect 6184 4088 6236 4140
rect 6644 4020 6696 4072
rect 8576 4020 8628 4072
rect 9588 4063 9640 4072
rect 9588 4029 9597 4063
rect 9597 4029 9631 4063
rect 9631 4029 9640 4063
rect 9588 4020 9640 4029
rect 9864 4063 9916 4072
rect 9864 4029 9873 4063
rect 9873 4029 9907 4063
rect 9907 4029 9916 4063
rect 9864 4020 9916 4029
rect 8208 3952 8260 4004
rect 2872 3884 2924 3936
rect 3240 3927 3292 3936
rect 3240 3893 3249 3927
rect 3249 3893 3283 3927
rect 3283 3893 3292 3927
rect 3240 3884 3292 3893
rect 6920 3884 6972 3936
rect 1839 3782 1891 3834
rect 1903 3782 1955 3834
rect 1967 3782 2019 3834
rect 2031 3782 2083 3834
rect 2095 3782 2147 3834
rect 5274 3782 5326 3834
rect 5338 3782 5390 3834
rect 5402 3782 5454 3834
rect 5466 3782 5518 3834
rect 5530 3782 5582 3834
rect 8708 3782 8760 3834
rect 8772 3782 8824 3834
rect 8836 3782 8888 3834
rect 8900 3782 8952 3834
rect 8964 3782 9016 3834
rect 1676 3680 1728 3732
rect 5172 3680 5224 3732
rect 5632 3680 5684 3732
rect 6276 3680 6328 3732
rect 9036 3680 9088 3732
rect 9128 3723 9180 3732
rect 9128 3689 9137 3723
rect 9137 3689 9171 3723
rect 9171 3689 9180 3723
rect 9128 3680 9180 3689
rect 4068 3544 4120 3596
rect 3056 3519 3108 3528
rect 2780 3408 2832 3460
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 4068 3408 4120 3460
rect 4620 3476 4672 3528
rect 5724 3476 5776 3528
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 6920 3519 6972 3528
rect 6920 3485 6929 3519
rect 6929 3485 6963 3519
rect 6963 3485 6972 3519
rect 6920 3476 6972 3485
rect 7380 3476 7432 3528
rect 8576 3476 8628 3528
rect 5080 3408 5132 3460
rect 2228 3340 2280 3392
rect 2688 3340 2740 3392
rect 3556 3238 3608 3290
rect 3620 3238 3672 3290
rect 3684 3238 3736 3290
rect 3748 3238 3800 3290
rect 3812 3238 3864 3290
rect 6991 3238 7043 3290
rect 7055 3238 7107 3290
rect 7119 3238 7171 3290
rect 7183 3238 7235 3290
rect 7247 3238 7299 3290
rect 1400 3136 1452 3188
rect 2872 3136 2924 3188
rect 5724 3136 5776 3188
rect 9864 3179 9916 3188
rect 9864 3145 9873 3179
rect 9873 3145 9907 3179
rect 9907 3145 9916 3179
rect 9864 3136 9916 3145
rect 6828 3068 6880 3120
rect 7840 3111 7892 3120
rect 7840 3077 7849 3111
rect 7849 3077 7883 3111
rect 7883 3077 7892 3111
rect 7840 3068 7892 3077
rect 572 3043 624 3052
rect 572 3009 581 3043
rect 581 3009 615 3043
rect 615 3009 624 3043
rect 572 3000 624 3009
rect 2688 3000 2740 3052
rect 3976 3000 4028 3052
rect 9680 3043 9732 3052
rect 3424 2932 3476 2984
rect 6184 2864 6236 2916
rect 6736 2796 6788 2848
rect 9680 3009 9689 3043
rect 9689 3009 9723 3043
rect 9723 3009 9732 3043
rect 9680 3000 9732 3009
rect 1839 2694 1891 2746
rect 1903 2694 1955 2746
rect 1967 2694 2019 2746
rect 2031 2694 2083 2746
rect 2095 2694 2147 2746
rect 5274 2694 5326 2746
rect 5338 2694 5390 2746
rect 5402 2694 5454 2746
rect 5466 2694 5518 2746
rect 5530 2694 5582 2746
rect 8708 2694 8760 2746
rect 8772 2694 8824 2746
rect 8836 2694 8888 2746
rect 8900 2694 8952 2746
rect 8964 2694 9016 2746
rect 6000 2592 6052 2644
rect 7380 2592 7432 2644
rect 6828 2524 6880 2576
rect 9496 2592 9548 2644
rect 9772 2592 9824 2644
rect 1400 2456 1452 2508
rect 3424 2499 3476 2508
rect 3424 2465 3433 2499
rect 3433 2465 3467 2499
rect 3467 2465 3476 2499
rect 3424 2456 3476 2465
rect 8392 2499 8444 2508
rect 8392 2465 8401 2499
rect 8401 2465 8435 2499
rect 8435 2465 8444 2499
rect 8392 2456 8444 2465
rect 572 2431 624 2440
rect 572 2397 581 2431
rect 581 2397 615 2431
rect 615 2397 624 2431
rect 572 2388 624 2397
rect 1492 2431 1544 2440
rect 1492 2397 1501 2431
rect 1501 2397 1535 2431
rect 1535 2397 1544 2431
rect 1492 2388 1544 2397
rect 5080 2388 5132 2440
rect 6184 2431 6236 2440
rect 6184 2397 6193 2431
rect 6193 2397 6227 2431
rect 6227 2397 6236 2431
rect 6184 2388 6236 2397
rect 7840 2388 7892 2440
rect 9496 2388 9548 2440
rect 1308 2252 1360 2304
rect 2688 2252 2740 2304
rect 6828 2252 6880 2304
rect 3556 2150 3608 2202
rect 3620 2150 3672 2202
rect 3684 2150 3736 2202
rect 3748 2150 3800 2202
rect 3812 2150 3864 2202
rect 6991 2150 7043 2202
rect 7055 2150 7107 2202
rect 7119 2150 7171 2202
rect 7183 2150 7235 2202
rect 7247 2150 7299 2202
<< metal2 >>
rect 1306 7485 1362 7885
rect 3974 7485 4030 7885
rect 6734 7485 6790 7885
rect 9402 7485 9458 7885
rect 570 6896 626 6905
rect 570 6831 626 6840
rect 664 6860 716 6866
rect 584 6322 612 6831
rect 664 6802 716 6808
rect 676 6458 704 6802
rect 1320 6474 1348 7485
rect 1839 7100 2147 7120
rect 1839 7098 1845 7100
rect 1901 7098 1925 7100
rect 1981 7098 2005 7100
rect 2061 7098 2085 7100
rect 2141 7098 2147 7100
rect 1901 7046 1903 7098
rect 2083 7046 2085 7098
rect 1839 7044 1845 7046
rect 1901 7044 1925 7046
rect 1981 7044 2005 7046
rect 2061 7044 2085 7046
rect 2141 7044 2147 7046
rect 1839 7024 2147 7044
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2320 6724 2372 6730
rect 2320 6666 2372 6672
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 1320 6458 1440 6474
rect 664 6452 716 6458
rect 1320 6452 1452 6458
rect 1320 6446 1400 6452
rect 664 6394 716 6400
rect 1400 6394 1452 6400
rect 2240 6322 2268 6598
rect 572 6316 624 6322
rect 572 6258 624 6264
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 848 6112 900 6118
rect 848 6054 900 6060
rect 860 5710 888 6054
rect 1839 6012 2147 6032
rect 1839 6010 1845 6012
rect 1901 6010 1925 6012
rect 1981 6010 2005 6012
rect 2061 6010 2085 6012
rect 2141 6010 2147 6012
rect 1901 5958 1903 6010
rect 2083 5958 2085 6010
rect 1839 5956 1845 5958
rect 1901 5956 1925 5958
rect 1981 5956 2005 5958
rect 2061 5956 2085 5958
rect 2141 5956 2147 5958
rect 1839 5936 2147 5956
rect 2240 5710 2268 6258
rect 848 5704 900 5710
rect 848 5646 900 5652
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 570 4992 626 5001
rect 570 4927 626 4936
rect 584 4622 612 4927
rect 572 4616 624 4622
rect 572 4558 624 4564
rect 1400 4480 1452 4486
rect 1400 4422 1452 4428
rect 1412 3194 1440 4422
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 572 3052 624 3058
rect 572 2994 624 3000
rect 584 2961 612 2994
rect 570 2952 626 2961
rect 570 2887 626 2896
rect 1412 2514 1440 3130
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1504 2446 1532 5510
rect 2056 5370 2084 5646
rect 2228 5568 2280 5574
rect 2332 5522 2360 6666
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2280 5516 2360 5522
rect 2228 5510 2360 5516
rect 2240 5494 2360 5510
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 1596 5234 1900 5250
rect 1584 5228 1912 5234
rect 1636 5222 1860 5228
rect 1584 5170 1636 5176
rect 1688 4282 1716 5222
rect 1860 5170 1912 5176
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 1780 4826 1808 5102
rect 1839 4924 2147 4944
rect 1839 4922 1845 4924
rect 1901 4922 1925 4924
rect 1981 4922 2005 4924
rect 2061 4922 2085 4924
rect 2141 4922 2147 4924
rect 1901 4870 1903 4922
rect 2083 4870 2085 4922
rect 1839 4868 1845 4870
rect 1901 4868 1925 4870
rect 1981 4868 2005 4870
rect 2061 4868 2085 4870
rect 2141 4868 2147 4870
rect 1839 4848 2147 4868
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 1768 4480 1820 4486
rect 1768 4422 1820 4428
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1780 4162 1808 4422
rect 1872 4214 1900 4558
rect 1688 4146 1808 4162
rect 1860 4208 1912 4214
rect 1860 4150 1912 4156
rect 1676 4140 1808 4146
rect 1728 4134 1808 4140
rect 1676 4082 1728 4088
rect 1688 3738 1716 4082
rect 1839 3836 2147 3856
rect 1839 3834 1845 3836
rect 1901 3834 1925 3836
rect 1981 3834 2005 3836
rect 2061 3834 2085 3836
rect 2141 3834 2147 3836
rect 1901 3782 1903 3834
rect 2083 3782 2085 3834
rect 1839 3780 1845 3782
rect 1901 3780 1925 3782
rect 1981 3780 2005 3782
rect 2061 3780 2085 3782
rect 2141 3780 2147 3782
rect 1839 3760 2147 3780
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 2240 3398 2268 5494
rect 2700 5370 2728 5578
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2332 4282 2360 4626
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2792 3466 2820 6734
rect 2884 6730 2912 6938
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2976 5914 3004 6258
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 3436 5710 3464 6802
rect 3556 6556 3864 6576
rect 3556 6554 3562 6556
rect 3618 6554 3642 6556
rect 3698 6554 3722 6556
rect 3778 6554 3802 6556
rect 3858 6554 3864 6556
rect 3618 6502 3620 6554
rect 3800 6502 3802 6554
rect 3556 6500 3562 6502
rect 3618 6500 3642 6502
rect 3698 6500 3722 6502
rect 3778 6500 3802 6502
rect 3858 6500 3864 6502
rect 3556 6480 3864 6500
rect 3988 6322 4016 7485
rect 5274 7100 5582 7120
rect 5274 7098 5280 7100
rect 5336 7098 5360 7100
rect 5416 7098 5440 7100
rect 5496 7098 5520 7100
rect 5576 7098 5582 7100
rect 5336 7046 5338 7098
rect 5518 7046 5520 7098
rect 5274 7044 5280 7046
rect 5336 7044 5360 7046
rect 5416 7044 5440 7046
rect 5496 7044 5520 7046
rect 5576 7044 5582 7046
rect 5274 7024 5582 7044
rect 6748 6798 6776 7485
rect 8708 7100 9016 7120
rect 8708 7098 8714 7100
rect 8770 7098 8794 7100
rect 8850 7098 8874 7100
rect 8930 7098 8954 7100
rect 9010 7098 9016 7100
rect 8770 7046 8772 7098
rect 8952 7046 8954 7098
rect 8708 7044 8714 7046
rect 8770 7044 8794 7046
rect 8850 7044 8874 7046
rect 8930 7044 8954 7046
rect 9010 7044 9016 7046
rect 8708 7024 9016 7044
rect 7840 6928 7892 6934
rect 7840 6870 7892 6876
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2884 3942 2912 5170
rect 2976 5098 3004 5646
rect 3436 5166 3464 5646
rect 3556 5468 3864 5488
rect 3556 5466 3562 5468
rect 3618 5466 3642 5468
rect 3698 5466 3722 5468
rect 3778 5466 3802 5468
rect 3858 5466 3864 5468
rect 3618 5414 3620 5466
rect 3800 5414 3802 5466
rect 3556 5412 3562 5414
rect 3618 5412 3642 5414
rect 3698 5412 3722 5414
rect 3778 5412 3802 5414
rect 3858 5412 3864 5414
rect 3556 5392 3864 5412
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 2964 5092 3016 5098
rect 2964 5034 3016 5040
rect 3620 4826 3648 5170
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3556 4380 3864 4400
rect 3556 4378 3562 4380
rect 3618 4378 3642 4380
rect 3698 4378 3722 4380
rect 3778 4378 3802 4380
rect 3858 4378 3864 4380
rect 3618 4326 3620 4378
rect 3800 4326 3802 4378
rect 3556 4324 3562 4326
rect 3618 4324 3642 4326
rect 3698 4324 3722 4326
rect 3778 4324 3802 4326
rect 3858 4324 3864 4326
rect 3556 4304 3864 4324
rect 4080 4146 4108 4626
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 3068 3534 3096 4082
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3252 3942 3280 4014
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 4080 3602 4108 4082
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 3056 3528 3108 3534
rect 4172 3482 4200 6190
rect 4540 5914 4568 6258
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 5184 5846 5212 6734
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5274 6012 5582 6032
rect 5274 6010 5280 6012
rect 5336 6010 5360 6012
rect 5416 6010 5440 6012
rect 5496 6010 5520 6012
rect 5576 6010 5582 6012
rect 5336 5958 5338 6010
rect 5518 5958 5520 6010
rect 5274 5956 5280 5958
rect 5336 5956 5360 5958
rect 5416 5956 5440 5958
rect 5496 5956 5520 5958
rect 5576 5956 5582 5958
rect 5274 5936 5582 5956
rect 5172 5840 5224 5846
rect 5172 5782 5224 5788
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4344 5296 4396 5302
rect 4344 5238 4396 5244
rect 4356 4826 4384 5238
rect 4448 4826 4476 5646
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 5092 5370 5120 5510
rect 5080 5364 5132 5370
rect 5644 5352 5672 6258
rect 5736 6186 5764 6734
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 5724 6180 5776 6186
rect 5724 6122 5776 6128
rect 5724 5364 5776 5370
rect 5644 5324 5724 5352
rect 5080 5306 5132 5312
rect 5724 5306 5776 5312
rect 5736 5234 5764 5306
rect 5920 5234 5948 6598
rect 6564 6322 6592 6598
rect 6991 6556 7299 6576
rect 6991 6554 6997 6556
rect 7053 6554 7077 6556
rect 7133 6554 7157 6556
rect 7213 6554 7237 6556
rect 7293 6554 7299 6556
rect 7053 6502 7055 6554
rect 7235 6502 7237 6554
rect 6991 6500 6997 6502
rect 7053 6500 7077 6502
rect 7133 6500 7157 6502
rect 7213 6500 7237 6502
rect 7293 6500 7299 6502
rect 6991 6480 7299 6500
rect 7392 6458 7420 6598
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 4724 5114 4752 5170
rect 4724 5086 4936 5114
rect 4908 5030 4936 5086
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4540 4282 4568 4558
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4632 3534 4660 4082
rect 4816 4078 4844 4966
rect 5274 4924 5582 4944
rect 5274 4922 5280 4924
rect 5336 4922 5360 4924
rect 5416 4922 5440 4924
rect 5496 4922 5520 4924
rect 5576 4922 5582 4924
rect 5336 4870 5338 4922
rect 5518 4870 5520 4922
rect 5274 4868 5280 4870
rect 5336 4868 5360 4870
rect 5416 4868 5440 4870
rect 5496 4868 5520 4870
rect 5576 4868 5582 4870
rect 5274 4848 5582 4868
rect 5644 4622 5672 5170
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5080 4548 5132 4554
rect 5080 4490 5132 4496
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 3056 3470 3108 3476
rect 4080 3466 4200 3482
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 5092 3466 5120 4490
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5184 3738 5212 4082
rect 5274 3836 5582 3856
rect 5274 3834 5280 3836
rect 5336 3834 5360 3836
rect 5416 3834 5440 3836
rect 5496 3834 5520 3836
rect 5576 3834 5582 3836
rect 5336 3782 5338 3834
rect 5518 3782 5520 3834
rect 5274 3780 5280 3782
rect 5336 3780 5360 3782
rect 5416 3780 5440 3782
rect 5496 3780 5520 3782
rect 5576 3780 5582 3782
rect 5274 3760 5582 3780
rect 5644 3738 5672 4558
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5736 3534 5764 5170
rect 5920 4214 5948 5170
rect 6012 5030 6040 5646
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6472 5030 6500 5510
rect 6564 5234 6592 6258
rect 6991 5468 7299 5488
rect 6991 5466 6997 5468
rect 7053 5466 7077 5468
rect 7133 5466 7157 5468
rect 7213 5466 7237 5468
rect 7293 5466 7299 5468
rect 7053 5414 7055 5466
rect 7235 5414 7237 5466
rect 6991 5412 6997 5414
rect 7053 5412 7077 5414
rect 7133 5412 7157 5414
rect 7213 5412 7237 5414
rect 7293 5412 7299 5414
rect 6991 5392 7299 5412
rect 7392 5370 7420 6258
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7576 5710 7604 6054
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7392 5234 7420 5306
rect 7576 5234 7604 5646
rect 7748 5296 7800 5302
rect 7748 5238 7800 5244
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 5908 4208 5960 4214
rect 5908 4150 5960 4156
rect 6196 4146 6224 4422
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6012 3534 6040 4082
rect 6288 3738 6316 4966
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6564 4214 6592 4626
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6656 4078 6684 4558
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6840 4214 6868 4422
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6932 3942 6960 4558
rect 6991 4380 7299 4400
rect 6991 4378 6997 4380
rect 7053 4378 7077 4380
rect 7133 4378 7157 4380
rect 7213 4378 7237 4380
rect 7293 4378 7299 4380
rect 7053 4326 7055 4378
rect 7235 4326 7237 4378
rect 6991 4324 6997 4326
rect 7053 4324 7077 4326
rect 7133 4324 7157 4326
rect 7213 4324 7237 4326
rect 7293 4324 7299 4326
rect 6991 4304 7299 4324
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6932 3534 6960 3878
rect 7392 3534 7420 4558
rect 7760 4486 7788 5238
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 2780 3460 2832 3466
rect 2780 3402 2832 3408
rect 4068 3460 4200 3466
rect 4120 3454 4200 3460
rect 5080 3460 5132 3466
rect 4068 3402 4120 3408
rect 5080 3402 5132 3408
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 2700 3058 2728 3334
rect 2792 3210 2820 3402
rect 3556 3292 3864 3312
rect 3556 3290 3562 3292
rect 3618 3290 3642 3292
rect 3698 3290 3722 3292
rect 3778 3290 3802 3292
rect 3858 3290 3864 3292
rect 3618 3238 3620 3290
rect 3800 3238 3802 3290
rect 3556 3236 3562 3238
rect 3618 3236 3642 3238
rect 3698 3236 3722 3238
rect 3778 3236 3802 3238
rect 3858 3236 3864 3238
rect 3556 3216 3864 3236
rect 2792 3194 2912 3210
rect 2792 3188 2924 3194
rect 2792 3182 2872 3188
rect 2872 3130 2924 3136
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 1839 2748 2147 2768
rect 1839 2746 1845 2748
rect 1901 2746 1925 2748
rect 1981 2746 2005 2748
rect 2061 2746 2085 2748
rect 2141 2746 2147 2748
rect 1901 2694 1903 2746
rect 2083 2694 2085 2746
rect 1839 2692 1845 2694
rect 1901 2692 1925 2694
rect 1981 2692 2005 2694
rect 2061 2692 2085 2694
rect 2141 2692 2147 2694
rect 1839 2672 2147 2692
rect 572 2440 624 2446
rect 572 2382 624 2388
rect 1492 2440 1544 2446
rect 1492 2382 1544 2388
rect 584 1657 612 2382
rect 2700 2310 2728 2994
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3436 2514 3464 2926
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 2688 2304 2740 2310
rect 2688 2246 2740 2252
rect 1320 1800 1348 2246
rect 3556 2204 3864 2224
rect 3556 2202 3562 2204
rect 3618 2202 3642 2204
rect 3698 2202 3722 2204
rect 3778 2202 3802 2204
rect 3858 2202 3864 2204
rect 3618 2150 3620 2202
rect 3800 2150 3802 2202
rect 3556 2148 3562 2150
rect 3618 2148 3642 2150
rect 3698 2148 3722 2150
rect 3778 2148 3802 2150
rect 3858 2148 3864 2150
rect 3556 2128 3864 2148
rect 3988 1800 4016 2994
rect 5092 2446 5120 3402
rect 5736 3194 5764 3470
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5274 2748 5582 2768
rect 5274 2746 5280 2748
rect 5336 2746 5360 2748
rect 5416 2746 5440 2748
rect 5496 2746 5520 2748
rect 5576 2746 5582 2748
rect 5336 2694 5338 2746
rect 5518 2694 5520 2746
rect 5274 2692 5280 2694
rect 5336 2692 5360 2694
rect 5416 2692 5440 2694
rect 5496 2692 5520 2694
rect 5576 2692 5582 2694
rect 5274 2672 5582 2692
rect 6012 2650 6040 3470
rect 6991 3292 7299 3312
rect 6991 3290 6997 3292
rect 7053 3290 7077 3292
rect 7133 3290 7157 3292
rect 7213 3290 7237 3292
rect 7293 3290 7299 3292
rect 7053 3238 7055 3290
rect 7235 3238 7237 3290
rect 6991 3236 6997 3238
rect 7053 3236 7077 3238
rect 7133 3236 7157 3238
rect 7213 3236 7237 3238
rect 7293 3236 7299 3238
rect 6991 3216 7299 3236
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 6184 2916 6236 2922
rect 6184 2858 6236 2864
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 6196 2446 6224 2858
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 6748 1800 6776 2790
rect 6840 2582 6868 3062
rect 7392 2650 7420 3470
rect 7852 3126 7880 6870
rect 9416 6798 9444 7485
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 8220 6458 8248 6734
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8036 4214 8064 6258
rect 8312 6225 8340 6258
rect 8298 6216 8354 6225
rect 8772 6186 8800 6734
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9036 6384 9088 6390
rect 9128 6384 9180 6390
rect 9088 6344 9128 6372
rect 9036 6326 9088 6332
rect 9128 6326 9180 6332
rect 9404 6384 9456 6390
rect 9404 6326 9456 6332
rect 8852 6316 8904 6322
rect 9312 6316 9364 6322
rect 8852 6258 8904 6264
rect 9232 6276 9312 6304
rect 8864 6186 8892 6258
rect 9232 6186 9260 6276
rect 9312 6258 9364 6264
rect 8298 6151 8354 6160
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 9220 6180 9272 6186
rect 9220 6122 9272 6128
rect 8708 6012 9016 6032
rect 8708 6010 8714 6012
rect 8770 6010 8794 6012
rect 8850 6010 8874 6012
rect 8930 6010 8954 6012
rect 9010 6010 9016 6012
rect 8770 5958 8772 6010
rect 8952 5958 8954 6010
rect 8708 5956 8714 5958
rect 8770 5956 8794 5958
rect 8850 5956 8874 5958
rect 8930 5956 8954 5958
rect 9010 5956 9016 5958
rect 8708 5936 9016 5956
rect 9232 5914 9260 6122
rect 9416 5914 9444 6326
rect 9494 6216 9550 6225
rect 9494 6151 9496 6160
rect 9548 6151 9550 6160
rect 9496 6122 9548 6128
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8128 5370 8156 5646
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8496 5166 8524 5782
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8588 5234 8616 5714
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9048 5234 9076 5646
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8312 4622 8340 5102
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 8024 4208 8076 4214
rect 8024 4150 8076 4156
rect 8220 4010 8248 4490
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 6828 2576 6880 2582
rect 6828 2518 6880 2524
rect 6840 2310 6868 2518
rect 7852 2446 7880 3062
rect 8404 2514 8432 5034
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8588 4622 8616 4966
rect 8708 4924 9016 4944
rect 8708 4922 8714 4924
rect 8770 4922 8794 4924
rect 8850 4922 8874 4924
rect 8930 4922 8954 4924
rect 9010 4922 9016 4924
rect 8770 4870 8772 4922
rect 8952 4870 8954 4922
rect 8708 4868 8714 4870
rect 8770 4868 8794 4870
rect 8850 4868 8874 4870
rect 8930 4868 8954 4870
rect 9010 4868 9016 4870
rect 8708 4848 9016 4868
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8588 3534 8616 4014
rect 8708 3836 9016 3856
rect 8708 3834 8714 3836
rect 8770 3834 8794 3836
rect 8850 3834 8874 3836
rect 8930 3834 8954 3836
rect 9010 3834 9016 3836
rect 8770 3782 8772 3834
rect 8952 3782 8954 3834
rect 8708 3780 8714 3782
rect 8770 3780 8794 3782
rect 8850 3780 8874 3782
rect 8930 3780 8954 3782
rect 9010 3780 9016 3782
rect 8708 3760 9016 3780
rect 9048 3738 9076 5170
rect 9140 4622 9168 5238
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9140 3738 9168 4558
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8708 2748 9016 2768
rect 8708 2746 8714 2748
rect 8770 2746 8794 2748
rect 8850 2746 8874 2748
rect 8930 2746 8954 2748
rect 9010 2746 9016 2748
rect 8770 2694 8772 2746
rect 8952 2694 8954 2746
rect 8708 2692 8714 2694
rect 8770 2692 8794 2694
rect 8850 2692 8874 2694
rect 8930 2692 8954 2694
rect 9010 2692 9016 2694
rect 8708 2672 9016 2692
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 6991 2204 7299 2224
rect 6991 2202 6997 2204
rect 7053 2202 7077 2204
rect 7133 2202 7157 2204
rect 7213 2202 7237 2204
rect 7293 2202 7299 2204
rect 7053 2150 7055 2202
rect 7235 2150 7237 2202
rect 6991 2148 6997 2150
rect 7053 2148 7077 2150
rect 7133 2148 7157 2150
rect 7213 2148 7237 2150
rect 7293 2148 7299 2150
rect 6991 2128 7299 2148
rect 9416 1800 9444 5170
rect 9508 4826 9536 5646
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9508 2650 9536 4218
rect 9600 4078 9628 6394
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9678 4040 9734 4049
rect 9678 3975 9734 3984
rect 9692 3058 9720 3975
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9784 2650 9812 6190
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9876 3194 9904 4014
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9508 2446 9536 2586
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 570 1648 626 1657
rect 570 1583 626 1592
rect 584 1574 612 1583
rect 1306 1400 1362 1800
rect 3974 1400 4030 1800
rect 6734 1400 6790 1800
rect 9402 1400 9458 1800
<< via2 >>
rect 570 6840 626 6896
rect 1845 7098 1901 7100
rect 1925 7098 1981 7100
rect 2005 7098 2061 7100
rect 2085 7098 2141 7100
rect 1845 7046 1891 7098
rect 1891 7046 1901 7098
rect 1925 7046 1955 7098
rect 1955 7046 1967 7098
rect 1967 7046 1981 7098
rect 2005 7046 2019 7098
rect 2019 7046 2031 7098
rect 2031 7046 2061 7098
rect 2085 7046 2095 7098
rect 2095 7046 2141 7098
rect 1845 7044 1901 7046
rect 1925 7044 1981 7046
rect 2005 7044 2061 7046
rect 2085 7044 2141 7046
rect 1845 6010 1901 6012
rect 1925 6010 1981 6012
rect 2005 6010 2061 6012
rect 2085 6010 2141 6012
rect 1845 5958 1891 6010
rect 1891 5958 1901 6010
rect 1925 5958 1955 6010
rect 1955 5958 1967 6010
rect 1967 5958 1981 6010
rect 2005 5958 2019 6010
rect 2019 5958 2031 6010
rect 2031 5958 2061 6010
rect 2085 5958 2095 6010
rect 2095 5958 2141 6010
rect 1845 5956 1901 5958
rect 1925 5956 1981 5958
rect 2005 5956 2061 5958
rect 2085 5956 2141 5958
rect 570 4936 626 4992
rect 570 2896 626 2952
rect 1845 4922 1901 4924
rect 1925 4922 1981 4924
rect 2005 4922 2061 4924
rect 2085 4922 2141 4924
rect 1845 4870 1891 4922
rect 1891 4870 1901 4922
rect 1925 4870 1955 4922
rect 1955 4870 1967 4922
rect 1967 4870 1981 4922
rect 2005 4870 2019 4922
rect 2019 4870 2031 4922
rect 2031 4870 2061 4922
rect 2085 4870 2095 4922
rect 2095 4870 2141 4922
rect 1845 4868 1901 4870
rect 1925 4868 1981 4870
rect 2005 4868 2061 4870
rect 2085 4868 2141 4870
rect 1845 3834 1901 3836
rect 1925 3834 1981 3836
rect 2005 3834 2061 3836
rect 2085 3834 2141 3836
rect 1845 3782 1891 3834
rect 1891 3782 1901 3834
rect 1925 3782 1955 3834
rect 1955 3782 1967 3834
rect 1967 3782 1981 3834
rect 2005 3782 2019 3834
rect 2019 3782 2031 3834
rect 2031 3782 2061 3834
rect 2085 3782 2095 3834
rect 2095 3782 2141 3834
rect 1845 3780 1901 3782
rect 1925 3780 1981 3782
rect 2005 3780 2061 3782
rect 2085 3780 2141 3782
rect 3562 6554 3618 6556
rect 3642 6554 3698 6556
rect 3722 6554 3778 6556
rect 3802 6554 3858 6556
rect 3562 6502 3608 6554
rect 3608 6502 3618 6554
rect 3642 6502 3672 6554
rect 3672 6502 3684 6554
rect 3684 6502 3698 6554
rect 3722 6502 3736 6554
rect 3736 6502 3748 6554
rect 3748 6502 3778 6554
rect 3802 6502 3812 6554
rect 3812 6502 3858 6554
rect 3562 6500 3618 6502
rect 3642 6500 3698 6502
rect 3722 6500 3778 6502
rect 3802 6500 3858 6502
rect 5280 7098 5336 7100
rect 5360 7098 5416 7100
rect 5440 7098 5496 7100
rect 5520 7098 5576 7100
rect 5280 7046 5326 7098
rect 5326 7046 5336 7098
rect 5360 7046 5390 7098
rect 5390 7046 5402 7098
rect 5402 7046 5416 7098
rect 5440 7046 5454 7098
rect 5454 7046 5466 7098
rect 5466 7046 5496 7098
rect 5520 7046 5530 7098
rect 5530 7046 5576 7098
rect 5280 7044 5336 7046
rect 5360 7044 5416 7046
rect 5440 7044 5496 7046
rect 5520 7044 5576 7046
rect 8714 7098 8770 7100
rect 8794 7098 8850 7100
rect 8874 7098 8930 7100
rect 8954 7098 9010 7100
rect 8714 7046 8760 7098
rect 8760 7046 8770 7098
rect 8794 7046 8824 7098
rect 8824 7046 8836 7098
rect 8836 7046 8850 7098
rect 8874 7046 8888 7098
rect 8888 7046 8900 7098
rect 8900 7046 8930 7098
rect 8954 7046 8964 7098
rect 8964 7046 9010 7098
rect 8714 7044 8770 7046
rect 8794 7044 8850 7046
rect 8874 7044 8930 7046
rect 8954 7044 9010 7046
rect 3562 5466 3618 5468
rect 3642 5466 3698 5468
rect 3722 5466 3778 5468
rect 3802 5466 3858 5468
rect 3562 5414 3608 5466
rect 3608 5414 3618 5466
rect 3642 5414 3672 5466
rect 3672 5414 3684 5466
rect 3684 5414 3698 5466
rect 3722 5414 3736 5466
rect 3736 5414 3748 5466
rect 3748 5414 3778 5466
rect 3802 5414 3812 5466
rect 3812 5414 3858 5466
rect 3562 5412 3618 5414
rect 3642 5412 3698 5414
rect 3722 5412 3778 5414
rect 3802 5412 3858 5414
rect 3562 4378 3618 4380
rect 3642 4378 3698 4380
rect 3722 4378 3778 4380
rect 3802 4378 3858 4380
rect 3562 4326 3608 4378
rect 3608 4326 3618 4378
rect 3642 4326 3672 4378
rect 3672 4326 3684 4378
rect 3684 4326 3698 4378
rect 3722 4326 3736 4378
rect 3736 4326 3748 4378
rect 3748 4326 3778 4378
rect 3802 4326 3812 4378
rect 3812 4326 3858 4378
rect 3562 4324 3618 4326
rect 3642 4324 3698 4326
rect 3722 4324 3778 4326
rect 3802 4324 3858 4326
rect 5280 6010 5336 6012
rect 5360 6010 5416 6012
rect 5440 6010 5496 6012
rect 5520 6010 5576 6012
rect 5280 5958 5326 6010
rect 5326 5958 5336 6010
rect 5360 5958 5390 6010
rect 5390 5958 5402 6010
rect 5402 5958 5416 6010
rect 5440 5958 5454 6010
rect 5454 5958 5466 6010
rect 5466 5958 5496 6010
rect 5520 5958 5530 6010
rect 5530 5958 5576 6010
rect 5280 5956 5336 5958
rect 5360 5956 5416 5958
rect 5440 5956 5496 5958
rect 5520 5956 5576 5958
rect 6997 6554 7053 6556
rect 7077 6554 7133 6556
rect 7157 6554 7213 6556
rect 7237 6554 7293 6556
rect 6997 6502 7043 6554
rect 7043 6502 7053 6554
rect 7077 6502 7107 6554
rect 7107 6502 7119 6554
rect 7119 6502 7133 6554
rect 7157 6502 7171 6554
rect 7171 6502 7183 6554
rect 7183 6502 7213 6554
rect 7237 6502 7247 6554
rect 7247 6502 7293 6554
rect 6997 6500 7053 6502
rect 7077 6500 7133 6502
rect 7157 6500 7213 6502
rect 7237 6500 7293 6502
rect 5280 4922 5336 4924
rect 5360 4922 5416 4924
rect 5440 4922 5496 4924
rect 5520 4922 5576 4924
rect 5280 4870 5326 4922
rect 5326 4870 5336 4922
rect 5360 4870 5390 4922
rect 5390 4870 5402 4922
rect 5402 4870 5416 4922
rect 5440 4870 5454 4922
rect 5454 4870 5466 4922
rect 5466 4870 5496 4922
rect 5520 4870 5530 4922
rect 5530 4870 5576 4922
rect 5280 4868 5336 4870
rect 5360 4868 5416 4870
rect 5440 4868 5496 4870
rect 5520 4868 5576 4870
rect 5280 3834 5336 3836
rect 5360 3834 5416 3836
rect 5440 3834 5496 3836
rect 5520 3834 5576 3836
rect 5280 3782 5326 3834
rect 5326 3782 5336 3834
rect 5360 3782 5390 3834
rect 5390 3782 5402 3834
rect 5402 3782 5416 3834
rect 5440 3782 5454 3834
rect 5454 3782 5466 3834
rect 5466 3782 5496 3834
rect 5520 3782 5530 3834
rect 5530 3782 5576 3834
rect 5280 3780 5336 3782
rect 5360 3780 5416 3782
rect 5440 3780 5496 3782
rect 5520 3780 5576 3782
rect 6997 5466 7053 5468
rect 7077 5466 7133 5468
rect 7157 5466 7213 5468
rect 7237 5466 7293 5468
rect 6997 5414 7043 5466
rect 7043 5414 7053 5466
rect 7077 5414 7107 5466
rect 7107 5414 7119 5466
rect 7119 5414 7133 5466
rect 7157 5414 7171 5466
rect 7171 5414 7183 5466
rect 7183 5414 7213 5466
rect 7237 5414 7247 5466
rect 7247 5414 7293 5466
rect 6997 5412 7053 5414
rect 7077 5412 7133 5414
rect 7157 5412 7213 5414
rect 7237 5412 7293 5414
rect 6997 4378 7053 4380
rect 7077 4378 7133 4380
rect 7157 4378 7213 4380
rect 7237 4378 7293 4380
rect 6997 4326 7043 4378
rect 7043 4326 7053 4378
rect 7077 4326 7107 4378
rect 7107 4326 7119 4378
rect 7119 4326 7133 4378
rect 7157 4326 7171 4378
rect 7171 4326 7183 4378
rect 7183 4326 7213 4378
rect 7237 4326 7247 4378
rect 7247 4326 7293 4378
rect 6997 4324 7053 4326
rect 7077 4324 7133 4326
rect 7157 4324 7213 4326
rect 7237 4324 7293 4326
rect 3562 3290 3618 3292
rect 3642 3290 3698 3292
rect 3722 3290 3778 3292
rect 3802 3290 3858 3292
rect 3562 3238 3608 3290
rect 3608 3238 3618 3290
rect 3642 3238 3672 3290
rect 3672 3238 3684 3290
rect 3684 3238 3698 3290
rect 3722 3238 3736 3290
rect 3736 3238 3748 3290
rect 3748 3238 3778 3290
rect 3802 3238 3812 3290
rect 3812 3238 3858 3290
rect 3562 3236 3618 3238
rect 3642 3236 3698 3238
rect 3722 3236 3778 3238
rect 3802 3236 3858 3238
rect 1845 2746 1901 2748
rect 1925 2746 1981 2748
rect 2005 2746 2061 2748
rect 2085 2746 2141 2748
rect 1845 2694 1891 2746
rect 1891 2694 1901 2746
rect 1925 2694 1955 2746
rect 1955 2694 1967 2746
rect 1967 2694 1981 2746
rect 2005 2694 2019 2746
rect 2019 2694 2031 2746
rect 2031 2694 2061 2746
rect 2085 2694 2095 2746
rect 2095 2694 2141 2746
rect 1845 2692 1901 2694
rect 1925 2692 1981 2694
rect 2005 2692 2061 2694
rect 2085 2692 2141 2694
rect 3562 2202 3618 2204
rect 3642 2202 3698 2204
rect 3722 2202 3778 2204
rect 3802 2202 3858 2204
rect 3562 2150 3608 2202
rect 3608 2150 3618 2202
rect 3642 2150 3672 2202
rect 3672 2150 3684 2202
rect 3684 2150 3698 2202
rect 3722 2150 3736 2202
rect 3736 2150 3748 2202
rect 3748 2150 3778 2202
rect 3802 2150 3812 2202
rect 3812 2150 3858 2202
rect 3562 2148 3618 2150
rect 3642 2148 3698 2150
rect 3722 2148 3778 2150
rect 3802 2148 3858 2150
rect 5280 2746 5336 2748
rect 5360 2746 5416 2748
rect 5440 2746 5496 2748
rect 5520 2746 5576 2748
rect 5280 2694 5326 2746
rect 5326 2694 5336 2746
rect 5360 2694 5390 2746
rect 5390 2694 5402 2746
rect 5402 2694 5416 2746
rect 5440 2694 5454 2746
rect 5454 2694 5466 2746
rect 5466 2694 5496 2746
rect 5520 2694 5530 2746
rect 5530 2694 5576 2746
rect 5280 2692 5336 2694
rect 5360 2692 5416 2694
rect 5440 2692 5496 2694
rect 5520 2692 5576 2694
rect 6997 3290 7053 3292
rect 7077 3290 7133 3292
rect 7157 3290 7213 3292
rect 7237 3290 7293 3292
rect 6997 3238 7043 3290
rect 7043 3238 7053 3290
rect 7077 3238 7107 3290
rect 7107 3238 7119 3290
rect 7119 3238 7133 3290
rect 7157 3238 7171 3290
rect 7171 3238 7183 3290
rect 7183 3238 7213 3290
rect 7237 3238 7247 3290
rect 7247 3238 7293 3290
rect 6997 3236 7053 3238
rect 7077 3236 7133 3238
rect 7157 3236 7213 3238
rect 7237 3236 7293 3238
rect 8298 6160 8354 6216
rect 8714 6010 8770 6012
rect 8794 6010 8850 6012
rect 8874 6010 8930 6012
rect 8954 6010 9010 6012
rect 8714 5958 8760 6010
rect 8760 5958 8770 6010
rect 8794 5958 8824 6010
rect 8824 5958 8836 6010
rect 8836 5958 8850 6010
rect 8874 5958 8888 6010
rect 8888 5958 8900 6010
rect 8900 5958 8930 6010
rect 8954 5958 8964 6010
rect 8964 5958 9010 6010
rect 8714 5956 8770 5958
rect 8794 5956 8850 5958
rect 8874 5956 8930 5958
rect 8954 5956 9010 5958
rect 9494 6180 9550 6216
rect 9494 6160 9496 6180
rect 9496 6160 9548 6180
rect 9548 6160 9550 6180
rect 8714 4922 8770 4924
rect 8794 4922 8850 4924
rect 8874 4922 8930 4924
rect 8954 4922 9010 4924
rect 8714 4870 8760 4922
rect 8760 4870 8770 4922
rect 8794 4870 8824 4922
rect 8824 4870 8836 4922
rect 8836 4870 8850 4922
rect 8874 4870 8888 4922
rect 8888 4870 8900 4922
rect 8900 4870 8930 4922
rect 8954 4870 8964 4922
rect 8964 4870 9010 4922
rect 8714 4868 8770 4870
rect 8794 4868 8850 4870
rect 8874 4868 8930 4870
rect 8954 4868 9010 4870
rect 8714 3834 8770 3836
rect 8794 3834 8850 3836
rect 8874 3834 8930 3836
rect 8954 3834 9010 3836
rect 8714 3782 8760 3834
rect 8760 3782 8770 3834
rect 8794 3782 8824 3834
rect 8824 3782 8836 3834
rect 8836 3782 8850 3834
rect 8874 3782 8888 3834
rect 8888 3782 8900 3834
rect 8900 3782 8930 3834
rect 8954 3782 8964 3834
rect 8964 3782 9010 3834
rect 8714 3780 8770 3782
rect 8794 3780 8850 3782
rect 8874 3780 8930 3782
rect 8954 3780 9010 3782
rect 8714 2746 8770 2748
rect 8794 2746 8850 2748
rect 8874 2746 8930 2748
rect 8954 2746 9010 2748
rect 8714 2694 8760 2746
rect 8760 2694 8770 2746
rect 8794 2694 8824 2746
rect 8824 2694 8836 2746
rect 8836 2694 8850 2746
rect 8874 2694 8888 2746
rect 8888 2694 8900 2746
rect 8900 2694 8930 2746
rect 8954 2694 8964 2746
rect 8964 2694 9010 2746
rect 8714 2692 8770 2694
rect 8794 2692 8850 2694
rect 8874 2692 8930 2694
rect 8954 2692 9010 2694
rect 6997 2202 7053 2204
rect 7077 2202 7133 2204
rect 7157 2202 7213 2204
rect 7237 2202 7293 2204
rect 6997 2150 7043 2202
rect 7043 2150 7053 2202
rect 7077 2150 7107 2202
rect 7107 2150 7119 2202
rect 7119 2150 7133 2202
rect 7157 2150 7171 2202
rect 7171 2150 7183 2202
rect 7183 2150 7213 2202
rect 7237 2150 7247 2202
rect 7247 2150 7293 2202
rect 6997 2148 7053 2150
rect 7077 2148 7133 2150
rect 7157 2148 7213 2150
rect 7237 2148 7293 2150
rect 9678 3984 9734 4040
rect 570 1592 626 1648
<< metal3 >>
rect 1833 7104 2153 7105
rect 1833 7040 1841 7104
rect 1905 7040 1921 7104
rect 1985 7040 2001 7104
rect 2065 7040 2081 7104
rect 2145 7040 2153 7104
rect 1833 7039 2153 7040
rect 5268 7104 5588 7105
rect 5268 7040 5276 7104
rect 5340 7040 5356 7104
rect 5420 7040 5436 7104
rect 5500 7040 5516 7104
rect 5580 7040 5588 7104
rect 5268 7039 5588 7040
rect 8702 7104 9022 7105
rect 8702 7040 8710 7104
rect 8774 7040 8790 7104
rect 8854 7040 8870 7104
rect 8934 7040 8950 7104
rect 9014 7040 9022 7104
rect 8702 7039 9022 7040
rect 0 6898 400 6928
rect 565 6898 631 6901
rect 0 6896 631 6898
rect 0 6840 570 6896
rect 626 6840 631 6896
rect 0 6838 631 6840
rect 0 6808 400 6838
rect 565 6835 631 6838
rect 3550 6560 3870 6561
rect 3550 6496 3558 6560
rect 3622 6496 3638 6560
rect 3702 6496 3718 6560
rect 3782 6496 3798 6560
rect 3862 6496 3870 6560
rect 3550 6495 3870 6496
rect 6985 6560 7305 6561
rect 6985 6496 6993 6560
rect 7057 6496 7073 6560
rect 7137 6496 7153 6560
rect 7217 6496 7233 6560
rect 7297 6496 7305 6560
rect 6985 6495 7305 6496
rect 8293 6218 8359 6221
rect 9489 6218 9555 6221
rect 8293 6216 9555 6218
rect 8293 6160 8298 6216
rect 8354 6160 9494 6216
rect 9550 6160 9555 6216
rect 8293 6158 9555 6160
rect 8293 6155 8359 6158
rect 9489 6155 9555 6158
rect 1833 6016 2153 6017
rect 1833 5952 1841 6016
rect 1905 5952 1921 6016
rect 1985 5952 2001 6016
rect 2065 5952 2081 6016
rect 2145 5952 2153 6016
rect 1833 5951 2153 5952
rect 5268 6016 5588 6017
rect 5268 5952 5276 6016
rect 5340 5952 5356 6016
rect 5420 5952 5436 6016
rect 5500 5952 5516 6016
rect 5580 5952 5588 6016
rect 5268 5951 5588 5952
rect 8702 6016 9022 6017
rect 8702 5952 8710 6016
rect 8774 5952 8790 6016
rect 8854 5952 8870 6016
rect 8934 5952 8950 6016
rect 9014 5952 9022 6016
rect 8702 5951 9022 5952
rect 3550 5472 3870 5473
rect 3550 5408 3558 5472
rect 3622 5408 3638 5472
rect 3702 5408 3718 5472
rect 3782 5408 3798 5472
rect 3862 5408 3870 5472
rect 3550 5407 3870 5408
rect 6985 5472 7305 5473
rect 6985 5408 6993 5472
rect 7057 5408 7073 5472
rect 7137 5408 7153 5472
rect 7217 5408 7233 5472
rect 7297 5408 7305 5472
rect 6985 5407 7305 5408
rect 0 4994 400 5024
rect 565 4994 631 4997
rect 0 4992 631 4994
rect 0 4936 570 4992
rect 626 4936 631 4992
rect 0 4934 631 4936
rect 0 4904 400 4934
rect 565 4931 631 4934
rect 1833 4928 2153 4929
rect 1833 4864 1841 4928
rect 1905 4864 1921 4928
rect 1985 4864 2001 4928
rect 2065 4864 2081 4928
rect 2145 4864 2153 4928
rect 1833 4863 2153 4864
rect 5268 4928 5588 4929
rect 5268 4864 5276 4928
rect 5340 4864 5356 4928
rect 5420 4864 5436 4928
rect 5500 4864 5516 4928
rect 5580 4864 5588 4928
rect 5268 4863 5588 4864
rect 8702 4928 9022 4929
rect 8702 4864 8710 4928
rect 8774 4864 8790 4928
rect 8854 4864 8870 4928
rect 8934 4864 8950 4928
rect 9014 4864 9022 4928
rect 8702 4863 9022 4864
rect 3550 4384 3870 4385
rect 3550 4320 3558 4384
rect 3622 4320 3638 4384
rect 3702 4320 3718 4384
rect 3782 4320 3798 4384
rect 3862 4320 3870 4384
rect 3550 4319 3870 4320
rect 6985 4384 7305 4385
rect 6985 4320 6993 4384
rect 7057 4320 7073 4384
rect 7137 4320 7153 4384
rect 7217 4320 7233 4384
rect 7297 4320 7305 4384
rect 6985 4319 7305 4320
rect 9673 4042 9739 4045
rect 10482 4042 10882 4072
rect 9673 4040 10882 4042
rect 9673 3984 9678 4040
rect 9734 3984 10882 4040
rect 9673 3982 10882 3984
rect 9673 3979 9739 3982
rect 10482 3952 10882 3982
rect 1833 3840 2153 3841
rect 1833 3776 1841 3840
rect 1905 3776 1921 3840
rect 1985 3776 2001 3840
rect 2065 3776 2081 3840
rect 2145 3776 2153 3840
rect 1833 3775 2153 3776
rect 5268 3840 5588 3841
rect 5268 3776 5276 3840
rect 5340 3776 5356 3840
rect 5420 3776 5436 3840
rect 5500 3776 5516 3840
rect 5580 3776 5588 3840
rect 5268 3775 5588 3776
rect 8702 3840 9022 3841
rect 8702 3776 8710 3840
rect 8774 3776 8790 3840
rect 8854 3776 8870 3840
rect 8934 3776 8950 3840
rect 9014 3776 9022 3840
rect 8702 3775 9022 3776
rect 3550 3296 3870 3297
rect 3550 3232 3558 3296
rect 3622 3232 3638 3296
rect 3702 3232 3718 3296
rect 3782 3232 3798 3296
rect 3862 3232 3870 3296
rect 3550 3231 3870 3232
rect 6985 3296 7305 3297
rect 6985 3232 6993 3296
rect 7057 3232 7073 3296
rect 7137 3232 7153 3296
rect 7217 3232 7233 3296
rect 7297 3232 7305 3296
rect 6985 3231 7305 3232
rect 0 2954 400 2984
rect 565 2954 631 2957
rect 0 2952 631 2954
rect 0 2896 570 2952
rect 626 2896 631 2952
rect 0 2894 631 2896
rect 0 2864 400 2894
rect 565 2891 631 2894
rect 1833 2752 2153 2753
rect 1833 2688 1841 2752
rect 1905 2688 1921 2752
rect 1985 2688 2001 2752
rect 2065 2688 2081 2752
rect 2145 2688 2153 2752
rect 1833 2687 2153 2688
rect 5268 2752 5588 2753
rect 5268 2688 5276 2752
rect 5340 2688 5356 2752
rect 5420 2688 5436 2752
rect 5500 2688 5516 2752
rect 5580 2688 5588 2752
rect 5268 2687 5588 2688
rect 8702 2752 9022 2753
rect 8702 2688 8710 2752
rect 8774 2688 8790 2752
rect 8854 2688 8870 2752
rect 8934 2688 8950 2752
rect 9014 2688 9022 2752
rect 8702 2687 9022 2688
rect 3550 2208 3870 2209
rect 3550 2144 3558 2208
rect 3622 2144 3638 2208
rect 3702 2144 3718 2208
rect 3782 2144 3798 2208
rect 3862 2144 3870 2208
rect 3550 2143 3870 2144
rect 6985 2208 7305 2209
rect 6985 2144 6993 2208
rect 7057 2144 7073 2208
rect 7137 2144 7153 2208
rect 7217 2144 7233 2208
rect 7297 2144 7305 2208
rect 6985 2143 7305 2144
rect 0 1650 400 1680
rect 565 1650 631 1653
rect 0 1648 631 1650
rect 0 1592 570 1648
rect 626 1592 631 1648
rect 0 1590 631 1592
rect 0 1560 400 1590
rect 565 1587 631 1590
<< via3 >>
rect 1841 7100 1905 7104
rect 1841 7044 1845 7100
rect 1845 7044 1901 7100
rect 1901 7044 1905 7100
rect 1841 7040 1905 7044
rect 1921 7100 1985 7104
rect 1921 7044 1925 7100
rect 1925 7044 1981 7100
rect 1981 7044 1985 7100
rect 1921 7040 1985 7044
rect 2001 7100 2065 7104
rect 2001 7044 2005 7100
rect 2005 7044 2061 7100
rect 2061 7044 2065 7100
rect 2001 7040 2065 7044
rect 2081 7100 2145 7104
rect 2081 7044 2085 7100
rect 2085 7044 2141 7100
rect 2141 7044 2145 7100
rect 2081 7040 2145 7044
rect 5276 7100 5340 7104
rect 5276 7044 5280 7100
rect 5280 7044 5336 7100
rect 5336 7044 5340 7100
rect 5276 7040 5340 7044
rect 5356 7100 5420 7104
rect 5356 7044 5360 7100
rect 5360 7044 5416 7100
rect 5416 7044 5420 7100
rect 5356 7040 5420 7044
rect 5436 7100 5500 7104
rect 5436 7044 5440 7100
rect 5440 7044 5496 7100
rect 5496 7044 5500 7100
rect 5436 7040 5500 7044
rect 5516 7100 5580 7104
rect 5516 7044 5520 7100
rect 5520 7044 5576 7100
rect 5576 7044 5580 7100
rect 5516 7040 5580 7044
rect 8710 7100 8774 7104
rect 8710 7044 8714 7100
rect 8714 7044 8770 7100
rect 8770 7044 8774 7100
rect 8710 7040 8774 7044
rect 8790 7100 8854 7104
rect 8790 7044 8794 7100
rect 8794 7044 8850 7100
rect 8850 7044 8854 7100
rect 8790 7040 8854 7044
rect 8870 7100 8934 7104
rect 8870 7044 8874 7100
rect 8874 7044 8930 7100
rect 8930 7044 8934 7100
rect 8870 7040 8934 7044
rect 8950 7100 9014 7104
rect 8950 7044 8954 7100
rect 8954 7044 9010 7100
rect 9010 7044 9014 7100
rect 8950 7040 9014 7044
rect 3558 6556 3622 6560
rect 3558 6500 3562 6556
rect 3562 6500 3618 6556
rect 3618 6500 3622 6556
rect 3558 6496 3622 6500
rect 3638 6556 3702 6560
rect 3638 6500 3642 6556
rect 3642 6500 3698 6556
rect 3698 6500 3702 6556
rect 3638 6496 3702 6500
rect 3718 6556 3782 6560
rect 3718 6500 3722 6556
rect 3722 6500 3778 6556
rect 3778 6500 3782 6556
rect 3718 6496 3782 6500
rect 3798 6556 3862 6560
rect 3798 6500 3802 6556
rect 3802 6500 3858 6556
rect 3858 6500 3862 6556
rect 3798 6496 3862 6500
rect 6993 6556 7057 6560
rect 6993 6500 6997 6556
rect 6997 6500 7053 6556
rect 7053 6500 7057 6556
rect 6993 6496 7057 6500
rect 7073 6556 7137 6560
rect 7073 6500 7077 6556
rect 7077 6500 7133 6556
rect 7133 6500 7137 6556
rect 7073 6496 7137 6500
rect 7153 6556 7217 6560
rect 7153 6500 7157 6556
rect 7157 6500 7213 6556
rect 7213 6500 7217 6556
rect 7153 6496 7217 6500
rect 7233 6556 7297 6560
rect 7233 6500 7237 6556
rect 7237 6500 7293 6556
rect 7293 6500 7297 6556
rect 7233 6496 7297 6500
rect 1841 6012 1905 6016
rect 1841 5956 1845 6012
rect 1845 5956 1901 6012
rect 1901 5956 1905 6012
rect 1841 5952 1905 5956
rect 1921 6012 1985 6016
rect 1921 5956 1925 6012
rect 1925 5956 1981 6012
rect 1981 5956 1985 6012
rect 1921 5952 1985 5956
rect 2001 6012 2065 6016
rect 2001 5956 2005 6012
rect 2005 5956 2061 6012
rect 2061 5956 2065 6012
rect 2001 5952 2065 5956
rect 2081 6012 2145 6016
rect 2081 5956 2085 6012
rect 2085 5956 2141 6012
rect 2141 5956 2145 6012
rect 2081 5952 2145 5956
rect 5276 6012 5340 6016
rect 5276 5956 5280 6012
rect 5280 5956 5336 6012
rect 5336 5956 5340 6012
rect 5276 5952 5340 5956
rect 5356 6012 5420 6016
rect 5356 5956 5360 6012
rect 5360 5956 5416 6012
rect 5416 5956 5420 6012
rect 5356 5952 5420 5956
rect 5436 6012 5500 6016
rect 5436 5956 5440 6012
rect 5440 5956 5496 6012
rect 5496 5956 5500 6012
rect 5436 5952 5500 5956
rect 5516 6012 5580 6016
rect 5516 5956 5520 6012
rect 5520 5956 5576 6012
rect 5576 5956 5580 6012
rect 5516 5952 5580 5956
rect 8710 6012 8774 6016
rect 8710 5956 8714 6012
rect 8714 5956 8770 6012
rect 8770 5956 8774 6012
rect 8710 5952 8774 5956
rect 8790 6012 8854 6016
rect 8790 5956 8794 6012
rect 8794 5956 8850 6012
rect 8850 5956 8854 6012
rect 8790 5952 8854 5956
rect 8870 6012 8934 6016
rect 8870 5956 8874 6012
rect 8874 5956 8930 6012
rect 8930 5956 8934 6012
rect 8870 5952 8934 5956
rect 8950 6012 9014 6016
rect 8950 5956 8954 6012
rect 8954 5956 9010 6012
rect 9010 5956 9014 6012
rect 8950 5952 9014 5956
rect 3558 5468 3622 5472
rect 3558 5412 3562 5468
rect 3562 5412 3618 5468
rect 3618 5412 3622 5468
rect 3558 5408 3622 5412
rect 3638 5468 3702 5472
rect 3638 5412 3642 5468
rect 3642 5412 3698 5468
rect 3698 5412 3702 5468
rect 3638 5408 3702 5412
rect 3718 5468 3782 5472
rect 3718 5412 3722 5468
rect 3722 5412 3778 5468
rect 3778 5412 3782 5468
rect 3718 5408 3782 5412
rect 3798 5468 3862 5472
rect 3798 5412 3802 5468
rect 3802 5412 3858 5468
rect 3858 5412 3862 5468
rect 3798 5408 3862 5412
rect 6993 5468 7057 5472
rect 6993 5412 6997 5468
rect 6997 5412 7053 5468
rect 7053 5412 7057 5468
rect 6993 5408 7057 5412
rect 7073 5468 7137 5472
rect 7073 5412 7077 5468
rect 7077 5412 7133 5468
rect 7133 5412 7137 5468
rect 7073 5408 7137 5412
rect 7153 5468 7217 5472
rect 7153 5412 7157 5468
rect 7157 5412 7213 5468
rect 7213 5412 7217 5468
rect 7153 5408 7217 5412
rect 7233 5468 7297 5472
rect 7233 5412 7237 5468
rect 7237 5412 7293 5468
rect 7293 5412 7297 5468
rect 7233 5408 7297 5412
rect 1841 4924 1905 4928
rect 1841 4868 1845 4924
rect 1845 4868 1901 4924
rect 1901 4868 1905 4924
rect 1841 4864 1905 4868
rect 1921 4924 1985 4928
rect 1921 4868 1925 4924
rect 1925 4868 1981 4924
rect 1981 4868 1985 4924
rect 1921 4864 1985 4868
rect 2001 4924 2065 4928
rect 2001 4868 2005 4924
rect 2005 4868 2061 4924
rect 2061 4868 2065 4924
rect 2001 4864 2065 4868
rect 2081 4924 2145 4928
rect 2081 4868 2085 4924
rect 2085 4868 2141 4924
rect 2141 4868 2145 4924
rect 2081 4864 2145 4868
rect 5276 4924 5340 4928
rect 5276 4868 5280 4924
rect 5280 4868 5336 4924
rect 5336 4868 5340 4924
rect 5276 4864 5340 4868
rect 5356 4924 5420 4928
rect 5356 4868 5360 4924
rect 5360 4868 5416 4924
rect 5416 4868 5420 4924
rect 5356 4864 5420 4868
rect 5436 4924 5500 4928
rect 5436 4868 5440 4924
rect 5440 4868 5496 4924
rect 5496 4868 5500 4924
rect 5436 4864 5500 4868
rect 5516 4924 5580 4928
rect 5516 4868 5520 4924
rect 5520 4868 5576 4924
rect 5576 4868 5580 4924
rect 5516 4864 5580 4868
rect 8710 4924 8774 4928
rect 8710 4868 8714 4924
rect 8714 4868 8770 4924
rect 8770 4868 8774 4924
rect 8710 4864 8774 4868
rect 8790 4924 8854 4928
rect 8790 4868 8794 4924
rect 8794 4868 8850 4924
rect 8850 4868 8854 4924
rect 8790 4864 8854 4868
rect 8870 4924 8934 4928
rect 8870 4868 8874 4924
rect 8874 4868 8930 4924
rect 8930 4868 8934 4924
rect 8870 4864 8934 4868
rect 8950 4924 9014 4928
rect 8950 4868 8954 4924
rect 8954 4868 9010 4924
rect 9010 4868 9014 4924
rect 8950 4864 9014 4868
rect 3558 4380 3622 4384
rect 3558 4324 3562 4380
rect 3562 4324 3618 4380
rect 3618 4324 3622 4380
rect 3558 4320 3622 4324
rect 3638 4380 3702 4384
rect 3638 4324 3642 4380
rect 3642 4324 3698 4380
rect 3698 4324 3702 4380
rect 3638 4320 3702 4324
rect 3718 4380 3782 4384
rect 3718 4324 3722 4380
rect 3722 4324 3778 4380
rect 3778 4324 3782 4380
rect 3718 4320 3782 4324
rect 3798 4380 3862 4384
rect 3798 4324 3802 4380
rect 3802 4324 3858 4380
rect 3858 4324 3862 4380
rect 3798 4320 3862 4324
rect 6993 4380 7057 4384
rect 6993 4324 6997 4380
rect 6997 4324 7053 4380
rect 7053 4324 7057 4380
rect 6993 4320 7057 4324
rect 7073 4380 7137 4384
rect 7073 4324 7077 4380
rect 7077 4324 7133 4380
rect 7133 4324 7137 4380
rect 7073 4320 7137 4324
rect 7153 4380 7217 4384
rect 7153 4324 7157 4380
rect 7157 4324 7213 4380
rect 7213 4324 7217 4380
rect 7153 4320 7217 4324
rect 7233 4380 7297 4384
rect 7233 4324 7237 4380
rect 7237 4324 7293 4380
rect 7293 4324 7297 4380
rect 7233 4320 7297 4324
rect 1841 3836 1905 3840
rect 1841 3780 1845 3836
rect 1845 3780 1901 3836
rect 1901 3780 1905 3836
rect 1841 3776 1905 3780
rect 1921 3836 1985 3840
rect 1921 3780 1925 3836
rect 1925 3780 1981 3836
rect 1981 3780 1985 3836
rect 1921 3776 1985 3780
rect 2001 3836 2065 3840
rect 2001 3780 2005 3836
rect 2005 3780 2061 3836
rect 2061 3780 2065 3836
rect 2001 3776 2065 3780
rect 2081 3836 2145 3840
rect 2081 3780 2085 3836
rect 2085 3780 2141 3836
rect 2141 3780 2145 3836
rect 2081 3776 2145 3780
rect 5276 3836 5340 3840
rect 5276 3780 5280 3836
rect 5280 3780 5336 3836
rect 5336 3780 5340 3836
rect 5276 3776 5340 3780
rect 5356 3836 5420 3840
rect 5356 3780 5360 3836
rect 5360 3780 5416 3836
rect 5416 3780 5420 3836
rect 5356 3776 5420 3780
rect 5436 3836 5500 3840
rect 5436 3780 5440 3836
rect 5440 3780 5496 3836
rect 5496 3780 5500 3836
rect 5436 3776 5500 3780
rect 5516 3836 5580 3840
rect 5516 3780 5520 3836
rect 5520 3780 5576 3836
rect 5576 3780 5580 3836
rect 5516 3776 5580 3780
rect 8710 3836 8774 3840
rect 8710 3780 8714 3836
rect 8714 3780 8770 3836
rect 8770 3780 8774 3836
rect 8710 3776 8774 3780
rect 8790 3836 8854 3840
rect 8790 3780 8794 3836
rect 8794 3780 8850 3836
rect 8850 3780 8854 3836
rect 8790 3776 8854 3780
rect 8870 3836 8934 3840
rect 8870 3780 8874 3836
rect 8874 3780 8930 3836
rect 8930 3780 8934 3836
rect 8870 3776 8934 3780
rect 8950 3836 9014 3840
rect 8950 3780 8954 3836
rect 8954 3780 9010 3836
rect 9010 3780 9014 3836
rect 8950 3776 9014 3780
rect 3558 3292 3622 3296
rect 3558 3236 3562 3292
rect 3562 3236 3618 3292
rect 3618 3236 3622 3292
rect 3558 3232 3622 3236
rect 3638 3292 3702 3296
rect 3638 3236 3642 3292
rect 3642 3236 3698 3292
rect 3698 3236 3702 3292
rect 3638 3232 3702 3236
rect 3718 3292 3782 3296
rect 3718 3236 3722 3292
rect 3722 3236 3778 3292
rect 3778 3236 3782 3292
rect 3718 3232 3782 3236
rect 3798 3292 3862 3296
rect 3798 3236 3802 3292
rect 3802 3236 3858 3292
rect 3858 3236 3862 3292
rect 3798 3232 3862 3236
rect 6993 3292 7057 3296
rect 6993 3236 6997 3292
rect 6997 3236 7053 3292
rect 7053 3236 7057 3292
rect 6993 3232 7057 3236
rect 7073 3292 7137 3296
rect 7073 3236 7077 3292
rect 7077 3236 7133 3292
rect 7133 3236 7137 3292
rect 7073 3232 7137 3236
rect 7153 3292 7217 3296
rect 7153 3236 7157 3292
rect 7157 3236 7213 3292
rect 7213 3236 7217 3292
rect 7153 3232 7217 3236
rect 7233 3292 7297 3296
rect 7233 3236 7237 3292
rect 7237 3236 7293 3292
rect 7293 3236 7297 3292
rect 7233 3232 7297 3236
rect 1841 2748 1905 2752
rect 1841 2692 1845 2748
rect 1845 2692 1901 2748
rect 1901 2692 1905 2748
rect 1841 2688 1905 2692
rect 1921 2748 1985 2752
rect 1921 2692 1925 2748
rect 1925 2692 1981 2748
rect 1981 2692 1985 2748
rect 1921 2688 1985 2692
rect 2001 2748 2065 2752
rect 2001 2692 2005 2748
rect 2005 2692 2061 2748
rect 2061 2692 2065 2748
rect 2001 2688 2065 2692
rect 2081 2748 2145 2752
rect 2081 2692 2085 2748
rect 2085 2692 2141 2748
rect 2141 2692 2145 2748
rect 2081 2688 2145 2692
rect 5276 2748 5340 2752
rect 5276 2692 5280 2748
rect 5280 2692 5336 2748
rect 5336 2692 5340 2748
rect 5276 2688 5340 2692
rect 5356 2748 5420 2752
rect 5356 2692 5360 2748
rect 5360 2692 5416 2748
rect 5416 2692 5420 2748
rect 5356 2688 5420 2692
rect 5436 2748 5500 2752
rect 5436 2692 5440 2748
rect 5440 2692 5496 2748
rect 5496 2692 5500 2748
rect 5436 2688 5500 2692
rect 5516 2748 5580 2752
rect 5516 2692 5520 2748
rect 5520 2692 5576 2748
rect 5576 2692 5580 2748
rect 5516 2688 5580 2692
rect 8710 2748 8774 2752
rect 8710 2692 8714 2748
rect 8714 2692 8770 2748
rect 8770 2692 8774 2748
rect 8710 2688 8774 2692
rect 8790 2748 8854 2752
rect 8790 2692 8794 2748
rect 8794 2692 8850 2748
rect 8850 2692 8854 2748
rect 8790 2688 8854 2692
rect 8870 2748 8934 2752
rect 8870 2692 8874 2748
rect 8874 2692 8930 2748
rect 8930 2692 8934 2748
rect 8870 2688 8934 2692
rect 8950 2748 9014 2752
rect 8950 2692 8954 2748
rect 8954 2692 9010 2748
rect 9010 2692 9014 2748
rect 8950 2688 9014 2692
rect 3558 2204 3622 2208
rect 3558 2148 3562 2204
rect 3562 2148 3618 2204
rect 3618 2148 3622 2204
rect 3558 2144 3622 2148
rect 3638 2204 3702 2208
rect 3638 2148 3642 2204
rect 3642 2148 3698 2204
rect 3698 2148 3702 2204
rect 3638 2144 3702 2148
rect 3718 2204 3782 2208
rect 3718 2148 3722 2204
rect 3722 2148 3778 2204
rect 3778 2148 3782 2204
rect 3718 2144 3782 2148
rect 3798 2204 3862 2208
rect 3798 2148 3802 2204
rect 3802 2148 3858 2204
rect 3858 2148 3862 2204
rect 3798 2144 3862 2148
rect 6993 2204 7057 2208
rect 6993 2148 6997 2204
rect 6997 2148 7053 2204
rect 7053 2148 7057 2204
rect 6993 2144 7057 2148
rect 7073 2204 7137 2208
rect 7073 2148 7077 2204
rect 7077 2148 7133 2204
rect 7133 2148 7137 2204
rect 7073 2144 7137 2148
rect 7153 2204 7217 2208
rect 7153 2148 7157 2204
rect 7157 2148 7213 2204
rect 7213 2148 7217 2204
rect 7153 2144 7217 2148
rect 7233 2204 7297 2208
rect 7233 2148 7237 2204
rect 7237 2148 7293 2204
rect 7293 2148 7297 2204
rect 7233 2144 7297 2148
<< metal4 >>
rect 1833 7104 2154 7120
rect 1833 7040 1841 7104
rect 1905 7040 1921 7104
rect 1985 7040 2001 7104
rect 2065 7040 2081 7104
rect 2145 7040 2154 7104
rect 1833 6016 2154 7040
rect 1833 5952 1841 6016
rect 1905 5952 1921 6016
rect 1985 5952 2001 6016
rect 2065 5952 2081 6016
rect 2145 5952 2154 6016
rect 1833 4928 2154 5952
rect 1833 4864 1841 4928
rect 1905 4864 1921 4928
rect 1985 4864 2001 4928
rect 2065 4864 2081 4928
rect 2145 4864 2154 4928
rect 1833 3840 2154 4864
rect 1833 3776 1841 3840
rect 1905 3776 1921 3840
rect 1985 3776 2001 3840
rect 2065 3776 2081 3840
rect 2145 3776 2154 3840
rect 1833 2752 2154 3776
rect 1833 2688 1841 2752
rect 1905 2688 1921 2752
rect 1985 2688 2001 2752
rect 2065 2688 2081 2752
rect 2145 2688 2154 2752
rect 1833 2128 2154 2688
rect 3550 6560 3870 7120
rect 3550 6496 3558 6560
rect 3622 6496 3638 6560
rect 3702 6496 3718 6560
rect 3782 6496 3798 6560
rect 3862 6496 3870 6560
rect 3550 5472 3870 6496
rect 3550 5408 3558 5472
rect 3622 5408 3638 5472
rect 3702 5408 3718 5472
rect 3782 5408 3798 5472
rect 3862 5408 3870 5472
rect 3550 4384 3870 5408
rect 3550 4320 3558 4384
rect 3622 4320 3638 4384
rect 3702 4320 3718 4384
rect 3782 4320 3798 4384
rect 3862 4320 3870 4384
rect 3550 3296 3870 4320
rect 3550 3232 3558 3296
rect 3622 3232 3638 3296
rect 3702 3232 3718 3296
rect 3782 3232 3798 3296
rect 3862 3232 3870 3296
rect 3550 2208 3870 3232
rect 3550 2144 3558 2208
rect 3622 2144 3638 2208
rect 3702 2144 3718 2208
rect 3782 2144 3798 2208
rect 3862 2144 3870 2208
rect 3550 2128 3870 2144
rect 5268 7104 5588 7120
rect 5268 7040 5276 7104
rect 5340 7040 5356 7104
rect 5420 7040 5436 7104
rect 5500 7040 5516 7104
rect 5580 7040 5588 7104
rect 5268 6016 5588 7040
rect 5268 5952 5276 6016
rect 5340 5952 5356 6016
rect 5420 5952 5436 6016
rect 5500 5952 5516 6016
rect 5580 5952 5588 6016
rect 5268 4928 5588 5952
rect 5268 4864 5276 4928
rect 5340 4864 5356 4928
rect 5420 4864 5436 4928
rect 5500 4864 5516 4928
rect 5580 4864 5588 4928
rect 5268 3840 5588 4864
rect 5268 3776 5276 3840
rect 5340 3776 5356 3840
rect 5420 3776 5436 3840
rect 5500 3776 5516 3840
rect 5580 3776 5588 3840
rect 5268 2752 5588 3776
rect 5268 2688 5276 2752
rect 5340 2688 5356 2752
rect 5420 2688 5436 2752
rect 5500 2688 5516 2752
rect 5580 2688 5588 2752
rect 5268 2128 5588 2688
rect 6985 6560 7305 7120
rect 6985 6496 6993 6560
rect 7057 6496 7073 6560
rect 7137 6496 7153 6560
rect 7217 6496 7233 6560
rect 7297 6496 7305 6560
rect 6985 5472 7305 6496
rect 6985 5408 6993 5472
rect 7057 5408 7073 5472
rect 7137 5408 7153 5472
rect 7217 5408 7233 5472
rect 7297 5408 7305 5472
rect 6985 4384 7305 5408
rect 6985 4320 6993 4384
rect 7057 4320 7073 4384
rect 7137 4320 7153 4384
rect 7217 4320 7233 4384
rect 7297 4320 7305 4384
rect 6985 3296 7305 4320
rect 6985 3232 6993 3296
rect 7057 3232 7073 3296
rect 7137 3232 7153 3296
rect 7217 3232 7233 3296
rect 7297 3232 7305 3296
rect 6985 2208 7305 3232
rect 6985 2144 6993 2208
rect 7057 2144 7073 2208
rect 7137 2144 7153 2208
rect 7217 2144 7233 2208
rect 7297 2144 7305 2208
rect 6985 2128 7305 2144
rect 8702 7104 9023 7120
rect 8702 7040 8710 7104
rect 8774 7040 8790 7104
rect 8854 7040 8870 7104
rect 8934 7040 8950 7104
rect 9014 7040 9023 7104
rect 8702 6016 9023 7040
rect 8702 5952 8710 6016
rect 8774 5952 8790 6016
rect 8854 5952 8870 6016
rect 8934 5952 8950 6016
rect 9014 5952 9023 6016
rect 8702 4928 9023 5952
rect 8702 4864 8710 4928
rect 8774 4864 8790 4928
rect 8854 4864 8870 4928
rect 8934 4864 8950 4928
rect 9014 4864 9023 4928
rect 8702 3840 9023 4864
rect 8702 3776 8710 3840
rect 8774 3776 8790 3840
rect 8854 3776 8870 3840
rect 8934 3776 8950 3840
rect 9014 3776 9023 3840
rect 8702 2752 9023 3776
rect 8702 2688 8710 2752
rect 8774 2688 8790 2752
rect 8854 2688 8870 2752
rect 8934 2688 8950 2752
rect 9014 2688 9023 2752
rect 8702 2128 9023 2688
use sky130_fd_sc_hd__decap_4  FILLER_0_9
timestamp 1626515363
transform 1 0 1104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6
timestamp 1626515363
transform 1 0 828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_10
timestamp 1626515363
transform 1 0 1196 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1626515363
transform 1 0 276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1626515363
transform 1 0 276 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1626515363
transform -1 0 828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input11
timestamp 1626515363
transform 1 0 552 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17
timestamp 1626515363
transform 1 0 1840 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1626515363
transform 1 0 1472 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _118_
timestamp 1626515363
transform 1 0 1288 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1626515363
transform 1 0 4048 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _116_
timestamp 1626515363
transform 1 0 3128 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_18
timestamp 1626515363
transform 1 0 2852 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25
timestamp 1626515363
transform 1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_39
timestamp 1626515363
transform 1 0 3864 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1626515363
transform 1 0 2944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_31
timestamp 1626515363
transform 1 0 3128 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _114_
timestamp 1626515363
transform -1 0 8188 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_6  _058_
timestamp 1626515363
transform -1 0 6348 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1626515363
transform 1 0 5428 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_19
timestamp 1626515363
transform 1 0 5428 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1626515363
transform 1 0 4324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1626515363
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1626515363
transform 1 0 5060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _112_
timestamp 1626515363
transform 1 0 8096 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _055_
timestamp 1626515363
transform 1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20
timestamp 1626515363
transform 1 0 8004 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1626515363
transform 1 0 7820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74
timestamp 1626515363
transform 1 0 7084 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70
timestamp 1626515363
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_86
timestamp 1626515363
transform 1 0 8188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66
timestamp 1626515363
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1626515363
transform 1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1626515363
transform -1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1626515363
transform -1 0 10580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1626515363
transform -1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_93
timestamp 1626515363
transform 1 0 8832 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_101
timestamp 1626515363
transform 1 0 9568 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_105
timestamp 1626515363
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_105
timestamp 1626515363
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _117_
timestamp 1626515363
transform -1 0 2484 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1626515363
transform 1 0 276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1626515363
transform 1 0 552 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _096_
timestamp 1626515363
transform -1 0 4416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _059_
timestamp 1626515363
transform 1 0 2944 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1626515363
transform 1 0 2852 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_38
timestamp 1626515363
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1626515363
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _094_
timestamp 1626515363
transform -1 0 5428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _069_
timestamp 1626515363
transform -1 0 6072 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_63
timestamp 1626515363
transform 1 0 6072 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_45
timestamp 1626515363
transform 1 0 4416 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_56
timestamp 1626515363
transform 1 0 5428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _057_
timestamp 1626515363
transform 1 0 6900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1626515363
transform 1 0 8004 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_75
timestamp 1626515363
transform 1 0 7176 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1626515363
transform 1 0 7912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_71
timestamp 1626515363
transform 1 0 6808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1626515363
transform 1 0 8096 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _079_
timestamp 1626515363
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _067_
timestamp 1626515363
transform -1 0 8740 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1626515363
transform -1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_107
timestamp 1626515363
transform 1 0 10120 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_99
timestamp 1626515363
transform 1 0 9384 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_92
timestamp 1626515363
transform 1 0 8740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _099_
timestamp 1626515363
transform 1 0 1656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1626515363
transform -1 0 1288 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1626515363
transform 1 0 276 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1626515363
transform 1 0 920 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_19
timestamp 1626515363
transform 1 0 2024 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_11
timestamp 1626515363
transform 1 0 1288 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1626515363
transform 1 0 552 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _107_
timestamp 1626515363
transform 1 0 2392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _056_
timestamp 1626515363
transform 1 0 3128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_42
timestamp 1626515363
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_34
timestamp 1626515363
transform 1 0 3404 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1626515363
transform 1 0 2760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _074_
timestamp 1626515363
transform -1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _095_
timestamp 1626515363
transform -1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1626515363
transform 1 0 5428 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_61
timestamp 1626515363
transform 1 0 5888 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_48
timestamp 1626515363
transform 1 0 4692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _119_
timestamp 1626515363
transform -1 0 9936 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__nand3_1  _072_
timestamp 1626515363
transform -1 0 7084 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_82
timestamp 1626515363
transform 1 0 7820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_74
timestamp 1626515363
transform 1 0 7084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_69
timestamp 1626515363
transform 1 0 6624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1626515363
transform -1 0 10580 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_105
timestamp 1626515363
transform 1 0 9936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1626515363
transform -1 0 828 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _097_
timestamp 1626515363
transform 1 0 1472 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1626515363
transform 1 0 276 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6
timestamp 1626515363
transform 1 0 828 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1626515363
transform 1 0 2024 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_12
timestamp 1626515363
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _078_
timestamp 1626515363
transform -1 0 4416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _060_
timestamp 1626515363
transform 1 0 3496 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1626515363
transform 1 0 2852 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_29
timestamp 1626515363
transform 1 0 2944 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1626515363
transform 1 0 2760 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_38
timestamp 1626515363
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _070_
timestamp 1626515363
transform -1 0 6348 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _089_
timestamp 1626515363
transform -1 0 5336 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_45
timestamp 1626515363
transform 1 0 4416 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_55
timestamp 1626515363
transform 1 0 5336 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _073_
timestamp 1626515363
transform 1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _071_
timestamp 1626515363
transform -1 0 6992 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _075_
timestamp 1626515363
transform 1 0 8096 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1626515363
transform 1 0 8004 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1626515363
transform 1 0 7636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_73
timestamp 1626515363
transform 1 0 6992 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_66
timestamp 1626515363
transform 1 0 6348 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _081_
timestamp 1626515363
transform -1 0 9936 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _080_
timestamp 1626515363
transform -1 0 9200 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1626515363
transform -1 0 10580 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_105
timestamp 1626515363
transform 1 0 9936 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_97
timestamp 1626515363
transform 1 0 9200 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_89
timestamp 1626515363
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _105_
timestamp 1626515363
transform 1 0 1012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _101_
timestamp 1626515363
transform 1 0 1656 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1626515363
transform 1 0 276 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1626515363
transform 1 0 920 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_19
timestamp 1626515363
transform 1 0 2024 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_11
timestamp 1626515363
transform 1 0 1288 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1626515363
transform 1 0 552 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _108_
timestamp 1626515363
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _061_
timestamp 1626515363
transform 1 0 3956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp 1626515363
transform -1 0 2668 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_43
timestamp 1626515363
transform 1 0 4232 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_33
timestamp 1626515363
transform 1 0 3312 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_39
timestamp 1626515363
transform 1 0 3864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_26
timestamp 1626515363
transform 1 0 2668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _098_
timestamp 1626515363
transform 1 0 4784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _076_
timestamp 1626515363
transform -1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1626515363
transform 1 0 5428 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1626515363
transform 1 0 5520 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1626515363
transform 1 0 5980 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1626515363
transform 1 0 5060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _065_
timestamp 1626515363
transform 1 0 6992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _100_
timestamp 1626515363
transform -1 0 8004 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _077_
timestamp 1626515363
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_84
timestamp 1626515363
transform 1 0 8004 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_76
timestamp 1626515363
transform 1 0 7268 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_69
timestamp 1626515363
transform 1 0 6624 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1626515363
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _066_
timestamp 1626515363
transform 1 0 8372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _087_
timestamp 1626515363
transform 1 0 9016 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1626515363
transform -1 0 10580 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_105
timestamp 1626515363
transform 1 0 9936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_98
timestamp 1626515363
transform 1 0 9292 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_91
timestamp 1626515363
transform 1 0 8648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1626515363
transform 1 0 552 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6
timestamp 1626515363
transform 1 0 828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1626515363
transform 1 0 276 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1626515363
transform 1 0 276 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _111_
timestamp 1626515363
transform -1 0 1012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1626515363
transform -1 0 828 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_8
timestamp 1626515363
transform 1 0 1012 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _110_
timestamp 1626515363
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1626515363
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp 1626515363
transform 1 0 1656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_16
timestamp 1626515363
transform 1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _109_
timestamp 1626515363
transform -1 0 2392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _103_
timestamp 1626515363
transform -1 0 2392 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1626515363
transform 1 0 4048 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _102_
timestamp 1626515363
transform 1 0 2944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1626515363
transform 1 0 2852 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_35
timestamp 1626515363
transform 1 0 3496 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_23
timestamp 1626515363
transform 1 0 2392 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1626515363
transform 1 0 3220 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1626515363
transform 1 0 2760 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1626515363
transform 1 0 2392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_48
timestamp 1626515363
transform 1 0 4692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1626515363
transform 1 0 4968 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_44
timestamp 1626515363
transform 1 0 4324 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _092_
timestamp 1626515363
transform -1 0 5428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _090_
timestamp 1626515363
transform 1 0 4416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_56
timestamp 1626515363
transform 1 0 5428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_61
timestamp 1626515363
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1626515363
transform 1 0 5336 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_65
timestamp 1626515363
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1626515363
transform 1 0 5428 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _091_
timestamp 1626515363
transform -1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _088_
timestamp 1626515363
transform -1 0 6072 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_63
timestamp 1626515363
transform 1 0 6072 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_69
timestamp 1626515363
transform 1 0 6624 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _062_
timestamp 1626515363
transform -1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _063_
timestamp 1626515363
transform 1 0 6992 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1626515363
transform 1 0 7636 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_76
timestamp 1626515363
transform 1 0 7268 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_75
timestamp 1626515363
transform 1 0 7176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _064_
timestamp 1626515363
transform -1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_84
timestamp 1626515363
transform 1 0 8004 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1626515363
transform 1 0 8004 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_1  _068_
timestamp 1626515363
transform -1 0 8648 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _085_
timestamp 1626515363
transform 1 0 8096 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_88
timestamp 1626515363
transform 1 0 8372 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_96
timestamp 1626515363
transform 1 0 9108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_91
timestamp 1626515363
transform 1 0 8648 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _083_
timestamp 1626515363
transform 1 0 8740 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_104
timestamp 1626515363
transform 1 0 9844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_97
timestamp 1626515363
transform 1 0 9200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_101
timestamp 1626515363
transform 1 0 9568 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _082_
timestamp 1626515363
transform -1 0 9568 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _084_
timestamp 1626515363
transform -1 0 9844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_108
timestamp 1626515363
transform 1 0 10212 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1626515363
transform -1 0 10580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1626515363
transform -1 0 10580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _113_
timestamp 1626515363
transform 1 0 644 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1626515363
transform 1 0 276 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1626515363
transform 1 0 552 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _115_
timestamp 1626515363
transform 1 0 3036 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1626515363
transform 1 0 2852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1626515363
transform 1 0 2944 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1626515363
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _093_
timestamp 1626515363
transform 1 0 5520 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1626515363
transform 1 0 5428 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_60
timestamp 1626515363
transform 1 0 5796 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_55
timestamp 1626515363
transform 1 0 5336 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_51
timestamp 1626515363
transform 1 0 4968 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1626515363
transform -1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _086_
timestamp 1626515363
transform 1 0 8096 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1626515363
transform 1 0 8004 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_68
timestamp 1626515363
transform 1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1626515363
transform 1 0 7820 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_74
timestamp 1626515363
transform 1 0 7084 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1626515363
transform 1 0 9476 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1626515363
transform -1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_103
timestamp 1626515363
transform 1 0 9752 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_88
timestamp 1626515363
transform 1 0 8372 0 1 6528
box -38 -48 1142 592
<< labels >>
rlabel metal4 s 3550 2128 3870 7120 6 VGND
port 0 nsew ground input
rlabel metal4 s 6985 2128 7305 7120 6 VGND
port 0 nsew ground input
rlabel metal4 s 1834 2128 2154 7120 6 VPWR
port 1 nsew power input
rlabel metal4 s 5268 2128 5588 7120 6 VPWR
port 1 nsew power input
rlabel metal4 s 8703 2128 9023 7120 6 VPWR
port 1 nsew power input
rlabel metal3 s 10482 3952 10882 4072 6 f_clk[0]
port 3 nsew signal input
rlabel metal3 s 0 2864 400 2984 6 f_clk[1]
port 4 nsew signal input
rlabel metal2 s 3974 7485 4030 7885 6 f_clk[2]
port 5 nsew signal input
rlabel metal3 s 0 4904 400 5024 6 f_clk[3]
port 6 nsew signal input
rlabel metal3 s 0 6808 400 6928 6 f_clk[6]
port 9 nsew signal input
rlabel metal2 s 6734 7485 6790 7885 6 f_clk[7]
port 10 nsew signal input
rlabel metal2 s 9402 7485 9458 7885 6 f_clk[8]
port 11 nsew signal input
rlabel metal2 s 1306 7485 1362 7885 6 sin_out
port 14 nsew signal tristate
rlabel metal2 s 1306 1400 1362 1800 6 cos_out
port 2 nsew signal tristate
rlabel metal2 s 3974 1400 4030 1800 6 f_clk[4]
port 7 nsew signal input
rlabel metal2 s 6734 1400 6790 1800 6 f_clk[5]
port 8 nsew signal input
rlabel metal2 s 9402 1400 9458 1800 6 f_clk[9]
port 12 nsew signal input
rlabel metal3 s 0 1560 400 1680 6 rstb
port 13 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 10882 7885
<< end >>
