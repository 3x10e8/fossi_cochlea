magic
tech sky130B
magscale 1 2
timestamp 1662948631
<< nwell >>
rect -204 204 302 417
<< nmos >>
rect -6 0 30 84
<< pmos >>
rect -6 240 30 366
rect 110 240 146 366
<< ndiff >>
rect -71 72 -6 84
rect -71 13 -63 72
rect -17 13 -6 72
rect -71 0 -6 13
rect 30 58 92 84
rect 30 24 48 58
rect 82 24 92 58
rect 30 0 92 24
<< pdiff >>
rect -84 354 -6 366
rect -84 259 -75 354
rect -17 259 -6 354
rect -84 240 -6 259
rect 30 354 110 366
rect 30 259 41 354
rect 99 259 110 354
rect 30 240 110 259
rect 146 353 254 366
rect 146 258 158 353
rect 216 258 254 353
rect 146 240 254 258
<< ndiffc >>
rect -63 13 -17 72
rect 48 24 82 58
<< pdiffc >>
rect -75 259 -17 354
rect 41 259 99 354
rect 158 258 216 353
<< psubdiff >>
rect -177 71 -71 84
rect -177 12 -153 71
rect -107 12 -71 71
rect -177 0 -71 12
<< nsubdiff >>
rect -168 350 -84 366
rect -168 261 -144 350
rect -109 261 -84 350
rect -168 240 -84 261
<< psubdiffcont >>
rect -153 12 -107 71
<< nsubdiffcont >>
rect -144 261 -109 350
<< poly >>
rect -6 392 146 424
rect -6 366 30 392
rect 110 366 146 392
rect -151 180 -95 189
rect -6 180 30 240
rect 110 214 146 240
rect -151 179 30 180
rect -157 145 -141 179
rect -107 145 30 179
rect -151 144 30 145
rect -151 135 -95 144
rect -6 84 30 144
rect -6 -26 30 0
<< polycont >>
rect -141 145 -107 179
<< locali >>
rect -276 447 -247 481
rect -213 447 -155 481
rect -121 447 -63 481
rect -29 447 29 481
rect 63 447 121 481
rect 155 447 213 481
rect 247 447 305 481
rect 339 447 368 481
rect -148 374 -38 447
rect -148 366 -10 374
rect -152 354 -10 366
rect -152 350 -75 354
rect -152 261 -144 350
rect -109 261 -75 350
rect -152 259 -75 261
rect -17 259 -10 354
rect -152 245 -10 259
rect 32 366 105 374
rect 164 373 200 447
rect 32 354 106 366
rect 32 259 41 354
rect 99 259 106 354
rect 32 245 106 259
rect 149 365 222 373
rect 149 353 223 365
rect 149 258 158 353
rect 216 258 223 353
rect -75 243 -17 245
rect 41 243 99 245
rect 149 244 223 258
rect -157 145 -141 179
rect -107 145 -91 179
rect -153 84 -107 87
rect -63 84 -17 89
rect 158 242 216 244
rect -153 83 -17 84
rect -153 72 -8 83
rect -153 71 -63 72
rect -107 13 -63 71
rect -17 13 -8 72
rect -107 12 -8 13
rect -153 1 -8 12
rect 32 58 92 84
rect 32 24 48 58
rect 82 24 92 58
rect -153 -3 -17 1
rect 32 0 92 24
rect -153 -4 -53 -3
rect -147 -63 -53 -4
rect -276 -97 -247 -63
rect -213 -97 -155 -63
rect -121 -97 -63 -63
rect -29 -97 29 -63
rect 63 -97 121 -63
rect 155 -97 213 -63
rect 247 -97 305 -63
rect 339 -97 368 -63
<< viali >>
rect -247 447 -213 481
rect -155 447 -121 481
rect -63 447 -29 481
rect 29 447 63 481
rect 121 447 155 481
rect 213 447 247 481
rect 305 447 339 481
rect -141 145 -107 179
rect 48 84 82 243
rect -247 -97 -213 -63
rect -155 -97 -121 -63
rect -63 -97 -29 -63
rect 29 -97 63 -63
rect 121 -97 155 -63
rect 213 -97 247 -63
rect 305 -97 339 -63
<< metal1 >>
rect -276 481 368 512
rect -276 447 -247 481
rect -213 447 -155 481
rect -121 447 -63 481
rect -29 447 29 481
rect 63 447 121 481
rect 155 447 213 481
rect 247 447 305 481
rect 339 447 368 481
rect -276 416 368 447
rect 39 243 90 256
rect -154 188 -91 189
rect -156 136 -150 188
rect -98 136 -91 188
rect -154 135 -91 136
rect 39 84 48 243
rect 82 84 90 243
rect 39 72 90 84
rect -276 -63 368 -32
rect -276 -97 -247 -63
rect -213 -97 -155 -63
rect -121 -97 -63 -63
rect -29 -97 29 -63
rect 63 -97 121 -63
rect 155 -97 213 -63
rect 247 -97 305 -63
rect 339 -97 368 -63
rect -276 -128 368 -97
<< via1 >>
rect -150 179 -98 188
rect -150 145 -141 179
rect -141 145 -107 179
rect -107 145 -98 179
rect -150 136 -98 145
<< metal2 >>
rect -156 136 -150 188
rect -98 136 -92 188
<< labels >>
flabel metal2 -141 145 -107 179 0 FreeSans 160 0 0 0 in
port 2 nsew default input
flabel viali 48 84 82 243 0 FreeSans 160 0 0 0 out
port 3 nsew default output
flabel metal1 -29 -128 29 -32 1 FreeSans 320 0 0 0 vss
port 4 n default bidirectional
flabel metal1 -10 416 84 512 1 FreeSans 320 0 0 0 vdd
port 5 n default bidirectional
<< end >>
