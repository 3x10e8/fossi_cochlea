magic
tech sky130A
magscale 1 2
timestamp 1654644553
<< viali >>
rect 1501 27557 1535 27591
rect 2881 27557 2915 27591
rect 9045 27557 9079 27591
rect 20177 27557 20211 27591
rect 24777 27557 24811 27591
rect 30113 27557 30147 27591
rect 33057 27557 33091 27591
rect 35633 27557 35667 27591
rect 52009 27557 52043 27591
rect 36185 27489 36219 27523
rect 1685 27421 1719 27455
rect 3065 27421 3099 27455
rect 9229 27421 9263 27455
rect 14105 27421 14139 27455
rect 14749 27421 14783 27455
rect 19533 27421 19567 27455
rect 19993 27421 20027 27455
rect 24593 27421 24627 27455
rect 28089 27421 28123 27455
rect 30297 27421 30331 27455
rect 34713 27421 34747 27455
rect 35449 27421 35483 27455
rect 40417 27421 40451 27455
rect 40877 27421 40911 27455
rect 45937 27421 45971 27455
rect 46397 27421 46431 27455
rect 51825 27421 51859 27455
rect 56885 27421 56919 27455
rect 57253 27421 57287 27455
rect 20637 27353 20671 27387
rect 27537 27353 27571 27387
rect 33517 27353 33551 27387
rect 34161 27353 34195 27387
rect 57897 27353 57931 27387
rect 58081 27353 58115 27387
rect 3893 27285 3927 27319
rect 9781 27285 9815 27319
rect 14289 27285 14323 27319
rect 19349 27285 19383 27319
rect 25789 27285 25823 27319
rect 26433 27285 26467 27319
rect 28549 27285 28583 27319
rect 31309 27285 31343 27319
rect 32505 27285 32539 27319
rect 34897 27285 34931 27319
rect 41061 27285 41095 27319
rect 46581 27285 46615 27319
rect 1501 27081 1535 27115
rect 20821 27081 20855 27115
rect 25789 27081 25823 27115
rect 34069 27081 34103 27115
rect 58081 27081 58115 27115
rect 57253 27013 57287 27047
rect 1685 26945 1719 26979
rect 21005 26945 21039 26979
rect 21833 26945 21867 26979
rect 30757 26945 30791 26979
rect 31585 26945 31619 26979
rect 57897 26945 57931 26979
rect 26433 26877 26467 26911
rect 34621 26877 34655 26911
rect 28917 26809 28951 26843
rect 35173 26809 35207 26843
rect 25237 26741 25271 26775
rect 27353 26741 27387 26775
rect 28365 26741 28399 26775
rect 29469 26741 29503 26775
rect 30297 26741 30331 26775
rect 30849 26741 30883 26775
rect 31493 26741 31527 26775
rect 32137 26741 32171 26775
rect 32689 26741 32723 26775
rect 33425 26741 33459 26775
rect 35725 26741 35759 26775
rect 36185 26741 36219 26775
rect 37381 26741 37415 26775
rect 30481 26537 30515 26571
rect 31217 26537 31251 26571
rect 58081 26537 58115 26571
rect 29561 26469 29595 26503
rect 30389 26469 30423 26503
rect 26433 26401 26467 26435
rect 30573 26401 30607 26435
rect 1685 26333 1719 26367
rect 27629 26333 27663 26367
rect 29745 26333 29779 26367
rect 30297 26333 30331 26367
rect 31217 26333 31251 26367
rect 31953 26333 31987 26367
rect 32413 26333 32447 26367
rect 32505 26333 32539 26367
rect 33241 26333 33275 26367
rect 36461 26333 36495 26367
rect 28273 26265 28307 26299
rect 33149 26265 33183 26299
rect 33793 26265 33827 26299
rect 34713 26265 34747 26299
rect 36921 26265 36955 26299
rect 38117 26265 38151 26299
rect 1501 26197 1535 26231
rect 24685 26197 24719 26231
rect 25145 26197 25179 26231
rect 25789 26197 25823 26231
rect 26985 26197 27019 26231
rect 29009 26197 29043 26231
rect 31769 26197 31803 26231
rect 35265 26197 35299 26231
rect 35817 26197 35851 26231
rect 37565 26197 37599 26231
rect 30481 25993 30515 26027
rect 37289 25993 37323 26027
rect 38393 25993 38427 26027
rect 38945 25993 38979 26027
rect 44373 25993 44407 26027
rect 23765 25925 23799 25959
rect 30941 25925 30975 25959
rect 32413 25925 32447 25959
rect 28825 25857 28859 25891
rect 29009 25857 29043 25891
rect 29837 25857 29871 25891
rect 31585 25857 31619 25891
rect 32137 25857 32171 25891
rect 33057 25857 33091 25891
rect 33701 25857 33735 25891
rect 44189 25857 44223 25891
rect 47593 25857 47627 25891
rect 58081 25857 58115 25891
rect 29745 25789 29779 25823
rect 27261 25721 27295 25755
rect 27813 25721 27847 25755
rect 30573 25721 30607 25755
rect 35357 25721 35391 25755
rect 36369 25721 36403 25755
rect 57897 25721 57931 25755
rect 23213 25653 23247 25687
rect 24409 25653 24443 25687
rect 24869 25653 24903 25687
rect 25421 25653 25455 25687
rect 26433 25653 26467 25687
rect 28273 25653 28307 25687
rect 28917 25653 28951 25687
rect 29469 25653 29503 25687
rect 31493 25653 31527 25687
rect 32965 25653 32999 25687
rect 33609 25653 33643 25687
rect 34253 25653 34287 25687
rect 34713 25653 34747 25687
rect 35909 25653 35943 25687
rect 37933 25653 37967 25687
rect 47777 25653 47811 25687
rect 23305 25449 23339 25483
rect 32413 25449 32447 25483
rect 34713 25449 34747 25483
rect 35357 25449 35391 25483
rect 37565 25449 37599 25483
rect 58173 25449 58207 25483
rect 14473 25381 14507 25415
rect 23857 25381 23891 25415
rect 27353 25381 27387 25415
rect 29561 25381 29595 25415
rect 25513 25313 25547 25347
rect 28825 25313 28859 25347
rect 30481 25313 30515 25347
rect 31401 25313 31435 25347
rect 27997 25245 28031 25279
rect 28641 25245 28675 25279
rect 29929 25245 29963 25279
rect 30573 25245 30607 25279
rect 31585 25245 31619 25279
rect 33057 25245 33091 25279
rect 33793 25245 33827 25279
rect 35449 25245 35483 25279
rect 37013 25245 37047 25279
rect 39221 25245 39255 25279
rect 14657 25177 14691 25211
rect 29745 25177 29779 25211
rect 31769 25177 31803 25211
rect 32229 25177 32263 25211
rect 32445 25177 32479 25211
rect 33885 25177 33919 25211
rect 24961 25109 24995 25143
rect 26065 25109 26099 25143
rect 26801 25109 26835 25143
rect 27905 25109 27939 25143
rect 28457 25109 28491 25143
rect 30941 25109 30975 25143
rect 32597 25109 32631 25143
rect 33241 25109 33275 25143
rect 35909 25109 35943 25143
rect 36553 25109 36587 25143
rect 38117 25109 38151 25143
rect 38761 25109 38795 25143
rect 32505 24905 32539 24939
rect 27905 24837 27939 24871
rect 28135 24803 28169 24837
rect 1685 24769 1719 24803
rect 11713 24769 11747 24803
rect 27261 24769 27295 24803
rect 27445 24769 27479 24803
rect 29101 24769 29135 24803
rect 30021 24769 30055 24803
rect 30665 24769 30699 24803
rect 31585 24769 31619 24803
rect 32137 24769 32171 24803
rect 32321 24769 32355 24803
rect 32413 24769 32447 24803
rect 33149 24769 33183 24803
rect 33977 24769 34011 24803
rect 34161 24769 34195 24803
rect 34805 24769 34839 24803
rect 35541 24769 35575 24803
rect 36185 24769 36219 24803
rect 36737 24769 36771 24803
rect 40601 24769 40635 24803
rect 25237 24701 25271 24735
rect 29009 24701 29043 24735
rect 29745 24701 29779 24735
rect 37841 24701 37875 24735
rect 11529 24633 11563 24667
rect 22201 24633 22235 24667
rect 27353 24633 27387 24667
rect 28273 24633 28307 24667
rect 32689 24633 32723 24667
rect 34621 24633 34655 24667
rect 38393 24633 38427 24667
rect 40141 24633 40175 24667
rect 1501 24565 1535 24599
rect 22753 24565 22787 24599
rect 23213 24565 23247 24599
rect 24225 24565 24259 24599
rect 24777 24565 24811 24599
rect 25789 24565 25823 24599
rect 26341 24565 26375 24599
rect 28089 24565 28123 24599
rect 28825 24565 28859 24599
rect 30849 24565 30883 24599
rect 31493 24565 31527 24599
rect 33149 24565 33183 24599
rect 35449 24565 35483 24599
rect 36093 24565 36127 24599
rect 37289 24565 37323 24599
rect 38945 24565 38979 24599
rect 39497 24565 39531 24599
rect 16681 24361 16715 24395
rect 17417 24361 17451 24395
rect 23857 24361 23891 24395
rect 33977 24361 34011 24395
rect 40509 24361 40543 24395
rect 14473 24293 14507 24327
rect 21649 24293 21683 24327
rect 22201 24293 22235 24327
rect 25605 24293 25639 24327
rect 34161 24293 34195 24327
rect 34897 24293 34931 24327
rect 36921 24293 36955 24327
rect 27905 24225 27939 24259
rect 29009 24225 29043 24259
rect 29653 24225 29687 24259
rect 32781 24225 32815 24259
rect 32965 24225 32999 24259
rect 33242 24225 33276 24259
rect 39221 24225 39255 24259
rect 16773 24157 16807 24191
rect 21097 24157 21131 24191
rect 23305 24157 23339 24191
rect 26065 24157 26099 24191
rect 26801 24157 26835 24191
rect 27735 24157 27769 24191
rect 28825 24157 28859 24191
rect 29745 24157 29779 24191
rect 32321 24157 32355 24191
rect 33057 24157 33091 24191
rect 33149 24157 33183 24191
rect 34713 24157 34747 24191
rect 35541 24157 35575 24191
rect 36185 24157 36219 24191
rect 36829 24157 36863 24191
rect 37473 24157 37507 24191
rect 58173 24157 58207 24191
rect 14657 24089 14691 24123
rect 25053 24089 25087 24123
rect 26709 24089 26743 24123
rect 28641 24089 28675 24123
rect 32045 24089 32079 24123
rect 33793 24089 33827 24123
rect 34009 24089 34043 24123
rect 37565 24089 37599 24123
rect 39865 24089 39899 24123
rect 40969 24089 41003 24123
rect 57897 24089 57931 24123
rect 22661 24021 22695 24055
rect 24501 24021 24535 24055
rect 26157 24021 26191 24055
rect 27445 24021 27479 24055
rect 28457 24021 28491 24055
rect 28733 24021 28767 24055
rect 30113 24021 30147 24055
rect 30573 24021 30607 24055
rect 35725 24021 35759 24055
rect 36277 24021 36311 24055
rect 38209 24021 38243 24055
rect 38669 24021 38703 24055
rect 25697 23817 25731 23851
rect 32137 23817 32171 23851
rect 35541 23817 35575 23851
rect 40785 23817 40819 23851
rect 58173 23817 58207 23851
rect 20177 23749 20211 23783
rect 20729 23749 20763 23783
rect 25513 23681 25547 23715
rect 25697 23681 25731 23715
rect 26157 23681 26191 23715
rect 26433 23681 26467 23715
rect 27445 23681 27479 23715
rect 28549 23681 28583 23715
rect 28825 23681 28859 23715
rect 29745 23681 29779 23715
rect 32965 23681 32999 23715
rect 33885 23681 33919 23715
rect 35081 23681 35115 23715
rect 35725 23681 35759 23715
rect 35817 23681 35851 23715
rect 36645 23681 36679 23715
rect 37289 23681 37323 23715
rect 38117 23681 38151 23715
rect 39221 23681 39255 23715
rect 21925 23613 21959 23647
rect 24593 23613 24627 23647
rect 24869 23613 24903 23647
rect 27353 23613 27387 23647
rect 30021 23613 30055 23647
rect 31493 23613 31527 23647
rect 32873 23613 32907 23647
rect 33977 23613 34011 23647
rect 34989 23613 35023 23647
rect 36369 23613 36403 23647
rect 22569 23545 22603 23579
rect 26341 23545 26375 23579
rect 26433 23545 26467 23579
rect 28365 23545 28399 23579
rect 28733 23545 28767 23579
rect 34253 23545 34287 23579
rect 37473 23545 37507 23579
rect 40325 23545 40359 23579
rect 21281 23477 21315 23511
rect 23121 23477 23155 23511
rect 27721 23477 27755 23511
rect 34713 23477 34747 23511
rect 35081 23477 35115 23511
rect 36461 23477 36495 23511
rect 36553 23477 36587 23511
rect 38025 23477 38059 23511
rect 38669 23477 38703 23511
rect 39681 23477 39715 23511
rect 41429 23477 41463 23511
rect 2237 23273 2271 23307
rect 20177 23273 20211 23307
rect 26893 23273 26927 23307
rect 30021 23273 30055 23307
rect 40969 23273 41003 23307
rect 19533 23205 19567 23239
rect 32229 23205 32263 23239
rect 38117 23205 38151 23239
rect 24593 23137 24627 23171
rect 26341 23137 26375 23171
rect 27445 23137 27479 23171
rect 28917 23137 28951 23171
rect 31493 23137 31527 23171
rect 34989 23137 35023 23171
rect 36001 23137 36035 23171
rect 36645 23137 36679 23171
rect 1685 23069 1719 23103
rect 21649 23069 21683 23103
rect 24501 23069 24535 23103
rect 24685 23069 24719 23103
rect 25237 23069 25271 23103
rect 26249 23069 26283 23103
rect 27261 23069 27295 23103
rect 27997 23069 28031 23103
rect 28181 23069 28215 23103
rect 31769 23069 31803 23103
rect 33977 23069 34011 23103
rect 34897 23069 34931 23103
rect 37381 23069 37415 23103
rect 38025 23069 38059 23103
rect 38669 23069 38703 23103
rect 25145 23001 25179 23035
rect 27077 23001 27111 23035
rect 33701 23001 33735 23035
rect 36093 23001 36127 23035
rect 38761 23001 38795 23035
rect 1501 22933 1535 22967
rect 20729 22933 20763 22967
rect 22201 22933 22235 22967
rect 22753 22933 22787 22967
rect 23305 22933 23339 22967
rect 23857 22933 23891 22967
rect 25881 22933 25915 22967
rect 27169 22933 27203 22967
rect 35265 22933 35299 22967
rect 37473 22933 37507 22967
rect 39865 22933 39899 22967
rect 40417 22933 40451 22967
rect 41521 22933 41555 22967
rect 42165 22933 42199 22967
rect 42625 22933 42659 22967
rect 18429 22729 18463 22763
rect 20085 22729 20119 22763
rect 21281 22729 21315 22763
rect 27445 22729 27479 22763
rect 32137 22729 32171 22763
rect 37289 22729 37323 22763
rect 37473 22729 37507 22763
rect 41429 22729 41463 22763
rect 42993 22729 43027 22763
rect 20545 22661 20579 22695
rect 24041 22661 24075 22695
rect 25605 22661 25639 22695
rect 26157 22661 26191 22695
rect 26249 22661 26283 22695
rect 26985 22661 27019 22695
rect 29101 22661 29135 22695
rect 38301 22661 38335 22695
rect 40785 22661 40819 22695
rect 23489 22593 23523 22627
rect 23949 22593 23983 22627
rect 24133 22593 24167 22627
rect 24961 22593 24995 22627
rect 27169 22593 27203 22627
rect 27261 22593 27295 22627
rect 28181 22593 28215 22627
rect 28825 22593 28859 22627
rect 35357 22593 35391 22627
rect 35725 22593 35759 22627
rect 36369 22593 36403 22627
rect 36737 22593 36771 22627
rect 37841 22593 37875 22627
rect 38577 22593 38611 22627
rect 39221 22593 39255 22627
rect 19533 22525 19567 22559
rect 25053 22525 25087 22559
rect 27905 22525 27939 22559
rect 31033 22525 31067 22559
rect 31309 22525 31343 22559
rect 33609 22525 33643 22559
rect 33885 22525 33919 22559
rect 34713 22525 34747 22559
rect 36461 22457 36495 22491
rect 39129 22457 39163 22491
rect 43545 22457 43579 22491
rect 18981 22389 19015 22423
rect 22109 22389 22143 22423
rect 22753 22389 22787 22423
rect 23397 22389 23431 22423
rect 24685 22389 24719 22423
rect 26985 22389 27019 22423
rect 29561 22389 29595 22423
rect 36553 22389 36587 22423
rect 36737 22389 36771 22423
rect 37473 22389 37507 22423
rect 39681 22389 39715 22423
rect 40233 22389 40267 22423
rect 42533 22389 42567 22423
rect 27524 22185 27558 22219
rect 31493 22185 31527 22219
rect 43269 22185 43303 22219
rect 43821 22185 43855 22219
rect 23857 22117 23891 22151
rect 25605 22117 25639 22151
rect 38577 22117 38611 22151
rect 39957 22117 39991 22151
rect 41061 22117 41095 22151
rect 18705 22049 18739 22083
rect 23029 22049 23063 22083
rect 25329 22049 25363 22083
rect 26249 22049 26283 22083
rect 30021 22049 30055 22083
rect 37657 22049 37691 22083
rect 38485 22049 38519 22083
rect 38669 22049 38703 22083
rect 44373 22049 44407 22083
rect 22293 21981 22327 22015
rect 22937 21981 22971 22015
rect 23121 21981 23155 22015
rect 24409 21981 24443 22015
rect 25237 21981 25271 22015
rect 26433 21981 26467 22015
rect 27261 21981 27295 22015
rect 29745 21981 29779 22015
rect 33701 21981 33735 22015
rect 37749 21981 37783 22015
rect 38393 21981 38427 22015
rect 39129 21981 39163 22015
rect 39313 21981 39347 22015
rect 39865 21981 39899 22015
rect 58173 21981 58207 22015
rect 20545 21913 20579 21947
rect 23673 21913 23707 21947
rect 24501 21913 24535 21947
rect 33425 21913 33459 21947
rect 36921 21913 36955 21947
rect 41613 21913 41647 21947
rect 57897 21913 57931 21947
rect 17509 21845 17543 21879
rect 18061 21845 18095 21879
rect 19441 21845 19475 21879
rect 19993 21845 20027 21879
rect 21005 21845 21039 21879
rect 21557 21845 21591 21879
rect 22109 21845 22143 21879
rect 26341 21845 26375 21879
rect 26801 21845 26835 21879
rect 29009 21845 29043 21879
rect 31953 21845 31987 21879
rect 35633 21845 35667 21879
rect 37381 21845 37415 21879
rect 39221 21845 39255 21879
rect 40509 21845 40543 21879
rect 42257 21845 42291 21879
rect 42809 21845 42843 21879
rect 17693 21641 17727 21675
rect 20729 21641 20763 21675
rect 38761 21641 38795 21675
rect 39681 21641 39715 21675
rect 41613 21641 41647 21675
rect 44097 21641 44131 21675
rect 58173 21641 58207 21675
rect 17141 21573 17175 21607
rect 22845 21573 22879 21607
rect 34621 21573 34655 21607
rect 39957 21573 39991 21607
rect 1685 21505 1719 21539
rect 22385 21505 22419 21539
rect 24317 21505 24351 21539
rect 24685 21505 24719 21539
rect 25237 21505 25271 21539
rect 25513 21505 25547 21539
rect 26157 21505 26191 21539
rect 26985 21505 27019 21539
rect 27629 21505 27663 21539
rect 32137 21505 32171 21539
rect 34345 21505 34379 21539
rect 36737 21505 36771 21539
rect 37565 21505 37599 21539
rect 39681 21505 39715 21539
rect 40601 21505 40635 21539
rect 41153 21505 41187 21539
rect 18245 21437 18279 21471
rect 19625 21437 19659 21471
rect 27905 21437 27939 21471
rect 29837 21437 29871 21471
rect 30113 21437 30147 21471
rect 32413 21437 32447 21471
rect 37289 21437 37323 21471
rect 39221 21437 39255 21471
rect 43085 21437 43119 21471
rect 36093 21369 36127 21403
rect 38853 21369 38887 21403
rect 39773 21369 39807 21403
rect 43545 21369 43579 21403
rect 1501 21301 1535 21335
rect 18705 21301 18739 21335
rect 20177 21301 20211 21335
rect 21281 21301 21315 21335
rect 22293 21301 22327 21335
rect 26341 21301 26375 21335
rect 27077 21301 27111 21335
rect 29377 21301 29411 21335
rect 31585 21301 31619 21335
rect 33885 21301 33919 21335
rect 36645 21301 36679 21335
rect 40509 21301 40543 21335
rect 42533 21301 42567 21335
rect 44741 21301 44775 21335
rect 45293 21301 45327 21335
rect 15761 21097 15795 21131
rect 21833 21097 21867 21131
rect 23765 21097 23799 21131
rect 24409 21097 24443 21131
rect 27261 21097 27295 21131
rect 32965 21097 32999 21131
rect 40049 21097 40083 21131
rect 42073 21097 42107 21131
rect 45017 21097 45051 21131
rect 34713 21029 34747 21063
rect 42625 21029 42659 21063
rect 17969 20961 18003 20995
rect 18705 20961 18739 20995
rect 22569 20961 22603 20995
rect 23397 20961 23431 20995
rect 24961 20961 24995 20995
rect 25605 20961 25639 20995
rect 28733 20961 28767 20995
rect 29009 20961 29043 20995
rect 30113 20961 30147 20995
rect 30941 20961 30975 20995
rect 32413 20961 32447 20995
rect 34069 20961 34103 20995
rect 19901 20893 19935 20927
rect 21189 20893 21223 20927
rect 21649 20893 21683 20927
rect 22477 20893 22511 20927
rect 23489 20893 23523 20927
rect 24869 20893 24903 20927
rect 25881 20893 25915 20927
rect 26525 20893 26559 20927
rect 29745 20893 29779 20927
rect 29837 20893 29871 20927
rect 30205 20893 30239 20927
rect 30665 20893 30699 20927
rect 33149 20893 33183 20927
rect 33793 20893 33827 20927
rect 36461 20893 36495 20927
rect 39313 20893 39347 20927
rect 40693 20893 40727 20927
rect 41337 20893 41371 20927
rect 41521 20893 41555 20927
rect 42165 20893 42199 20927
rect 43821 20893 43855 20927
rect 21097 20825 21131 20859
rect 26801 20825 26835 20859
rect 29561 20825 29595 20859
rect 36185 20825 36219 20859
rect 36921 20825 36955 20859
rect 38669 20825 38703 20859
rect 39957 20825 39991 20859
rect 40877 20825 40911 20859
rect 44373 20825 44407 20859
rect 16221 20757 16255 20791
rect 16773 20757 16807 20791
rect 17417 20757 17451 20791
rect 19441 20757 19475 20791
rect 20545 20757 20579 20791
rect 22845 20757 22879 20791
rect 24777 20757 24811 20791
rect 30021 20757 30055 20791
rect 39221 20757 39255 20791
rect 41429 20757 41463 20791
rect 43177 20757 43211 20791
rect 45661 20757 45695 20791
rect 46213 20757 46247 20791
rect 16129 20553 16163 20587
rect 17049 20553 17083 20587
rect 18153 20553 18187 20587
rect 21005 20553 21039 20587
rect 32137 20553 32171 20587
rect 36645 20553 36679 20587
rect 40877 20553 40911 20587
rect 43177 20553 43211 20587
rect 45385 20553 45419 20587
rect 46489 20553 46523 20587
rect 19809 20485 19843 20519
rect 24041 20485 24075 20519
rect 24133 20485 24167 20519
rect 29469 20485 29503 20519
rect 33609 20485 33643 20519
rect 39037 20485 39071 20519
rect 40969 20485 41003 20519
rect 44281 20485 44315 20519
rect 19901 20417 19935 20451
rect 20545 20417 20579 20451
rect 21281 20417 21315 20451
rect 21833 20417 21867 20451
rect 22661 20417 22695 20451
rect 26433 20417 26467 20451
rect 26985 20417 27019 20451
rect 31585 20417 31619 20451
rect 33885 20417 33919 20451
rect 36093 20417 36127 20451
rect 36737 20417 36771 20451
rect 37657 20417 37691 20451
rect 37933 20417 37967 20451
rect 40049 20417 40083 20451
rect 40325 20417 40359 20451
rect 41705 20417 41739 20451
rect 42625 20417 42659 20451
rect 43269 20417 43303 20451
rect 21005 20349 21039 20383
rect 22569 20349 22603 20383
rect 23673 20349 23707 20383
rect 26157 20349 26191 20383
rect 27261 20349 27295 20383
rect 29193 20349 29227 20383
rect 35817 20349 35851 20383
rect 37381 20349 37415 20383
rect 38945 20349 38979 20383
rect 39221 20349 39255 20383
rect 40141 20349 40175 20383
rect 43729 20349 43763 20383
rect 15577 20281 15611 20315
rect 20453 20281 20487 20315
rect 23029 20281 23063 20315
rect 24685 20281 24719 20315
rect 14933 20213 14967 20247
rect 17509 20213 17543 20247
rect 18613 20213 18647 20247
rect 19165 20213 19199 20247
rect 21189 20213 21223 20247
rect 21925 20213 21959 20247
rect 28733 20213 28767 20247
rect 30941 20213 30975 20247
rect 31493 20213 31527 20247
rect 34345 20213 34379 20247
rect 40233 20213 40267 20247
rect 41613 20213 41647 20247
rect 42533 20213 42567 20247
rect 44833 20213 44867 20247
rect 46029 20213 46063 20247
rect 15393 20009 15427 20043
rect 17601 20009 17635 20043
rect 20085 20009 20119 20043
rect 22109 20009 22143 20043
rect 29009 20009 29043 20043
rect 38669 20009 38703 20043
rect 39865 20009 39899 20043
rect 40785 20009 40819 20043
rect 41797 20009 41831 20043
rect 44281 20009 44315 20043
rect 46673 20009 46707 20043
rect 12265 19941 12299 19975
rect 17049 19941 17083 19975
rect 21189 19941 21223 19975
rect 24501 19941 24535 19975
rect 26801 19941 26835 19975
rect 29561 19941 29595 19975
rect 40049 19941 40083 19975
rect 40877 19941 40911 19975
rect 20729 19873 20763 19907
rect 21925 19873 21959 19907
rect 22661 19873 22695 19907
rect 25329 19873 25363 19907
rect 27261 19873 27295 19907
rect 27537 19873 27571 19907
rect 30205 19873 30239 19907
rect 32597 19873 32631 19907
rect 34713 19873 34747 19907
rect 34989 19873 35023 19907
rect 36921 19873 36955 19907
rect 43085 19873 43119 19907
rect 1685 19805 1719 19839
rect 12449 19805 12483 19839
rect 18613 19805 18647 19839
rect 19533 19805 19567 19839
rect 19993 19805 20027 19839
rect 20821 19805 20855 19839
rect 21833 19805 21867 19839
rect 22937 19805 22971 19839
rect 23581 19805 23615 19839
rect 24409 19805 24443 19839
rect 25053 19805 25087 19839
rect 30757 19805 30791 19839
rect 33701 19805 33735 19839
rect 34069 19805 34103 19839
rect 39129 19805 39163 19839
rect 39221 19805 39255 19839
rect 41889 19805 41923 19839
rect 42533 19805 42567 19839
rect 43177 19805 43211 19839
rect 47317 19805 47351 19839
rect 58173 19805 58207 19839
rect 15945 19737 15979 19771
rect 19441 19737 19475 19771
rect 23857 19737 23891 19771
rect 32413 19737 32447 19771
rect 33057 19737 33091 19771
rect 37197 19737 37231 19771
rect 40325 19737 40359 19771
rect 41245 19737 41279 19771
rect 57897 19737 57931 19771
rect 1501 19669 1535 19703
rect 14197 19669 14231 19703
rect 14841 19669 14875 19703
rect 16405 19669 16439 19703
rect 18061 19669 18095 19703
rect 29929 19669 29963 19703
rect 30021 19669 30055 19703
rect 36461 19669 36495 19703
rect 42441 19669 42475 19703
rect 43729 19669 43763 19703
rect 45017 19669 45051 19703
rect 45661 19669 45695 19703
rect 46213 19669 46247 19703
rect 47777 19669 47811 19703
rect 12081 19465 12115 19499
rect 16129 19465 16163 19499
rect 20729 19465 20763 19499
rect 20913 19465 20947 19499
rect 21005 19465 21039 19499
rect 22293 19465 22327 19499
rect 22569 19465 22603 19499
rect 26433 19465 26467 19499
rect 27077 19465 27111 19499
rect 39037 19465 39071 19499
rect 46673 19465 46707 19499
rect 58173 19465 58207 19499
rect 17325 19397 17359 19431
rect 18521 19397 18555 19431
rect 29745 19397 29779 19431
rect 31401 19397 31435 19431
rect 33793 19397 33827 19431
rect 37565 19397 37599 19431
rect 43913 19397 43947 19431
rect 12265 19329 12299 19363
rect 17785 19329 17819 19363
rect 18429 19329 18463 19363
rect 19065 19329 19099 19363
rect 19901 19329 19935 19363
rect 21097 19329 21131 19363
rect 22201 19329 22235 19363
rect 22410 19329 22444 19363
rect 23305 19329 23339 19363
rect 23949 19329 23983 19363
rect 24225 19329 24259 19363
rect 24685 19329 24719 19363
rect 27537 19329 27571 19363
rect 31585 19329 31619 19363
rect 33977 19329 34011 19363
rect 36185 19329 36219 19363
rect 37289 19329 37323 19363
rect 39865 19329 39899 19363
rect 40141 19329 40175 19363
rect 41521 19329 41555 19363
rect 42717 19329 42751 19363
rect 43177 19329 43211 19363
rect 43269 19329 43303 19363
rect 43821 19329 43855 19363
rect 44557 19329 44591 19363
rect 12725 19261 12759 19295
rect 13553 19261 13587 19295
rect 15577 19261 15611 19295
rect 19165 19261 19199 19295
rect 19993 19261 20027 19295
rect 21925 19261 21959 19295
rect 23029 19261 23063 19295
rect 24961 19261 24995 19295
rect 27813 19261 27847 19295
rect 33425 19261 33459 19295
rect 35909 19261 35943 19295
rect 36645 19261 36679 19295
rect 39497 19261 39531 19295
rect 48145 19261 48179 19295
rect 48697 19261 48731 19295
rect 14473 19193 14507 19227
rect 16773 19193 16807 19227
rect 17877 19193 17911 19227
rect 21281 19193 21315 19227
rect 41153 19193 41187 19227
rect 42533 19193 42567 19227
rect 45569 19193 45603 19227
rect 47685 19193 47719 19227
rect 15025 19125 15059 19159
rect 20177 19125 20211 19159
rect 29285 19125 29319 19159
rect 34437 19125 34471 19159
rect 41061 19125 41095 19159
rect 45017 19125 45051 19159
rect 46213 19125 46247 19159
rect 12449 18921 12483 18955
rect 13001 18921 13035 18955
rect 17601 18921 17635 18955
rect 20453 18921 20487 18955
rect 26801 18921 26835 18955
rect 29009 18921 29043 18955
rect 41613 18921 41647 18955
rect 49433 18921 49467 18955
rect 14749 18853 14783 18887
rect 38669 18853 38703 18887
rect 42441 18853 42475 18887
rect 47869 18853 47903 18887
rect 14197 18785 14231 18819
rect 18429 18785 18463 18819
rect 20085 18785 20119 18819
rect 21189 18785 21223 18819
rect 21649 18785 21683 18819
rect 23857 18785 23891 18819
rect 32229 18785 32263 18819
rect 34989 18785 35023 18819
rect 36921 18785 36955 18819
rect 39865 18785 39899 18819
rect 40141 18785 40175 18819
rect 42073 18785 42107 18819
rect 42993 18785 43027 18819
rect 43177 18785 43211 18819
rect 46121 18785 46155 18819
rect 48329 18785 48363 18819
rect 48881 18785 48915 18819
rect 13553 18717 13587 18751
rect 16865 18717 16899 18751
rect 17517 18717 17551 18751
rect 18337 18717 18371 18751
rect 20177 18717 20211 18751
rect 21005 18717 21039 18751
rect 21281 18717 21315 18751
rect 22109 18717 22143 18751
rect 24593 18717 24627 18751
rect 25053 18717 25087 18751
rect 27261 18717 27295 18751
rect 29929 18717 29963 18751
rect 30297 18717 30331 18751
rect 34713 18717 34747 18751
rect 39129 18717 39163 18751
rect 43269 18717 43303 18751
rect 43729 18717 43763 18751
rect 46673 18717 46707 18751
rect 58173 18717 58207 18751
rect 15209 18649 15243 18683
rect 19349 18649 19383 18683
rect 22385 18649 22419 18683
rect 24501 18649 24535 18683
rect 25329 18649 25363 18683
rect 27537 18649 27571 18683
rect 32413 18649 32447 18683
rect 34069 18649 34103 18683
rect 37197 18649 37231 18683
rect 47225 18649 47259 18683
rect 57897 18649 57931 18683
rect 15761 18581 15795 18615
rect 16313 18581 16347 18615
rect 16957 18581 16991 18615
rect 18705 18581 18739 18615
rect 19441 18581 19475 18615
rect 21373 18581 21407 18615
rect 21557 18581 21591 18615
rect 31723 18581 31757 18615
rect 36461 18581 36495 18615
rect 39221 18581 39255 18615
rect 42533 18581 42567 18615
rect 42993 18581 43027 18615
rect 43821 18581 43855 18615
rect 44465 18581 44499 18615
rect 45109 18581 45143 18615
rect 45661 18581 45695 18615
rect 13185 18377 13219 18411
rect 17601 18377 17635 18411
rect 19625 18377 19659 18411
rect 39037 18377 39071 18411
rect 41797 18377 41831 18411
rect 43545 18377 43579 18411
rect 45017 18377 45051 18411
rect 45569 18377 45603 18411
rect 46121 18377 46155 18411
rect 48145 18377 48179 18411
rect 48697 18377 48731 18411
rect 58173 18377 58207 18411
rect 12725 18309 12759 18343
rect 13921 18309 13955 18343
rect 17325 18309 17359 18343
rect 22753 18309 22787 18343
rect 24961 18309 24995 18343
rect 29101 18309 29135 18343
rect 30021 18309 30055 18343
rect 37565 18309 37599 18343
rect 40969 18309 41003 18343
rect 46673 18309 46707 18343
rect 1685 18241 1719 18275
rect 13369 18241 13403 18275
rect 16681 18241 16715 18275
rect 17509 18241 17543 18275
rect 17601 18241 17635 18275
rect 18245 18241 18279 18275
rect 19257 18241 19291 18275
rect 20361 18241 20395 18275
rect 21005 18241 21039 18275
rect 21281 18241 21315 18275
rect 21833 18241 21867 18275
rect 22477 18241 22511 18275
rect 33977 18241 34011 18275
rect 37289 18241 37323 18275
rect 41245 18241 41279 18275
rect 41889 18241 41923 18275
rect 42809 18241 42843 18275
rect 43545 18241 43579 18275
rect 44465 18241 44499 18275
rect 45109 18241 45143 18275
rect 49801 18241 49835 18275
rect 18153 18173 18187 18207
rect 19165 18173 19199 18207
rect 20085 18173 20119 18207
rect 24685 18173 24719 18207
rect 28825 18173 28859 18207
rect 29285 18173 29319 18207
rect 29745 18173 29779 18207
rect 31493 18173 31527 18207
rect 33425 18173 33459 18207
rect 33793 18173 33827 18207
rect 34713 18173 34747 18207
rect 36093 18173 36127 18207
rect 36277 18173 36311 18207
rect 42901 18173 42935 18207
rect 44189 18173 44223 18207
rect 47593 18173 47627 18207
rect 15577 18105 15611 18139
rect 16773 18105 16807 18139
rect 50445 18105 50479 18139
rect 1501 18037 1535 18071
rect 11621 18037 11655 18071
rect 12173 18037 12207 18071
rect 14381 18037 14415 18071
rect 15025 18037 15059 18071
rect 16129 18037 16163 18071
rect 18521 18037 18555 18071
rect 21925 18037 21959 18071
rect 24225 18037 24259 18071
rect 26433 18037 26467 18071
rect 39497 18037 39531 18071
rect 42441 18037 42475 18071
rect 49341 18037 49375 18071
rect 13001 17833 13035 17867
rect 15945 17833 15979 17867
rect 16589 17833 16623 17867
rect 18705 17833 18739 17867
rect 19993 17833 20027 17867
rect 21557 17833 21591 17867
rect 24501 17833 24535 17867
rect 31493 17833 31527 17867
rect 44373 17833 44407 17867
rect 45109 17833 45143 17867
rect 46489 17833 46523 17867
rect 49249 17833 49283 17867
rect 14841 17765 14875 17799
rect 24961 17765 24995 17799
rect 33793 17765 33827 17799
rect 39221 17765 39255 17799
rect 43269 17765 43303 17799
rect 47593 17765 47627 17799
rect 13553 17697 13587 17731
rect 17417 17697 17451 17731
rect 18245 17697 18279 17731
rect 18337 17697 18371 17731
rect 18429 17697 18463 17731
rect 20453 17697 20487 17731
rect 22385 17697 22419 17731
rect 26709 17697 26743 17731
rect 27169 17697 27203 17731
rect 28825 17697 28859 17731
rect 29009 17697 29043 17731
rect 36553 17697 36587 17731
rect 37013 17697 37047 17731
rect 37289 17697 37323 17731
rect 42533 17697 42567 17731
rect 42717 17697 42751 17731
rect 43729 17697 43763 17731
rect 16037 17629 16071 17663
rect 16497 17629 16531 17663
rect 17325 17629 17359 17663
rect 18521 17629 18555 17663
rect 19441 17629 19475 17663
rect 19533 17629 19567 17663
rect 19717 17629 19751 17663
rect 19809 17629 19843 17663
rect 20729 17629 20763 17663
rect 21373 17629 21407 17663
rect 22109 17629 22143 17663
rect 29745 17629 29779 17663
rect 32045 17629 32079 17663
rect 41606 17629 41640 17663
rect 43637 17629 43671 17663
rect 44281 17629 44315 17663
rect 45293 17629 45327 17663
rect 45937 17629 45971 17663
rect 46581 17629 46615 17663
rect 48697 17629 48731 17663
rect 14289 17561 14323 17595
rect 26433 17561 26467 17595
rect 30021 17561 30055 17595
rect 32321 17561 32355 17595
rect 34713 17561 34747 17595
rect 36369 17561 36403 17595
rect 41337 17561 41371 17595
rect 11345 17493 11379 17527
rect 11805 17493 11839 17527
rect 12449 17493 12483 17527
rect 15393 17493 15427 17527
rect 17693 17493 17727 17527
rect 23857 17493 23891 17527
rect 38761 17493 38795 17527
rect 39865 17493 39899 17527
rect 42073 17493 42107 17527
rect 42441 17493 42475 17527
rect 45845 17493 45879 17527
rect 47041 17493 47075 17527
rect 48237 17493 48271 17527
rect 50169 17493 50203 17527
rect 12081 17289 12115 17323
rect 28825 17289 28859 17323
rect 41337 17289 41371 17323
rect 43729 17289 43763 17323
rect 50353 17289 50387 17323
rect 19349 17221 19383 17255
rect 22753 17221 22787 17255
rect 24961 17221 24995 17255
rect 27353 17221 27387 17255
rect 37473 17221 37507 17255
rect 39865 17221 39899 17255
rect 49249 17221 49283 17255
rect 49801 17221 49835 17255
rect 10977 17153 11011 17187
rect 13277 17153 13311 17187
rect 15209 17153 15243 17187
rect 16129 17153 16163 17187
rect 17219 17153 17253 17187
rect 18153 17153 18187 17187
rect 20361 17153 20395 17187
rect 21005 17153 21039 17187
rect 21833 17153 21867 17187
rect 24685 17153 24719 17187
rect 27077 17153 27111 17187
rect 31217 17153 31251 17187
rect 39589 17153 39623 17187
rect 42717 17153 42751 17187
rect 44097 17153 44131 17187
rect 45017 17153 45051 17187
rect 45661 17153 45695 17187
rect 45753 17153 45787 17187
rect 45937 17153 45971 17187
rect 46581 17153 46615 17187
rect 15853 17085 15887 17119
rect 17141 17085 17175 17119
rect 18245 17085 18279 17119
rect 18981 17085 19015 17119
rect 19257 17085 19291 17119
rect 19466 17085 19500 17119
rect 21281 17085 21315 17119
rect 22477 17085 22511 17119
rect 24225 17085 24259 17119
rect 30941 17085 30975 17119
rect 32137 17085 32171 17119
rect 32413 17085 32447 17119
rect 34437 17085 34471 17119
rect 34621 17085 34655 17119
rect 34989 17085 35023 17119
rect 37289 17085 37323 17119
rect 39129 17085 39163 17119
rect 42441 17085 42475 17119
rect 44005 17085 44039 17119
rect 44741 17085 44775 17119
rect 47593 17085 47627 17119
rect 17509 17017 17543 17051
rect 18521 17017 18555 17051
rect 21925 17017 21959 17051
rect 48145 17017 48179 17051
rect 12633 16949 12667 16983
rect 13093 16949 13127 16983
rect 14105 16949 14139 16983
rect 14657 16949 14691 16983
rect 15301 16949 15335 16983
rect 15945 16949 15979 16983
rect 16037 16949 16071 16983
rect 19625 16949 19659 16983
rect 20177 16949 20211 16983
rect 26433 16949 26467 16983
rect 29469 16949 29503 16983
rect 33885 16949 33919 16983
rect 41797 16949 41831 16983
rect 44833 16949 44867 16983
rect 45201 16949 45235 16983
rect 45661 16949 45695 16983
rect 46489 16949 46523 16983
rect 48789 16949 48823 16983
rect 11897 16745 11931 16779
rect 12449 16745 12483 16779
rect 14841 16745 14875 16779
rect 15393 16745 15427 16779
rect 16589 16745 16623 16779
rect 33977 16745 34011 16779
rect 42165 16745 42199 16779
rect 44281 16745 44315 16779
rect 47501 16745 47535 16779
rect 48697 16745 48731 16779
rect 50169 16745 50203 16779
rect 13001 16677 13035 16711
rect 14289 16677 14323 16711
rect 17693 16677 17727 16711
rect 18705 16677 18739 16711
rect 39221 16677 39255 16711
rect 39865 16677 39899 16711
rect 43085 16677 43119 16711
rect 46949 16677 46983 16711
rect 13553 16609 13587 16643
rect 17233 16609 17267 16643
rect 18429 16609 18463 16643
rect 19926 16609 19960 16643
rect 21649 16609 21683 16643
rect 24961 16609 24995 16643
rect 32229 16609 32263 16643
rect 34713 16609 34747 16643
rect 35173 16609 35207 16643
rect 37289 16609 37323 16643
rect 41337 16609 41371 16643
rect 42349 16609 42383 16643
rect 43361 16609 43395 16643
rect 44373 16609 44407 16643
rect 45017 16609 45051 16643
rect 46397 16609 46431 16643
rect 48053 16609 48087 16643
rect 1685 16541 1719 16575
rect 15853 16541 15887 16575
rect 15945 16541 15979 16575
rect 16497 16541 16531 16575
rect 17325 16541 17359 16575
rect 18337 16541 18371 16575
rect 19441 16541 19475 16575
rect 19717 16541 19751 16575
rect 20821 16541 20855 16575
rect 21189 16541 21223 16575
rect 22109 16541 22143 16575
rect 24501 16541 24535 16575
rect 27169 16541 27203 16575
rect 29009 16541 29043 16575
rect 29929 16541 29963 16575
rect 30297 16541 30331 16575
rect 31723 16541 31757 16575
rect 37013 16541 37047 16575
rect 41613 16541 41647 16575
rect 42441 16541 42475 16575
rect 43453 16541 43487 16575
rect 44465 16541 44499 16575
rect 45109 16541 45143 16575
rect 45937 16541 45971 16575
rect 58173 16541 58207 16575
rect 22385 16473 22419 16507
rect 25237 16473 25271 16507
rect 28825 16473 28859 16507
rect 32505 16473 32539 16507
rect 34897 16473 34931 16507
rect 57897 16473 57931 16507
rect 1501 16405 1535 16439
rect 19809 16405 19843 16439
rect 20085 16405 20119 16439
rect 23857 16405 23891 16439
rect 26709 16405 26743 16439
rect 38761 16405 38795 16439
rect 44097 16405 44131 16439
rect 45845 16405 45879 16439
rect 49157 16405 49191 16439
rect 12265 16201 12299 16235
rect 14473 16201 14507 16235
rect 39497 16201 39531 16235
rect 41291 16201 41325 16235
rect 46581 16201 46615 16235
rect 47593 16201 47627 16235
rect 48237 16201 48271 16235
rect 58173 16201 58207 16235
rect 13369 16133 13403 16167
rect 15577 16133 15611 16167
rect 18061 16133 18095 16167
rect 20913 16133 20947 16167
rect 26157 16133 26191 16167
rect 49249 16133 49283 16167
rect 13921 16065 13955 16099
rect 17233 16065 17267 16099
rect 17417 16065 17451 16099
rect 17877 16065 17911 16099
rect 18153 16065 18187 16099
rect 18797 16065 18831 16099
rect 19809 16065 19843 16099
rect 20637 16065 20671 16099
rect 21833 16065 21867 16099
rect 26433 16065 26467 16099
rect 27261 16065 27295 16099
rect 29653 16065 29687 16099
rect 30205 16065 30239 16099
rect 32137 16065 32171 16099
rect 34437 16065 34471 16099
rect 39037 16065 39071 16099
rect 39865 16065 39899 16099
rect 40141 16065 40175 16099
rect 42625 16065 42659 16099
rect 42809 16065 42843 16099
rect 42901 16065 42935 16099
rect 43361 16065 43395 16099
rect 43453 16065 43487 16099
rect 44373 16065 44407 16099
rect 45017 16065 45051 16099
rect 48697 16065 48731 16099
rect 49801 16065 49835 16099
rect 12817 15997 12851 16031
rect 17325 15997 17359 16031
rect 18705 15997 18739 16031
rect 19165 15997 19199 16031
rect 19717 15997 19751 16031
rect 21005 15997 21039 16031
rect 21122 15997 21156 16031
rect 22477 15997 22511 16031
rect 22753 15997 22787 16031
rect 24685 15997 24719 16031
rect 28917 15997 28951 16031
rect 29101 15997 29135 16031
rect 32321 15997 32355 16031
rect 33977 15997 34011 16031
rect 34621 15997 34655 16031
rect 34897 15997 34931 16031
rect 38761 15997 38795 16031
rect 41061 15997 41095 16031
rect 43637 15997 43671 16031
rect 44097 15997 44131 16031
rect 21281 15929 21315 15963
rect 24225 15929 24259 15963
rect 15025 15861 15059 15895
rect 16129 15861 16163 15895
rect 16681 15861 16715 15895
rect 18153 15861 18187 15895
rect 20085 15861 20119 15895
rect 21925 15861 21959 15895
rect 31493 15861 31527 15895
rect 37289 15861 37323 15895
rect 42441 15861 42475 15895
rect 43545 15861 43579 15895
rect 44189 15861 44223 15895
rect 44281 15861 44315 15895
rect 44925 15861 44959 15895
rect 45569 15861 45603 15895
rect 46029 15861 46063 15895
rect 15117 15657 15151 15691
rect 15669 15657 15703 15691
rect 16221 15657 16255 15691
rect 21925 15657 21959 15691
rect 24409 15657 24443 15691
rect 25053 15657 25087 15691
rect 39221 15657 39255 15691
rect 41705 15657 41739 15691
rect 42533 15657 42567 15691
rect 43361 15657 43395 15691
rect 45017 15657 45051 15691
rect 45569 15657 45603 15691
rect 47317 15657 47351 15691
rect 47777 15657 47811 15691
rect 48881 15657 48915 15691
rect 49433 15657 49467 15691
rect 13553 15589 13587 15623
rect 16773 15589 16807 15623
rect 20361 15589 20395 15623
rect 29009 15589 29043 15623
rect 38669 15589 38703 15623
rect 42625 15589 42659 15623
rect 43269 15589 43303 15623
rect 19625 15521 19659 15555
rect 20913 15521 20947 15555
rect 26801 15521 26835 15555
rect 27537 15521 27571 15555
rect 31861 15521 31895 15555
rect 36921 15521 36955 15555
rect 41061 15521 41095 15555
rect 46121 15521 46155 15555
rect 11437 15453 11471 15487
rect 14565 15453 14599 15487
rect 17785 15453 17819 15487
rect 19533 15453 19567 15487
rect 20637 15453 20671 15487
rect 20729 15453 20763 15487
rect 21373 15453 21407 15487
rect 21649 15453 21683 15487
rect 21793 15453 21827 15487
rect 23121 15453 23155 15487
rect 23765 15453 23799 15487
rect 24593 15453 24627 15487
rect 27261 15453 27295 15487
rect 32321 15453 32355 15487
rect 36461 15453 36495 15487
rect 39129 15453 39163 15487
rect 40141 15453 40175 15487
rect 40785 15453 40819 15487
rect 41981 15453 42015 15487
rect 42717 15453 42751 15487
rect 43177 15453 43211 15487
rect 44097 15453 44131 15487
rect 58173 15453 58207 15487
rect 11989 15385 12023 15419
rect 18521 15385 18555 15419
rect 21557 15385 21591 15419
rect 26525 15385 26559 15419
rect 31585 15385 31619 15419
rect 32505 15385 32539 15419
rect 34161 15385 34195 15419
rect 36185 15385 36219 15419
rect 37197 15385 37231 15419
rect 39865 15385 39899 15419
rect 42441 15385 42475 15419
rect 43453 15385 43487 15419
rect 57897 15385 57931 15419
rect 11253 15317 11287 15351
rect 13001 15317 13035 15351
rect 17325 15317 17359 15351
rect 17877 15317 17911 15351
rect 18613 15317 18647 15351
rect 19901 15317 19935 15351
rect 20545 15317 20579 15351
rect 22937 15317 22971 15351
rect 30113 15317 30147 15351
rect 34713 15317 34747 15351
rect 41521 15317 41555 15351
rect 44005 15317 44039 15351
rect 46673 15317 46707 15351
rect 48329 15317 48363 15351
rect 13829 15113 13863 15147
rect 15025 15113 15059 15147
rect 16129 15113 16163 15147
rect 21281 15113 21315 15147
rect 22477 15113 22511 15147
rect 27077 15113 27111 15147
rect 43545 15113 43579 15147
rect 44189 15113 44223 15147
rect 46397 15113 46431 15147
rect 47593 15113 47627 15147
rect 14473 15045 14507 15079
rect 17969 15045 18003 15079
rect 19165 15045 19199 15079
rect 29009 15045 29043 15079
rect 29929 15045 29963 15079
rect 32321 15045 32355 15079
rect 42865 15045 42899 15079
rect 46949 15045 46983 15079
rect 58173 15045 58207 15079
rect 1685 14977 1719 15011
rect 17325 14977 17359 15011
rect 18429 14977 18463 15011
rect 19073 14977 19107 15011
rect 19257 14977 19291 15011
rect 19901 14977 19935 15011
rect 20991 14977 21025 15011
rect 22569 14977 22603 15011
rect 23673 14977 23707 15011
rect 29285 14977 29319 15011
rect 32137 14977 32171 15011
rect 34437 14977 34471 15011
rect 37565 14977 37599 15011
rect 38209 14977 38243 15011
rect 39221 14977 39255 15011
rect 39865 14977 39899 15011
rect 40141 14977 40175 15011
rect 40969 14977 41003 15011
rect 41613 14977 41647 15011
rect 43729 14977 43763 15011
rect 44741 14977 44775 15011
rect 45845 14977 45879 15011
rect 16865 14909 16899 14943
rect 18521 14909 18555 14943
rect 19993 14909 20027 14943
rect 20821 14909 20855 14943
rect 22385 14909 22419 14943
rect 23397 14909 23431 14943
rect 24685 14909 24719 14943
rect 24961 14909 24995 14943
rect 29745 14909 29779 14943
rect 30389 14909 30423 14943
rect 32597 14909 32631 14943
rect 34713 14909 34747 14943
rect 37289 14909 37323 14943
rect 38945 14909 38979 14943
rect 40877 14909 40911 14943
rect 41705 14909 41739 14943
rect 41889 14909 41923 14943
rect 1501 14841 1535 14875
rect 15577 14841 15611 14875
rect 45293 14841 45327 14875
rect 20177 14773 20211 14807
rect 22937 14773 22971 14807
rect 26433 14773 26467 14807
rect 27537 14773 27571 14807
rect 36185 14773 36219 14807
rect 36645 14773 36679 14807
rect 38393 14773 38427 14807
rect 40693 14773 40727 14807
rect 41797 14773 41831 14807
rect 42993 14773 43027 14807
rect 48145 14773 48179 14807
rect 14289 14569 14323 14603
rect 15393 14569 15427 14603
rect 15853 14569 15887 14603
rect 17601 14569 17635 14603
rect 19717 14569 19751 14603
rect 24501 14569 24535 14603
rect 38669 14569 38703 14603
rect 41061 14569 41095 14603
rect 42901 14569 42935 14603
rect 45017 14569 45051 14603
rect 46673 14569 46707 14603
rect 18705 14501 18739 14535
rect 20361 14501 20395 14535
rect 20453 14501 20487 14535
rect 23259 14501 23293 14535
rect 26801 14501 26835 14535
rect 27261 14501 27295 14535
rect 36461 14501 36495 14535
rect 39865 14501 39899 14535
rect 43545 14501 43579 14535
rect 20269 14433 20303 14467
rect 21097 14433 21131 14467
rect 22293 14433 22327 14467
rect 22569 14433 22603 14467
rect 25329 14433 25363 14467
rect 29009 14433 29043 14467
rect 30849 14433 30883 14467
rect 31033 14433 31067 14467
rect 33701 14433 33735 14467
rect 39037 14433 39071 14467
rect 40785 14433 40819 14467
rect 44005 14433 44039 14467
rect 10793 14365 10827 14399
rect 19625 14365 19659 14399
rect 20544 14365 20578 14399
rect 21267 14365 21301 14399
rect 22201 14365 22235 14399
rect 23029 14365 23063 14399
rect 24593 14365 24627 14399
rect 25053 14365 25087 14399
rect 29561 14365 29595 14399
rect 29837 14365 29871 14399
rect 32689 14365 32723 14399
rect 33977 14365 34011 14399
rect 34713 14365 34747 14399
rect 36921 14365 36955 14399
rect 37197 14365 37231 14399
rect 37841 14365 37875 14399
rect 38867 14365 38901 14399
rect 40049 14365 40083 14399
rect 40141 14365 40175 14399
rect 40233 14365 40267 14399
rect 40969 14365 41003 14399
rect 41061 14365 41095 14399
rect 41705 14365 41739 14399
rect 42257 14365 42291 14399
rect 18153 14297 18187 14331
rect 28733 14297 28767 14331
rect 34989 14297 35023 14331
rect 38117 14297 38151 14331
rect 47225 14297 47259 14331
rect 47777 14297 47811 14331
rect 10609 14229 10643 14263
rect 11345 14229 11379 14263
rect 14841 14229 14875 14263
rect 16405 14229 16439 14263
rect 17049 14229 17083 14263
rect 21557 14229 21591 14263
rect 41613 14229 41647 14263
rect 42349 14229 42383 14263
rect 45569 14229 45603 14263
rect 46121 14229 46155 14263
rect 16129 14025 16163 14059
rect 17785 14025 17819 14059
rect 18337 14025 18371 14059
rect 19441 14025 19475 14059
rect 21833 14025 21867 14059
rect 29653 14025 29687 14059
rect 36737 14025 36771 14059
rect 39957 14025 39991 14059
rect 42993 14025 43027 14059
rect 44189 14025 44223 14059
rect 46305 14025 46339 14059
rect 17233 13957 17267 13991
rect 18889 13957 18923 13991
rect 21281 13957 21315 13991
rect 27721 13957 27755 13991
rect 34621 13957 34655 13991
rect 45201 13957 45235 13991
rect 45845 13957 45879 13991
rect 1685 13889 1719 13923
rect 15577 13889 15611 13923
rect 20545 13889 20579 13923
rect 21005 13889 21039 13923
rect 22201 13889 22235 13923
rect 22845 13889 22879 13923
rect 23857 13889 23891 13923
rect 23949 13889 23983 13923
rect 24133 13889 24167 13923
rect 24225 13889 24259 13923
rect 24685 13889 24719 13923
rect 27445 13889 27479 13923
rect 34345 13889 34379 13923
rect 36553 13889 36587 13923
rect 37565 13889 37599 13923
rect 38209 13889 38243 13923
rect 39313 13889 39347 13923
rect 40233 13889 40267 13923
rect 40785 13889 40819 13923
rect 40969 13889 41003 13923
rect 41613 13889 41647 13923
rect 43637 13889 43671 13923
rect 20453 13821 20487 13855
rect 21281 13821 21315 13855
rect 22109 13821 22143 13855
rect 22753 13821 22787 13855
rect 23213 13821 23247 13855
rect 26433 13821 26467 13855
rect 29193 13821 29227 13855
rect 31401 13821 31435 13855
rect 32137 13821 32171 13855
rect 33885 13821 33919 13855
rect 37289 13821 37323 13855
rect 38945 13821 38979 13855
rect 39221 13821 39255 13855
rect 39957 13821 39991 13855
rect 41521 13821 41555 13855
rect 44649 13821 44683 13855
rect 23673 13753 23707 13787
rect 36093 13753 36127 13787
rect 1501 13685 1535 13719
rect 21097 13685 21131 13719
rect 22109 13685 22143 13719
rect 24942 13685 24976 13719
rect 31143 13685 31177 13719
rect 32394 13685 32428 13719
rect 38393 13685 38427 13719
rect 40141 13685 40175 13719
rect 42533 13685 42567 13719
rect 46857 13685 46891 13719
rect 12081 13481 12115 13515
rect 16681 13481 16715 13515
rect 19625 13481 19659 13515
rect 21281 13481 21315 13515
rect 24777 13481 24811 13515
rect 33793 13481 33827 13515
rect 40601 13481 40635 13515
rect 41245 13481 41279 13515
rect 42809 13481 42843 13515
rect 43913 13481 43947 13515
rect 46213 13481 46247 13515
rect 16037 13413 16071 13447
rect 17141 13413 17175 13447
rect 17785 13413 17819 13447
rect 27261 13413 27295 13447
rect 38025 13413 38059 13447
rect 39957 13413 39991 13447
rect 45569 13413 45603 13447
rect 23581 13345 23615 13379
rect 25421 13345 25455 13379
rect 26249 13345 26283 13379
rect 30113 13345 30147 13379
rect 32321 13345 32355 13379
rect 36369 13345 36403 13379
rect 38301 13345 38335 13379
rect 45109 13345 45143 13379
rect 11529 13277 11563 13311
rect 20177 13277 20211 13311
rect 21373 13277 21407 13311
rect 23857 13277 23891 13311
rect 25973 13277 26007 13311
rect 29009 13277 29043 13311
rect 29837 13277 29871 13311
rect 32045 13277 32079 13311
rect 34713 13277 34747 13311
rect 34989 13277 35023 13311
rect 35633 13277 35667 13311
rect 36645 13277 36679 13311
rect 37289 13277 37323 13311
rect 38393 13277 38427 13311
rect 40049 13277 40083 13311
rect 40693 13277 40727 13311
rect 43361 13277 43395 13311
rect 58173 13277 58207 13311
rect 20637 13209 20671 13243
rect 21833 13209 21867 13243
rect 25237 13209 25271 13243
rect 28733 13209 28767 13243
rect 35909 13209 35943 13243
rect 37565 13209 37599 13243
rect 39221 13209 39255 13243
rect 41705 13209 41739 13243
rect 57897 13209 57931 13243
rect 11345 13141 11379 13175
rect 18245 13141 18279 13175
rect 25145 13141 25179 13175
rect 31585 13141 31619 13175
rect 39129 13141 39163 13175
rect 42257 13141 42291 13175
rect 18521 12937 18555 12971
rect 20085 12937 20119 12971
rect 21281 12937 21315 12971
rect 22385 12937 22419 12971
rect 26433 12937 26467 12971
rect 29101 12937 29135 12971
rect 31309 12937 31343 12971
rect 37289 12937 37323 12971
rect 38485 12937 38519 12971
rect 39773 12937 39807 12971
rect 41061 12937 41095 12971
rect 41613 12937 41647 12971
rect 42533 12937 42567 12971
rect 58173 12937 58207 12971
rect 17969 12869 18003 12903
rect 19625 12869 19659 12903
rect 23121 12869 23155 12903
rect 32413 12869 32447 12903
rect 39129 12869 39163 12903
rect 43545 12869 43579 12903
rect 20729 12801 20763 12835
rect 22477 12801 22511 12835
rect 22937 12801 22971 12835
rect 23213 12801 23247 12835
rect 23857 12801 23891 12835
rect 25053 12801 25087 12835
rect 25697 12801 25731 12835
rect 25881 12801 25915 12835
rect 26182 12801 26216 12835
rect 34621 12801 34655 12835
rect 35265 12801 35299 12835
rect 36277 12801 36311 12835
rect 36553 12801 36587 12835
rect 37657 12801 37691 12835
rect 38301 12801 38335 12835
rect 38577 12801 38611 12835
rect 39037 12801 39071 12835
rect 39865 12801 39899 12835
rect 40509 12801 40543 12835
rect 18981 12733 19015 12767
rect 23765 12733 23799 12767
rect 24961 12733 24995 12767
rect 27353 12733 27387 12767
rect 27629 12733 27663 12767
rect 29561 12733 29595 12767
rect 29837 12733 29871 12767
rect 32137 12733 32171 12767
rect 33885 12733 33919 12767
rect 34345 12733 34379 12767
rect 36461 12733 36495 12767
rect 37565 12733 37599 12767
rect 42993 12733 43027 12767
rect 24685 12665 24719 12699
rect 25973 12665 26007 12699
rect 36093 12665 36127 12699
rect 38301 12665 38335 12699
rect 44189 12665 44223 12699
rect 16865 12597 16899 12631
rect 17417 12597 17451 12631
rect 23213 12597 23247 12631
rect 24133 12597 24167 12631
rect 26065 12597 26099 12631
rect 35449 12597 35483 12631
rect 36277 12597 36311 12631
rect 44649 12597 44683 12631
rect 45201 12597 45235 12631
rect 12909 12393 12943 12427
rect 18705 12393 18739 12427
rect 19717 12393 19751 12427
rect 20913 12393 20947 12427
rect 21925 12393 21959 12427
rect 25789 12393 25823 12427
rect 26801 12393 26835 12427
rect 29009 12393 29043 12427
rect 36277 12393 36311 12427
rect 36461 12393 36495 12427
rect 37933 12393 37967 12427
rect 41521 12393 41555 12427
rect 43269 12393 43303 12427
rect 20361 12325 20395 12359
rect 22385 12325 22419 12359
rect 24777 12325 24811 12359
rect 31493 12325 31527 12359
rect 39865 12325 39899 12359
rect 40417 12325 40451 12359
rect 42717 12325 42751 12359
rect 23029 12257 23063 12291
rect 24593 12257 24627 12291
rect 25513 12257 25547 12291
rect 26341 12257 26375 12291
rect 36093 12257 36127 12291
rect 1685 12189 1719 12223
rect 12357 12189 12391 12223
rect 22937 12189 22971 12223
rect 23121 12189 23155 12223
rect 23581 12189 23615 12223
rect 24409 12189 24443 12223
rect 24501 12189 24535 12223
rect 24777 12189 24811 12223
rect 25421 12189 25455 12223
rect 26433 12189 26467 12223
rect 27261 12189 27295 12223
rect 29745 12189 29779 12223
rect 31953 12189 31987 12223
rect 34713 12189 34747 12223
rect 34989 12189 35023 12223
rect 36277 12189 36311 12223
rect 37197 12189 37231 12223
rect 37933 12189 37967 12223
rect 38669 12189 38703 12223
rect 27537 12121 27571 12155
rect 30021 12121 30055 12155
rect 32229 12121 32263 12155
rect 36001 12121 36035 12155
rect 1501 12053 1535 12087
rect 12173 12053 12207 12087
rect 18153 12053 18187 12087
rect 23765 12053 23799 12087
rect 33701 12053 33735 12087
rect 37105 12053 37139 12087
rect 38577 12053 38611 12087
rect 39129 12053 39163 12087
rect 40969 12053 41003 12087
rect 42073 12053 42107 12087
rect 43729 12053 43763 12087
rect 44373 12053 44407 12087
rect 21925 11849 21959 11883
rect 23029 11849 23063 11883
rect 36093 11849 36127 11883
rect 36645 11849 36679 11883
rect 38025 11849 38059 11883
rect 38761 11849 38795 11883
rect 39313 11849 39347 11883
rect 40325 11849 40359 11883
rect 40877 11849 40911 11883
rect 41429 11849 41463 11883
rect 42533 11849 42567 11883
rect 20545 11781 20579 11815
rect 23673 11781 23707 11815
rect 32413 11781 32447 11815
rect 20453 11713 20487 11747
rect 22477 11713 22511 11747
rect 23581 11713 23615 11747
rect 23765 11713 23799 11747
rect 24409 11713 24443 11747
rect 25053 11713 25087 11747
rect 26065 11713 26099 11747
rect 27997 11713 28031 11747
rect 28733 11713 28767 11747
rect 29837 11713 29871 11747
rect 32137 11713 32171 11747
rect 34621 11713 34655 11747
rect 35633 11713 35667 11747
rect 35909 11713 35943 11747
rect 36737 11713 36771 11747
rect 37289 11713 37323 11747
rect 37473 11713 37507 11747
rect 38117 11713 38151 11747
rect 42993 11713 43027 11747
rect 43545 11713 43579 11747
rect 19809 11645 19843 11679
rect 25145 11645 25179 11679
rect 25973 11645 26007 11679
rect 30113 11645 30147 11679
rect 34345 11645 34379 11679
rect 35725 11645 35759 11679
rect 26433 11577 26467 11611
rect 39865 11577 39899 11611
rect 18613 11509 18647 11543
rect 19257 11509 19291 11543
rect 21005 11509 21039 11543
rect 24225 11509 24259 11543
rect 25421 11509 25455 11543
rect 29285 11509 29319 11543
rect 31585 11509 31619 11543
rect 33885 11509 33919 11543
rect 35633 11509 35667 11543
rect 37381 11509 37415 11543
rect 19901 11305 19935 11339
rect 21557 11305 21591 11339
rect 22201 11305 22235 11339
rect 22753 11305 22787 11339
rect 23857 11305 23891 11339
rect 25605 11305 25639 11339
rect 27261 11305 27295 11339
rect 27445 11305 27479 11339
rect 28825 11305 28859 11339
rect 34805 11305 34839 11339
rect 35817 11305 35851 11339
rect 36645 11305 36679 11339
rect 38301 11305 38335 11339
rect 38853 11305 38887 11339
rect 39865 11305 39899 11339
rect 42717 11305 42751 11339
rect 20453 11237 20487 11271
rect 26801 11237 26835 11271
rect 27813 11237 27847 11271
rect 28273 11237 28307 11271
rect 37749 11237 37783 11271
rect 26341 11169 26375 11203
rect 30297 11169 30331 11203
rect 30573 11169 30607 11203
rect 34161 11169 34195 11203
rect 35173 11169 35207 11203
rect 41521 11169 41555 11203
rect 19349 11101 19383 11135
rect 23305 11101 23339 11135
rect 25053 11101 25087 11135
rect 26433 11101 26467 11135
rect 28549 11101 28583 11135
rect 28641 11101 28675 11135
rect 28733 11101 28767 11135
rect 29009 11101 29043 11135
rect 31033 11101 31067 11135
rect 33885 11101 33919 11135
rect 34713 11101 34747 11135
rect 34989 11101 35023 11135
rect 36461 11101 36495 11135
rect 37297 11103 37331 11137
rect 40417 11101 40451 11135
rect 41061 11101 41095 11135
rect 58173 11101 58207 11135
rect 21097 11033 21131 11067
rect 24961 11033 24995 11067
rect 25697 11033 25731 11067
rect 27445 11033 27479 11067
rect 31309 11033 31343 11067
rect 35633 11033 35667 11067
rect 37197 11033 37231 11067
rect 42073 11033 42107 11067
rect 57897 11033 57931 11067
rect 32781 10965 32815 10999
rect 35833 10965 35867 10999
rect 36001 10965 36035 10999
rect 20729 10761 20763 10795
rect 21281 10761 21315 10795
rect 22661 10761 22695 10795
rect 23213 10761 23247 10795
rect 23765 10761 23799 10795
rect 28917 10761 28951 10795
rect 36277 10761 36311 10795
rect 37841 10761 37875 10795
rect 40693 10761 40727 10795
rect 41245 10761 41279 10795
rect 41797 10761 41831 10795
rect 58173 10761 58207 10795
rect 24317 10693 24351 10727
rect 25605 10693 25639 10727
rect 31309 10693 31343 10727
rect 33333 10693 33367 10727
rect 35081 10693 35115 10727
rect 38393 10693 38427 10727
rect 40141 10693 40175 10727
rect 34851 10659 34885 10693
rect 1685 10625 1719 10659
rect 11713 10625 11747 10659
rect 24777 10625 24811 10659
rect 24961 10625 24995 10659
rect 26341 10625 26375 10659
rect 27629 10625 27663 10659
rect 30205 10625 30239 10659
rect 31585 10625 31619 10659
rect 32413 10625 32447 10659
rect 33057 10625 33091 10659
rect 33977 10625 34011 10659
rect 34253 10625 34287 10659
rect 35725 10625 35759 10659
rect 36369 10625 36403 10659
rect 38945 10625 38979 10659
rect 12265 10557 12299 10591
rect 25421 10557 25455 10591
rect 27721 10557 27755 10591
rect 32137 10557 32171 10591
rect 34069 10557 34103 10591
rect 37289 10557 37323 10591
rect 22109 10489 22143 10523
rect 26157 10489 26191 10523
rect 27997 10489 28031 10523
rect 30849 10489 30883 10523
rect 33793 10489 33827 10523
rect 34713 10489 34747 10523
rect 35541 10489 35575 10523
rect 1501 10421 1535 10455
rect 11529 10421 11563 10455
rect 20177 10421 20211 10455
rect 24869 10421 24903 10455
rect 33977 10421 34011 10455
rect 34897 10421 34931 10455
rect 39497 10421 39531 10455
rect 21005 10217 21039 10251
rect 21557 10217 21591 10251
rect 22201 10217 22235 10251
rect 23765 10217 23799 10251
rect 24593 10217 24627 10251
rect 26249 10217 26283 10251
rect 27077 10217 27111 10251
rect 28457 10217 28491 10251
rect 38393 10217 38427 10251
rect 39957 10217 39991 10251
rect 41061 10217 41095 10251
rect 25329 10149 25363 10183
rect 27813 10149 27847 10183
rect 27997 10149 28031 10183
rect 34989 10149 35023 10183
rect 23213 10081 23247 10115
rect 27629 10081 27663 10115
rect 28733 10081 28767 10115
rect 29745 10081 29779 10115
rect 30021 10081 30055 10115
rect 31953 10081 31987 10115
rect 36185 10081 36219 10115
rect 38945 10081 38979 10115
rect 26249 10013 26283 10047
rect 26893 10013 26927 10047
rect 27721 10013 27755 10047
rect 28825 10013 28859 10047
rect 32229 10013 32263 10047
rect 32873 10013 32907 10047
rect 33885 10013 33919 10047
rect 34805 10013 34839 10047
rect 35449 10013 35483 10047
rect 35633 10013 35667 10047
rect 36277 10013 36311 10047
rect 37841 10013 37875 10047
rect 58081 10013 58115 10047
rect 22753 9945 22787 9979
rect 27997 9945 28031 9979
rect 33149 9945 33183 9979
rect 33609 9945 33643 9979
rect 57529 9945 57563 9979
rect 31493 9877 31527 9911
rect 33793 9877 33827 9911
rect 33977 9877 34011 9911
rect 34161 9877 34195 9911
rect 35449 9877 35483 9911
rect 36829 9877 36863 9911
rect 37289 9877 37323 9911
rect 40417 9877 40451 9911
rect 24685 9673 24719 9707
rect 28273 9673 28307 9707
rect 28457 9673 28491 9707
rect 28641 9673 28675 9707
rect 58173 9673 58207 9707
rect 11621 9605 11655 9639
rect 22753 9605 22787 9639
rect 27445 9605 27479 9639
rect 27629 9605 27663 9639
rect 32321 9605 32355 9639
rect 32505 9605 32539 9639
rect 33609 9605 33643 9639
rect 33793 9605 33827 9639
rect 35725 9605 35759 9639
rect 36369 9605 36403 9639
rect 10609 9537 10643 9571
rect 26157 9537 26191 9571
rect 26249 9537 26283 9571
rect 28089 9537 28123 9571
rect 28365 9537 28399 9571
rect 29285 9537 29319 9571
rect 30113 9537 30147 9571
rect 31125 9537 31159 9571
rect 32413 9537 32447 9571
rect 33977 9537 34011 9571
rect 34437 9537 34471 9571
rect 34621 9537 34655 9571
rect 35265 9537 35299 9571
rect 25145 9469 25179 9503
rect 29101 9469 29135 9503
rect 30021 9469 30055 9503
rect 31033 9469 31067 9503
rect 30481 9401 30515 9435
rect 31493 9401 31527 9435
rect 32689 9401 32723 9435
rect 39497 9401 39531 9435
rect 40049 9401 40083 9435
rect 10425 9333 10459 9367
rect 22201 9333 22235 9367
rect 23305 9333 23339 9367
rect 24133 9333 24167 9367
rect 29469 9333 29503 9367
rect 32137 9333 32171 9367
rect 34529 9333 34563 9367
rect 35173 9333 35207 9367
rect 37289 9333 37323 9367
rect 37933 9333 37967 9367
rect 38485 9333 38519 9367
rect 38945 9333 38979 9367
rect 24961 9129 24995 9163
rect 26525 9129 26559 9163
rect 27721 9129 27755 9163
rect 28825 9129 28859 9163
rect 29745 9129 29779 9163
rect 31585 9129 31619 9163
rect 32505 9129 32539 9163
rect 33333 9129 33367 9163
rect 33977 9129 34011 9163
rect 35265 9129 35299 9163
rect 37473 9129 37507 9163
rect 26065 9061 26099 9095
rect 30941 9061 30975 9095
rect 38025 9061 38059 9095
rect 28273 8993 28307 9027
rect 30665 8993 30699 9027
rect 31769 8993 31803 9027
rect 33149 8993 33183 9027
rect 34713 8993 34747 9027
rect 35909 8993 35943 9027
rect 1685 8925 1719 8959
rect 25421 8925 25455 8959
rect 27169 8925 27203 8959
rect 28825 8925 28859 8959
rect 30573 8925 30607 8959
rect 31592 8925 31626 8959
rect 31861 8925 31895 8959
rect 32321 8925 32355 8959
rect 33425 8925 33459 8959
rect 34069 8925 34103 8959
rect 29791 8891 29825 8925
rect 29561 8857 29595 8891
rect 36369 8857 36403 8891
rect 36921 8857 36955 8891
rect 38577 8857 38611 8891
rect 39129 8857 39163 8891
rect 1501 8789 1535 8823
rect 22753 8789 22787 8823
rect 23305 8789 23339 8823
rect 23857 8789 23891 8823
rect 29929 8789 29963 8823
rect 31401 8789 31435 8823
rect 33149 8789 33183 8823
rect 24593 8585 24627 8619
rect 25145 8585 25179 8619
rect 26341 8585 26375 8619
rect 27077 8585 27111 8619
rect 27629 8585 27663 8619
rect 28181 8585 28215 8619
rect 28733 8585 28767 8619
rect 32321 8585 32355 8619
rect 33609 8585 33643 8619
rect 34161 8585 34195 8619
rect 35173 8585 35207 8619
rect 36369 8585 36403 8619
rect 37381 8585 37415 8619
rect 31125 8517 31159 8551
rect 31341 8517 31375 8551
rect 35725 8517 35759 8551
rect 38485 8517 38519 8551
rect 25789 8449 25823 8483
rect 28825 8449 28859 8483
rect 29469 8449 29503 8483
rect 30297 8449 30331 8483
rect 32137 8449 32171 8483
rect 32873 8449 32907 8483
rect 24041 8381 24075 8415
rect 29377 8381 29411 8415
rect 29837 8381 29871 8415
rect 30389 8381 30423 8415
rect 30665 8313 30699 8347
rect 31493 8313 31527 8347
rect 32965 8313 32999 8347
rect 30481 8245 30515 8279
rect 31309 8245 31343 8279
rect 34713 8245 34747 8279
rect 37841 8245 37875 8279
rect 24869 8041 24903 8075
rect 25973 8041 26007 8075
rect 26525 8041 26559 8075
rect 27261 8041 27295 8075
rect 27905 8041 27939 8075
rect 29653 8041 29687 8075
rect 31217 8041 31251 8075
rect 32965 8041 32999 8075
rect 33609 8041 33643 8075
rect 28365 7973 28399 8007
rect 30389 7973 30423 8007
rect 35909 7973 35943 8007
rect 30297 7905 30331 7939
rect 31861 7905 31895 7939
rect 34161 7905 34195 7939
rect 57897 7905 57931 7939
rect 29837 7837 29871 7871
rect 30481 7837 30515 7871
rect 30572 7847 30606 7881
rect 31125 7837 31159 7871
rect 31769 7837 31803 7871
rect 58173 7837 58207 7871
rect 14473 7769 14507 7803
rect 14657 7769 14691 7803
rect 32413 7769 32447 7803
rect 34713 7769 34747 7803
rect 35265 7769 35299 7803
rect 37473 7769 37507 7803
rect 15301 7701 15335 7735
rect 25513 7701 25547 7735
rect 29009 7701 29043 7735
rect 36369 7701 36403 7735
rect 36921 7701 36955 7735
rect 25881 7497 25915 7531
rect 27353 7497 27387 7531
rect 27905 7497 27939 7531
rect 28549 7497 28583 7531
rect 29101 7497 29135 7531
rect 30389 7497 30423 7531
rect 31033 7497 31067 7531
rect 32137 7497 32171 7531
rect 32689 7497 32723 7531
rect 33885 7497 33919 7531
rect 34989 7497 35023 7531
rect 36093 7497 36127 7531
rect 58173 7497 58207 7531
rect 29745 7429 29779 7463
rect 33241 7429 33275 7463
rect 1685 7361 1719 7395
rect 29837 7361 29871 7395
rect 30297 7361 30331 7395
rect 31125 7361 31159 7395
rect 36553 7225 36587 7259
rect 1501 7157 1535 7191
rect 26433 7157 26467 7191
rect 34437 7157 34471 7191
rect 35449 7157 35483 7191
rect 31033 6953 31067 6987
rect 31585 6953 31619 6987
rect 32689 6953 32723 6987
rect 30481 6817 30515 6851
rect 33885 6817 33919 6851
rect 34713 6817 34747 6851
rect 29009 6749 29043 6783
rect 32229 6749 32263 6783
rect 27261 6681 27295 6715
rect 27905 6681 27939 6715
rect 29929 6681 29963 6715
rect 26249 6613 26283 6647
rect 26801 6613 26835 6647
rect 33333 6613 33367 6647
rect 35357 6613 35391 6647
rect 35909 6613 35943 6647
rect 28273 6409 28307 6443
rect 30205 6409 30239 6443
rect 30665 6409 30699 6443
rect 32137 6409 32171 6443
rect 32781 6409 32815 6443
rect 34437 6409 34471 6443
rect 34989 6409 35023 6443
rect 28733 6341 28767 6375
rect 29285 6341 29319 6375
rect 33241 6273 33275 6307
rect 33793 6273 33827 6307
rect 35449 6273 35483 6307
rect 31217 6137 31251 6171
rect 27353 6069 27387 6103
rect 28457 5865 28491 5899
rect 29009 5865 29043 5899
rect 29653 5865 29687 5899
rect 30205 5865 30239 5899
rect 30665 5865 30699 5899
rect 31217 5865 31251 5899
rect 32413 5865 32447 5899
rect 32873 5797 32907 5831
rect 33517 5797 33551 5831
rect 34069 5797 34103 5831
rect 31861 5729 31895 5763
rect 1685 5661 1719 5695
rect 13553 5661 13587 5695
rect 58173 5661 58207 5695
rect 57897 5593 57931 5627
rect 1501 5525 1535 5559
rect 13369 5525 13403 5559
rect 14197 5525 14231 5559
rect 29469 5321 29503 5355
rect 30481 5321 30515 5355
rect 58173 5321 58207 5355
rect 32229 5253 32263 5287
rect 28917 5185 28951 5219
rect 30021 5185 30055 5219
rect 29561 4777 29595 4811
rect 58081 4573 58115 4607
rect 57529 4505 57563 4539
rect 58173 4233 58207 4267
rect 1685 4097 1719 4131
rect 2237 3961 2271 3995
rect 1501 3893 1535 3927
rect 40049 3621 40083 3655
rect 39865 3485 39899 3519
rect 40509 3485 40543 3519
rect 1593 3009 1627 3043
rect 37749 3009 37783 3043
rect 37933 2873 37967 2907
rect 1409 2805 1443 2839
rect 4537 2465 4571 2499
rect 7205 2465 7239 2499
rect 1685 2397 1719 2431
rect 3985 2397 4019 2431
rect 6653 2397 6687 2431
rect 18337 2397 18371 2431
rect 30021 2397 30055 2431
rect 30665 2397 30699 2431
rect 37565 2397 37599 2431
rect 42441 2397 42475 2431
rect 54033 2397 54067 2431
rect 57345 2397 57379 2431
rect 19349 2329 19383 2363
rect 56149 2329 56183 2363
rect 1501 2261 1535 2295
rect 3801 2261 3835 2295
rect 6469 2261 6503 2295
rect 18153 2261 18187 2295
rect 30205 2261 30239 2295
rect 42625 2261 42659 2295
rect 54217 2261 54251 2295
rect 57897 2261 57931 2295
<< metal1 >>
rect 17218 28160 17224 28212
rect 17276 28200 17282 28212
rect 32306 28200 32312 28212
rect 17276 28172 32312 28200
rect 17276 28160 17282 28172
rect 32306 28160 32312 28172
rect 32364 28160 32370 28212
rect 14642 28092 14648 28144
rect 14700 28132 14706 28144
rect 38194 28132 38200 28144
rect 14700 28104 38200 28132
rect 14700 28092 14706 28104
rect 38194 28092 38200 28104
rect 38252 28132 38258 28144
rect 41414 28132 41420 28144
rect 38252 28104 41420 28132
rect 38252 28092 38258 28104
rect 41414 28092 41420 28104
rect 41472 28092 41478 28144
rect 18782 28024 18788 28076
rect 18840 28064 18846 28076
rect 32858 28064 32864 28076
rect 18840 28036 32864 28064
rect 18840 28024 18846 28036
rect 32858 28024 32864 28036
rect 32916 28024 32922 28076
rect 19058 27956 19064 28008
rect 19116 27996 19122 28008
rect 37458 27996 37464 28008
rect 19116 27968 37464 27996
rect 19116 27956 19122 27968
rect 37458 27956 37464 27968
rect 37516 27956 37522 28008
rect 23934 27888 23940 27940
rect 23992 27928 23998 27940
rect 44266 27928 44272 27940
rect 23992 27900 44272 27928
rect 23992 27888 23998 27900
rect 44266 27888 44272 27900
rect 44324 27888 44330 27940
rect 14090 27820 14096 27872
rect 14148 27860 14154 27872
rect 37366 27860 37372 27872
rect 14148 27832 37372 27860
rect 14148 27820 14154 27832
rect 37366 27820 37372 27832
rect 37424 27820 37430 27872
rect 1104 27770 58880 27792
rect 1104 27718 10582 27770
rect 10634 27718 10646 27770
rect 10698 27718 10710 27770
rect 10762 27718 10774 27770
rect 10826 27718 10838 27770
rect 10890 27718 29846 27770
rect 29898 27718 29910 27770
rect 29962 27718 29974 27770
rect 30026 27718 30038 27770
rect 30090 27718 30102 27770
rect 30154 27718 49110 27770
rect 49162 27718 49174 27770
rect 49226 27718 49238 27770
rect 49290 27718 49302 27770
rect 49354 27718 49366 27770
rect 49418 27718 58880 27770
rect 1104 27696 58880 27718
rect 30282 27616 30288 27668
rect 30340 27656 30346 27668
rect 39850 27656 39856 27668
rect 30340 27628 39856 27656
rect 30340 27616 30346 27628
rect 39850 27616 39856 27628
rect 39908 27616 39914 27668
rect 1486 27588 1492 27600
rect 1447 27560 1492 27588
rect 1486 27548 1492 27560
rect 1544 27548 1550 27600
rect 2774 27548 2780 27600
rect 2832 27588 2838 27600
rect 2869 27591 2927 27597
rect 2869 27588 2881 27591
rect 2832 27560 2881 27588
rect 2832 27548 2838 27560
rect 2869 27557 2881 27560
rect 2915 27557 2927 27591
rect 2869 27551 2927 27557
rect 8294 27548 8300 27600
rect 8352 27588 8358 27600
rect 9033 27591 9091 27597
rect 9033 27588 9045 27591
rect 8352 27560 9045 27588
rect 8352 27548 8358 27560
rect 9033 27557 9045 27560
rect 9079 27557 9091 27591
rect 9033 27551 9091 27557
rect 20165 27591 20223 27597
rect 20165 27557 20177 27591
rect 20211 27557 20223 27591
rect 20165 27551 20223 27557
rect 14366 27520 14372 27532
rect 6886 27492 14372 27520
rect 1673 27455 1731 27461
rect 1673 27421 1685 27455
rect 1719 27421 1731 27455
rect 1673 27415 1731 27421
rect 3053 27455 3111 27461
rect 3053 27421 3065 27455
rect 3099 27452 3111 27455
rect 3878 27452 3884 27464
rect 3099 27424 3884 27452
rect 3099 27421 3111 27424
rect 3053 27415 3111 27421
rect 1688 27384 1716 27415
rect 3878 27412 3884 27424
rect 3936 27412 3942 27464
rect 6886 27384 6914 27492
rect 14366 27480 14372 27492
rect 14424 27480 14430 27532
rect 9217 27455 9275 27461
rect 9217 27421 9229 27455
rect 9263 27452 9275 27455
rect 9263 27424 9812 27452
rect 9263 27421 9275 27424
rect 9217 27415 9275 27421
rect 1688 27356 6914 27384
rect 9784 27328 9812 27424
rect 13814 27412 13820 27464
rect 13872 27452 13878 27464
rect 14093 27455 14151 27461
rect 14093 27452 14105 27455
rect 13872 27424 14105 27452
rect 13872 27412 13878 27424
rect 14093 27421 14105 27424
rect 14139 27452 14151 27455
rect 14737 27455 14795 27461
rect 14737 27452 14749 27455
rect 14139 27424 14749 27452
rect 14139 27421 14151 27424
rect 14093 27415 14151 27421
rect 14737 27421 14749 27424
rect 14783 27421 14795 27455
rect 19518 27452 19524 27464
rect 19479 27424 19524 27452
rect 14737 27415 14795 27421
rect 19518 27412 19524 27424
rect 19576 27412 19582 27464
rect 19978 27452 19984 27464
rect 19939 27424 19984 27452
rect 19978 27412 19984 27424
rect 20036 27412 20042 27464
rect 20180 27452 20208 27551
rect 24486 27548 24492 27600
rect 24544 27588 24550 27600
rect 24765 27591 24823 27597
rect 24765 27588 24777 27591
rect 24544 27560 24777 27588
rect 24544 27548 24550 27560
rect 24765 27557 24777 27560
rect 24811 27557 24823 27591
rect 24765 27551 24823 27557
rect 30101 27591 30159 27597
rect 30101 27557 30113 27591
rect 30147 27588 30159 27591
rect 30190 27588 30196 27600
rect 30147 27560 30196 27588
rect 30147 27557 30159 27560
rect 30101 27551 30159 27557
rect 30190 27548 30196 27560
rect 30248 27548 30254 27600
rect 30742 27548 30748 27600
rect 30800 27588 30806 27600
rect 33045 27591 33103 27597
rect 33045 27588 33057 27591
rect 30800 27560 33057 27588
rect 30800 27548 30806 27560
rect 33045 27557 33057 27560
rect 33091 27588 33103 27591
rect 35342 27588 35348 27600
rect 33091 27560 35348 27588
rect 33091 27557 33103 27560
rect 33045 27551 33103 27557
rect 35342 27548 35348 27560
rect 35400 27548 35406 27600
rect 35618 27588 35624 27600
rect 35579 27560 35624 27588
rect 35618 27548 35624 27560
rect 35676 27548 35682 27600
rect 51994 27588 52000 27600
rect 51955 27560 52000 27588
rect 51994 27548 52000 27560
rect 52052 27548 52058 27600
rect 33502 27520 33508 27532
rect 26896 27492 33508 27520
rect 24581 27455 24639 27461
rect 24581 27452 24593 27455
rect 20180 27424 24593 27452
rect 24581 27421 24593 27424
rect 24627 27421 24639 27455
rect 24581 27415 24639 27421
rect 18414 27344 18420 27396
rect 18472 27384 18478 27396
rect 19996 27384 20024 27412
rect 20622 27384 20628 27396
rect 18472 27356 19472 27384
rect 19996 27356 20628 27384
rect 18472 27344 18478 27356
rect 3878 27316 3884 27328
rect 3839 27288 3884 27316
rect 3878 27276 3884 27288
rect 3936 27276 3942 27328
rect 9766 27316 9772 27328
rect 9727 27288 9772 27316
rect 9766 27276 9772 27288
rect 9824 27276 9830 27328
rect 14274 27316 14280 27328
rect 14235 27288 14280 27316
rect 14274 27276 14280 27288
rect 14332 27276 14338 27328
rect 19334 27316 19340 27328
rect 19295 27288 19340 27316
rect 19334 27276 19340 27288
rect 19392 27276 19398 27328
rect 19444 27316 19472 27356
rect 20622 27344 20628 27356
rect 20680 27344 20686 27396
rect 26896 27384 26924 27492
rect 33502 27480 33508 27492
rect 33560 27480 33566 27532
rect 36173 27523 36231 27529
rect 36173 27520 36185 27523
rect 34716 27492 36185 27520
rect 28077 27455 28135 27461
rect 28077 27421 28089 27455
rect 28123 27452 28135 27455
rect 28626 27452 28632 27464
rect 28123 27424 28632 27452
rect 28123 27421 28135 27424
rect 28077 27415 28135 27421
rect 28626 27412 28632 27424
rect 28684 27412 28690 27464
rect 30285 27455 30343 27461
rect 30285 27421 30297 27455
rect 30331 27452 30343 27455
rect 30374 27452 30380 27464
rect 30331 27424 30380 27452
rect 30331 27421 30343 27424
rect 30285 27415 30343 27421
rect 30374 27412 30380 27424
rect 30432 27452 30438 27464
rect 34716 27461 34744 27492
rect 36173 27489 36185 27492
rect 36219 27489 36231 27523
rect 36173 27483 36231 27489
rect 34701 27455 34759 27461
rect 34701 27452 34713 27455
rect 30432 27424 34713 27452
rect 30432 27412 30438 27424
rect 34701 27421 34713 27424
rect 34747 27421 34759 27455
rect 35437 27455 35495 27461
rect 35437 27452 35449 27455
rect 34701 27415 34759 27421
rect 34900 27424 35449 27452
rect 20732 27356 26924 27384
rect 27525 27387 27583 27393
rect 20732 27316 20760 27356
rect 27525 27353 27537 27387
rect 27571 27384 27583 27387
rect 29638 27384 29644 27396
rect 27571 27356 29644 27384
rect 27571 27353 27583 27356
rect 27525 27347 27583 27353
rect 29638 27344 29644 27356
rect 29696 27344 29702 27396
rect 32122 27344 32128 27396
rect 32180 27384 32186 27396
rect 33505 27387 33563 27393
rect 33505 27384 33517 27387
rect 32180 27356 33517 27384
rect 32180 27344 32186 27356
rect 33505 27353 33517 27356
rect 33551 27353 33563 27387
rect 34146 27384 34152 27396
rect 34107 27356 34152 27384
rect 33505 27347 33563 27353
rect 34146 27344 34152 27356
rect 34204 27344 34210 27396
rect 25774 27316 25780 27328
rect 19444 27288 20760 27316
rect 25735 27288 25780 27316
rect 25774 27276 25780 27288
rect 25832 27276 25838 27328
rect 26418 27316 26424 27328
rect 26379 27288 26424 27316
rect 26418 27276 26424 27288
rect 26476 27276 26482 27328
rect 28534 27316 28540 27328
rect 28495 27288 28540 27316
rect 28534 27276 28540 27288
rect 28592 27276 28598 27328
rect 31297 27319 31355 27325
rect 31297 27285 31309 27319
rect 31343 27316 31355 27319
rect 31570 27316 31576 27328
rect 31343 27288 31576 27316
rect 31343 27285 31355 27288
rect 31297 27279 31355 27285
rect 31570 27276 31576 27288
rect 31628 27276 31634 27328
rect 32493 27319 32551 27325
rect 32493 27285 32505 27319
rect 32539 27316 32551 27319
rect 32858 27316 32864 27328
rect 32539 27288 32864 27316
rect 32539 27285 32551 27288
rect 32493 27279 32551 27285
rect 32858 27276 32864 27288
rect 32916 27316 32922 27328
rect 33134 27316 33140 27328
rect 32916 27288 33140 27316
rect 32916 27276 32922 27288
rect 33134 27276 33140 27288
rect 33192 27276 33198 27328
rect 34900 27325 34928 27424
rect 35437 27421 35449 27424
rect 35483 27421 35495 27455
rect 35437 27415 35495 27421
rect 40405 27455 40463 27461
rect 40405 27421 40417 27455
rect 40451 27452 40463 27455
rect 40862 27452 40868 27464
rect 40451 27424 40868 27452
rect 40451 27421 40463 27424
rect 40405 27415 40463 27421
rect 40862 27412 40868 27424
rect 40920 27412 40926 27464
rect 45925 27455 45983 27461
rect 45925 27421 45937 27455
rect 45971 27452 45983 27455
rect 46382 27452 46388 27464
rect 45971 27424 46388 27452
rect 45971 27421 45983 27424
rect 45925 27415 45983 27421
rect 46382 27412 46388 27424
rect 46440 27412 46446 27464
rect 46474 27412 46480 27464
rect 46532 27452 46538 27464
rect 51813 27455 51871 27461
rect 51813 27452 51825 27455
rect 46532 27424 51825 27452
rect 46532 27412 46538 27424
rect 51813 27421 51825 27424
rect 51859 27421 51871 27455
rect 51813 27415 51871 27421
rect 52454 27412 52460 27464
rect 52512 27452 52518 27464
rect 56873 27455 56931 27461
rect 56873 27452 56885 27455
rect 52512 27424 56885 27452
rect 52512 27412 52518 27424
rect 56873 27421 56885 27424
rect 56919 27421 56931 27455
rect 57238 27452 57244 27464
rect 57199 27424 57244 27452
rect 56873 27415 56931 27421
rect 57238 27412 57244 27424
rect 57296 27412 57302 27464
rect 57882 27384 57888 27396
rect 57843 27356 57888 27384
rect 57882 27344 57888 27356
rect 57940 27344 57946 27396
rect 58066 27384 58072 27396
rect 58027 27356 58072 27384
rect 58066 27344 58072 27356
rect 58124 27344 58130 27396
rect 34885 27319 34943 27325
rect 34885 27285 34897 27319
rect 34931 27285 34943 27319
rect 41046 27316 41052 27328
rect 41007 27288 41052 27316
rect 34885 27279 34943 27285
rect 41046 27276 41052 27288
rect 41104 27276 41110 27328
rect 46290 27276 46296 27328
rect 46348 27316 46354 27328
rect 46569 27319 46627 27325
rect 46569 27316 46581 27319
rect 46348 27288 46581 27316
rect 46348 27276 46354 27288
rect 46569 27285 46581 27288
rect 46615 27285 46627 27319
rect 46569 27279 46627 27285
rect 1104 27226 58880 27248
rect 1104 27174 20214 27226
rect 20266 27174 20278 27226
rect 20330 27174 20342 27226
rect 20394 27174 20406 27226
rect 20458 27174 20470 27226
rect 20522 27174 39478 27226
rect 39530 27174 39542 27226
rect 39594 27174 39606 27226
rect 39658 27174 39670 27226
rect 39722 27174 39734 27226
rect 39786 27174 58880 27226
rect 1104 27152 58880 27174
rect 1394 27072 1400 27124
rect 1452 27112 1458 27124
rect 1489 27115 1547 27121
rect 1489 27112 1501 27115
rect 1452 27084 1501 27112
rect 1452 27072 1458 27084
rect 1489 27081 1501 27084
rect 1535 27081 1547 27115
rect 1489 27075 1547 27081
rect 9766 27072 9772 27124
rect 9824 27112 9830 27124
rect 9824 27084 19472 27112
rect 9824 27072 9830 27084
rect 1673 26979 1731 26985
rect 1673 26945 1685 26979
rect 1719 26976 1731 26979
rect 14458 26976 14464 26988
rect 1719 26948 14464 26976
rect 1719 26945 1731 26948
rect 1673 26939 1731 26945
rect 14458 26936 14464 26948
rect 14516 26936 14522 26988
rect 19444 26976 19472 27084
rect 19518 27072 19524 27124
rect 19576 27112 19582 27124
rect 20809 27115 20867 27121
rect 20809 27112 20821 27115
rect 19576 27084 20821 27112
rect 19576 27072 19582 27084
rect 20809 27081 20821 27084
rect 20855 27081 20867 27115
rect 25774 27112 25780 27124
rect 25735 27084 25780 27112
rect 20809 27075 20867 27081
rect 25774 27072 25780 27084
rect 25832 27072 25838 27124
rect 34054 27112 34060 27124
rect 34015 27084 34060 27112
rect 34054 27072 34060 27084
rect 34112 27072 34118 27124
rect 57146 27072 57152 27124
rect 57204 27112 57210 27124
rect 58069 27115 58127 27121
rect 58069 27112 58081 27115
rect 57204 27084 58081 27112
rect 57204 27072 57210 27084
rect 58069 27081 58081 27084
rect 58115 27081 58127 27115
rect 58069 27075 58127 27081
rect 28626 27004 28632 27056
rect 28684 27044 28690 27056
rect 33042 27044 33048 27056
rect 28684 27016 33048 27044
rect 28684 27004 28690 27016
rect 33042 27004 33048 27016
rect 33100 27004 33106 27056
rect 33134 27004 33140 27056
rect 33192 27044 33198 27056
rect 44174 27044 44180 27056
rect 33192 27016 44180 27044
rect 33192 27004 33198 27016
rect 44174 27004 44180 27016
rect 44232 27004 44238 27056
rect 57238 27044 57244 27056
rect 57199 27016 57244 27044
rect 57238 27004 57244 27016
rect 57296 27004 57302 27056
rect 20993 26979 21051 26985
rect 20993 26976 21005 26979
rect 19444 26948 21005 26976
rect 20993 26945 21005 26948
rect 21039 26976 21051 26979
rect 21821 26979 21879 26985
rect 21821 26976 21833 26979
rect 21039 26948 21833 26976
rect 21039 26945 21051 26948
rect 20993 26939 21051 26945
rect 21821 26945 21833 26948
rect 21867 26976 21879 26979
rect 21910 26976 21916 26988
rect 21867 26948 21916 26976
rect 21867 26945 21879 26948
rect 21821 26939 21879 26945
rect 21910 26936 21916 26948
rect 21968 26936 21974 26988
rect 30745 26979 30803 26985
rect 30745 26976 30757 26979
rect 28184 26948 30757 26976
rect 14274 26868 14280 26920
rect 14332 26908 14338 26920
rect 22830 26908 22836 26920
rect 14332 26880 22836 26908
rect 14332 26868 14338 26880
rect 22830 26868 22836 26880
rect 22888 26868 22894 26920
rect 26421 26911 26479 26917
rect 26421 26877 26433 26911
rect 26467 26908 26479 26911
rect 27522 26908 27528 26920
rect 26467 26880 27528 26908
rect 26467 26877 26479 26880
rect 26421 26871 26479 26877
rect 27522 26868 27528 26880
rect 27580 26868 27586 26920
rect 3878 26800 3884 26852
rect 3936 26840 3942 26852
rect 19978 26840 19984 26852
rect 3936 26812 19984 26840
rect 3936 26800 3942 26812
rect 19978 26800 19984 26812
rect 20036 26800 20042 26852
rect 28184 26840 28212 26948
rect 30745 26945 30757 26948
rect 30791 26945 30803 26979
rect 30745 26939 30803 26945
rect 31573 26979 31631 26985
rect 31573 26945 31585 26979
rect 31619 26976 31631 26979
rect 32030 26976 32036 26988
rect 31619 26948 32036 26976
rect 31619 26945 31631 26948
rect 31573 26939 31631 26945
rect 30760 26908 30788 26939
rect 32030 26936 32036 26948
rect 32088 26936 32094 26988
rect 32306 26936 32312 26988
rect 32364 26976 32370 26988
rect 32364 26948 34652 26976
rect 32364 26936 32370 26948
rect 33226 26908 33232 26920
rect 30760 26880 33232 26908
rect 33226 26868 33232 26880
rect 33284 26868 33290 26920
rect 34624 26917 34652 26948
rect 56594 26936 56600 26988
rect 56652 26976 56658 26988
rect 57885 26979 57943 26985
rect 57885 26976 57897 26979
rect 56652 26948 57897 26976
rect 56652 26936 56658 26948
rect 57885 26945 57897 26948
rect 57931 26945 57943 26979
rect 57885 26939 57943 26945
rect 34609 26911 34667 26917
rect 34609 26877 34621 26911
rect 34655 26908 34667 26911
rect 37090 26908 37096 26920
rect 34655 26880 37096 26908
rect 34655 26877 34667 26880
rect 34609 26871 34667 26877
rect 37090 26868 37096 26880
rect 37148 26868 37154 26920
rect 20088 26812 28212 26840
rect 28905 26843 28963 26849
rect 17402 26732 17408 26784
rect 17460 26772 17466 26784
rect 20088 26772 20116 26812
rect 28905 26809 28917 26843
rect 28951 26840 28963 26843
rect 30190 26840 30196 26852
rect 28951 26812 30196 26840
rect 28951 26809 28963 26812
rect 28905 26803 28963 26809
rect 30190 26800 30196 26812
rect 30248 26800 30254 26852
rect 33042 26800 33048 26852
rect 33100 26840 33106 26852
rect 35161 26843 35219 26849
rect 35161 26840 35173 26843
rect 33100 26812 35173 26840
rect 33100 26800 33106 26812
rect 35161 26809 35173 26812
rect 35207 26840 35219 26843
rect 41598 26840 41604 26852
rect 35207 26812 41604 26840
rect 35207 26809 35219 26812
rect 35161 26803 35219 26809
rect 41598 26800 41604 26812
rect 41656 26800 41662 26852
rect 17460 26744 20116 26772
rect 17460 26732 17466 26744
rect 25130 26732 25136 26784
rect 25188 26772 25194 26784
rect 25225 26775 25283 26781
rect 25225 26772 25237 26775
rect 25188 26744 25237 26772
rect 25188 26732 25194 26744
rect 25225 26741 25237 26744
rect 25271 26741 25283 26775
rect 27338 26772 27344 26784
rect 27299 26744 27344 26772
rect 25225 26735 25283 26741
rect 27338 26732 27344 26744
rect 27396 26732 27402 26784
rect 28350 26772 28356 26784
rect 28311 26744 28356 26772
rect 28350 26732 28356 26744
rect 28408 26732 28414 26784
rect 29454 26772 29460 26784
rect 29415 26744 29460 26772
rect 29454 26732 29460 26744
rect 29512 26732 29518 26784
rect 30285 26775 30343 26781
rect 30285 26741 30297 26775
rect 30331 26772 30343 26775
rect 30558 26772 30564 26784
rect 30331 26744 30564 26772
rect 30331 26741 30343 26744
rect 30285 26735 30343 26741
rect 30558 26732 30564 26744
rect 30616 26732 30622 26784
rect 30834 26772 30840 26784
rect 30795 26744 30840 26772
rect 30834 26732 30840 26744
rect 30892 26732 30898 26784
rect 31478 26772 31484 26784
rect 31439 26744 31484 26772
rect 31478 26732 31484 26744
rect 31536 26732 31542 26784
rect 31662 26732 31668 26784
rect 31720 26772 31726 26784
rect 32125 26775 32183 26781
rect 32125 26772 32137 26775
rect 31720 26744 32137 26772
rect 31720 26732 31726 26744
rect 32125 26741 32137 26744
rect 32171 26741 32183 26775
rect 32125 26735 32183 26741
rect 32582 26732 32588 26784
rect 32640 26772 32646 26784
rect 32677 26775 32735 26781
rect 32677 26772 32689 26775
rect 32640 26744 32689 26772
rect 32640 26732 32646 26744
rect 32677 26741 32689 26744
rect 32723 26741 32735 26775
rect 32677 26735 32735 26741
rect 33318 26732 33324 26784
rect 33376 26772 33382 26784
rect 33413 26775 33471 26781
rect 33413 26772 33425 26775
rect 33376 26744 33425 26772
rect 33376 26732 33382 26744
rect 33413 26741 33425 26744
rect 33459 26741 33471 26775
rect 35710 26772 35716 26784
rect 35671 26744 35716 26772
rect 33413 26735 33471 26741
rect 35710 26732 35716 26744
rect 35768 26732 35774 26784
rect 35894 26732 35900 26784
rect 35952 26772 35958 26784
rect 36173 26775 36231 26781
rect 36173 26772 36185 26775
rect 35952 26744 36185 26772
rect 35952 26732 35958 26744
rect 36173 26741 36185 26744
rect 36219 26741 36231 26775
rect 36173 26735 36231 26741
rect 37369 26775 37427 26781
rect 37369 26741 37381 26775
rect 37415 26772 37427 26775
rect 37550 26772 37556 26784
rect 37415 26744 37556 26772
rect 37415 26741 37427 26744
rect 37369 26735 37427 26741
rect 37550 26732 37556 26744
rect 37608 26732 37614 26784
rect 1104 26682 58880 26704
rect 1104 26630 10582 26682
rect 10634 26630 10646 26682
rect 10698 26630 10710 26682
rect 10762 26630 10774 26682
rect 10826 26630 10838 26682
rect 10890 26630 29846 26682
rect 29898 26630 29910 26682
rect 29962 26630 29974 26682
rect 30026 26630 30038 26682
rect 30090 26630 30102 26682
rect 30154 26630 49110 26682
rect 49162 26630 49174 26682
rect 49226 26630 49238 26682
rect 49290 26630 49302 26682
rect 49354 26630 49366 26682
rect 49418 26630 58880 26682
rect 1104 26608 58880 26630
rect 30466 26568 30472 26580
rect 30427 26540 30472 26568
rect 30466 26528 30472 26540
rect 30524 26528 30530 26580
rect 31202 26568 31208 26580
rect 31163 26540 31208 26568
rect 31202 26528 31208 26540
rect 31260 26528 31266 26580
rect 36906 26528 36912 26580
rect 36964 26568 36970 26580
rect 46566 26568 46572 26580
rect 36964 26540 46572 26568
rect 36964 26528 36970 26540
rect 46566 26528 46572 26540
rect 46624 26528 46630 26580
rect 58066 26568 58072 26580
rect 58027 26540 58072 26568
rect 58066 26528 58072 26540
rect 58124 26528 58130 26580
rect 23198 26460 23204 26512
rect 23256 26500 23262 26512
rect 29546 26500 29552 26512
rect 23256 26472 28948 26500
rect 29507 26472 29552 26500
rect 23256 26460 23262 26472
rect 23382 26392 23388 26444
rect 23440 26432 23446 26444
rect 26421 26435 26479 26441
rect 26421 26432 26433 26435
rect 23440 26404 26433 26432
rect 23440 26392 23446 26404
rect 26421 26401 26433 26404
rect 26467 26432 26479 26435
rect 28810 26432 28816 26444
rect 26467 26404 28816 26432
rect 26467 26401 26479 26404
rect 26421 26395 26479 26401
rect 28810 26392 28816 26404
rect 28868 26392 28874 26444
rect 28920 26432 28948 26472
rect 29546 26460 29552 26472
rect 29604 26460 29610 26512
rect 30377 26503 30435 26509
rect 30377 26469 30389 26503
rect 30423 26500 30435 26503
rect 35434 26500 35440 26512
rect 30423 26472 35440 26500
rect 30423 26469 30435 26472
rect 30377 26463 30435 26469
rect 35434 26460 35440 26472
rect 35492 26460 35498 26512
rect 35802 26460 35808 26512
rect 35860 26500 35866 26512
rect 45002 26500 45008 26512
rect 35860 26472 45008 26500
rect 35860 26460 35866 26472
rect 45002 26460 45008 26472
rect 45060 26460 45066 26512
rect 30561 26435 30619 26441
rect 28920 26404 30328 26432
rect 1673 26367 1731 26373
rect 1673 26333 1685 26367
rect 1719 26364 1731 26367
rect 8570 26364 8576 26376
rect 1719 26336 8576 26364
rect 1719 26333 1731 26336
rect 1673 26327 1731 26333
rect 8570 26324 8576 26336
rect 8628 26324 8634 26376
rect 27617 26367 27675 26373
rect 27617 26333 27629 26367
rect 27663 26364 27675 26367
rect 27706 26364 27712 26376
rect 27663 26336 27712 26364
rect 27663 26333 27675 26336
rect 27617 26327 27675 26333
rect 27706 26324 27712 26336
rect 27764 26364 27770 26376
rect 28350 26364 28356 26376
rect 27764 26336 28356 26364
rect 27764 26324 27770 26336
rect 28350 26324 28356 26336
rect 28408 26324 28414 26376
rect 29730 26364 29736 26376
rect 29691 26336 29736 26364
rect 29730 26324 29736 26336
rect 29788 26324 29794 26376
rect 30300 26373 30328 26404
rect 30561 26401 30573 26435
rect 30607 26432 30619 26435
rect 30742 26432 30748 26444
rect 30607 26404 30748 26432
rect 30607 26401 30619 26404
rect 30561 26395 30619 26401
rect 30742 26392 30748 26404
rect 30800 26392 30806 26444
rect 33962 26392 33968 26444
rect 34020 26432 34026 26444
rect 34238 26432 34244 26444
rect 34020 26404 34244 26432
rect 34020 26392 34026 26404
rect 34238 26392 34244 26404
rect 34296 26432 34302 26444
rect 37550 26432 37556 26444
rect 34296 26404 37556 26432
rect 34296 26392 34302 26404
rect 37550 26392 37556 26404
rect 37608 26432 37614 26444
rect 43530 26432 43536 26444
rect 37608 26404 43536 26432
rect 37608 26392 37614 26404
rect 43530 26392 43536 26404
rect 43588 26392 43594 26444
rect 30285 26367 30343 26373
rect 30285 26333 30297 26367
rect 30331 26333 30343 26367
rect 31202 26364 31208 26376
rect 31163 26336 31208 26364
rect 30285 26327 30343 26333
rect 31202 26324 31208 26336
rect 31260 26324 31266 26376
rect 31938 26364 31944 26376
rect 31899 26336 31944 26364
rect 31938 26324 31944 26336
rect 31996 26324 32002 26376
rect 32401 26367 32459 26373
rect 32401 26364 32413 26367
rect 32048 26336 32413 26364
rect 28258 26296 28264 26308
rect 28219 26268 28264 26296
rect 28258 26256 28264 26268
rect 28316 26256 28322 26308
rect 31846 26256 31852 26308
rect 31904 26296 31910 26308
rect 32048 26296 32076 26336
rect 32401 26333 32413 26336
rect 32447 26333 32459 26367
rect 32401 26327 32459 26333
rect 32490 26324 32496 26376
rect 32548 26364 32554 26376
rect 33226 26364 33232 26376
rect 32548 26336 32593 26364
rect 33139 26336 33232 26364
rect 32548 26324 32554 26336
rect 33226 26324 33232 26336
rect 33284 26364 33290 26376
rect 35710 26364 35716 26376
rect 33284 26336 35716 26364
rect 33284 26324 33290 26336
rect 35710 26324 35716 26336
rect 35768 26364 35774 26376
rect 36449 26367 36507 26373
rect 36449 26364 36461 26367
rect 35768 26336 36461 26364
rect 35768 26324 35774 26336
rect 36449 26333 36461 26336
rect 36495 26364 36507 26367
rect 45554 26364 45560 26376
rect 36495 26336 45560 26364
rect 36495 26333 36507 26336
rect 36449 26327 36507 26333
rect 45554 26324 45560 26336
rect 45612 26324 45618 26376
rect 33134 26296 33140 26308
rect 31904 26268 32076 26296
rect 33095 26268 33140 26296
rect 31904 26256 31910 26268
rect 33134 26256 33140 26268
rect 33192 26256 33198 26308
rect 33778 26296 33784 26308
rect 33739 26268 33784 26296
rect 33778 26256 33784 26268
rect 33836 26256 33842 26308
rect 34054 26256 34060 26308
rect 34112 26296 34118 26308
rect 34701 26299 34759 26305
rect 34701 26296 34713 26299
rect 34112 26268 34713 26296
rect 34112 26256 34118 26268
rect 34701 26265 34713 26268
rect 34747 26265 34759 26299
rect 34701 26259 34759 26265
rect 36170 26256 36176 26308
rect 36228 26296 36234 26308
rect 36906 26296 36912 26308
rect 36228 26268 36912 26296
rect 36228 26256 36234 26268
rect 36906 26256 36912 26268
rect 36964 26256 36970 26308
rect 38105 26299 38163 26305
rect 38105 26265 38117 26299
rect 38151 26296 38163 26299
rect 40954 26296 40960 26308
rect 38151 26268 40960 26296
rect 38151 26265 38163 26268
rect 38105 26259 38163 26265
rect 40954 26256 40960 26268
rect 41012 26256 41018 26308
rect 1486 26228 1492 26240
rect 1447 26200 1492 26228
rect 1486 26188 1492 26200
rect 1544 26188 1550 26240
rect 18966 26188 18972 26240
rect 19024 26228 19030 26240
rect 19334 26228 19340 26240
rect 19024 26200 19340 26228
rect 19024 26188 19030 26200
rect 19334 26188 19340 26200
rect 19392 26188 19398 26240
rect 24670 26228 24676 26240
rect 24631 26200 24676 26228
rect 24670 26188 24676 26200
rect 24728 26188 24734 26240
rect 25130 26228 25136 26240
rect 25091 26200 25136 26228
rect 25130 26188 25136 26200
rect 25188 26188 25194 26240
rect 25406 26188 25412 26240
rect 25464 26228 25470 26240
rect 25777 26231 25835 26237
rect 25777 26228 25789 26231
rect 25464 26200 25789 26228
rect 25464 26188 25470 26200
rect 25777 26197 25789 26200
rect 25823 26197 25835 26231
rect 25777 26191 25835 26197
rect 26973 26231 27031 26237
rect 26973 26197 26985 26231
rect 27019 26228 27031 26231
rect 28074 26228 28080 26240
rect 27019 26200 28080 26228
rect 27019 26197 27031 26200
rect 26973 26191 27031 26197
rect 28074 26188 28080 26200
rect 28132 26188 28138 26240
rect 28997 26231 29055 26237
rect 28997 26197 29009 26231
rect 29043 26228 29055 26231
rect 29086 26228 29092 26240
rect 29043 26200 29092 26228
rect 29043 26197 29055 26200
rect 28997 26191 29055 26197
rect 29086 26188 29092 26200
rect 29144 26188 29150 26240
rect 31478 26188 31484 26240
rect 31536 26228 31542 26240
rect 31757 26231 31815 26237
rect 31757 26228 31769 26231
rect 31536 26200 31769 26228
rect 31536 26188 31542 26200
rect 31757 26197 31769 26200
rect 31803 26197 31815 26231
rect 31757 26191 31815 26197
rect 32674 26188 32680 26240
rect 32732 26228 32738 26240
rect 35253 26231 35311 26237
rect 35253 26228 35265 26231
rect 32732 26200 35265 26228
rect 32732 26188 32738 26200
rect 35253 26197 35265 26200
rect 35299 26197 35311 26231
rect 35253 26191 35311 26197
rect 35618 26188 35624 26240
rect 35676 26228 35682 26240
rect 35802 26228 35808 26240
rect 35676 26200 35808 26228
rect 35676 26188 35682 26200
rect 35802 26188 35808 26200
rect 35860 26188 35866 26240
rect 37553 26231 37611 26237
rect 37553 26197 37565 26231
rect 37599 26228 37611 26231
rect 38378 26228 38384 26240
rect 37599 26200 38384 26228
rect 37599 26197 37611 26200
rect 37553 26191 37611 26197
rect 38378 26188 38384 26200
rect 38436 26188 38442 26240
rect 1104 26138 58880 26160
rect 1104 26086 20214 26138
rect 20266 26086 20278 26138
rect 20330 26086 20342 26138
rect 20394 26086 20406 26138
rect 20458 26086 20470 26138
rect 20522 26086 39478 26138
rect 39530 26086 39542 26138
rect 39594 26086 39606 26138
rect 39658 26086 39670 26138
rect 39722 26086 39734 26138
rect 39786 26086 58880 26138
rect 1104 26064 58880 26086
rect 25406 25984 25412 26036
rect 25464 26024 25470 26036
rect 30466 26024 30472 26036
rect 25464 25996 29592 26024
rect 30427 25996 30472 26024
rect 25464 25984 25470 25996
rect 23753 25959 23811 25965
rect 23753 25925 23765 25959
rect 23799 25956 23811 25959
rect 24670 25956 24676 25968
rect 23799 25928 24676 25956
rect 23799 25925 23811 25928
rect 23753 25919 23811 25925
rect 24670 25916 24676 25928
rect 24728 25956 24734 25968
rect 27798 25956 27804 25968
rect 24728 25928 27804 25956
rect 24728 25916 24734 25928
rect 27798 25916 27804 25928
rect 27856 25916 27862 25968
rect 28350 25916 28356 25968
rect 28408 25956 28414 25968
rect 28408 25928 29040 25956
rect 28408 25916 28414 25928
rect 26786 25848 26792 25900
rect 26844 25888 26850 25900
rect 29012 25897 29040 25928
rect 28813 25891 28871 25897
rect 28813 25888 28825 25891
rect 26844 25860 28825 25888
rect 26844 25848 26850 25860
rect 28813 25857 28825 25860
rect 28859 25857 28871 25891
rect 28813 25851 28871 25857
rect 28997 25891 29055 25897
rect 28997 25857 29009 25891
rect 29043 25888 29055 25891
rect 29362 25888 29368 25900
rect 29043 25860 29368 25888
rect 29043 25857 29055 25860
rect 28997 25851 29055 25857
rect 29362 25848 29368 25860
rect 29420 25848 29426 25900
rect 29564 25888 29592 25996
rect 30466 25984 30472 25996
rect 30524 25984 30530 26036
rect 32490 26024 32496 26036
rect 30944 25996 32496 26024
rect 29914 25916 29920 25968
rect 29972 25956 29978 25968
rect 30944 25965 30972 25996
rect 32490 25984 32496 25996
rect 32548 25984 32554 26036
rect 33502 25984 33508 26036
rect 33560 26024 33566 26036
rect 37274 26024 37280 26036
rect 33560 25996 37280 26024
rect 33560 25984 33566 25996
rect 37274 25984 37280 25996
rect 37332 25984 37338 26036
rect 38378 26024 38384 26036
rect 38339 25996 38384 26024
rect 38378 25984 38384 25996
rect 38436 26024 38442 26036
rect 38933 26027 38991 26033
rect 38933 26024 38945 26027
rect 38436 25996 38945 26024
rect 38436 25984 38442 25996
rect 38933 25993 38945 25996
rect 38979 26024 38991 26027
rect 40586 26024 40592 26036
rect 38979 25996 40592 26024
rect 38979 25993 38991 25996
rect 38933 25987 38991 25993
rect 40586 25984 40592 25996
rect 40644 25984 40650 26036
rect 44361 26027 44419 26033
rect 44361 25993 44373 26027
rect 44407 26024 44419 26027
rect 46474 26024 46480 26036
rect 44407 25996 46480 26024
rect 44407 25993 44419 25996
rect 44361 25987 44419 25993
rect 46474 25984 46480 25996
rect 46532 25984 46538 26036
rect 30929 25959 30987 25965
rect 30929 25956 30941 25959
rect 29972 25928 30941 25956
rect 29972 25916 29978 25928
rect 30929 25925 30941 25928
rect 30975 25925 30987 25959
rect 30929 25919 30987 25925
rect 32401 25959 32459 25965
rect 32401 25925 32413 25959
rect 32447 25956 32459 25959
rect 37734 25956 37740 25968
rect 32447 25928 37740 25956
rect 32447 25925 32459 25928
rect 32401 25919 32459 25925
rect 37734 25916 37740 25928
rect 37792 25916 37798 25968
rect 29825 25891 29883 25897
rect 29825 25888 29837 25891
rect 29564 25860 29837 25888
rect 29825 25857 29837 25860
rect 29871 25888 29883 25891
rect 31570 25888 31576 25900
rect 29871 25860 30972 25888
rect 31531 25860 31576 25888
rect 29871 25857 29883 25860
rect 29825 25851 29883 25857
rect 30944 25832 30972 25860
rect 31570 25848 31576 25860
rect 31628 25848 31634 25900
rect 32125 25891 32183 25897
rect 32125 25857 32137 25891
rect 32171 25857 32183 25891
rect 32125 25851 32183 25857
rect 33045 25891 33103 25897
rect 33045 25857 33057 25891
rect 33091 25857 33103 25891
rect 33686 25888 33692 25900
rect 33599 25860 33692 25888
rect 33045 25851 33103 25857
rect 29638 25780 29644 25832
rect 29696 25820 29702 25832
rect 29733 25823 29791 25829
rect 29733 25820 29745 25823
rect 29696 25792 29745 25820
rect 29696 25780 29702 25792
rect 29733 25789 29745 25792
rect 29779 25820 29791 25823
rect 29779 25792 30696 25820
rect 29779 25789 29791 25792
rect 29733 25783 29791 25789
rect 2222 25712 2228 25764
rect 2280 25752 2286 25764
rect 22002 25752 22008 25764
rect 2280 25724 22008 25752
rect 2280 25712 2286 25724
rect 22002 25712 22008 25724
rect 22060 25712 22066 25764
rect 23014 25712 23020 25764
rect 23072 25752 23078 25764
rect 27246 25752 27252 25764
rect 23072 25724 27252 25752
rect 23072 25712 23078 25724
rect 27246 25712 27252 25724
rect 27304 25712 27310 25764
rect 27801 25755 27859 25761
rect 27801 25721 27813 25755
rect 27847 25752 27859 25755
rect 28534 25752 28540 25764
rect 27847 25724 28540 25752
rect 27847 25721 27859 25724
rect 27801 25715 27859 25721
rect 28534 25712 28540 25724
rect 28592 25712 28598 25764
rect 28718 25712 28724 25764
rect 28776 25752 28782 25764
rect 29914 25752 29920 25764
rect 28776 25724 29920 25752
rect 28776 25712 28782 25724
rect 29914 25712 29920 25724
rect 29972 25712 29978 25764
rect 30374 25712 30380 25764
rect 30432 25752 30438 25764
rect 30561 25755 30619 25761
rect 30561 25752 30573 25755
rect 30432 25724 30573 25752
rect 30432 25712 30438 25724
rect 30561 25721 30573 25724
rect 30607 25721 30619 25755
rect 30668 25752 30696 25792
rect 30926 25780 30932 25832
rect 30984 25780 30990 25832
rect 31386 25780 31392 25832
rect 31444 25820 31450 25832
rect 32140 25820 32168 25851
rect 31444 25792 32168 25820
rect 31444 25780 31450 25792
rect 32950 25780 32956 25832
rect 33008 25780 33014 25832
rect 33060 25820 33088 25851
rect 33686 25848 33692 25860
rect 33744 25888 33750 25900
rect 34422 25888 34428 25900
rect 33744 25860 34428 25888
rect 33744 25848 33750 25860
rect 34422 25848 34428 25860
rect 34480 25848 34486 25900
rect 36630 25848 36636 25900
rect 36688 25888 36694 25900
rect 44177 25891 44235 25897
rect 44177 25888 44189 25891
rect 36688 25860 44189 25888
rect 36688 25848 36694 25860
rect 44177 25857 44189 25860
rect 44223 25857 44235 25891
rect 47581 25891 47639 25897
rect 47581 25888 47593 25891
rect 44177 25851 44235 25857
rect 45526 25860 47593 25888
rect 35250 25820 35256 25832
rect 33060 25792 35256 25820
rect 35250 25780 35256 25792
rect 35308 25780 35314 25832
rect 39206 25780 39212 25832
rect 39264 25820 39270 25832
rect 45526 25820 45554 25860
rect 47581 25857 47593 25860
rect 47627 25857 47639 25891
rect 47581 25851 47639 25857
rect 58069 25891 58127 25897
rect 58069 25857 58081 25891
rect 58115 25888 58127 25891
rect 58158 25888 58164 25900
rect 58115 25860 58164 25888
rect 58115 25857 58127 25860
rect 58069 25851 58127 25857
rect 58158 25848 58164 25860
rect 58216 25848 58222 25900
rect 39264 25792 45554 25820
rect 39264 25780 39270 25792
rect 32582 25752 32588 25764
rect 30668 25724 32588 25752
rect 30561 25715 30619 25721
rect 32582 25712 32588 25724
rect 32640 25712 32646 25764
rect 32968 25752 32996 25780
rect 35345 25755 35403 25761
rect 35345 25752 35357 25755
rect 32968 25724 35357 25752
rect 35345 25721 35357 25724
rect 35391 25752 35403 25755
rect 35526 25752 35532 25764
rect 35391 25724 35532 25752
rect 35391 25721 35403 25724
rect 35345 25715 35403 25721
rect 35526 25712 35532 25724
rect 35584 25712 35590 25764
rect 35710 25712 35716 25764
rect 35768 25752 35774 25764
rect 36357 25755 36415 25761
rect 36357 25752 36369 25755
rect 35768 25724 36369 25752
rect 35768 25712 35774 25724
rect 36357 25721 36369 25724
rect 36403 25721 36415 25755
rect 57882 25752 57888 25764
rect 57843 25724 57888 25752
rect 36357 25715 36415 25721
rect 57882 25712 57888 25724
rect 57940 25712 57946 25764
rect 20714 25644 20720 25696
rect 20772 25684 20778 25696
rect 23201 25687 23259 25693
rect 23201 25684 23213 25687
rect 20772 25656 23213 25684
rect 20772 25644 20778 25656
rect 23201 25653 23213 25656
rect 23247 25653 23259 25687
rect 24394 25684 24400 25696
rect 24355 25656 24400 25684
rect 23201 25647 23259 25653
rect 24394 25644 24400 25656
rect 24452 25644 24458 25696
rect 24854 25684 24860 25696
rect 24815 25656 24860 25684
rect 24854 25644 24860 25656
rect 24912 25644 24918 25696
rect 25038 25644 25044 25696
rect 25096 25684 25102 25696
rect 25406 25684 25412 25696
rect 25096 25656 25412 25684
rect 25096 25644 25102 25656
rect 25406 25644 25412 25656
rect 25464 25644 25470 25696
rect 26421 25687 26479 25693
rect 26421 25653 26433 25687
rect 26467 25684 26479 25687
rect 27154 25684 27160 25696
rect 26467 25656 27160 25684
rect 26467 25653 26479 25656
rect 26421 25647 26479 25653
rect 27154 25644 27160 25656
rect 27212 25644 27218 25696
rect 28074 25644 28080 25696
rect 28132 25684 28138 25696
rect 28261 25687 28319 25693
rect 28261 25684 28273 25687
rect 28132 25656 28273 25684
rect 28132 25644 28138 25656
rect 28261 25653 28273 25656
rect 28307 25653 28319 25687
rect 28902 25684 28908 25696
rect 28863 25656 28908 25684
rect 28261 25647 28319 25653
rect 28902 25644 28908 25656
rect 28960 25644 28966 25696
rect 29454 25684 29460 25696
rect 29415 25656 29460 25684
rect 29454 25644 29460 25656
rect 29512 25644 29518 25696
rect 30834 25644 30840 25696
rect 30892 25684 30898 25696
rect 31481 25687 31539 25693
rect 31481 25684 31493 25687
rect 30892 25656 31493 25684
rect 30892 25644 30898 25656
rect 31481 25653 31493 25656
rect 31527 25653 31539 25687
rect 31481 25647 31539 25653
rect 31754 25644 31760 25696
rect 31812 25684 31818 25696
rect 32306 25684 32312 25696
rect 31812 25656 32312 25684
rect 31812 25644 31818 25656
rect 32306 25644 32312 25656
rect 32364 25644 32370 25696
rect 32398 25644 32404 25696
rect 32456 25684 32462 25696
rect 32953 25687 33011 25693
rect 32953 25684 32965 25687
rect 32456 25656 32965 25684
rect 32456 25644 32462 25656
rect 32953 25653 32965 25656
rect 32999 25653 33011 25687
rect 33594 25684 33600 25696
rect 33555 25656 33600 25684
rect 32953 25647 33011 25653
rect 33594 25644 33600 25656
rect 33652 25644 33658 25696
rect 34241 25687 34299 25693
rect 34241 25653 34253 25687
rect 34287 25684 34299 25687
rect 34330 25684 34336 25696
rect 34287 25656 34336 25684
rect 34287 25653 34299 25656
rect 34241 25647 34299 25653
rect 34330 25644 34336 25656
rect 34388 25644 34394 25696
rect 34698 25684 34704 25696
rect 34659 25656 34704 25684
rect 34698 25644 34704 25656
rect 34756 25644 34762 25696
rect 35897 25687 35955 25693
rect 35897 25653 35909 25687
rect 35943 25684 35955 25687
rect 36446 25684 36452 25696
rect 35943 25656 36452 25684
rect 35943 25653 35955 25656
rect 35897 25647 35955 25653
rect 36446 25644 36452 25656
rect 36504 25644 36510 25696
rect 37921 25687 37979 25693
rect 37921 25653 37933 25687
rect 37967 25684 37979 25687
rect 38286 25684 38292 25696
rect 37967 25656 38292 25684
rect 37967 25653 37979 25656
rect 37921 25647 37979 25653
rect 38286 25644 38292 25656
rect 38344 25644 38350 25696
rect 47765 25687 47823 25693
rect 47765 25653 47777 25687
rect 47811 25684 47823 25687
rect 56594 25684 56600 25696
rect 47811 25656 56600 25684
rect 47811 25653 47823 25656
rect 47765 25647 47823 25653
rect 56594 25644 56600 25656
rect 56652 25644 56658 25696
rect 1104 25594 58880 25616
rect 1104 25542 10582 25594
rect 10634 25542 10646 25594
rect 10698 25542 10710 25594
rect 10762 25542 10774 25594
rect 10826 25542 10838 25594
rect 10890 25542 29846 25594
rect 29898 25542 29910 25594
rect 29962 25542 29974 25594
rect 30026 25542 30038 25594
rect 30090 25542 30102 25594
rect 30154 25542 49110 25594
rect 49162 25542 49174 25594
rect 49226 25542 49238 25594
rect 49290 25542 49302 25594
rect 49354 25542 49366 25594
rect 49418 25542 58880 25594
rect 1104 25520 58880 25542
rect 23293 25483 23351 25489
rect 23293 25449 23305 25483
rect 23339 25480 23351 25483
rect 25774 25480 25780 25492
rect 23339 25452 25780 25480
rect 23339 25449 23351 25452
rect 23293 25443 23351 25449
rect 14458 25412 14464 25424
rect 14419 25384 14464 25412
rect 14458 25372 14464 25384
rect 14516 25372 14522 25424
rect 21634 25372 21640 25424
rect 21692 25412 21698 25424
rect 23308 25412 23336 25443
rect 25774 25440 25780 25452
rect 25832 25440 25838 25492
rect 26418 25440 26424 25492
rect 26476 25480 26482 25492
rect 31570 25480 31576 25492
rect 26476 25452 31576 25480
rect 26476 25440 26482 25452
rect 31570 25440 31576 25452
rect 31628 25440 31634 25492
rect 32401 25483 32459 25489
rect 32401 25449 32413 25483
rect 32447 25480 32459 25483
rect 33042 25480 33048 25492
rect 32447 25452 33048 25480
rect 32447 25449 32459 25452
rect 32401 25443 32459 25449
rect 33042 25440 33048 25452
rect 33100 25440 33106 25492
rect 34606 25440 34612 25492
rect 34664 25480 34670 25492
rect 34701 25483 34759 25489
rect 34701 25480 34713 25483
rect 34664 25452 34713 25480
rect 34664 25440 34670 25452
rect 34701 25449 34713 25452
rect 34747 25480 34759 25483
rect 34790 25480 34796 25492
rect 34747 25452 34796 25480
rect 34747 25449 34759 25452
rect 34701 25443 34759 25449
rect 34790 25440 34796 25452
rect 34848 25440 34854 25492
rect 34974 25440 34980 25492
rect 35032 25480 35038 25492
rect 35345 25483 35403 25489
rect 35345 25480 35357 25483
rect 35032 25452 35357 25480
rect 35032 25440 35038 25452
rect 35345 25449 35357 25452
rect 35391 25449 35403 25483
rect 35345 25443 35403 25449
rect 37366 25440 37372 25492
rect 37424 25480 37430 25492
rect 37550 25480 37556 25492
rect 37424 25452 37556 25480
rect 37424 25440 37430 25452
rect 37550 25440 37556 25452
rect 37608 25440 37614 25492
rect 46934 25480 46940 25492
rect 39224 25452 46940 25480
rect 21692 25384 23336 25412
rect 23845 25415 23903 25421
rect 21692 25372 21698 25384
rect 23845 25381 23857 25415
rect 23891 25412 23903 25415
rect 23934 25412 23940 25424
rect 23891 25384 23940 25412
rect 23891 25381 23903 25384
rect 23845 25375 23903 25381
rect 23934 25372 23940 25384
rect 23992 25412 23998 25424
rect 25222 25412 25228 25424
rect 23992 25384 25228 25412
rect 23992 25372 23998 25384
rect 25222 25372 25228 25384
rect 25280 25372 25286 25424
rect 26234 25372 26240 25424
rect 26292 25412 26298 25424
rect 27341 25415 27399 25421
rect 27341 25412 27353 25415
rect 26292 25384 27353 25412
rect 26292 25372 26298 25384
rect 27341 25381 27353 25384
rect 27387 25412 27399 25415
rect 28718 25412 28724 25424
rect 27387 25384 28724 25412
rect 27387 25381 27399 25384
rect 27341 25375 27399 25381
rect 28718 25372 28724 25384
rect 28776 25372 28782 25424
rect 29549 25415 29607 25421
rect 29549 25381 29561 25415
rect 29595 25412 29607 25415
rect 35526 25412 35532 25424
rect 29595 25384 35532 25412
rect 29595 25381 29607 25384
rect 29549 25375 29607 25381
rect 35526 25372 35532 25384
rect 35584 25372 35590 25424
rect 35618 25372 35624 25424
rect 35676 25412 35682 25424
rect 38286 25412 38292 25424
rect 35676 25384 38292 25412
rect 35676 25372 35682 25384
rect 38286 25372 38292 25384
rect 38344 25372 38350 25424
rect 25501 25347 25559 25353
rect 25501 25313 25513 25347
rect 25547 25344 25559 25347
rect 25774 25344 25780 25356
rect 25547 25316 25780 25344
rect 25547 25313 25559 25316
rect 25501 25307 25559 25313
rect 25774 25304 25780 25316
rect 25832 25344 25838 25356
rect 27706 25344 27712 25356
rect 25832 25316 27712 25344
rect 25832 25304 25838 25316
rect 27706 25304 27712 25316
rect 27764 25304 27770 25356
rect 28810 25344 28816 25356
rect 28771 25316 28816 25344
rect 28810 25304 28816 25316
rect 28868 25304 28874 25356
rect 28994 25304 29000 25356
rect 29052 25344 29058 25356
rect 30469 25347 30527 25353
rect 30469 25344 30481 25347
rect 29052 25316 30481 25344
rect 29052 25304 29058 25316
rect 30469 25313 30481 25316
rect 30515 25344 30527 25347
rect 31389 25347 31447 25353
rect 30515 25316 31340 25344
rect 30515 25313 30527 25316
rect 30469 25307 30527 25313
rect 21450 25236 21456 25288
rect 21508 25276 21514 25288
rect 26878 25276 26884 25288
rect 21508 25248 26884 25276
rect 21508 25236 21514 25248
rect 26878 25236 26884 25248
rect 26936 25236 26942 25288
rect 27985 25279 28043 25285
rect 27985 25245 27997 25279
rect 28031 25276 28043 25279
rect 28166 25276 28172 25288
rect 28031 25248 28172 25276
rect 28031 25245 28043 25248
rect 27985 25239 28043 25245
rect 28166 25236 28172 25248
rect 28224 25236 28230 25288
rect 28626 25276 28632 25288
rect 28587 25248 28632 25276
rect 28626 25236 28632 25248
rect 28684 25236 28690 25288
rect 29917 25279 29975 25285
rect 29917 25245 29929 25279
rect 29963 25276 29975 25279
rect 30282 25276 30288 25288
rect 29963 25248 30288 25276
rect 29963 25245 29975 25248
rect 29917 25239 29975 25245
rect 30282 25236 30288 25248
rect 30340 25236 30346 25288
rect 30558 25276 30564 25288
rect 30519 25248 30564 25276
rect 30558 25236 30564 25248
rect 30616 25236 30622 25288
rect 14645 25211 14703 25217
rect 14645 25177 14657 25211
rect 14691 25208 14703 25211
rect 21082 25208 21088 25220
rect 14691 25180 21088 25208
rect 14691 25177 14703 25180
rect 14645 25171 14703 25177
rect 21082 25168 21088 25180
rect 21140 25168 21146 25220
rect 23842 25168 23848 25220
rect 23900 25208 23906 25220
rect 29178 25208 29184 25220
rect 23900 25180 29184 25208
rect 23900 25168 23906 25180
rect 29178 25168 29184 25180
rect 29236 25168 29242 25220
rect 29730 25208 29736 25220
rect 29691 25180 29736 25208
rect 29730 25168 29736 25180
rect 29788 25168 29794 25220
rect 24946 25140 24952 25152
rect 24907 25112 24952 25140
rect 24946 25100 24952 25112
rect 25004 25100 25010 25152
rect 26053 25143 26111 25149
rect 26053 25109 26065 25143
rect 26099 25140 26111 25143
rect 26142 25140 26148 25152
rect 26099 25112 26148 25140
rect 26099 25109 26111 25112
rect 26053 25103 26111 25109
rect 26142 25100 26148 25112
rect 26200 25100 26206 25152
rect 26789 25143 26847 25149
rect 26789 25109 26801 25143
rect 26835 25140 26847 25143
rect 27154 25140 27160 25152
rect 26835 25112 27160 25140
rect 26835 25109 26847 25112
rect 26789 25103 26847 25109
rect 27154 25100 27160 25112
rect 27212 25100 27218 25152
rect 27890 25140 27896 25152
rect 27851 25112 27896 25140
rect 27890 25100 27896 25112
rect 27948 25100 27954 25152
rect 28442 25140 28448 25152
rect 28403 25112 28448 25140
rect 28442 25100 28448 25112
rect 28500 25100 28506 25152
rect 30929 25143 30987 25149
rect 30929 25109 30941 25143
rect 30975 25140 30987 25143
rect 31110 25140 31116 25152
rect 30975 25112 31116 25140
rect 30975 25109 30987 25112
rect 30929 25103 30987 25109
rect 31110 25100 31116 25112
rect 31168 25100 31174 25152
rect 31312 25140 31340 25316
rect 31389 25313 31401 25347
rect 31435 25344 31447 25347
rect 37182 25344 37188 25356
rect 31435 25316 37188 25344
rect 31435 25313 31447 25316
rect 31389 25307 31447 25313
rect 37182 25304 37188 25316
rect 37240 25304 37246 25356
rect 31570 25276 31576 25288
rect 31531 25248 31576 25276
rect 31570 25236 31576 25248
rect 31628 25236 31634 25288
rect 32030 25236 32036 25288
rect 32088 25276 32094 25288
rect 33042 25276 33048 25288
rect 32088 25248 32352 25276
rect 33003 25248 33048 25276
rect 32088 25236 32094 25248
rect 31478 25168 31484 25220
rect 31536 25208 31542 25220
rect 31757 25211 31815 25217
rect 31757 25208 31769 25211
rect 31536 25180 31769 25208
rect 31536 25168 31542 25180
rect 31757 25177 31769 25180
rect 31803 25177 31815 25211
rect 32214 25208 32220 25220
rect 32175 25180 32220 25208
rect 31757 25171 31815 25177
rect 32214 25168 32220 25180
rect 32272 25168 32278 25220
rect 32324 25208 32352 25248
rect 33042 25236 33048 25248
rect 33100 25236 33106 25288
rect 33502 25236 33508 25288
rect 33560 25276 33566 25288
rect 33781 25279 33839 25285
rect 33781 25276 33793 25279
rect 33560 25248 33793 25276
rect 33560 25236 33566 25248
rect 33781 25245 33793 25248
rect 33827 25245 33839 25279
rect 33781 25239 33839 25245
rect 35437 25279 35495 25285
rect 35437 25245 35449 25279
rect 35483 25276 35495 25279
rect 35618 25276 35624 25288
rect 35483 25248 35624 25276
rect 35483 25245 35495 25248
rect 35437 25239 35495 25245
rect 35618 25236 35624 25248
rect 35676 25236 35682 25288
rect 35710 25236 35716 25288
rect 35768 25276 35774 25288
rect 37001 25279 37059 25285
rect 37001 25276 37013 25279
rect 35768 25248 37013 25276
rect 35768 25236 35774 25248
rect 37001 25245 37013 25248
rect 37047 25245 37059 25279
rect 37001 25239 37059 25245
rect 37274 25236 37280 25288
rect 37332 25276 37338 25288
rect 39224 25285 39252 25452
rect 46934 25440 46940 25452
rect 46992 25440 46998 25492
rect 58158 25480 58164 25492
rect 58119 25452 58164 25480
rect 58158 25440 58164 25452
rect 58216 25440 58222 25492
rect 39209 25279 39267 25285
rect 39209 25276 39221 25279
rect 37332 25248 39221 25276
rect 37332 25236 37338 25248
rect 39209 25245 39221 25248
rect 39255 25245 39267 25279
rect 39209 25239 39267 25245
rect 32433 25211 32491 25217
rect 32433 25208 32445 25211
rect 32324 25180 32445 25208
rect 32433 25177 32445 25180
rect 32479 25208 32491 25211
rect 33873 25211 33931 25217
rect 32479 25180 33456 25208
rect 32479 25177 32491 25180
rect 32433 25171 32491 25177
rect 32030 25140 32036 25152
rect 31312 25112 32036 25140
rect 32030 25100 32036 25112
rect 32088 25100 32094 25152
rect 32582 25140 32588 25152
rect 32543 25112 32588 25140
rect 32582 25100 32588 25112
rect 32640 25100 32646 25152
rect 33226 25140 33232 25152
rect 33187 25112 33232 25140
rect 33226 25100 33232 25112
rect 33284 25100 33290 25152
rect 33428 25140 33456 25180
rect 33873 25177 33885 25211
rect 33919 25208 33931 25211
rect 36354 25208 36360 25220
rect 33919 25180 36360 25208
rect 33919 25177 33931 25180
rect 33873 25171 33931 25177
rect 36354 25168 36360 25180
rect 36412 25168 36418 25220
rect 35618 25140 35624 25152
rect 33428 25112 35624 25140
rect 35618 25100 35624 25112
rect 35676 25100 35682 25152
rect 35894 25140 35900 25152
rect 35855 25112 35900 25140
rect 35894 25100 35900 25112
rect 35952 25100 35958 25152
rect 36538 25140 36544 25152
rect 36499 25112 36544 25140
rect 36538 25100 36544 25112
rect 36596 25100 36602 25152
rect 38102 25140 38108 25152
rect 38063 25112 38108 25140
rect 38102 25100 38108 25112
rect 38160 25100 38166 25152
rect 38746 25140 38752 25152
rect 38707 25112 38752 25140
rect 38746 25100 38752 25112
rect 38804 25100 38810 25152
rect 1104 25050 58880 25072
rect 1104 24998 20214 25050
rect 20266 24998 20278 25050
rect 20330 24998 20342 25050
rect 20394 24998 20406 25050
rect 20458 24998 20470 25050
rect 20522 24998 39478 25050
rect 39530 24998 39542 25050
rect 39594 24998 39606 25050
rect 39658 24998 39670 25050
rect 39722 24998 39734 25050
rect 39786 24998 58880 25050
rect 1104 24976 58880 24998
rect 25498 24896 25504 24948
rect 25556 24936 25562 24948
rect 25556 24908 27936 24936
rect 25556 24896 25562 24908
rect 27706 24868 27712 24880
rect 27448 24840 27712 24868
rect 1673 24803 1731 24809
rect 1673 24769 1685 24803
rect 1719 24800 1731 24803
rect 9122 24800 9128 24812
rect 1719 24772 9128 24800
rect 1719 24769 1731 24772
rect 1673 24763 1731 24769
rect 9122 24760 9128 24772
rect 9180 24760 9186 24812
rect 11701 24803 11759 24809
rect 11701 24769 11713 24803
rect 11747 24800 11759 24803
rect 22186 24800 22192 24812
rect 11747 24772 22192 24800
rect 11747 24769 11759 24772
rect 11701 24763 11759 24769
rect 22186 24760 22192 24772
rect 22244 24760 22250 24812
rect 27448 24809 27476 24840
rect 27706 24828 27712 24840
rect 27764 24828 27770 24880
rect 27908 24877 27936 24908
rect 31754 24896 31760 24948
rect 31812 24936 31818 24948
rect 32214 24936 32220 24948
rect 31812 24908 32220 24936
rect 31812 24896 31818 24908
rect 32214 24896 32220 24908
rect 32272 24896 32278 24948
rect 32306 24896 32312 24948
rect 32364 24936 32370 24948
rect 32493 24939 32551 24945
rect 32493 24936 32505 24939
rect 32364 24908 32505 24936
rect 32364 24896 32370 24908
rect 32493 24905 32505 24908
rect 32539 24905 32551 24939
rect 32493 24899 32551 24905
rect 32582 24896 32588 24948
rect 32640 24936 32646 24948
rect 32640 24908 41414 24936
rect 32640 24896 32646 24908
rect 27893 24871 27951 24877
rect 27893 24837 27905 24871
rect 27939 24837 27951 24871
rect 27893 24831 27951 24837
rect 28123 24837 28181 24843
rect 28123 24834 28135 24837
rect 27249 24803 27307 24809
rect 27249 24800 27261 24803
rect 22296 24772 27261 24800
rect 19794 24692 19800 24744
rect 19852 24732 19858 24744
rect 22296 24732 22324 24772
rect 27249 24769 27261 24772
rect 27295 24769 27307 24803
rect 27249 24763 27307 24769
rect 27433 24803 27491 24809
rect 27433 24769 27445 24803
rect 27479 24769 27491 24803
rect 27433 24763 27491 24769
rect 27522 24760 27528 24812
rect 27580 24800 27586 24812
rect 28108 24803 28135 24834
rect 28169 24803 28181 24837
rect 28442 24828 28448 24880
rect 28500 24868 28506 24880
rect 33226 24868 33232 24880
rect 28500 24840 33232 24868
rect 28500 24828 28506 24840
rect 33226 24828 33232 24840
rect 33284 24828 33290 24880
rect 38654 24868 38660 24880
rect 36740 24840 38660 24868
rect 36740 24812 36768 24840
rect 38654 24828 38660 24840
rect 38712 24828 38718 24880
rect 41386 24868 41414 24908
rect 42886 24868 42892 24880
rect 41386 24840 42892 24868
rect 42886 24828 42892 24840
rect 42944 24828 42950 24880
rect 28108 24800 28181 24803
rect 27580 24797 28181 24800
rect 27580 24772 28136 24797
rect 27580 24760 27586 24772
rect 28534 24760 28540 24812
rect 28592 24800 28598 24812
rect 29089 24803 29147 24809
rect 29089 24800 29101 24803
rect 28592 24772 29101 24800
rect 28592 24760 28598 24772
rect 29089 24769 29101 24772
rect 29135 24769 29147 24803
rect 29089 24763 29147 24769
rect 29914 24760 29920 24812
rect 29972 24800 29978 24812
rect 30009 24803 30067 24809
rect 30009 24800 30021 24803
rect 29972 24772 30021 24800
rect 29972 24760 29978 24772
rect 30009 24769 30021 24772
rect 30055 24769 30067 24803
rect 30650 24800 30656 24812
rect 30611 24772 30656 24800
rect 30009 24763 30067 24769
rect 30650 24760 30656 24772
rect 30708 24760 30714 24812
rect 31570 24760 31576 24812
rect 31628 24800 31634 24812
rect 32122 24800 32128 24812
rect 31628 24772 31673 24800
rect 32083 24772 32128 24800
rect 31628 24760 31634 24772
rect 32122 24760 32128 24772
rect 32180 24760 32186 24812
rect 32214 24760 32220 24812
rect 32272 24800 32278 24812
rect 32309 24803 32367 24809
rect 32309 24800 32321 24803
rect 32272 24772 32321 24800
rect 32272 24760 32278 24772
rect 32309 24769 32321 24772
rect 32355 24769 32367 24803
rect 32309 24763 32367 24769
rect 32401 24803 32459 24809
rect 32401 24769 32413 24803
rect 32447 24800 32459 24803
rect 32674 24800 32680 24812
rect 32447 24772 32680 24800
rect 32447 24769 32459 24772
rect 32401 24763 32459 24769
rect 32674 24760 32680 24772
rect 32732 24760 32738 24812
rect 33137 24803 33195 24809
rect 33137 24800 33149 24803
rect 32876 24772 33149 24800
rect 19852 24704 22324 24732
rect 25225 24735 25283 24741
rect 19852 24692 19858 24704
rect 25225 24701 25237 24735
rect 25271 24732 25283 24735
rect 25498 24732 25504 24744
rect 25271 24704 25504 24732
rect 25271 24701 25283 24704
rect 25225 24695 25283 24701
rect 25498 24692 25504 24704
rect 25556 24692 25562 24744
rect 25682 24692 25688 24744
rect 25740 24732 25746 24744
rect 28997 24735 29055 24741
rect 28997 24732 29009 24735
rect 25740 24704 29009 24732
rect 25740 24692 25746 24704
rect 28997 24701 29009 24704
rect 29043 24701 29055 24735
rect 28997 24695 29055 24701
rect 29178 24692 29184 24744
rect 29236 24732 29242 24744
rect 29638 24732 29644 24744
rect 29236 24704 29644 24732
rect 29236 24692 29242 24704
rect 29638 24692 29644 24704
rect 29696 24732 29702 24744
rect 29733 24735 29791 24741
rect 29733 24732 29745 24735
rect 29696 24704 29745 24732
rect 29696 24692 29702 24704
rect 29733 24701 29745 24704
rect 29779 24701 29791 24735
rect 29733 24695 29791 24701
rect 30558 24692 30564 24744
rect 30616 24732 30622 24744
rect 31846 24732 31852 24744
rect 30616 24704 31852 24732
rect 30616 24692 30622 24704
rect 31846 24692 31852 24704
rect 31904 24692 31910 24744
rect 32030 24692 32036 24744
rect 32088 24732 32094 24744
rect 32876 24732 32904 24772
rect 33137 24769 33149 24772
rect 33183 24769 33195 24803
rect 33962 24800 33968 24812
rect 33923 24772 33968 24800
rect 33137 24763 33195 24769
rect 33962 24760 33968 24772
rect 34020 24760 34026 24812
rect 34149 24803 34207 24809
rect 34149 24769 34161 24803
rect 34195 24800 34207 24803
rect 34606 24800 34612 24812
rect 34195 24772 34612 24800
rect 34195 24769 34207 24772
rect 34149 24763 34207 24769
rect 34606 24760 34612 24772
rect 34664 24760 34670 24812
rect 34793 24803 34851 24809
rect 34793 24769 34805 24803
rect 34839 24800 34851 24803
rect 35158 24800 35164 24812
rect 34839 24772 35164 24800
rect 34839 24769 34851 24772
rect 34793 24763 34851 24769
rect 35158 24760 35164 24772
rect 35216 24760 35222 24812
rect 35529 24803 35587 24809
rect 35529 24769 35541 24803
rect 35575 24800 35587 24803
rect 35618 24800 35624 24812
rect 35575 24772 35624 24800
rect 35575 24769 35587 24772
rect 35529 24763 35587 24769
rect 35618 24760 35624 24772
rect 35676 24800 35682 24812
rect 35802 24800 35808 24812
rect 35676 24772 35808 24800
rect 35676 24760 35682 24772
rect 35802 24760 35808 24772
rect 35860 24760 35866 24812
rect 36170 24800 36176 24812
rect 36131 24772 36176 24800
rect 36170 24760 36176 24772
rect 36228 24760 36234 24812
rect 36722 24800 36728 24812
rect 36635 24772 36728 24800
rect 36722 24760 36728 24772
rect 36780 24760 36786 24812
rect 40586 24800 40592 24812
rect 40547 24772 40592 24800
rect 40586 24760 40592 24772
rect 40644 24760 40650 24812
rect 35986 24732 35992 24744
rect 32088 24704 32904 24732
rect 34348 24704 35992 24732
rect 32088 24692 32094 24704
rect 8570 24624 8576 24676
rect 8628 24664 8634 24676
rect 11517 24667 11575 24673
rect 11517 24664 11529 24667
rect 8628 24636 11529 24664
rect 8628 24624 8634 24636
rect 11517 24633 11529 24636
rect 11563 24633 11575 24667
rect 11517 24627 11575 24633
rect 12342 24624 12348 24676
rect 12400 24664 12406 24676
rect 22189 24667 22247 24673
rect 12400 24636 22094 24664
rect 12400 24624 12406 24636
rect 1486 24596 1492 24608
rect 1447 24568 1492 24596
rect 1486 24556 1492 24568
rect 1544 24556 1550 24608
rect 22066 24596 22094 24636
rect 22189 24633 22201 24667
rect 22235 24664 22247 24667
rect 22278 24664 22284 24676
rect 22235 24636 22284 24664
rect 22235 24633 22247 24636
rect 22189 24627 22247 24633
rect 22278 24624 22284 24636
rect 22336 24664 22342 24676
rect 24118 24664 24124 24676
rect 22336 24636 24124 24664
rect 22336 24624 22342 24636
rect 24118 24624 24124 24636
rect 24176 24624 24182 24676
rect 25314 24624 25320 24676
rect 25372 24664 25378 24676
rect 27341 24667 27399 24673
rect 27341 24664 27353 24667
rect 25372 24636 27353 24664
rect 25372 24624 25378 24636
rect 27341 24633 27353 24636
rect 27387 24633 27399 24667
rect 27341 24627 27399 24633
rect 27706 24624 27712 24676
rect 27764 24664 27770 24676
rect 28261 24667 28319 24673
rect 27764 24636 28212 24664
rect 27764 24624 27770 24636
rect 22738 24596 22744 24608
rect 22066 24568 22744 24596
rect 22738 24556 22744 24568
rect 22796 24556 22802 24608
rect 23106 24556 23112 24608
rect 23164 24596 23170 24608
rect 23201 24599 23259 24605
rect 23201 24596 23213 24599
rect 23164 24568 23213 24596
rect 23164 24556 23170 24568
rect 23201 24565 23213 24568
rect 23247 24565 23259 24599
rect 23201 24559 23259 24565
rect 24213 24599 24271 24605
rect 24213 24565 24225 24599
rect 24259 24596 24271 24599
rect 24394 24596 24400 24608
rect 24259 24568 24400 24596
rect 24259 24565 24271 24568
rect 24213 24559 24271 24565
rect 24394 24556 24400 24568
rect 24452 24556 24458 24608
rect 24765 24599 24823 24605
rect 24765 24565 24777 24599
rect 24811 24596 24823 24599
rect 25406 24596 25412 24608
rect 24811 24568 25412 24596
rect 24811 24565 24823 24568
rect 24765 24559 24823 24565
rect 25406 24556 25412 24568
rect 25464 24556 25470 24608
rect 25590 24556 25596 24608
rect 25648 24596 25654 24608
rect 25777 24599 25835 24605
rect 25777 24596 25789 24599
rect 25648 24568 25789 24596
rect 25648 24556 25654 24568
rect 25777 24565 25789 24568
rect 25823 24565 25835 24599
rect 25777 24559 25835 24565
rect 26142 24556 26148 24608
rect 26200 24596 26206 24608
rect 26326 24596 26332 24608
rect 26200 24568 26332 24596
rect 26200 24556 26206 24568
rect 26326 24556 26332 24568
rect 26384 24556 26390 24608
rect 26510 24556 26516 24608
rect 26568 24596 26574 24608
rect 28077 24599 28135 24605
rect 28077 24596 28089 24599
rect 26568 24568 28089 24596
rect 26568 24556 26574 24568
rect 28077 24565 28089 24568
rect 28123 24565 28135 24599
rect 28184 24596 28212 24636
rect 28261 24633 28273 24667
rect 28307 24664 28319 24667
rect 31754 24664 31760 24676
rect 28307 24636 28994 24664
rect 28307 24633 28319 24636
rect 28261 24627 28319 24633
rect 28813 24599 28871 24605
rect 28813 24596 28825 24599
rect 28184 24568 28825 24596
rect 28077 24559 28135 24565
rect 28813 24565 28825 24568
rect 28859 24565 28871 24599
rect 28966 24596 28994 24636
rect 30760 24636 31760 24664
rect 30760 24596 30788 24636
rect 31754 24624 31760 24636
rect 31812 24624 31818 24676
rect 32677 24667 32735 24673
rect 32677 24633 32689 24667
rect 32723 24664 32735 24667
rect 34348 24664 34376 24704
rect 35986 24692 35992 24704
rect 36044 24692 36050 24744
rect 36446 24692 36452 24744
rect 36504 24732 36510 24744
rect 37829 24735 37887 24741
rect 37829 24732 37841 24735
rect 36504 24704 37841 24732
rect 36504 24692 36510 24704
rect 37829 24701 37841 24704
rect 37875 24701 37887 24735
rect 37829 24695 37887 24701
rect 32723 24636 34376 24664
rect 32723 24633 32735 24636
rect 32677 24627 32735 24633
rect 34422 24624 34428 24676
rect 34480 24664 34486 24676
rect 34609 24667 34667 24673
rect 34609 24664 34621 24667
rect 34480 24636 34621 24664
rect 34480 24624 34486 24636
rect 34609 24633 34621 24636
rect 34655 24633 34667 24667
rect 34609 24627 34667 24633
rect 36170 24624 36176 24676
rect 36228 24664 36234 24676
rect 38381 24667 38439 24673
rect 38381 24664 38393 24667
rect 36228 24636 38393 24664
rect 36228 24624 36234 24636
rect 38381 24633 38393 24636
rect 38427 24633 38439 24667
rect 38381 24627 38439 24633
rect 40129 24667 40187 24673
rect 40129 24633 40141 24667
rect 40175 24664 40187 24667
rect 44542 24664 44548 24676
rect 40175 24636 44548 24664
rect 40175 24633 40187 24636
rect 40129 24627 40187 24633
rect 44542 24624 44548 24636
rect 44600 24624 44606 24676
rect 28966 24568 30788 24596
rect 30837 24599 30895 24605
rect 28813 24559 28871 24565
rect 30837 24565 30849 24599
rect 30883 24596 30895 24599
rect 31294 24596 31300 24608
rect 30883 24568 31300 24596
rect 30883 24565 30895 24568
rect 30837 24559 30895 24565
rect 31294 24556 31300 24568
rect 31352 24556 31358 24608
rect 31478 24596 31484 24608
rect 31439 24568 31484 24596
rect 31478 24556 31484 24568
rect 31536 24556 31542 24608
rect 32030 24556 32036 24608
rect 32088 24596 32094 24608
rect 32398 24596 32404 24608
rect 32088 24568 32404 24596
rect 32088 24556 32094 24568
rect 32398 24556 32404 24568
rect 32456 24556 32462 24608
rect 33134 24596 33140 24608
rect 33095 24568 33140 24596
rect 33134 24556 33140 24568
rect 33192 24556 33198 24608
rect 34514 24556 34520 24608
rect 34572 24596 34578 24608
rect 35437 24599 35495 24605
rect 35437 24596 35449 24599
rect 34572 24568 35449 24596
rect 34572 24556 34578 24568
rect 35437 24565 35449 24568
rect 35483 24565 35495 24599
rect 36078 24596 36084 24608
rect 36039 24568 36084 24596
rect 35437 24559 35495 24565
rect 36078 24556 36084 24568
rect 36136 24556 36142 24608
rect 37274 24596 37280 24608
rect 37235 24568 37280 24596
rect 37274 24556 37280 24568
rect 37332 24556 37338 24608
rect 38562 24556 38568 24608
rect 38620 24596 38626 24608
rect 38933 24599 38991 24605
rect 38933 24596 38945 24599
rect 38620 24568 38945 24596
rect 38620 24556 38626 24568
rect 38933 24565 38945 24568
rect 38979 24565 38991 24599
rect 39482 24596 39488 24608
rect 39443 24568 39488 24596
rect 38933 24559 38991 24565
rect 39482 24556 39488 24568
rect 39540 24556 39546 24608
rect 1104 24506 58880 24528
rect 1104 24454 10582 24506
rect 10634 24454 10646 24506
rect 10698 24454 10710 24506
rect 10762 24454 10774 24506
rect 10826 24454 10838 24506
rect 10890 24454 29846 24506
rect 29898 24454 29910 24506
rect 29962 24454 29974 24506
rect 30026 24454 30038 24506
rect 30090 24454 30102 24506
rect 30154 24454 49110 24506
rect 49162 24454 49174 24506
rect 49226 24454 49238 24506
rect 49290 24454 49302 24506
rect 49354 24454 49366 24506
rect 49418 24454 58880 24506
rect 1104 24432 58880 24454
rect 9122 24352 9128 24404
rect 9180 24392 9186 24404
rect 16669 24395 16727 24401
rect 16669 24392 16681 24395
rect 9180 24364 16681 24392
rect 9180 24352 9186 24364
rect 16669 24361 16681 24364
rect 16715 24361 16727 24395
rect 16669 24355 16727 24361
rect 17405 24395 17463 24401
rect 17405 24361 17417 24395
rect 17451 24392 17463 24395
rect 23382 24392 23388 24404
rect 17451 24364 23388 24392
rect 17451 24361 17463 24364
rect 17405 24355 17463 24361
rect 14366 24284 14372 24336
rect 14424 24324 14430 24336
rect 14461 24327 14519 24333
rect 14461 24324 14473 24327
rect 14424 24296 14473 24324
rect 14424 24284 14430 24296
rect 14461 24293 14473 24296
rect 14507 24293 14519 24327
rect 14461 24287 14519 24293
rect 16761 24191 16819 24197
rect 16761 24157 16773 24191
rect 16807 24188 16819 24191
rect 17420 24188 17448 24355
rect 23382 24352 23388 24364
rect 23440 24352 23446 24404
rect 23845 24395 23903 24401
rect 23845 24361 23857 24395
rect 23891 24392 23903 24395
rect 27154 24392 27160 24404
rect 23891 24364 27160 24392
rect 23891 24361 23903 24364
rect 23845 24355 23903 24361
rect 27154 24352 27160 24364
rect 27212 24352 27218 24404
rect 27246 24352 27252 24404
rect 27304 24392 27310 24404
rect 32766 24392 32772 24404
rect 27304 24364 32772 24392
rect 27304 24352 27310 24364
rect 32766 24352 32772 24364
rect 32824 24352 32830 24404
rect 33502 24352 33508 24404
rect 33560 24392 33566 24404
rect 33965 24395 34023 24401
rect 33965 24392 33977 24395
rect 33560 24364 33977 24392
rect 33560 24352 33566 24364
rect 33965 24361 33977 24364
rect 34011 24392 34023 24395
rect 34698 24392 34704 24404
rect 34011 24364 34704 24392
rect 34011 24361 34023 24364
rect 33965 24355 34023 24361
rect 34698 24352 34704 24364
rect 34756 24352 34762 24404
rect 36262 24392 36268 24404
rect 34808 24364 36268 24392
rect 19242 24284 19248 24336
rect 19300 24324 19306 24336
rect 21634 24324 21640 24336
rect 19300 24284 19334 24324
rect 21595 24296 21640 24324
rect 21634 24284 21640 24296
rect 21692 24284 21698 24336
rect 22189 24327 22247 24333
rect 22189 24293 22201 24327
rect 22235 24324 22247 24327
rect 23566 24324 23572 24336
rect 22235 24296 23572 24324
rect 22235 24293 22247 24296
rect 22189 24287 22247 24293
rect 23566 24284 23572 24296
rect 23624 24284 23630 24336
rect 25593 24327 25651 24333
rect 25593 24293 25605 24327
rect 25639 24324 25651 24327
rect 27430 24324 27436 24336
rect 25639 24296 27436 24324
rect 25639 24293 25651 24296
rect 25593 24287 25651 24293
rect 27430 24284 27436 24296
rect 27488 24324 27494 24336
rect 30558 24324 30564 24336
rect 27488 24296 27614 24324
rect 27488 24284 27494 24296
rect 16807 24160 17448 24188
rect 19306 24188 19334 24284
rect 22002 24216 22008 24268
rect 22060 24256 22066 24268
rect 25222 24256 25228 24268
rect 22060 24228 25228 24256
rect 22060 24216 22066 24228
rect 25222 24216 25228 24228
rect 25280 24256 25286 24268
rect 27586 24256 27614 24296
rect 27908 24296 30564 24324
rect 27908 24265 27936 24296
rect 30558 24284 30564 24296
rect 30616 24284 30622 24336
rect 33870 24324 33876 24336
rect 33245 24296 33876 24324
rect 27893 24259 27951 24265
rect 25280 24228 26832 24256
rect 27586 24228 27844 24256
rect 25280 24216 25286 24228
rect 21085 24191 21143 24197
rect 21085 24188 21097 24191
rect 19306 24160 21097 24188
rect 16807 24157 16819 24160
rect 16761 24151 16819 24157
rect 21085 24157 21097 24160
rect 21131 24188 21143 24191
rect 22278 24188 22284 24200
rect 21131 24160 22284 24188
rect 21131 24157 21143 24160
rect 21085 24151 21143 24157
rect 22278 24148 22284 24160
rect 22336 24148 22342 24200
rect 22922 24148 22928 24200
rect 22980 24188 22986 24200
rect 23293 24191 23351 24197
rect 23293 24188 23305 24191
rect 22980 24160 23305 24188
rect 22980 24148 22986 24160
rect 23293 24157 23305 24160
rect 23339 24188 23351 24191
rect 23339 24160 25912 24188
rect 23339 24157 23351 24160
rect 23293 24151 23351 24157
rect 14645 24123 14703 24129
rect 14645 24089 14657 24123
rect 14691 24120 14703 24123
rect 23658 24120 23664 24132
rect 14691 24092 23664 24120
rect 14691 24089 14703 24092
rect 14645 24083 14703 24089
rect 23658 24080 23664 24092
rect 23716 24080 23722 24132
rect 25041 24123 25099 24129
rect 24412 24092 24716 24120
rect 22002 24012 22008 24064
rect 22060 24052 22066 24064
rect 22649 24055 22707 24061
rect 22649 24052 22661 24055
rect 22060 24024 22661 24052
rect 22060 24012 22066 24024
rect 22649 24021 22661 24024
rect 22695 24021 22707 24055
rect 22649 24015 22707 24021
rect 23566 24012 23572 24064
rect 23624 24052 23630 24064
rect 24412 24052 24440 24092
rect 23624 24024 24440 24052
rect 24489 24055 24547 24061
rect 23624 24012 23630 24024
rect 24489 24021 24501 24055
rect 24535 24052 24547 24055
rect 24578 24052 24584 24064
rect 24535 24024 24584 24052
rect 24535 24021 24547 24024
rect 24489 24015 24547 24021
rect 24578 24012 24584 24024
rect 24636 24012 24642 24064
rect 24688 24052 24716 24092
rect 25041 24089 25053 24123
rect 25087 24120 25099 24123
rect 25406 24120 25412 24132
rect 25087 24092 25412 24120
rect 25087 24089 25099 24092
rect 25041 24083 25099 24089
rect 25406 24080 25412 24092
rect 25464 24080 25470 24132
rect 25884 24120 25912 24160
rect 25958 24148 25964 24200
rect 26016 24188 26022 24200
rect 26804 24197 26832 24228
rect 26053 24191 26111 24197
rect 26053 24188 26065 24191
rect 26016 24160 26065 24188
rect 26016 24148 26022 24160
rect 26053 24157 26065 24160
rect 26099 24157 26111 24191
rect 26053 24151 26111 24157
rect 26789 24191 26847 24197
rect 26789 24157 26801 24191
rect 26835 24157 26847 24191
rect 27246 24188 27252 24200
rect 26789 24151 26847 24157
rect 26896 24160 27252 24188
rect 26694 24120 26700 24132
rect 25884 24092 26280 24120
rect 26655 24092 26700 24120
rect 25866 24052 25872 24064
rect 24688 24024 25872 24052
rect 25866 24012 25872 24024
rect 25924 24012 25930 24064
rect 26142 24052 26148 24064
rect 26103 24024 26148 24052
rect 26142 24012 26148 24024
rect 26200 24012 26206 24064
rect 26252 24052 26280 24092
rect 26694 24080 26700 24092
rect 26752 24080 26758 24132
rect 26896 24120 26924 24160
rect 27246 24148 27252 24160
rect 27304 24148 27310 24200
rect 27338 24148 27344 24200
rect 27396 24188 27402 24200
rect 27723 24191 27781 24197
rect 27723 24188 27735 24191
rect 27396 24160 27735 24188
rect 27396 24148 27402 24160
rect 27723 24157 27735 24160
rect 27769 24157 27781 24191
rect 27816 24188 27844 24228
rect 27893 24225 27905 24259
rect 27939 24225 27951 24259
rect 27893 24219 27951 24225
rect 28074 24216 28080 24268
rect 28132 24256 28138 24268
rect 28718 24256 28724 24268
rect 28132 24228 28724 24256
rect 28132 24216 28138 24228
rect 28718 24216 28724 24228
rect 28776 24256 28782 24268
rect 28997 24259 29055 24265
rect 28997 24256 29009 24259
rect 28776 24228 29009 24256
rect 28776 24216 28782 24228
rect 28997 24225 29009 24228
rect 29043 24256 29055 24259
rect 29638 24256 29644 24268
rect 29043 24228 29500 24256
rect 29599 24228 29644 24256
rect 29043 24225 29055 24228
rect 28997 24219 29055 24225
rect 28813 24191 28871 24197
rect 28813 24188 28825 24191
rect 27816 24160 28825 24188
rect 27723 24151 27781 24157
rect 28813 24157 28825 24160
rect 28859 24157 28871 24191
rect 28813 24151 28871 24157
rect 26804 24092 26924 24120
rect 26804 24052 26832 24092
rect 26970 24080 26976 24132
rect 27028 24120 27034 24132
rect 28258 24120 28264 24132
rect 27028 24092 28264 24120
rect 27028 24080 27034 24092
rect 28258 24080 28264 24092
rect 28316 24120 28322 24132
rect 28629 24123 28687 24129
rect 28629 24120 28641 24123
rect 28316 24092 28641 24120
rect 28316 24080 28322 24092
rect 28629 24089 28641 24092
rect 28675 24089 28687 24123
rect 29472 24120 29500 24228
rect 29638 24216 29644 24228
rect 29696 24216 29702 24268
rect 30484 24228 32476 24256
rect 29733 24191 29791 24197
rect 29733 24157 29745 24191
rect 29779 24188 29791 24191
rect 30374 24188 30380 24200
rect 29779 24160 30380 24188
rect 29779 24157 29791 24160
rect 29733 24151 29791 24157
rect 30374 24148 30380 24160
rect 30432 24148 30438 24200
rect 30484 24120 30512 24228
rect 32306 24148 32312 24200
rect 32364 24188 32370 24200
rect 32448 24188 32476 24228
rect 32582 24216 32588 24268
rect 32640 24256 32646 24268
rect 32769 24259 32827 24265
rect 32769 24256 32781 24259
rect 32640 24228 32781 24256
rect 32640 24216 32646 24228
rect 32769 24225 32781 24228
rect 32815 24225 32827 24259
rect 32769 24219 32827 24225
rect 32950 24216 32956 24268
rect 33008 24256 33014 24268
rect 33245 24265 33273 24296
rect 33870 24284 33876 24296
rect 33928 24284 33934 24336
rect 34146 24324 34152 24336
rect 34107 24296 34152 24324
rect 34146 24284 34152 24296
rect 34204 24284 34210 24336
rect 34238 24284 34244 24336
rect 34296 24324 34302 24336
rect 34808 24324 34836 24364
rect 36262 24352 36268 24364
rect 36320 24352 36326 24404
rect 38378 24352 38384 24404
rect 38436 24392 38442 24404
rect 39298 24392 39304 24404
rect 38436 24364 39304 24392
rect 38436 24352 38442 24364
rect 39298 24352 39304 24364
rect 39356 24352 39362 24404
rect 40497 24395 40555 24401
rect 40497 24361 40509 24395
rect 40543 24392 40555 24395
rect 40586 24392 40592 24404
rect 40543 24364 40592 24392
rect 40543 24361 40555 24364
rect 40497 24355 40555 24361
rect 40586 24352 40592 24364
rect 40644 24352 40650 24404
rect 34296 24296 34836 24324
rect 34885 24327 34943 24333
rect 34296 24284 34302 24296
rect 34885 24293 34897 24327
rect 34931 24324 34943 24327
rect 36814 24324 36820 24336
rect 34931 24296 36820 24324
rect 34931 24293 34943 24296
rect 34885 24287 34943 24293
rect 36814 24284 36820 24296
rect 36872 24284 36878 24336
rect 36909 24327 36967 24333
rect 36909 24293 36921 24327
rect 36955 24324 36967 24327
rect 41690 24324 41696 24336
rect 36955 24296 41696 24324
rect 36955 24293 36967 24296
rect 36909 24287 36967 24293
rect 41690 24284 41696 24296
rect 41748 24284 41754 24336
rect 33230 24259 33288 24265
rect 33008 24228 33053 24256
rect 33008 24216 33014 24228
rect 33230 24225 33242 24259
rect 33276 24225 33288 24259
rect 33230 24219 33288 24225
rect 34422 24216 34428 24268
rect 34480 24256 34486 24268
rect 34480 24228 37504 24256
rect 34480 24216 34486 24228
rect 33045 24191 33103 24197
rect 32364 24160 32409 24188
rect 32448 24160 32812 24188
rect 32364 24148 32370 24160
rect 29472 24092 30512 24120
rect 28629 24083 28687 24089
rect 31478 24080 31484 24132
rect 31536 24080 31542 24132
rect 32030 24120 32036 24132
rect 31991 24092 32036 24120
rect 32030 24080 32036 24092
rect 32088 24080 32094 24132
rect 26252 24024 26832 24052
rect 26878 24012 26884 24064
rect 26936 24052 26942 24064
rect 27433 24055 27491 24061
rect 27433 24052 27445 24055
rect 26936 24024 27445 24052
rect 26936 24012 26942 24024
rect 27433 24021 27445 24024
rect 27479 24021 27491 24055
rect 27433 24015 27491 24021
rect 27982 24012 27988 24064
rect 28040 24052 28046 24064
rect 28445 24055 28503 24061
rect 28445 24052 28457 24055
rect 28040 24024 28457 24052
rect 28040 24012 28046 24024
rect 28445 24021 28457 24024
rect 28491 24021 28503 24055
rect 28445 24015 28503 24021
rect 28534 24012 28540 24064
rect 28592 24052 28598 24064
rect 28721 24055 28779 24061
rect 28721 24052 28733 24055
rect 28592 24024 28733 24052
rect 28592 24012 28598 24024
rect 28721 24021 28733 24024
rect 28767 24021 28779 24055
rect 28721 24015 28779 24021
rect 28810 24012 28816 24064
rect 28868 24052 28874 24064
rect 29086 24052 29092 24064
rect 28868 24024 29092 24052
rect 28868 24012 28874 24024
rect 29086 24012 29092 24024
rect 29144 24012 29150 24064
rect 30098 24052 30104 24064
rect 30059 24024 30104 24052
rect 30098 24012 30104 24024
rect 30156 24012 30162 24064
rect 30561 24055 30619 24061
rect 30561 24021 30573 24055
rect 30607 24052 30619 24055
rect 32122 24052 32128 24064
rect 30607 24024 32128 24052
rect 30607 24021 30619 24024
rect 30561 24015 30619 24021
rect 32122 24012 32128 24024
rect 32180 24012 32186 24064
rect 32784 24052 32812 24160
rect 33045 24157 33057 24191
rect 33091 24157 33103 24191
rect 33045 24151 33103 24157
rect 33137 24191 33195 24197
rect 33137 24157 33149 24191
rect 33183 24190 33195 24191
rect 33318 24190 33324 24200
rect 33183 24162 33324 24190
rect 33183 24157 33195 24162
rect 33137 24151 33195 24157
rect 32858 24080 32864 24132
rect 32916 24120 32922 24132
rect 33060 24120 33088 24151
rect 33318 24148 33324 24162
rect 33376 24188 33382 24200
rect 33686 24188 33692 24200
rect 33376 24160 33692 24188
rect 33376 24148 33382 24160
rect 33686 24148 33692 24160
rect 33744 24148 33750 24200
rect 33870 24148 33876 24200
rect 33928 24188 33934 24200
rect 34701 24191 34759 24197
rect 34701 24188 34713 24191
rect 33928 24160 34713 24188
rect 33928 24148 33934 24160
rect 34701 24157 34713 24160
rect 34747 24188 34759 24191
rect 34882 24188 34888 24200
rect 34747 24160 34888 24188
rect 34747 24157 34759 24160
rect 34701 24151 34759 24157
rect 34882 24148 34888 24160
rect 34940 24148 34946 24200
rect 35526 24188 35532 24200
rect 35487 24160 35532 24188
rect 35526 24148 35532 24160
rect 35584 24148 35590 24200
rect 36170 24188 36176 24200
rect 36131 24160 36176 24188
rect 36170 24148 36176 24160
rect 36228 24148 36234 24200
rect 36262 24148 36268 24200
rect 36320 24188 36326 24200
rect 36817 24191 36875 24197
rect 36817 24188 36829 24191
rect 36320 24160 36829 24188
rect 36320 24148 36326 24160
rect 36817 24157 36829 24160
rect 36863 24188 36875 24191
rect 37366 24188 37372 24200
rect 36863 24160 37372 24188
rect 36863 24157 36875 24160
rect 36817 24151 36875 24157
rect 37366 24148 37372 24160
rect 37424 24148 37430 24200
rect 37476 24197 37504 24228
rect 39114 24216 39120 24268
rect 39172 24256 39178 24268
rect 39209 24259 39267 24265
rect 39209 24256 39221 24259
rect 39172 24228 39221 24256
rect 39172 24216 39178 24228
rect 39209 24225 39221 24228
rect 39255 24225 39267 24259
rect 39209 24219 39267 24225
rect 37461 24191 37519 24197
rect 37461 24157 37473 24191
rect 37507 24157 37519 24191
rect 37461 24151 37519 24157
rect 38286 24148 38292 24200
rect 38344 24188 38350 24200
rect 40770 24188 40776 24200
rect 38344 24160 40776 24188
rect 38344 24148 38350 24160
rect 40770 24148 40776 24160
rect 40828 24148 40834 24200
rect 58158 24188 58164 24200
rect 58119 24160 58164 24188
rect 58158 24148 58164 24160
rect 58216 24148 58222 24200
rect 32916 24092 33088 24120
rect 32916 24080 32922 24092
rect 33410 24080 33416 24132
rect 33468 24120 33474 24132
rect 33778 24120 33784 24132
rect 33468 24092 33784 24120
rect 33468 24080 33474 24092
rect 33778 24080 33784 24092
rect 33836 24080 33842 24132
rect 34054 24129 34060 24132
rect 33997 24123 34060 24129
rect 33997 24089 34009 24123
rect 34043 24089 34060 24123
rect 33997 24083 34060 24089
rect 34054 24080 34060 24083
rect 34112 24080 34118 24132
rect 35618 24080 35624 24132
rect 35676 24120 35682 24132
rect 37553 24123 37611 24129
rect 37553 24120 37565 24123
rect 35676 24092 37565 24120
rect 35676 24080 35682 24092
rect 37553 24089 37565 24092
rect 37599 24089 37611 24123
rect 37553 24083 37611 24089
rect 38102 24080 38108 24132
rect 38160 24120 38166 24132
rect 38746 24120 38752 24132
rect 38160 24092 38752 24120
rect 38160 24080 38166 24092
rect 38746 24080 38752 24092
rect 38804 24120 38810 24132
rect 39853 24123 39911 24129
rect 39853 24120 39865 24123
rect 38804 24092 39865 24120
rect 38804 24080 38810 24092
rect 39853 24089 39865 24092
rect 39899 24120 39911 24123
rect 40957 24123 41015 24129
rect 40957 24120 40969 24123
rect 39899 24092 40969 24120
rect 39899 24089 39911 24092
rect 39853 24083 39911 24089
rect 40957 24089 40969 24092
rect 41003 24120 41015 24123
rect 41003 24092 41414 24120
rect 41003 24089 41015 24092
rect 40957 24083 41015 24089
rect 35526 24052 35532 24064
rect 32784 24024 35532 24052
rect 35526 24012 35532 24024
rect 35584 24012 35590 24064
rect 35713 24055 35771 24061
rect 35713 24021 35725 24055
rect 35759 24052 35771 24055
rect 35986 24052 35992 24064
rect 35759 24024 35992 24052
rect 35759 24021 35771 24024
rect 35713 24015 35771 24021
rect 35986 24012 35992 24024
rect 36044 24012 36050 24064
rect 36262 24052 36268 24064
rect 36223 24024 36268 24052
rect 36262 24012 36268 24024
rect 36320 24012 36326 24064
rect 36906 24012 36912 24064
rect 36964 24052 36970 24064
rect 38197 24055 38255 24061
rect 38197 24052 38209 24055
rect 36964 24024 38209 24052
rect 36964 24012 36970 24024
rect 38197 24021 38209 24024
rect 38243 24052 38255 24055
rect 38378 24052 38384 24064
rect 38243 24024 38384 24052
rect 38243 24021 38255 24024
rect 38197 24015 38255 24021
rect 38378 24012 38384 24024
rect 38436 24012 38442 24064
rect 38657 24055 38715 24061
rect 38657 24021 38669 24055
rect 38703 24052 38715 24055
rect 38838 24052 38844 24064
rect 38703 24024 38844 24052
rect 38703 24021 38715 24024
rect 38657 24015 38715 24021
rect 38838 24012 38844 24024
rect 38896 24012 38902 24064
rect 41386 24052 41414 24092
rect 49694 24080 49700 24132
rect 49752 24120 49758 24132
rect 57885 24123 57943 24129
rect 57885 24120 57897 24123
rect 49752 24092 57897 24120
rect 49752 24080 49758 24092
rect 57885 24089 57897 24092
rect 57931 24089 57943 24123
rect 57885 24083 57943 24089
rect 42702 24052 42708 24064
rect 41386 24024 42708 24052
rect 42702 24012 42708 24024
rect 42760 24012 42766 24064
rect 1104 23962 58880 23984
rect 1104 23910 20214 23962
rect 20266 23910 20278 23962
rect 20330 23910 20342 23962
rect 20394 23910 20406 23962
rect 20458 23910 20470 23962
rect 20522 23910 39478 23962
rect 39530 23910 39542 23962
rect 39594 23910 39606 23962
rect 39658 23910 39670 23962
rect 39722 23910 39734 23962
rect 39786 23910 58880 23962
rect 1104 23888 58880 23910
rect 18598 23808 18604 23860
rect 18656 23848 18662 23860
rect 25682 23848 25688 23860
rect 18656 23820 25544 23848
rect 25643 23820 25688 23848
rect 18656 23808 18662 23820
rect 19978 23740 19984 23792
rect 20036 23780 20042 23792
rect 20165 23783 20223 23789
rect 20165 23780 20177 23783
rect 20036 23752 20177 23780
rect 20036 23740 20042 23752
rect 20165 23749 20177 23752
rect 20211 23780 20223 23783
rect 20714 23780 20720 23792
rect 20211 23752 20720 23780
rect 20211 23749 20223 23752
rect 20165 23743 20223 23749
rect 20714 23740 20720 23752
rect 20772 23740 20778 23792
rect 24118 23740 24124 23792
rect 24176 23780 24182 23792
rect 25130 23780 25136 23792
rect 24176 23752 25136 23780
rect 24176 23740 24182 23752
rect 25130 23740 25136 23752
rect 25188 23740 25194 23792
rect 25516 23721 25544 23820
rect 25682 23808 25688 23820
rect 25740 23808 25746 23860
rect 25866 23808 25872 23860
rect 25924 23848 25930 23860
rect 28810 23848 28816 23860
rect 25924 23820 28816 23848
rect 25924 23808 25930 23820
rect 28810 23808 28816 23820
rect 28868 23848 28874 23860
rect 28868 23820 29040 23848
rect 28868 23808 28874 23820
rect 26326 23780 26332 23792
rect 25608 23752 26332 23780
rect 25608 23724 25636 23752
rect 25501 23715 25559 23721
rect 25501 23681 25513 23715
rect 25547 23681 25559 23715
rect 25501 23675 25559 23681
rect 25590 23672 25596 23724
rect 25648 23672 25654 23724
rect 25685 23715 25743 23721
rect 25685 23681 25697 23715
rect 25731 23712 25743 23715
rect 25774 23712 25780 23724
rect 25731 23684 25780 23712
rect 25731 23681 25743 23684
rect 25685 23675 25743 23681
rect 25774 23672 25780 23684
rect 25832 23672 25838 23724
rect 26160 23721 26188 23752
rect 26326 23740 26332 23752
rect 26384 23740 26390 23792
rect 28902 23780 28908 23792
rect 27172 23752 28908 23780
rect 26145 23715 26203 23721
rect 26145 23681 26157 23715
rect 26191 23681 26203 23715
rect 26145 23675 26203 23681
rect 26421 23715 26479 23721
rect 26421 23681 26433 23715
rect 26467 23712 26479 23715
rect 26602 23712 26608 23724
rect 26467 23684 26608 23712
rect 26467 23681 26479 23684
rect 26421 23675 26479 23681
rect 26602 23672 26608 23684
rect 26660 23672 26666 23724
rect 20530 23604 20536 23656
rect 20588 23644 20594 23656
rect 21913 23647 21971 23653
rect 21913 23644 21925 23647
rect 20588 23616 21925 23644
rect 20588 23604 20594 23616
rect 21913 23613 21925 23616
rect 21959 23644 21971 23647
rect 22002 23644 22008 23656
rect 21959 23616 22008 23644
rect 21959 23613 21971 23616
rect 21913 23607 21971 23613
rect 22002 23604 22008 23616
rect 22060 23604 22066 23656
rect 22830 23604 22836 23656
rect 22888 23644 22894 23656
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 22888 23616 24593 23644
rect 22888 23604 22894 23616
rect 24581 23613 24593 23616
rect 24627 23613 24639 23647
rect 24854 23644 24860 23656
rect 24767 23616 24860 23644
rect 24581 23607 24639 23613
rect 24854 23604 24860 23616
rect 24912 23644 24918 23656
rect 25866 23644 25872 23656
rect 24912 23616 25872 23644
rect 24912 23604 24918 23616
rect 25866 23604 25872 23616
rect 25924 23604 25930 23656
rect 27172 23644 27200 23752
rect 28902 23740 28908 23752
rect 28960 23740 28966 23792
rect 27246 23672 27252 23724
rect 27304 23712 27310 23724
rect 27433 23715 27491 23721
rect 27433 23712 27445 23715
rect 27304 23684 27445 23712
rect 27304 23672 27310 23684
rect 27433 23681 27445 23684
rect 27479 23681 27491 23715
rect 27433 23675 27491 23681
rect 27614 23672 27620 23724
rect 27672 23712 27678 23724
rect 28537 23715 28595 23721
rect 28537 23712 28549 23715
rect 27672 23684 28549 23712
rect 27672 23672 27678 23684
rect 28537 23681 28549 23684
rect 28583 23681 28595 23715
rect 28537 23675 28595 23681
rect 28813 23715 28871 23721
rect 28813 23681 28825 23715
rect 28859 23712 28871 23715
rect 29012 23712 29040 23820
rect 29086 23808 29092 23860
rect 29144 23848 29150 23860
rect 32125 23851 32183 23857
rect 32125 23848 32137 23851
rect 29144 23820 32137 23848
rect 29144 23808 29150 23820
rect 32125 23817 32137 23820
rect 32171 23817 32183 23851
rect 32125 23811 32183 23817
rect 35434 23808 35440 23860
rect 35492 23848 35498 23860
rect 35529 23851 35587 23857
rect 35529 23848 35541 23851
rect 35492 23820 35541 23848
rect 35492 23808 35498 23820
rect 35529 23817 35541 23820
rect 35575 23817 35587 23851
rect 35529 23811 35587 23817
rect 35894 23808 35900 23860
rect 35952 23848 35958 23860
rect 35952 23820 36675 23848
rect 35952 23808 35958 23820
rect 30282 23780 30288 23792
rect 29748 23752 30288 23780
rect 29546 23712 29552 23724
rect 28859 23684 29552 23712
rect 28859 23681 28871 23684
rect 28813 23675 28871 23681
rect 29546 23672 29552 23684
rect 29604 23672 29610 23724
rect 29748 23721 29776 23752
rect 30282 23740 30288 23752
rect 30340 23740 30346 23792
rect 30742 23740 30748 23792
rect 30800 23740 30806 23792
rect 32766 23740 32772 23792
rect 32824 23780 32830 23792
rect 36446 23780 36452 23792
rect 32824 23752 36452 23780
rect 32824 23740 32830 23752
rect 29733 23715 29791 23721
rect 29733 23681 29745 23715
rect 29779 23681 29791 23715
rect 32953 23715 33011 23721
rect 32953 23712 32965 23715
rect 29733 23675 29791 23681
rect 32508 23684 32965 23712
rect 27338 23644 27344 23656
rect 27080 23616 27200 23644
rect 27299 23616 27344 23644
rect 22557 23579 22615 23585
rect 22557 23545 22569 23579
rect 22603 23576 22615 23579
rect 23290 23576 23296 23588
rect 22603 23548 23296 23576
rect 22603 23545 22615 23548
rect 22557 23539 22615 23545
rect 23290 23536 23296 23548
rect 23348 23536 23354 23588
rect 26329 23579 26387 23585
rect 26329 23545 26341 23579
rect 26375 23545 26387 23579
rect 26329 23539 26387 23545
rect 26421 23579 26479 23585
rect 26421 23545 26433 23579
rect 26467 23576 26479 23579
rect 27080 23576 27108 23616
rect 27338 23604 27344 23616
rect 27396 23604 27402 23656
rect 27798 23604 27804 23656
rect 27856 23644 27862 23656
rect 29178 23644 29184 23656
rect 27856 23616 29184 23644
rect 27856 23604 27862 23616
rect 29178 23604 29184 23616
rect 29236 23604 29242 23656
rect 30006 23644 30012 23656
rect 29967 23616 30012 23644
rect 30006 23604 30012 23616
rect 30064 23604 30070 23656
rect 30650 23604 30656 23656
rect 30708 23644 30714 23656
rect 31481 23647 31539 23653
rect 31481 23644 31493 23647
rect 30708 23616 31493 23644
rect 30708 23604 30714 23616
rect 31481 23613 31493 23616
rect 31527 23613 31539 23647
rect 32508 23644 32536 23684
rect 32953 23681 32965 23684
rect 32999 23712 33011 23715
rect 33042 23712 33048 23724
rect 32999 23684 33048 23712
rect 32999 23681 33011 23684
rect 32953 23675 33011 23681
rect 33042 23672 33048 23684
rect 33100 23672 33106 23724
rect 33870 23712 33876 23724
rect 33831 23684 33876 23712
rect 33870 23672 33876 23684
rect 33928 23672 33934 23724
rect 34790 23672 34796 23724
rect 34848 23712 34854 23724
rect 35066 23712 35072 23724
rect 34848 23684 35072 23712
rect 34848 23672 34854 23684
rect 35066 23672 35072 23684
rect 35124 23672 35130 23724
rect 35710 23712 35716 23724
rect 35671 23684 35716 23712
rect 35710 23672 35716 23684
rect 35768 23672 35774 23724
rect 35820 23721 35848 23752
rect 35805 23715 35863 23721
rect 35805 23681 35817 23715
rect 35851 23681 35863 23715
rect 35805 23675 35863 23681
rect 36188 23656 36216 23752
rect 36446 23740 36452 23752
rect 36504 23740 36510 23792
rect 36647 23780 36675 23820
rect 36998 23808 37004 23860
rect 37056 23848 37062 23860
rect 40218 23848 40224 23860
rect 37056 23820 40224 23848
rect 37056 23808 37062 23820
rect 40218 23808 40224 23820
rect 40276 23808 40282 23860
rect 40586 23808 40592 23860
rect 40644 23848 40650 23860
rect 40773 23851 40831 23857
rect 40773 23848 40785 23851
rect 40644 23820 40785 23848
rect 40644 23808 40650 23820
rect 40773 23817 40785 23820
rect 40819 23817 40831 23851
rect 58158 23848 58164 23860
rect 58119 23820 58164 23848
rect 40773 23811 40831 23817
rect 58158 23808 58164 23820
rect 58216 23808 58222 23860
rect 42058 23780 42064 23792
rect 36647 23752 42064 23780
rect 42058 23740 42064 23752
rect 42116 23740 42122 23792
rect 36633 23715 36691 23721
rect 36633 23681 36645 23715
rect 36679 23712 36691 23715
rect 36679 23684 37136 23712
rect 36679 23681 36691 23684
rect 36633 23675 36691 23681
rect 32858 23644 32864 23656
rect 31481 23607 31539 23613
rect 31726 23616 32536 23644
rect 32819 23616 32864 23644
rect 26467 23548 27108 23576
rect 26467 23545 26479 23548
rect 26421 23539 26479 23545
rect 21266 23508 21272 23520
rect 21227 23480 21272 23508
rect 21266 23468 21272 23480
rect 21324 23468 21330 23520
rect 21726 23468 21732 23520
rect 21784 23508 21790 23520
rect 23109 23511 23167 23517
rect 23109 23508 23121 23511
rect 21784 23480 23121 23508
rect 21784 23468 21790 23480
rect 23109 23477 23121 23480
rect 23155 23508 23167 23511
rect 26344 23508 26372 23539
rect 27154 23536 27160 23588
rect 27212 23576 27218 23588
rect 28353 23579 28411 23585
rect 28353 23576 28365 23579
rect 27212 23548 28365 23576
rect 27212 23536 27218 23548
rect 28353 23545 28365 23548
rect 28399 23545 28411 23579
rect 28718 23576 28724 23588
rect 28679 23548 28724 23576
rect 28353 23539 28411 23545
rect 28718 23536 28724 23548
rect 28776 23536 28782 23588
rect 31726 23576 31754 23616
rect 32858 23604 32864 23616
rect 32916 23604 32922 23656
rect 33962 23644 33968 23656
rect 33923 23616 33968 23644
rect 33962 23604 33968 23616
rect 34020 23604 34026 23656
rect 34977 23647 35035 23653
rect 34977 23644 34989 23647
rect 34072 23616 34989 23644
rect 31036 23548 31754 23576
rect 26510 23508 26516 23520
rect 23155 23480 26516 23508
rect 23155 23477 23167 23480
rect 23109 23471 23167 23477
rect 26510 23468 26516 23480
rect 26568 23468 26574 23520
rect 27338 23468 27344 23520
rect 27396 23508 27402 23520
rect 27614 23508 27620 23520
rect 27396 23480 27620 23508
rect 27396 23468 27402 23480
rect 27614 23468 27620 23480
rect 27672 23468 27678 23520
rect 27709 23511 27767 23517
rect 27709 23477 27721 23511
rect 27755 23508 27767 23511
rect 28258 23508 28264 23520
rect 27755 23480 28264 23508
rect 27755 23477 27767 23480
rect 27709 23471 27767 23477
rect 28258 23468 28264 23480
rect 28316 23468 28322 23520
rect 30190 23468 30196 23520
rect 30248 23508 30254 23520
rect 31036 23508 31064 23548
rect 31938 23536 31944 23588
rect 31996 23576 32002 23588
rect 34072 23576 34100 23616
rect 34977 23613 34989 23616
rect 35023 23644 35035 23647
rect 35894 23644 35900 23656
rect 35023 23616 35900 23644
rect 35023 23613 35035 23616
rect 34977 23607 35035 23613
rect 35894 23604 35900 23616
rect 35952 23604 35958 23656
rect 36170 23604 36176 23656
rect 36228 23604 36234 23656
rect 36357 23647 36415 23653
rect 36357 23613 36369 23647
rect 36403 23644 36415 23647
rect 36906 23644 36912 23656
rect 36403 23616 36912 23644
rect 36403 23613 36415 23616
rect 36357 23607 36415 23613
rect 36906 23604 36912 23616
rect 36964 23604 36970 23656
rect 37108 23644 37136 23684
rect 37182 23672 37188 23724
rect 37240 23712 37246 23724
rect 37277 23715 37335 23721
rect 37277 23712 37289 23715
rect 37240 23684 37289 23712
rect 37240 23672 37246 23684
rect 37277 23681 37289 23684
rect 37323 23681 37335 23715
rect 37277 23675 37335 23681
rect 37366 23672 37372 23724
rect 37424 23712 37430 23724
rect 38102 23712 38108 23724
rect 37424 23684 38108 23712
rect 37424 23672 37430 23684
rect 38102 23672 38108 23684
rect 38160 23672 38166 23724
rect 39209 23715 39267 23721
rect 38948 23684 39160 23712
rect 38948 23644 38976 23684
rect 37108 23616 38976 23644
rect 39132 23644 39160 23684
rect 39209 23681 39221 23715
rect 39255 23712 39267 23715
rect 40494 23712 40500 23724
rect 39255 23684 40500 23712
rect 39255 23681 39267 23684
rect 39209 23675 39267 23681
rect 40494 23672 40500 23684
rect 40552 23672 40558 23724
rect 40770 23672 40776 23724
rect 40828 23712 40834 23724
rect 49694 23712 49700 23724
rect 40828 23684 49700 23712
rect 40828 23672 40834 23684
rect 49694 23672 49700 23684
rect 49752 23672 49758 23724
rect 40678 23644 40684 23656
rect 39132 23616 40684 23644
rect 40678 23604 40684 23616
rect 40736 23604 40742 23656
rect 34238 23576 34244 23588
rect 31996 23548 34100 23576
rect 34199 23548 34244 23576
rect 31996 23536 32002 23548
rect 34238 23536 34244 23548
rect 34296 23536 34302 23588
rect 34422 23536 34428 23588
rect 34480 23576 34486 23588
rect 36722 23576 36728 23588
rect 34480 23548 34560 23576
rect 34480 23536 34486 23548
rect 30248 23480 31064 23508
rect 34532 23508 34560 23548
rect 35084 23548 36728 23576
rect 35084 23517 35112 23548
rect 36722 23536 36728 23548
rect 36780 23536 36786 23588
rect 37461 23579 37519 23585
rect 37461 23545 37473 23579
rect 37507 23576 37519 23579
rect 38930 23576 38936 23588
rect 37507 23548 38936 23576
rect 37507 23545 37519 23548
rect 37461 23539 37519 23545
rect 38930 23536 38936 23548
rect 38988 23536 38994 23588
rect 40313 23579 40371 23585
rect 40313 23545 40325 23579
rect 40359 23576 40371 23579
rect 41230 23576 41236 23588
rect 40359 23548 41236 23576
rect 40359 23545 40371 23548
rect 40313 23539 40371 23545
rect 41230 23536 41236 23548
rect 41288 23536 41294 23588
rect 34701 23511 34759 23517
rect 34701 23508 34713 23511
rect 34532 23480 34713 23508
rect 30248 23468 30254 23480
rect 34701 23477 34713 23480
rect 34747 23477 34759 23511
rect 34701 23471 34759 23477
rect 35069 23511 35127 23517
rect 35069 23477 35081 23511
rect 35115 23477 35127 23511
rect 36446 23508 36452 23520
rect 36407 23480 36452 23508
rect 35069 23471 35127 23477
rect 36446 23468 36452 23480
rect 36504 23468 36510 23520
rect 36538 23468 36544 23520
rect 36596 23508 36602 23520
rect 38010 23508 38016 23520
rect 36596 23480 36641 23508
rect 37971 23480 38016 23508
rect 36596 23468 36602 23480
rect 38010 23468 38016 23480
rect 38068 23468 38074 23520
rect 38657 23511 38715 23517
rect 38657 23477 38669 23511
rect 38703 23508 38715 23511
rect 39022 23508 39028 23520
rect 38703 23480 39028 23508
rect 38703 23477 38715 23480
rect 38657 23471 38715 23477
rect 39022 23468 39028 23480
rect 39080 23468 39086 23520
rect 39390 23468 39396 23520
rect 39448 23508 39454 23520
rect 39669 23511 39727 23517
rect 39669 23508 39681 23511
rect 39448 23480 39681 23508
rect 39448 23468 39454 23480
rect 39669 23477 39681 23480
rect 39715 23477 39727 23511
rect 39669 23471 39727 23477
rect 41417 23511 41475 23517
rect 41417 23477 41429 23511
rect 41463 23508 41475 23511
rect 41598 23508 41604 23520
rect 41463 23480 41604 23508
rect 41463 23477 41475 23480
rect 41417 23471 41475 23477
rect 41598 23468 41604 23480
rect 41656 23508 41662 23520
rect 41782 23508 41788 23520
rect 41656 23480 41788 23508
rect 41656 23468 41662 23480
rect 41782 23468 41788 23480
rect 41840 23468 41846 23520
rect 1104 23418 58880 23440
rect 1104 23366 10582 23418
rect 10634 23366 10646 23418
rect 10698 23366 10710 23418
rect 10762 23366 10774 23418
rect 10826 23366 10838 23418
rect 10890 23366 29846 23418
rect 29898 23366 29910 23418
rect 29962 23366 29974 23418
rect 30026 23366 30038 23418
rect 30090 23366 30102 23418
rect 30154 23366 49110 23418
rect 49162 23366 49174 23418
rect 49226 23366 49238 23418
rect 49290 23366 49302 23418
rect 49354 23366 49366 23418
rect 49418 23366 58880 23418
rect 1104 23344 58880 23366
rect 2222 23304 2228 23316
rect 2183 23276 2228 23304
rect 2222 23264 2228 23276
rect 2280 23264 2286 23316
rect 19334 23264 19340 23316
rect 19392 23304 19398 23316
rect 20165 23307 20223 23313
rect 20165 23304 20177 23307
rect 19392 23276 20177 23304
rect 19392 23264 19398 23276
rect 20165 23273 20177 23276
rect 20211 23304 20223 23307
rect 21634 23304 21640 23316
rect 20211 23276 21640 23304
rect 20211 23273 20223 23276
rect 20165 23267 20223 23273
rect 21634 23264 21640 23276
rect 21692 23264 21698 23316
rect 22002 23264 22008 23316
rect 22060 23304 22066 23316
rect 26881 23307 26939 23313
rect 26881 23304 26893 23307
rect 22060 23276 26893 23304
rect 22060 23264 22066 23276
rect 26881 23273 26893 23276
rect 26927 23304 26939 23307
rect 26927 23276 27476 23304
rect 26927 23273 26939 23276
rect 26881 23267 26939 23273
rect 19242 23196 19248 23248
rect 19300 23236 19306 23248
rect 19521 23239 19579 23245
rect 19521 23236 19533 23239
rect 19300 23208 19533 23236
rect 19300 23196 19306 23208
rect 19521 23205 19533 23208
rect 19567 23205 19579 23239
rect 19521 23199 19579 23205
rect 23290 23196 23296 23248
rect 23348 23236 23354 23248
rect 23348 23208 24716 23236
rect 23348 23196 23354 23208
rect 22554 23128 22560 23180
rect 22612 23168 22618 23180
rect 24581 23171 24639 23177
rect 24581 23168 24593 23171
rect 22612 23140 24593 23168
rect 22612 23128 22618 23140
rect 24581 23137 24593 23140
rect 24627 23137 24639 23171
rect 24581 23131 24639 23137
rect 24688 23112 24716 23208
rect 24854 23196 24860 23248
rect 24912 23236 24918 23248
rect 26050 23236 26056 23248
rect 24912 23208 26056 23236
rect 24912 23196 24918 23208
rect 26050 23196 26056 23208
rect 26108 23236 26114 23248
rect 27448 23236 27476 23276
rect 27982 23264 27988 23316
rect 28040 23264 28046 23316
rect 28902 23264 28908 23316
rect 28960 23304 28966 23316
rect 28960 23264 28994 23304
rect 29546 23264 29552 23316
rect 29604 23304 29610 23316
rect 30009 23307 30067 23313
rect 29604 23276 29776 23304
rect 29604 23264 29610 23276
rect 28000 23236 28028 23264
rect 26108 23208 26832 23236
rect 27448 23208 28028 23236
rect 28966 23236 28994 23264
rect 29638 23236 29644 23248
rect 28966 23208 29644 23236
rect 26108 23196 26114 23208
rect 24762 23128 24768 23180
rect 24820 23168 24826 23180
rect 25774 23168 25780 23180
rect 24820 23140 25780 23168
rect 24820 23128 24826 23140
rect 25774 23128 25780 23140
rect 25832 23128 25838 23180
rect 26326 23168 26332 23180
rect 26287 23140 26332 23168
rect 26326 23128 26332 23140
rect 26384 23128 26390 23180
rect 1673 23103 1731 23109
rect 1673 23069 1685 23103
rect 1719 23100 1731 23103
rect 2222 23100 2228 23112
rect 1719 23072 2228 23100
rect 1719 23069 1731 23072
rect 1673 23063 1731 23069
rect 2222 23060 2228 23072
rect 2280 23060 2286 23112
rect 21637 23103 21695 23109
rect 21637 23069 21649 23103
rect 21683 23100 21695 23103
rect 24118 23100 24124 23112
rect 21683 23072 24124 23100
rect 21683 23069 21695 23072
rect 21637 23063 21695 23069
rect 24118 23060 24124 23072
rect 24176 23060 24182 23112
rect 24486 23100 24492 23112
rect 24447 23072 24492 23100
rect 24486 23060 24492 23072
rect 24544 23060 24550 23112
rect 24670 23060 24676 23112
rect 24728 23100 24734 23112
rect 25222 23100 25228 23112
rect 24728 23072 24821 23100
rect 25183 23072 25228 23100
rect 24728 23060 24734 23072
rect 25222 23060 25228 23072
rect 25280 23060 25286 23112
rect 26237 23103 26295 23109
rect 26237 23069 26249 23103
rect 26283 23100 26295 23103
rect 26694 23100 26700 23112
rect 26283 23072 26700 23100
rect 26283 23069 26295 23072
rect 26237 23063 26295 23069
rect 26694 23060 26700 23072
rect 26752 23060 26758 23112
rect 26804 23100 26832 23208
rect 29638 23196 29644 23208
rect 29696 23196 29702 23248
rect 29748 23236 29776 23276
rect 30009 23273 30021 23307
rect 30055 23304 30067 23307
rect 30190 23304 30196 23316
rect 30055 23276 30196 23304
rect 30055 23273 30067 23276
rect 30009 23267 30067 23273
rect 30190 23264 30196 23276
rect 30248 23264 30254 23316
rect 31938 23304 31944 23316
rect 30300 23276 31944 23304
rect 30300 23236 30328 23276
rect 31938 23264 31944 23276
rect 31996 23264 32002 23316
rect 32122 23264 32128 23316
rect 32180 23304 32186 23316
rect 34330 23304 34336 23316
rect 32180 23276 34336 23304
rect 32180 23264 32186 23276
rect 34330 23264 34336 23276
rect 34388 23264 34394 23316
rect 34440 23276 40448 23304
rect 29748 23208 30328 23236
rect 31846 23196 31852 23248
rect 31904 23236 31910 23248
rect 32217 23239 32275 23245
rect 32217 23236 32229 23239
rect 31904 23208 32229 23236
rect 31904 23196 31910 23208
rect 32217 23205 32229 23208
rect 32263 23205 32275 23239
rect 32217 23199 32275 23205
rect 34146 23196 34152 23248
rect 34204 23236 34210 23248
rect 34440 23236 34468 23276
rect 38105 23239 38163 23245
rect 38105 23236 38117 23239
rect 34204 23208 34468 23236
rect 34716 23208 38117 23236
rect 34204 23196 34210 23208
rect 27433 23171 27491 23177
rect 27433 23137 27445 23171
rect 27479 23168 27491 23171
rect 27614 23168 27620 23180
rect 27479 23140 27620 23168
rect 27479 23137 27491 23140
rect 27433 23131 27491 23137
rect 27614 23128 27620 23140
rect 27672 23128 27678 23180
rect 28902 23168 28908 23180
rect 28863 23140 28908 23168
rect 28902 23128 28908 23140
rect 28960 23128 28966 23180
rect 29178 23128 29184 23180
rect 29236 23168 29242 23180
rect 31386 23168 31392 23180
rect 29236 23140 31392 23168
rect 29236 23128 29242 23140
rect 31386 23128 31392 23140
rect 31444 23128 31450 23180
rect 31481 23171 31539 23177
rect 31481 23137 31493 23171
rect 31527 23168 31539 23171
rect 34716 23168 34744 23208
rect 38105 23205 38117 23208
rect 38151 23205 38163 23239
rect 40420 23236 40448 23276
rect 40586 23264 40592 23316
rect 40644 23304 40650 23316
rect 40957 23307 41015 23313
rect 40957 23304 40969 23307
rect 40644 23276 40969 23304
rect 40644 23264 40650 23276
rect 40957 23273 40969 23276
rect 41003 23304 41015 23307
rect 42978 23304 42984 23316
rect 41003 23276 42984 23304
rect 41003 23273 41015 23276
rect 40957 23267 41015 23273
rect 42978 23264 42984 23276
rect 43036 23264 43042 23316
rect 41046 23236 41052 23248
rect 40420 23208 41052 23236
rect 38105 23199 38163 23205
rect 41046 23196 41052 23208
rect 41104 23236 41110 23248
rect 41104 23208 41414 23236
rect 41104 23196 41110 23208
rect 31527 23140 34744 23168
rect 34977 23171 35035 23177
rect 31527 23137 31539 23140
rect 31481 23131 31539 23137
rect 34977 23137 34989 23171
rect 35023 23168 35035 23171
rect 35066 23168 35072 23180
rect 35023 23140 35072 23168
rect 35023 23137 35035 23140
rect 34977 23131 35035 23137
rect 35066 23128 35072 23140
rect 35124 23168 35130 23180
rect 35250 23168 35256 23180
rect 35124 23140 35256 23168
rect 35124 23128 35130 23140
rect 35250 23128 35256 23140
rect 35308 23128 35314 23180
rect 35986 23168 35992 23180
rect 35947 23140 35992 23168
rect 35986 23128 35992 23140
rect 36044 23128 36050 23180
rect 36630 23168 36636 23180
rect 36591 23140 36636 23168
rect 36630 23128 36636 23140
rect 36688 23128 36694 23180
rect 38746 23128 38752 23180
rect 38804 23128 38810 23180
rect 27249 23103 27307 23109
rect 26804 23072 27016 23100
rect 23474 22992 23480 23044
rect 23532 23032 23538 23044
rect 25133 23035 25191 23041
rect 25133 23032 25145 23035
rect 23532 23004 25145 23032
rect 23532 22992 23538 23004
rect 25133 23001 25145 23004
rect 25179 23001 25191 23035
rect 25133 22995 25191 23001
rect 25406 22992 25412 23044
rect 25464 23032 25470 23044
rect 25464 23004 26096 23032
rect 25464 22992 25470 23004
rect 1486 22964 1492 22976
rect 1447 22936 1492 22964
rect 1486 22924 1492 22936
rect 1544 22924 1550 22976
rect 20717 22967 20775 22973
rect 20717 22933 20729 22967
rect 20763 22964 20775 22967
rect 20806 22964 20812 22976
rect 20763 22936 20812 22964
rect 20763 22933 20775 22936
rect 20717 22927 20775 22933
rect 20806 22924 20812 22936
rect 20864 22924 20870 22976
rect 22189 22967 22247 22973
rect 22189 22933 22201 22967
rect 22235 22964 22247 22967
rect 22370 22964 22376 22976
rect 22235 22936 22376 22964
rect 22235 22933 22247 22936
rect 22189 22927 22247 22933
rect 22370 22924 22376 22936
rect 22428 22924 22434 22976
rect 22738 22964 22744 22976
rect 22699 22936 22744 22964
rect 22738 22924 22744 22936
rect 22796 22924 22802 22976
rect 23290 22964 23296 22976
rect 23251 22936 23296 22964
rect 23290 22924 23296 22936
rect 23348 22924 23354 22976
rect 23845 22967 23903 22973
rect 23845 22933 23857 22967
rect 23891 22964 23903 22967
rect 23934 22964 23940 22976
rect 23891 22936 23940 22964
rect 23891 22933 23903 22936
rect 23845 22927 23903 22933
rect 23934 22924 23940 22936
rect 23992 22924 23998 22976
rect 24026 22924 24032 22976
rect 24084 22964 24090 22976
rect 25869 22967 25927 22973
rect 25869 22964 25881 22967
rect 24084 22936 25881 22964
rect 24084 22924 24090 22936
rect 25869 22933 25881 22936
rect 25915 22933 25927 22967
rect 26068 22964 26096 23004
rect 26878 22992 26884 23044
rect 26936 22992 26942 23044
rect 26988 23032 27016 23072
rect 27249 23069 27261 23103
rect 27295 23094 27307 23103
rect 27982 23100 27988 23112
rect 27295 23069 27476 23094
rect 27943 23072 27988 23100
rect 27249 23066 27476 23069
rect 27249 23063 27307 23066
rect 27065 23035 27123 23041
rect 27065 23032 27077 23035
rect 26988 23004 27077 23032
rect 27065 23001 27077 23004
rect 27111 23001 27123 23035
rect 27065 22995 27123 23001
rect 26896 22964 26924 22992
rect 27157 22967 27215 22973
rect 27157 22964 27169 22967
rect 26068 22936 27169 22964
rect 25869 22927 25927 22933
rect 27157 22933 27169 22936
rect 27203 22933 27215 22967
rect 27448 22964 27476 23066
rect 27982 23060 27988 23072
rect 28040 23060 28046 23112
rect 28166 23100 28172 23112
rect 28127 23072 28172 23100
rect 28166 23060 28172 23072
rect 28224 23060 28230 23112
rect 29270 23060 29276 23112
rect 29328 23100 29334 23112
rect 29546 23100 29552 23112
rect 29328 23072 29552 23100
rect 29328 23060 29334 23072
rect 29546 23060 29552 23072
rect 29604 23060 29610 23112
rect 31757 23103 31815 23109
rect 31757 23069 31769 23103
rect 31803 23100 31815 23103
rect 33965 23103 34023 23109
rect 31803 23072 32444 23100
rect 31803 23069 31815 23072
rect 31757 23063 31815 23069
rect 27614 22992 27620 23044
rect 27672 23032 27678 23044
rect 30098 23032 30104 23044
rect 27672 23004 30104 23032
rect 27672 22992 27678 23004
rect 30098 22992 30104 23004
rect 30156 22992 30162 23044
rect 30742 22992 30748 23044
rect 30800 22992 30806 23044
rect 28074 22964 28080 22976
rect 27448 22936 28080 22964
rect 27157 22927 27215 22933
rect 28074 22924 28080 22936
rect 28132 22924 28138 22976
rect 28258 22924 28264 22976
rect 28316 22964 28322 22976
rect 32122 22964 32128 22976
rect 28316 22936 32128 22964
rect 28316 22924 28322 22936
rect 32122 22924 32128 22936
rect 32180 22924 32186 22976
rect 32416 22964 32444 23072
rect 33965 23069 33977 23103
rect 34011 23100 34023 23103
rect 34054 23100 34060 23112
rect 34011 23072 34060 23100
rect 34011 23069 34023 23072
rect 33965 23063 34023 23069
rect 34054 23060 34060 23072
rect 34112 23060 34118 23112
rect 34882 23100 34888 23112
rect 34843 23072 34888 23100
rect 34882 23060 34888 23072
rect 34940 23060 34946 23112
rect 37366 23100 37372 23112
rect 37327 23072 37372 23100
rect 37366 23060 37372 23072
rect 37424 23060 37430 23112
rect 37458 23060 37464 23112
rect 37516 23100 37522 23112
rect 37826 23100 37832 23112
rect 37516 23072 37832 23100
rect 37516 23060 37522 23072
rect 37826 23060 37832 23072
rect 37884 23060 37890 23112
rect 38013 23103 38071 23109
rect 38013 23069 38025 23103
rect 38059 23069 38071 23103
rect 38013 23063 38071 23069
rect 38657 23103 38715 23109
rect 38657 23069 38669 23103
rect 38703 23100 38715 23103
rect 38764 23100 38792 23128
rect 38703 23072 38792 23100
rect 38703 23069 38715 23072
rect 38657 23063 38715 23069
rect 33594 23032 33600 23044
rect 33258 23004 33600 23032
rect 33594 22992 33600 23004
rect 33652 22992 33658 23044
rect 33686 22992 33692 23044
rect 33744 23032 33750 23044
rect 33744 23004 33789 23032
rect 33744 22992 33750 23004
rect 34238 22992 34244 23044
rect 34296 23032 34302 23044
rect 36081 23035 36139 23041
rect 36081 23032 36093 23035
rect 34296 23004 36093 23032
rect 34296 22992 34302 23004
rect 36081 23001 36093 23004
rect 36127 23001 36139 23035
rect 36081 22995 36139 23001
rect 37090 22992 37096 23044
rect 37148 23032 37154 23044
rect 38028 23032 38056 23063
rect 37148 23004 38056 23032
rect 37148 22992 37154 23004
rect 38378 22992 38384 23044
rect 38436 23032 38442 23044
rect 38749 23035 38807 23041
rect 38749 23032 38761 23035
rect 38436 23004 38761 23032
rect 38436 22992 38442 23004
rect 38749 23001 38761 23004
rect 38795 23001 38807 23035
rect 38749 22995 38807 23001
rect 41386 22976 41414 23208
rect 34514 22964 34520 22976
rect 32416 22936 34520 22964
rect 34514 22924 34520 22936
rect 34572 22924 34578 22976
rect 34698 22924 34704 22976
rect 34756 22964 34762 22976
rect 34882 22964 34888 22976
rect 34756 22936 34888 22964
rect 34756 22924 34762 22936
rect 34882 22924 34888 22936
rect 34940 22924 34946 22976
rect 35253 22967 35311 22973
rect 35253 22933 35265 22967
rect 35299 22964 35311 22967
rect 36814 22964 36820 22976
rect 35299 22936 36820 22964
rect 35299 22933 35311 22936
rect 35253 22927 35311 22933
rect 36814 22924 36820 22936
rect 36872 22924 36878 22976
rect 37182 22924 37188 22976
rect 37240 22964 37246 22976
rect 37461 22967 37519 22973
rect 37461 22964 37473 22967
rect 37240 22936 37473 22964
rect 37240 22924 37246 22936
rect 37461 22933 37473 22936
rect 37507 22933 37519 22967
rect 37461 22927 37519 22933
rect 38838 22924 38844 22976
rect 38896 22964 38902 22976
rect 39853 22967 39911 22973
rect 39853 22964 39865 22967
rect 38896 22936 39865 22964
rect 38896 22924 38902 22936
rect 39853 22933 39865 22936
rect 39899 22933 39911 22967
rect 40402 22964 40408 22976
rect 40363 22936 40408 22964
rect 39853 22927 39911 22933
rect 40402 22924 40408 22936
rect 40460 22924 40466 22976
rect 41322 22924 41328 22976
rect 41380 22964 41414 22976
rect 41509 22967 41567 22973
rect 41509 22964 41521 22967
rect 41380 22936 41521 22964
rect 41380 22924 41386 22936
rect 41509 22933 41521 22936
rect 41555 22933 41567 22967
rect 41509 22927 41567 22933
rect 42153 22967 42211 22973
rect 42153 22933 42165 22967
rect 42199 22964 42211 22967
rect 42334 22964 42340 22976
rect 42199 22936 42340 22964
rect 42199 22933 42211 22936
rect 42153 22927 42211 22933
rect 42334 22924 42340 22936
rect 42392 22924 42398 22976
rect 42610 22964 42616 22976
rect 42571 22936 42616 22964
rect 42610 22924 42616 22936
rect 42668 22924 42674 22976
rect 1104 22874 58880 22896
rect 1104 22822 20214 22874
rect 20266 22822 20278 22874
rect 20330 22822 20342 22874
rect 20394 22822 20406 22874
rect 20458 22822 20470 22874
rect 20522 22822 39478 22874
rect 39530 22822 39542 22874
rect 39594 22822 39606 22874
rect 39658 22822 39670 22874
rect 39722 22822 39734 22874
rect 39786 22822 58880 22874
rect 1104 22800 58880 22822
rect 17954 22720 17960 22772
rect 18012 22760 18018 22772
rect 18417 22763 18475 22769
rect 18417 22760 18429 22763
rect 18012 22732 18429 22760
rect 18012 22720 18018 22732
rect 18417 22729 18429 22732
rect 18463 22760 18475 22763
rect 19242 22760 19248 22772
rect 18463 22732 19248 22760
rect 18463 22729 18475 22732
rect 18417 22723 18475 22729
rect 19242 22720 19248 22732
rect 19300 22720 19306 22772
rect 20070 22760 20076 22772
rect 20031 22732 20076 22760
rect 20070 22720 20076 22732
rect 20128 22720 20134 22772
rect 21082 22720 21088 22772
rect 21140 22760 21146 22772
rect 21269 22763 21327 22769
rect 21269 22760 21281 22763
rect 21140 22732 21281 22760
rect 21140 22720 21146 22732
rect 21269 22729 21281 22732
rect 21315 22760 21327 22763
rect 21450 22760 21456 22772
rect 21315 22732 21456 22760
rect 21315 22729 21327 22732
rect 21269 22723 21327 22729
rect 21450 22720 21456 22732
rect 21508 22720 21514 22772
rect 23290 22720 23296 22772
rect 23348 22760 23354 22772
rect 25682 22760 25688 22772
rect 23348 22732 25688 22760
rect 23348 22720 23354 22732
rect 25682 22720 25688 22732
rect 25740 22760 25746 22772
rect 27246 22760 27252 22772
rect 25740 22732 27252 22760
rect 25740 22720 25746 22732
rect 27246 22720 27252 22732
rect 27304 22720 27310 22772
rect 27433 22763 27491 22769
rect 27433 22729 27445 22763
rect 27479 22760 27491 22763
rect 27614 22760 27620 22772
rect 27479 22732 27620 22760
rect 27479 22729 27491 22732
rect 27433 22723 27491 22729
rect 27614 22720 27620 22732
rect 27672 22720 27678 22772
rect 27982 22720 27988 22772
rect 28040 22760 28046 22772
rect 30834 22760 30840 22772
rect 28040 22732 28764 22760
rect 28040 22720 28046 22732
rect 19886 22652 19892 22704
rect 19944 22692 19950 22704
rect 20533 22695 20591 22701
rect 20533 22692 20545 22695
rect 19944 22664 20545 22692
rect 19944 22652 19950 22664
rect 20533 22661 20545 22664
rect 20579 22661 20591 22695
rect 20533 22655 20591 22661
rect 24029 22695 24087 22701
rect 24029 22661 24041 22695
rect 24075 22692 24087 22695
rect 24210 22692 24216 22704
rect 24075 22664 24216 22692
rect 24075 22661 24087 22664
rect 24029 22655 24087 22661
rect 24210 22652 24216 22664
rect 24268 22652 24274 22704
rect 25590 22692 25596 22704
rect 25551 22664 25596 22692
rect 25590 22652 25596 22664
rect 25648 22652 25654 22704
rect 25774 22652 25780 22704
rect 25832 22692 25838 22704
rect 26145 22695 26203 22701
rect 26145 22692 26157 22695
rect 25832 22664 26157 22692
rect 25832 22652 25838 22664
rect 26145 22661 26157 22664
rect 26191 22661 26203 22695
rect 26145 22655 26203 22661
rect 26237 22695 26295 22701
rect 26237 22661 26249 22695
rect 26283 22692 26295 22695
rect 26283 22664 26464 22692
rect 26283 22661 26295 22664
rect 26237 22655 26295 22661
rect 26436 22636 26464 22664
rect 26878 22652 26884 22704
rect 26936 22692 26942 22704
rect 26973 22695 27031 22701
rect 26973 22692 26985 22695
rect 26936 22664 26985 22692
rect 26936 22652 26942 22664
rect 26973 22661 26985 22664
rect 27019 22661 27031 22695
rect 27522 22692 27528 22704
rect 26973 22655 27031 22661
rect 27172 22664 27528 22692
rect 27172 22636 27200 22664
rect 27522 22652 27528 22664
rect 27580 22692 27586 22704
rect 27580 22664 28580 22692
rect 27580 22652 27586 22664
rect 23477 22627 23535 22633
rect 23477 22593 23489 22627
rect 23523 22624 23535 22627
rect 23842 22624 23848 22636
rect 23523 22596 23848 22624
rect 23523 22593 23535 22596
rect 23477 22587 23535 22593
rect 23842 22584 23848 22596
rect 23900 22584 23906 22636
rect 23937 22627 23995 22633
rect 23937 22593 23949 22627
rect 23983 22593 23995 22627
rect 24118 22624 24124 22636
rect 24079 22596 24124 22624
rect 23937 22587 23995 22593
rect 19242 22516 19248 22568
rect 19300 22556 19306 22568
rect 19521 22559 19579 22565
rect 19521 22556 19533 22559
rect 19300 22528 19533 22556
rect 19300 22516 19306 22528
rect 19521 22525 19533 22528
rect 19567 22556 19579 22559
rect 22830 22556 22836 22568
rect 19567 22528 22836 22556
rect 19567 22525 19579 22528
rect 19521 22519 19579 22525
rect 22830 22516 22836 22528
rect 22888 22516 22894 22568
rect 23566 22516 23572 22568
rect 23624 22556 23630 22568
rect 23750 22556 23756 22568
rect 23624 22528 23756 22556
rect 23624 22516 23630 22528
rect 23750 22516 23756 22528
rect 23808 22516 23814 22568
rect 23952 22556 23980 22587
rect 24118 22584 24124 22596
rect 24176 22584 24182 22636
rect 24946 22624 24952 22636
rect 24907 22596 24952 22624
rect 24946 22584 24952 22596
rect 25004 22584 25010 22636
rect 26418 22584 26424 22636
rect 26476 22584 26482 22636
rect 27154 22624 27160 22636
rect 27115 22596 27160 22624
rect 27154 22584 27160 22596
rect 27212 22584 27218 22636
rect 27246 22584 27252 22636
rect 27304 22624 27310 22636
rect 28169 22627 28227 22633
rect 28169 22624 28181 22627
rect 27304 22596 27349 22624
rect 27448 22596 28181 22624
rect 27304 22584 27310 22596
rect 24394 22556 24400 22568
rect 23952 22528 24400 22556
rect 24394 22516 24400 22528
rect 24452 22556 24458 22568
rect 25038 22556 25044 22568
rect 24452 22528 24808 22556
rect 24999 22528 25044 22556
rect 24452 22516 24458 22528
rect 21450 22448 21456 22500
rect 21508 22488 21514 22500
rect 24780 22488 24808 22528
rect 25038 22516 25044 22528
rect 25096 22516 25102 22568
rect 25130 22516 25136 22568
rect 25188 22556 25194 22568
rect 25590 22556 25596 22568
rect 25188 22528 25596 22556
rect 25188 22516 25194 22528
rect 25590 22516 25596 22528
rect 25648 22516 25654 22568
rect 27448 22556 27476 22596
rect 28169 22593 28181 22596
rect 28215 22624 28227 22627
rect 28258 22624 28264 22636
rect 28215 22596 28264 22624
rect 28215 22593 28227 22596
rect 28169 22587 28227 22593
rect 28258 22584 28264 22596
rect 28316 22584 28322 22636
rect 25700 22528 27476 22556
rect 25700 22500 25728 22528
rect 27798 22516 27804 22568
rect 27856 22556 27862 22568
rect 27893 22559 27951 22565
rect 27893 22556 27905 22559
rect 27856 22528 27905 22556
rect 27856 22516 27862 22528
rect 27893 22525 27905 22528
rect 27939 22525 27951 22559
rect 28552 22556 28580 22664
rect 28552 22528 28672 22556
rect 27893 22519 27951 22525
rect 25406 22488 25412 22500
rect 21508 22460 24716 22488
rect 24780 22460 25412 22488
rect 21508 22448 21514 22460
rect 18969 22423 19027 22429
rect 18969 22389 18981 22423
rect 19015 22420 19027 22423
rect 19978 22420 19984 22432
rect 19015 22392 19984 22420
rect 19015 22389 19027 22392
rect 18969 22383 19027 22389
rect 19978 22380 19984 22392
rect 20036 22380 20042 22432
rect 22002 22380 22008 22432
rect 22060 22420 22066 22432
rect 22097 22423 22155 22429
rect 22097 22420 22109 22423
rect 22060 22392 22109 22420
rect 22060 22380 22066 22392
rect 22097 22389 22109 22392
rect 22143 22389 22155 22423
rect 22097 22383 22155 22389
rect 22741 22423 22799 22429
rect 22741 22389 22753 22423
rect 22787 22420 22799 22423
rect 22830 22420 22836 22432
rect 22787 22392 22836 22420
rect 22787 22389 22799 22392
rect 22741 22383 22799 22389
rect 22830 22380 22836 22392
rect 22888 22380 22894 22432
rect 23382 22420 23388 22432
rect 23343 22392 23388 22420
rect 23382 22380 23388 22392
rect 23440 22380 23446 22432
rect 24688 22429 24716 22460
rect 25406 22448 25412 22460
rect 25464 22448 25470 22500
rect 25682 22448 25688 22500
rect 25740 22448 25746 22500
rect 25774 22448 25780 22500
rect 25832 22488 25838 22500
rect 28644 22488 28672 22528
rect 28736 22544 28764 22732
rect 28966 22732 30840 22760
rect 28813 22627 28871 22633
rect 28813 22593 28825 22627
rect 28859 22614 28871 22627
rect 28966 22614 28994 22732
rect 30834 22720 30840 22732
rect 30892 22720 30898 22772
rect 32125 22763 32183 22769
rect 32125 22729 32137 22763
rect 32171 22760 32183 22763
rect 32766 22760 32772 22772
rect 32171 22732 32772 22760
rect 32171 22729 32183 22732
rect 32125 22723 32183 22729
rect 32766 22720 32772 22732
rect 32824 22720 32830 22772
rect 32858 22720 32864 22772
rect 32916 22760 32922 22772
rect 37090 22760 37096 22772
rect 32916 22732 37096 22760
rect 32916 22720 32922 22732
rect 37090 22720 37096 22732
rect 37148 22720 37154 22772
rect 37274 22760 37280 22772
rect 37235 22732 37280 22760
rect 37274 22720 37280 22732
rect 37332 22720 37338 22772
rect 37461 22763 37519 22769
rect 37461 22729 37473 22763
rect 37507 22760 37519 22763
rect 39390 22760 39396 22772
rect 37507 22732 39396 22760
rect 37507 22729 37519 22732
rect 37461 22723 37519 22729
rect 39390 22720 39396 22732
rect 39448 22720 39454 22772
rect 41414 22760 41420 22772
rect 41375 22732 41420 22760
rect 41414 22720 41420 22732
rect 41472 22720 41478 22772
rect 42978 22760 42984 22772
rect 42939 22732 42984 22760
rect 42978 22720 42984 22732
rect 43036 22720 43042 22772
rect 29089 22695 29147 22701
rect 29089 22661 29101 22695
rect 29135 22692 29147 22695
rect 29178 22692 29184 22704
rect 29135 22664 29184 22692
rect 29135 22661 29147 22664
rect 29089 22655 29147 22661
rect 29178 22652 29184 22664
rect 29236 22652 29242 22704
rect 30852 22692 30880 22720
rect 30590 22664 30880 22692
rect 32950 22652 32956 22704
rect 33008 22652 33014 22704
rect 33686 22652 33692 22704
rect 33744 22692 33750 22704
rect 38289 22695 38347 22701
rect 38289 22692 38301 22695
rect 33744 22664 38301 22692
rect 33744 22652 33750 22664
rect 38289 22661 38301 22664
rect 38335 22661 38347 22695
rect 40773 22695 40831 22701
rect 40773 22692 40785 22695
rect 38289 22655 38347 22661
rect 39132 22664 40785 22692
rect 28859 22593 28994 22614
rect 28813 22587 28994 22593
rect 35345 22627 35403 22633
rect 35345 22593 35357 22627
rect 35391 22593 35403 22627
rect 35345 22587 35403 22593
rect 35713 22627 35771 22633
rect 35713 22593 35725 22627
rect 35759 22624 35771 22627
rect 35894 22624 35900 22636
rect 35759 22596 35900 22624
rect 35759 22593 35771 22596
rect 35713 22587 35771 22593
rect 28828 22586 28994 22587
rect 31021 22559 31079 22565
rect 31021 22556 31033 22559
rect 28920 22544 31033 22556
rect 28736 22528 31033 22544
rect 28736 22516 28948 22528
rect 31021 22525 31033 22528
rect 31067 22525 31079 22559
rect 31297 22559 31355 22565
rect 31297 22556 31309 22559
rect 31021 22519 31079 22525
rect 31220 22528 31309 22556
rect 25832 22460 28028 22488
rect 28644 22460 29592 22488
rect 25832 22448 25838 22460
rect 28000 22432 28028 22460
rect 24673 22423 24731 22429
rect 24673 22389 24685 22423
rect 24719 22420 24731 22423
rect 26418 22420 26424 22432
rect 24719 22392 26424 22420
rect 24719 22389 24731 22392
rect 24673 22383 24731 22389
rect 26418 22380 26424 22392
rect 26476 22380 26482 22432
rect 26510 22380 26516 22432
rect 26568 22420 26574 22432
rect 26973 22423 27031 22429
rect 26973 22420 26985 22423
rect 26568 22392 26985 22420
rect 26568 22380 26574 22392
rect 26973 22389 26985 22392
rect 27019 22420 27031 22423
rect 27522 22420 27528 22432
rect 27019 22392 27528 22420
rect 27019 22389 27031 22392
rect 26973 22383 27031 22389
rect 27522 22380 27528 22392
rect 27580 22380 27586 22432
rect 27982 22380 27988 22432
rect 28040 22380 28046 22432
rect 28626 22380 28632 22432
rect 28684 22420 28690 22432
rect 29178 22420 29184 22432
rect 28684 22392 29184 22420
rect 28684 22380 28690 22392
rect 29178 22380 29184 22392
rect 29236 22380 29242 22432
rect 29564 22429 29592 22460
rect 31220 22432 31248 22528
rect 31297 22525 31309 22528
rect 31343 22525 31355 22559
rect 31297 22519 31355 22525
rect 31846 22516 31852 22568
rect 31904 22556 31910 22568
rect 32858 22556 32864 22568
rect 31904 22528 32864 22556
rect 31904 22516 31910 22528
rect 32858 22516 32864 22528
rect 32916 22516 32922 22568
rect 33134 22516 33140 22568
rect 33192 22556 33198 22568
rect 33597 22559 33655 22565
rect 33597 22556 33609 22559
rect 33192 22528 33609 22556
rect 33192 22516 33198 22528
rect 33597 22525 33609 22528
rect 33643 22525 33655 22559
rect 33870 22556 33876 22568
rect 33831 22528 33876 22556
rect 33597 22519 33655 22525
rect 33870 22516 33876 22528
rect 33928 22516 33934 22568
rect 34698 22556 34704 22568
rect 34659 22528 34704 22556
rect 34698 22516 34704 22528
rect 34756 22516 34762 22568
rect 31386 22448 31392 22500
rect 31444 22488 31450 22500
rect 32398 22488 32404 22500
rect 31444 22460 32404 22488
rect 31444 22448 31450 22460
rect 32398 22448 32404 22460
rect 32456 22448 32462 22500
rect 35360 22488 35388 22587
rect 35894 22584 35900 22596
rect 35952 22584 35958 22636
rect 36170 22584 36176 22636
rect 36228 22624 36234 22636
rect 36357 22627 36415 22633
rect 36357 22624 36369 22627
rect 36228 22596 36369 22624
rect 36228 22584 36234 22596
rect 36357 22593 36369 22596
rect 36403 22593 36415 22627
rect 36722 22624 36728 22636
rect 36683 22596 36728 22624
rect 36357 22587 36415 22593
rect 36722 22584 36728 22596
rect 36780 22584 36786 22636
rect 37829 22627 37887 22633
rect 37829 22593 37841 22627
rect 37875 22624 37887 22627
rect 38194 22624 38200 22636
rect 37875 22596 38200 22624
rect 37875 22593 37887 22596
rect 37829 22587 37887 22593
rect 38194 22584 38200 22596
rect 38252 22584 38258 22636
rect 38562 22624 38568 22636
rect 38523 22596 38568 22624
rect 38562 22584 38568 22596
rect 38620 22584 38626 22636
rect 36814 22516 36820 22568
rect 36872 22556 36878 22568
rect 36872 22528 38056 22556
rect 36872 22516 36878 22528
rect 33796 22460 35388 22488
rect 36449 22491 36507 22497
rect 29549 22423 29607 22429
rect 29549 22389 29561 22423
rect 29595 22389 29607 22423
rect 29549 22383 29607 22389
rect 30466 22380 30472 22432
rect 30524 22420 30530 22432
rect 31202 22420 31208 22432
rect 30524 22392 31208 22420
rect 30524 22380 30530 22392
rect 31202 22380 31208 22392
rect 31260 22380 31266 22432
rect 31570 22380 31576 22432
rect 31628 22420 31634 22432
rect 33796 22420 33824 22460
rect 36449 22457 36461 22491
rect 36495 22488 36507 22491
rect 36998 22488 37004 22500
rect 36495 22460 37004 22488
rect 36495 22457 36507 22460
rect 36449 22451 36507 22457
rect 36998 22448 37004 22460
rect 37056 22448 37062 22500
rect 38028 22488 38056 22528
rect 38102 22516 38108 22568
rect 38160 22556 38166 22568
rect 39132 22556 39160 22664
rect 40773 22661 40785 22664
rect 40819 22692 40831 22695
rect 43898 22692 43904 22704
rect 40819 22664 43904 22692
rect 40819 22661 40831 22664
rect 40773 22655 40831 22661
rect 43898 22652 43904 22664
rect 43956 22652 43962 22704
rect 39209 22627 39267 22633
rect 39209 22593 39221 22627
rect 39255 22624 39267 22627
rect 41230 22624 41236 22636
rect 39255 22596 41236 22624
rect 39255 22593 39267 22596
rect 39209 22587 39267 22593
rect 41230 22584 41236 22596
rect 41288 22584 41294 22636
rect 45462 22556 45468 22568
rect 38160 22528 39160 22556
rect 39684 22528 45468 22556
rect 38160 22516 38166 22528
rect 38194 22488 38200 22500
rect 38028 22460 38200 22488
rect 38194 22448 38200 22460
rect 38252 22448 38258 22500
rect 39117 22491 39175 22497
rect 39117 22457 39129 22491
rect 39163 22488 39175 22491
rect 39574 22488 39580 22500
rect 39163 22460 39580 22488
rect 39163 22457 39175 22460
rect 39117 22451 39175 22457
rect 39574 22448 39580 22460
rect 39632 22448 39638 22500
rect 31628 22392 33824 22420
rect 31628 22380 31634 22392
rect 35986 22380 35992 22432
rect 36044 22420 36050 22432
rect 36541 22423 36599 22429
rect 36541 22420 36553 22423
rect 36044 22392 36553 22420
rect 36044 22380 36050 22392
rect 36541 22389 36553 22392
rect 36587 22389 36599 22423
rect 36722 22420 36728 22432
rect 36683 22392 36728 22420
rect 36541 22383 36599 22389
rect 36722 22380 36728 22392
rect 36780 22380 36786 22432
rect 37461 22423 37519 22429
rect 37461 22389 37473 22423
rect 37507 22420 37519 22423
rect 37550 22420 37556 22432
rect 37507 22392 37556 22420
rect 37507 22389 37519 22392
rect 37461 22383 37519 22389
rect 37550 22380 37556 22392
rect 37608 22380 37614 22432
rect 37642 22380 37648 22432
rect 37700 22420 37706 22432
rect 37918 22420 37924 22432
rect 37700 22392 37924 22420
rect 37700 22380 37706 22392
rect 37918 22380 37924 22392
rect 37976 22380 37982 22432
rect 38746 22380 38752 22432
rect 38804 22420 38810 22432
rect 39684 22429 39712 22528
rect 45462 22516 45468 22528
rect 45520 22516 45526 22568
rect 42794 22448 42800 22500
rect 42852 22488 42858 22500
rect 43530 22488 43536 22500
rect 42852 22460 43536 22488
rect 42852 22448 42858 22460
rect 43530 22448 43536 22460
rect 43588 22448 43594 22500
rect 39669 22423 39727 22429
rect 39669 22420 39681 22423
rect 38804 22392 39681 22420
rect 38804 22380 38810 22392
rect 39669 22389 39681 22392
rect 39715 22389 39727 22423
rect 39669 22383 39727 22389
rect 39850 22380 39856 22432
rect 39908 22420 39914 22432
rect 40221 22423 40279 22429
rect 40221 22420 40233 22423
rect 39908 22392 40233 22420
rect 39908 22380 39914 22392
rect 40221 22389 40233 22392
rect 40267 22389 40279 22423
rect 40221 22383 40279 22389
rect 41322 22380 41328 22432
rect 41380 22420 41386 22432
rect 42521 22423 42579 22429
rect 42521 22420 42533 22423
rect 41380 22392 42533 22420
rect 41380 22380 41386 22392
rect 42521 22389 42533 22392
rect 42567 22420 42579 22423
rect 45370 22420 45376 22432
rect 42567 22392 45376 22420
rect 42567 22389 42579 22392
rect 42521 22383 42579 22389
rect 45370 22380 45376 22392
rect 45428 22380 45434 22432
rect 1104 22330 58880 22352
rect 1104 22278 10582 22330
rect 10634 22278 10646 22330
rect 10698 22278 10710 22330
rect 10762 22278 10774 22330
rect 10826 22278 10838 22330
rect 10890 22278 29846 22330
rect 29898 22278 29910 22330
rect 29962 22278 29974 22330
rect 30026 22278 30038 22330
rect 30090 22278 30102 22330
rect 30154 22278 49110 22330
rect 49162 22278 49174 22330
rect 49226 22278 49238 22330
rect 49290 22278 49302 22330
rect 49354 22278 49366 22330
rect 49418 22278 58880 22330
rect 1104 22256 58880 22278
rect 20714 22176 20720 22228
rect 20772 22216 20778 22228
rect 22738 22216 22744 22228
rect 20772 22188 22744 22216
rect 20772 22176 20778 22188
rect 22738 22176 22744 22188
rect 22796 22216 22802 22228
rect 23566 22216 23572 22228
rect 22796 22188 23572 22216
rect 22796 22176 22802 22188
rect 23566 22176 23572 22188
rect 23624 22176 23630 22228
rect 24118 22176 24124 22228
rect 24176 22216 24182 22228
rect 26234 22216 26240 22228
rect 24176 22188 26240 22216
rect 24176 22176 24182 22188
rect 26234 22176 26240 22188
rect 26292 22176 26298 22228
rect 26510 22176 26516 22228
rect 26568 22216 26574 22228
rect 26970 22216 26976 22228
rect 26568 22188 26976 22216
rect 26568 22176 26574 22188
rect 26970 22176 26976 22188
rect 27028 22176 27034 22228
rect 27512 22219 27570 22225
rect 27512 22185 27524 22219
rect 27558 22216 27570 22219
rect 27890 22216 27896 22228
rect 27558 22188 27896 22216
rect 27558 22185 27570 22188
rect 27512 22179 27570 22185
rect 27890 22176 27896 22188
rect 27948 22176 27954 22228
rect 28258 22176 28264 22228
rect 28316 22216 28322 22228
rect 29730 22216 29736 22228
rect 28316 22188 29736 22216
rect 28316 22176 28322 22188
rect 29730 22176 29736 22188
rect 29788 22176 29794 22228
rect 31481 22219 31539 22225
rect 31481 22185 31493 22219
rect 31527 22216 31539 22219
rect 31570 22216 31576 22228
rect 31527 22188 31576 22216
rect 31527 22185 31539 22188
rect 31481 22179 31539 22185
rect 31570 22176 31576 22188
rect 31628 22176 31634 22228
rect 33870 22216 33876 22228
rect 31726 22188 33876 22216
rect 19518 22108 19524 22160
rect 19576 22148 19582 22160
rect 23845 22151 23903 22157
rect 23845 22148 23857 22151
rect 19576 22120 23857 22148
rect 19576 22108 19582 22120
rect 23845 22117 23857 22120
rect 23891 22148 23903 22151
rect 25498 22148 25504 22160
rect 23891 22120 25504 22148
rect 23891 22117 23903 22120
rect 23845 22111 23903 22117
rect 25498 22108 25504 22120
rect 25556 22108 25562 22160
rect 25593 22151 25651 22157
rect 25593 22117 25605 22151
rect 25639 22148 25651 22151
rect 25774 22148 25780 22160
rect 25639 22120 25780 22148
rect 25639 22117 25651 22120
rect 25593 22111 25651 22117
rect 25774 22108 25780 22120
rect 25832 22108 25838 22160
rect 26602 22148 26608 22160
rect 26160 22120 26608 22148
rect 18693 22083 18751 22089
rect 18693 22049 18705 22083
rect 18739 22080 18751 22083
rect 19334 22080 19340 22092
rect 18739 22052 19340 22080
rect 18739 22049 18751 22052
rect 18693 22043 18751 22049
rect 19334 22040 19340 22052
rect 19392 22040 19398 22092
rect 23017 22083 23075 22089
rect 23017 22049 23029 22083
rect 23063 22080 23075 22083
rect 23198 22080 23204 22092
rect 23063 22052 23204 22080
rect 23063 22049 23075 22052
rect 23017 22043 23075 22049
rect 23198 22040 23204 22052
rect 23256 22040 23262 22092
rect 24210 22040 24216 22092
rect 24268 22080 24274 22092
rect 24486 22080 24492 22092
rect 24268 22052 24492 22080
rect 24268 22040 24274 22052
rect 24486 22040 24492 22052
rect 24544 22040 24550 22092
rect 25314 22080 25320 22092
rect 25275 22052 25320 22080
rect 25314 22040 25320 22052
rect 25372 22040 25378 22092
rect 22094 21972 22100 22024
rect 22152 22012 22158 22024
rect 22281 22015 22339 22021
rect 22281 22012 22293 22015
rect 22152 21984 22293 22012
rect 22152 21972 22158 21984
rect 22281 21981 22293 21984
rect 22327 21981 22339 22015
rect 22281 21975 22339 21981
rect 22738 21972 22744 22024
rect 22796 22012 22802 22024
rect 22922 22012 22928 22024
rect 22796 21984 22928 22012
rect 22796 21972 22802 21984
rect 22922 21972 22928 21984
rect 22980 21972 22986 22024
rect 23106 22012 23112 22024
rect 23067 21984 23112 22012
rect 23106 21972 23112 21984
rect 23164 21972 23170 22024
rect 23934 21972 23940 22024
rect 23992 22012 23998 22024
rect 24397 22015 24455 22021
rect 24397 22012 24409 22015
rect 23992 21984 24409 22012
rect 23992 21972 23998 21984
rect 24397 21981 24409 21984
rect 24443 21981 24455 22015
rect 25222 22012 25228 22024
rect 25183 21984 25228 22012
rect 24397 21975 24455 21981
rect 25222 21972 25228 21984
rect 25280 22012 25286 22024
rect 26160 22012 26188 22120
rect 26602 22108 26608 22120
rect 26660 22148 26666 22160
rect 27154 22148 27160 22160
rect 26660 22120 27160 22148
rect 26660 22108 26666 22120
rect 27154 22108 27160 22120
rect 27212 22108 27218 22160
rect 31202 22108 31208 22160
rect 31260 22148 31266 22160
rect 31726 22148 31754 22188
rect 33870 22176 33876 22188
rect 33928 22176 33934 22228
rect 35066 22176 35072 22228
rect 35124 22216 35130 22228
rect 35894 22216 35900 22228
rect 35124 22188 35900 22216
rect 35124 22176 35130 22188
rect 35894 22176 35900 22188
rect 35952 22176 35958 22228
rect 36170 22176 36176 22228
rect 36228 22216 36234 22228
rect 36630 22216 36636 22228
rect 36228 22188 36636 22216
rect 36228 22176 36234 22188
rect 36630 22176 36636 22188
rect 36688 22176 36694 22228
rect 42610 22216 42616 22228
rect 36924 22188 42616 22216
rect 31260 22120 31754 22148
rect 31260 22108 31266 22120
rect 34514 22108 34520 22160
rect 34572 22148 34578 22160
rect 36924 22148 36952 22188
rect 42610 22176 42616 22188
rect 42668 22176 42674 22228
rect 42978 22176 42984 22228
rect 43036 22216 43042 22228
rect 43257 22219 43315 22225
rect 43257 22216 43269 22219
rect 43036 22188 43269 22216
rect 43036 22176 43042 22188
rect 43257 22185 43269 22188
rect 43303 22216 43315 22219
rect 43809 22219 43867 22225
rect 43809 22216 43821 22219
rect 43303 22188 43821 22216
rect 43303 22185 43315 22188
rect 43257 22179 43315 22185
rect 43809 22185 43821 22188
rect 43855 22185 43867 22219
rect 43809 22179 43867 22185
rect 38562 22148 38568 22160
rect 34572 22120 36952 22148
rect 38523 22120 38568 22148
rect 34572 22108 34578 22120
rect 38562 22108 38568 22120
rect 38620 22108 38626 22160
rect 39298 22148 39304 22160
rect 38672 22120 39304 22148
rect 26234 22040 26240 22092
rect 26292 22080 26298 22092
rect 26292 22052 26337 22080
rect 26292 22040 26298 22052
rect 27522 22040 27528 22092
rect 27580 22080 27586 22092
rect 29178 22080 29184 22092
rect 27580 22052 29184 22080
rect 27580 22040 27586 22052
rect 29178 22040 29184 22052
rect 29236 22040 29242 22092
rect 29546 22040 29552 22092
rect 29604 22080 29610 22092
rect 30009 22083 30067 22089
rect 30009 22080 30021 22083
rect 29604 22052 30021 22080
rect 29604 22040 29610 22052
rect 30009 22049 30021 22052
rect 30055 22049 30067 22083
rect 30009 22043 30067 22049
rect 30374 22040 30380 22092
rect 30432 22080 30438 22092
rect 36078 22080 36084 22092
rect 30432 22052 36084 22080
rect 30432 22040 30438 22052
rect 36078 22040 36084 22052
rect 36136 22040 36142 22092
rect 36446 22040 36452 22092
rect 36504 22080 36510 22092
rect 37645 22083 37703 22089
rect 37645 22080 37657 22083
rect 36504 22052 37657 22080
rect 36504 22040 36510 22052
rect 37645 22049 37657 22052
rect 37691 22049 37703 22083
rect 38102 22080 38108 22092
rect 37645 22043 37703 22049
rect 37752 22052 38108 22080
rect 25280 21984 26188 22012
rect 25280 21972 25286 21984
rect 26326 21972 26332 22024
rect 26384 22012 26390 22024
rect 26421 22015 26479 22021
rect 26421 22012 26433 22015
rect 26384 21984 26433 22012
rect 26384 21972 26390 21984
rect 26421 21981 26433 21984
rect 26467 21981 26479 22015
rect 26421 21975 26479 21981
rect 26602 21972 26608 22024
rect 26660 22012 26666 22024
rect 27249 22015 27307 22021
rect 27249 22012 27261 22015
rect 26660 21984 27261 22012
rect 26660 21972 26666 21984
rect 27249 21981 27261 21984
rect 27295 21981 27307 22015
rect 27249 21975 27307 21981
rect 28902 21972 28908 22024
rect 28960 22012 28966 22024
rect 29733 22015 29791 22021
rect 29733 22012 29745 22015
rect 28960 21984 29745 22012
rect 28960 21972 28966 21984
rect 29733 21981 29745 21984
rect 29779 21981 29791 22015
rect 29733 21975 29791 21981
rect 32306 21972 32312 22024
rect 32364 21972 32370 22024
rect 33686 21972 33692 22024
rect 33744 22012 33750 22024
rect 33744 21984 33789 22012
rect 33744 21972 33750 21984
rect 34330 21972 34336 22024
rect 34388 22012 34394 22024
rect 37366 22012 37372 22024
rect 34388 21984 37372 22012
rect 34388 21972 34394 21984
rect 37366 21972 37372 21984
rect 37424 21972 37430 22024
rect 37550 21972 37556 22024
rect 37608 22012 37614 22024
rect 37752 22021 37780 22052
rect 38102 22040 38108 22052
rect 38160 22040 38166 22092
rect 38470 22080 38476 22092
rect 38431 22052 38476 22080
rect 38470 22040 38476 22052
rect 38528 22040 38534 22092
rect 38672 22089 38700 22120
rect 39298 22108 39304 22120
rect 39356 22148 39362 22160
rect 39850 22148 39856 22160
rect 39356 22120 39856 22148
rect 39356 22108 39362 22120
rect 39850 22108 39856 22120
rect 39908 22108 39914 22160
rect 39945 22151 40003 22157
rect 39945 22117 39957 22151
rect 39991 22148 40003 22151
rect 40034 22148 40040 22160
rect 39991 22120 40040 22148
rect 39991 22117 40003 22120
rect 39945 22111 40003 22117
rect 40034 22108 40040 22120
rect 40092 22108 40098 22160
rect 40218 22108 40224 22160
rect 40276 22148 40282 22160
rect 41049 22151 41107 22157
rect 41049 22148 41061 22151
rect 40276 22120 41061 22148
rect 40276 22108 40282 22120
rect 41049 22117 41061 22120
rect 41095 22117 41107 22151
rect 41049 22111 41107 22117
rect 38657 22083 38715 22089
rect 38657 22049 38669 22083
rect 38703 22080 38715 22083
rect 41690 22080 41696 22092
rect 38703 22052 38805 22080
rect 39316 22052 41696 22080
rect 38703 22049 38715 22052
rect 38657 22043 38715 22049
rect 37737 22015 37795 22021
rect 37737 22012 37749 22015
rect 37608 21984 37749 22012
rect 37608 21972 37614 21984
rect 37737 21981 37749 21984
rect 37783 21981 37795 22015
rect 37737 21975 37795 21981
rect 37918 21972 37924 22024
rect 37976 22012 37982 22024
rect 38381 22015 38439 22021
rect 38381 22012 38393 22015
rect 37976 21984 38393 22012
rect 37976 21972 37982 21984
rect 38381 21981 38393 21984
rect 38427 21981 38439 22015
rect 38381 21975 38439 21981
rect 20533 21947 20591 21953
rect 20533 21913 20545 21947
rect 20579 21944 20591 21947
rect 21174 21944 21180 21956
rect 20579 21916 21180 21944
rect 20579 21913 20591 21916
rect 20533 21907 20591 21913
rect 21174 21904 21180 21916
rect 21232 21904 21238 21956
rect 23290 21944 23296 21956
rect 21560 21916 23296 21944
rect 15010 21836 15016 21888
rect 15068 21876 15074 21888
rect 17497 21879 17555 21885
rect 17497 21876 17509 21879
rect 15068 21848 17509 21876
rect 15068 21836 15074 21848
rect 17497 21845 17509 21848
rect 17543 21876 17555 21879
rect 18046 21876 18052 21888
rect 17543 21848 18052 21876
rect 17543 21845 17555 21848
rect 17497 21839 17555 21845
rect 18046 21836 18052 21848
rect 18104 21836 18110 21888
rect 19426 21876 19432 21888
rect 19387 21848 19432 21876
rect 19426 21836 19432 21848
rect 19484 21836 19490 21888
rect 19981 21879 20039 21885
rect 19981 21845 19993 21879
rect 20027 21876 20039 21879
rect 20070 21876 20076 21888
rect 20027 21848 20076 21876
rect 20027 21845 20039 21848
rect 19981 21839 20039 21845
rect 20070 21836 20076 21848
rect 20128 21836 20134 21888
rect 20898 21836 20904 21888
rect 20956 21876 20962 21888
rect 20993 21879 21051 21885
rect 20993 21876 21005 21879
rect 20956 21848 21005 21876
rect 20956 21836 20962 21848
rect 20993 21845 21005 21848
rect 21039 21845 21051 21879
rect 20993 21839 21051 21845
rect 21266 21836 21272 21888
rect 21324 21876 21330 21888
rect 21560 21885 21588 21916
rect 23290 21904 23296 21916
rect 23348 21944 23354 21956
rect 23661 21947 23719 21953
rect 23661 21944 23673 21947
rect 23348 21916 23673 21944
rect 23348 21904 23354 21916
rect 23661 21913 23673 21916
rect 23707 21913 23719 21947
rect 23661 21907 23719 21913
rect 24489 21947 24547 21953
rect 24489 21913 24501 21947
rect 24535 21944 24547 21947
rect 24535 21916 27936 21944
rect 24535 21913 24547 21916
rect 24489 21907 24547 21913
rect 21545 21879 21603 21885
rect 21545 21876 21557 21879
rect 21324 21848 21557 21876
rect 21324 21836 21330 21848
rect 21545 21845 21557 21848
rect 21591 21845 21603 21879
rect 21545 21839 21603 21845
rect 22097 21879 22155 21885
rect 22097 21845 22109 21879
rect 22143 21876 22155 21879
rect 22186 21876 22192 21888
rect 22143 21848 22192 21876
rect 22143 21845 22155 21848
rect 22097 21839 22155 21845
rect 22186 21836 22192 21848
rect 22244 21836 22250 21888
rect 22370 21836 22376 21888
rect 22428 21876 22434 21888
rect 25406 21876 25412 21888
rect 22428 21848 25412 21876
rect 22428 21836 22434 21848
rect 25406 21836 25412 21848
rect 25464 21876 25470 21888
rect 26050 21876 26056 21888
rect 25464 21848 26056 21876
rect 25464 21836 25470 21848
rect 26050 21836 26056 21848
rect 26108 21836 26114 21888
rect 26326 21876 26332 21888
rect 26239 21848 26332 21876
rect 26326 21836 26332 21848
rect 26384 21876 26390 21888
rect 26510 21876 26516 21888
rect 26384 21848 26516 21876
rect 26384 21836 26390 21848
rect 26510 21836 26516 21848
rect 26568 21836 26574 21888
rect 26789 21879 26847 21885
rect 26789 21845 26801 21879
rect 26835 21876 26847 21879
rect 26878 21876 26884 21888
rect 26835 21848 26884 21876
rect 26835 21845 26847 21848
rect 26789 21839 26847 21845
rect 26878 21836 26884 21848
rect 26936 21836 26942 21888
rect 27908 21876 27936 21916
rect 28166 21904 28172 21956
rect 28224 21904 28230 21956
rect 33413 21947 33471 21953
rect 28828 21916 30498 21944
rect 28828 21876 28856 21916
rect 33413 21913 33425 21947
rect 33459 21944 33471 21947
rect 33502 21944 33508 21956
rect 33459 21916 33508 21944
rect 33459 21913 33471 21916
rect 33413 21907 33471 21913
rect 33502 21904 33508 21916
rect 33560 21904 33566 21956
rect 33962 21904 33968 21956
rect 34020 21944 34026 21956
rect 36078 21944 36084 21956
rect 34020 21916 36084 21944
rect 34020 21904 34026 21916
rect 36078 21904 36084 21916
rect 36136 21904 36142 21956
rect 36909 21947 36967 21953
rect 36909 21913 36921 21947
rect 36955 21944 36967 21947
rect 36955 21916 37228 21944
rect 36955 21913 36967 21916
rect 36909 21907 36967 21913
rect 37200 21888 37228 21916
rect 37826 21904 37832 21956
rect 37884 21944 37890 21956
rect 38672 21944 38700 22043
rect 39114 22012 39120 22024
rect 39075 21984 39120 22012
rect 39114 21972 39120 21984
rect 39172 21972 39178 22024
rect 39316 22021 39344 22052
rect 41690 22040 41696 22052
rect 41748 22040 41754 22092
rect 43824 22080 43852 22179
rect 43898 22108 43904 22160
rect 43956 22148 43962 22160
rect 48682 22148 48688 22160
rect 43956 22120 48688 22148
rect 43956 22108 43962 22120
rect 48682 22108 48688 22120
rect 48740 22108 48746 22160
rect 44082 22080 44088 22092
rect 43824 22052 44088 22080
rect 44082 22040 44088 22052
rect 44140 22080 44146 22092
rect 44361 22083 44419 22089
rect 44361 22080 44373 22083
rect 44140 22052 44373 22080
rect 44140 22040 44146 22052
rect 44361 22049 44373 22052
rect 44407 22049 44419 22083
rect 44361 22043 44419 22049
rect 39301 22015 39359 22021
rect 39301 21981 39313 22015
rect 39347 21981 39359 22015
rect 39301 21975 39359 21981
rect 39853 22015 39911 22021
rect 39853 21981 39865 22015
rect 39899 22012 39911 22015
rect 40126 22012 40132 22024
rect 39899 21984 40132 22012
rect 39899 21981 39911 21984
rect 39853 21975 39911 21981
rect 40126 21972 40132 21984
rect 40184 21972 40190 22024
rect 58158 22012 58164 22024
rect 58119 21984 58164 22012
rect 58158 21972 58164 21984
rect 58216 21972 58222 22024
rect 37884 21916 38700 21944
rect 37884 21904 37890 21916
rect 41138 21904 41144 21956
rect 41196 21944 41202 21956
rect 41601 21947 41659 21953
rect 41601 21944 41613 21947
rect 41196 21916 41613 21944
rect 41196 21904 41202 21916
rect 41601 21913 41613 21916
rect 41647 21913 41659 21947
rect 41601 21907 41659 21913
rect 47854 21904 47860 21956
rect 47912 21944 47918 21956
rect 57885 21947 57943 21953
rect 57885 21944 57897 21947
rect 47912 21916 57897 21944
rect 47912 21904 47918 21916
rect 57885 21913 57897 21916
rect 57931 21913 57943 21947
rect 57885 21907 57943 21913
rect 27908 21848 28856 21876
rect 28997 21879 29055 21885
rect 28997 21845 29009 21879
rect 29043 21876 29055 21879
rect 29546 21876 29552 21888
rect 29043 21848 29552 21876
rect 29043 21845 29055 21848
rect 28997 21839 29055 21845
rect 29546 21836 29552 21848
rect 29604 21836 29610 21888
rect 31938 21876 31944 21888
rect 31899 21848 31944 21876
rect 31938 21836 31944 21848
rect 31996 21836 32002 21888
rect 32674 21836 32680 21888
rect 32732 21876 32738 21888
rect 33134 21876 33140 21888
rect 32732 21848 33140 21876
rect 32732 21836 32738 21848
rect 33134 21836 33140 21848
rect 33192 21836 33198 21888
rect 35158 21836 35164 21888
rect 35216 21876 35222 21888
rect 35621 21879 35679 21885
rect 35621 21876 35633 21879
rect 35216 21848 35633 21876
rect 35216 21836 35222 21848
rect 35621 21845 35633 21848
rect 35667 21876 35679 21879
rect 36998 21876 37004 21888
rect 35667 21848 37004 21876
rect 35667 21845 35679 21848
rect 35621 21839 35679 21845
rect 36998 21836 37004 21848
rect 37056 21836 37062 21888
rect 37182 21836 37188 21888
rect 37240 21836 37246 21888
rect 37274 21836 37280 21888
rect 37332 21876 37338 21888
rect 37369 21879 37427 21885
rect 37369 21876 37381 21879
rect 37332 21848 37381 21876
rect 37332 21836 37338 21848
rect 37369 21845 37381 21848
rect 37415 21845 37427 21879
rect 37369 21839 37427 21845
rect 39209 21879 39267 21885
rect 39209 21845 39221 21879
rect 39255 21876 39267 21879
rect 39298 21876 39304 21888
rect 39255 21848 39304 21876
rect 39255 21845 39267 21848
rect 39209 21839 39267 21845
rect 39298 21836 39304 21848
rect 39356 21836 39362 21888
rect 40402 21836 40408 21888
rect 40460 21876 40466 21888
rect 40497 21879 40555 21885
rect 40497 21876 40509 21879
rect 40460 21848 40509 21876
rect 40460 21836 40466 21848
rect 40497 21845 40509 21848
rect 40543 21845 40555 21879
rect 40497 21839 40555 21845
rect 41322 21836 41328 21888
rect 41380 21876 41386 21888
rect 42058 21876 42064 21888
rect 41380 21848 42064 21876
rect 41380 21836 41386 21848
rect 42058 21836 42064 21848
rect 42116 21876 42122 21888
rect 42245 21879 42303 21885
rect 42245 21876 42257 21879
rect 42116 21848 42257 21876
rect 42116 21836 42122 21848
rect 42245 21845 42257 21848
rect 42291 21876 42303 21879
rect 42426 21876 42432 21888
rect 42291 21848 42432 21876
rect 42291 21845 42303 21848
rect 42245 21839 42303 21845
rect 42426 21836 42432 21848
rect 42484 21836 42490 21888
rect 42702 21836 42708 21888
rect 42760 21876 42766 21888
rect 42797 21879 42855 21885
rect 42797 21876 42809 21879
rect 42760 21848 42809 21876
rect 42760 21836 42766 21848
rect 42797 21845 42809 21848
rect 42843 21876 42855 21879
rect 43254 21876 43260 21888
rect 42843 21848 43260 21876
rect 42843 21845 42855 21848
rect 42797 21839 42855 21845
rect 43254 21836 43260 21848
rect 43312 21836 43318 21888
rect 1104 21786 58880 21808
rect 1104 21734 20214 21786
rect 20266 21734 20278 21786
rect 20330 21734 20342 21786
rect 20394 21734 20406 21786
rect 20458 21734 20470 21786
rect 20522 21734 39478 21786
rect 39530 21734 39542 21786
rect 39594 21734 39606 21786
rect 39658 21734 39670 21786
rect 39722 21734 39734 21786
rect 39786 21734 58880 21786
rect 1104 21712 58880 21734
rect 16114 21632 16120 21684
rect 16172 21672 16178 21684
rect 17681 21675 17739 21681
rect 17681 21672 17693 21675
rect 16172 21644 17693 21672
rect 16172 21632 16178 21644
rect 17681 21641 17693 21644
rect 17727 21672 17739 21675
rect 19334 21672 19340 21684
rect 17727 21644 19340 21672
rect 17727 21641 17739 21644
rect 17681 21635 17739 21641
rect 19334 21632 19340 21644
rect 19392 21632 19398 21684
rect 20714 21672 20720 21684
rect 20675 21644 20720 21672
rect 20714 21632 20720 21644
rect 20772 21632 20778 21684
rect 21174 21632 21180 21684
rect 21232 21672 21238 21684
rect 26326 21672 26332 21684
rect 21232 21644 26332 21672
rect 21232 21632 21238 21644
rect 26326 21632 26332 21644
rect 26384 21632 26390 21684
rect 27614 21632 27620 21684
rect 27672 21672 27678 21684
rect 27798 21672 27804 21684
rect 27672 21644 27804 21672
rect 27672 21632 27678 21644
rect 27798 21632 27804 21644
rect 27856 21632 27862 21684
rect 27890 21632 27896 21684
rect 27948 21672 27954 21684
rect 29546 21672 29552 21684
rect 27948 21644 29552 21672
rect 27948 21632 27954 21644
rect 29546 21632 29552 21644
rect 29604 21632 29610 21684
rect 30190 21632 30196 21684
rect 30248 21672 30254 21684
rect 30466 21672 30472 21684
rect 30248 21644 30472 21672
rect 30248 21632 30254 21644
rect 30466 21632 30472 21644
rect 30524 21632 30530 21684
rect 30834 21632 30840 21684
rect 30892 21672 30898 21684
rect 30892 21644 31432 21672
rect 30892 21632 30898 21644
rect 15746 21564 15752 21616
rect 15804 21604 15810 21616
rect 17129 21607 17187 21613
rect 17129 21604 17141 21607
rect 15804 21576 17141 21604
rect 15804 21564 15810 21576
rect 17129 21573 17141 21576
rect 17175 21604 17187 21607
rect 19610 21604 19616 21616
rect 17175 21576 19616 21604
rect 17175 21573 17187 21576
rect 17129 21567 17187 21573
rect 19610 21564 19616 21576
rect 19668 21604 19674 21616
rect 19978 21604 19984 21616
rect 19668 21576 19984 21604
rect 19668 21564 19674 21576
rect 19978 21564 19984 21576
rect 20036 21564 20042 21616
rect 20622 21564 20628 21616
rect 20680 21604 20686 21616
rect 21192 21604 21220 21632
rect 22830 21604 22836 21616
rect 20680 21576 21220 21604
rect 22791 21576 22836 21604
rect 20680 21564 20686 21576
rect 22830 21564 22836 21576
rect 22888 21564 22894 21616
rect 22922 21564 22928 21616
rect 22980 21604 22986 21616
rect 23198 21604 23204 21616
rect 22980 21576 23204 21604
rect 22980 21564 22986 21576
rect 23198 21564 23204 21576
rect 23256 21604 23262 21616
rect 24118 21604 24124 21616
rect 23256 21576 24124 21604
rect 23256 21564 23262 21576
rect 24118 21564 24124 21576
rect 24176 21564 24182 21616
rect 24578 21604 24584 21616
rect 24320 21576 24584 21604
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 12250 21536 12256 21548
rect 1719 21508 12256 21536
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 12250 21496 12256 21508
rect 12308 21496 12314 21548
rect 17862 21496 17868 21548
rect 17920 21536 17926 21548
rect 17920 21508 22094 21536
rect 17920 21496 17926 21508
rect 18233 21471 18291 21477
rect 18233 21437 18245 21471
rect 18279 21468 18291 21471
rect 18322 21468 18328 21480
rect 18279 21440 18328 21468
rect 18279 21437 18291 21440
rect 18233 21431 18291 21437
rect 18322 21428 18328 21440
rect 18380 21428 18386 21480
rect 19613 21471 19671 21477
rect 19613 21437 19625 21471
rect 19659 21468 19671 21471
rect 21174 21468 21180 21480
rect 19659 21440 21180 21468
rect 19659 21437 19671 21440
rect 19613 21431 19671 21437
rect 21174 21428 21180 21440
rect 21232 21428 21238 21480
rect 22066 21468 22094 21508
rect 22278 21496 22284 21548
rect 22336 21536 22342 21548
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 22336 21508 22385 21536
rect 22336 21496 22342 21508
rect 22373 21505 22385 21508
rect 22419 21536 22431 21539
rect 23382 21536 23388 21548
rect 22419 21508 23388 21536
rect 22419 21505 22431 21508
rect 22373 21499 22431 21505
rect 23382 21496 23388 21508
rect 23440 21496 23446 21548
rect 24320 21545 24348 21576
rect 24578 21564 24584 21576
rect 24636 21564 24642 21616
rect 24946 21564 24952 21616
rect 25004 21604 25010 21616
rect 25004 21576 26464 21604
rect 25004 21564 25010 21576
rect 24305 21539 24363 21545
rect 24305 21505 24317 21539
rect 24351 21505 24363 21539
rect 24305 21499 24363 21505
rect 24673 21539 24731 21545
rect 24673 21505 24685 21539
rect 24719 21536 24731 21539
rect 24762 21536 24768 21548
rect 24719 21508 24768 21536
rect 24719 21505 24731 21508
rect 24673 21499 24731 21505
rect 24762 21496 24768 21508
rect 24820 21496 24826 21548
rect 25225 21539 25283 21545
rect 25225 21505 25237 21539
rect 25271 21536 25283 21539
rect 25406 21536 25412 21548
rect 25271 21508 25412 21536
rect 25271 21505 25283 21508
rect 25225 21499 25283 21505
rect 25406 21496 25412 21508
rect 25464 21496 25470 21548
rect 25501 21539 25559 21545
rect 25501 21505 25513 21539
rect 25547 21536 25559 21539
rect 25682 21536 25688 21548
rect 25547 21508 25688 21536
rect 25547 21505 25559 21508
rect 25501 21499 25559 21505
rect 25682 21496 25688 21508
rect 25740 21496 25746 21548
rect 26145 21539 26203 21545
rect 26145 21505 26157 21539
rect 26191 21536 26203 21539
rect 26326 21536 26332 21548
rect 26191 21508 26332 21536
rect 26191 21505 26203 21508
rect 26145 21499 26203 21505
rect 26326 21496 26332 21508
rect 26384 21496 26390 21548
rect 26436 21536 26464 21576
rect 26510 21564 26516 21616
rect 26568 21604 26574 21616
rect 27982 21604 27988 21616
rect 26568 21576 27988 21604
rect 26568 21564 26574 21576
rect 27982 21564 27988 21576
rect 28040 21564 28046 21616
rect 30374 21604 30380 21616
rect 29118 21576 30380 21604
rect 30374 21564 30380 21576
rect 30432 21564 30438 21616
rect 31404 21604 31432 21644
rect 32600 21644 34008 21672
rect 31570 21604 31576 21616
rect 31326 21576 31576 21604
rect 31570 21564 31576 21576
rect 31628 21564 31634 21616
rect 32600 21604 32628 21644
rect 32140 21576 32628 21604
rect 26973 21539 27031 21545
rect 26973 21536 26985 21539
rect 26436 21508 26985 21536
rect 26973 21505 26985 21508
rect 27019 21505 27031 21539
rect 27614 21536 27620 21548
rect 27575 21508 27620 21536
rect 26973 21499 27031 21505
rect 27614 21496 27620 21508
rect 27672 21496 27678 21548
rect 32140 21545 32168 21576
rect 32950 21564 32956 21616
rect 33008 21564 33014 21616
rect 32125 21539 32183 21545
rect 32125 21505 32137 21539
rect 32171 21505 32183 21539
rect 32125 21499 32183 21505
rect 22738 21468 22744 21480
rect 22066 21440 22744 21468
rect 22738 21428 22744 21440
rect 22796 21428 22802 21480
rect 26050 21428 26056 21480
rect 26108 21468 26114 21480
rect 27522 21468 27528 21480
rect 26108 21440 27528 21468
rect 26108 21428 26114 21440
rect 27522 21428 27528 21440
rect 27580 21428 27586 21480
rect 27893 21471 27951 21477
rect 27893 21437 27905 21471
rect 27939 21468 27951 21471
rect 28442 21468 28448 21480
rect 27939 21440 28448 21468
rect 27939 21437 27951 21440
rect 27893 21431 27951 21437
rect 28442 21428 28448 21440
rect 28500 21428 28506 21480
rect 29546 21468 29552 21480
rect 28966 21440 29552 21468
rect 19978 21360 19984 21412
rect 20036 21400 20042 21412
rect 20036 21372 25360 21400
rect 20036 21360 20042 21372
rect 1486 21332 1492 21344
rect 1447 21304 1492 21332
rect 1486 21292 1492 21304
rect 1544 21292 1550 21344
rect 18690 21332 18696 21344
rect 18651 21304 18696 21332
rect 18690 21292 18696 21304
rect 18748 21292 18754 21344
rect 20162 21332 20168 21344
rect 20123 21304 20168 21332
rect 20162 21292 20168 21304
rect 20220 21292 20226 21344
rect 20714 21292 20720 21344
rect 20772 21332 20778 21344
rect 20898 21332 20904 21344
rect 20772 21304 20904 21332
rect 20772 21292 20778 21304
rect 20898 21292 20904 21304
rect 20956 21292 20962 21344
rect 21269 21335 21327 21341
rect 21269 21301 21281 21335
rect 21315 21332 21327 21335
rect 21542 21332 21548 21344
rect 21315 21304 21548 21332
rect 21315 21301 21327 21304
rect 21269 21295 21327 21301
rect 21542 21292 21548 21304
rect 21600 21332 21606 21344
rect 21818 21332 21824 21344
rect 21600 21304 21824 21332
rect 21600 21292 21606 21304
rect 21818 21292 21824 21304
rect 21876 21292 21882 21344
rect 22278 21332 22284 21344
rect 22191 21304 22284 21332
rect 22278 21292 22284 21304
rect 22336 21332 22342 21344
rect 22922 21332 22928 21344
rect 22336 21304 22928 21332
rect 22336 21292 22342 21304
rect 22922 21292 22928 21304
rect 22980 21292 22986 21344
rect 23934 21292 23940 21344
rect 23992 21332 23998 21344
rect 24118 21332 24124 21344
rect 23992 21304 24124 21332
rect 23992 21292 23998 21304
rect 24118 21292 24124 21304
rect 24176 21292 24182 21344
rect 24210 21292 24216 21344
rect 24268 21332 24274 21344
rect 24486 21332 24492 21344
rect 24268 21304 24492 21332
rect 24268 21292 24274 21304
rect 24486 21292 24492 21304
rect 24544 21292 24550 21344
rect 24762 21292 24768 21344
rect 24820 21332 24826 21344
rect 24946 21332 24952 21344
rect 24820 21304 24952 21332
rect 24820 21292 24826 21304
rect 24946 21292 24952 21304
rect 25004 21292 25010 21344
rect 25332 21332 25360 21372
rect 25866 21360 25872 21412
rect 25924 21400 25930 21412
rect 25924 21372 27752 21400
rect 25924 21360 25930 21372
rect 26234 21332 26240 21344
rect 25332 21304 26240 21332
rect 26234 21292 26240 21304
rect 26292 21292 26298 21344
rect 26329 21335 26387 21341
rect 26329 21301 26341 21335
rect 26375 21332 26387 21335
rect 26786 21332 26792 21344
rect 26375 21304 26792 21332
rect 26375 21301 26387 21304
rect 26329 21295 26387 21301
rect 26786 21292 26792 21304
rect 26844 21292 26850 21344
rect 27062 21332 27068 21344
rect 27023 21304 27068 21332
rect 27062 21292 27068 21304
rect 27120 21292 27126 21344
rect 27724 21332 27752 21372
rect 28966 21332 28994 21440
rect 29546 21428 29552 21440
rect 29604 21468 29610 21480
rect 29825 21471 29883 21477
rect 29825 21468 29837 21471
rect 29604 21440 29837 21468
rect 29604 21428 29610 21440
rect 29825 21437 29837 21440
rect 29871 21437 29883 21471
rect 30101 21471 30159 21477
rect 30101 21468 30113 21471
rect 29825 21431 29883 21437
rect 29932 21440 30113 21468
rect 29178 21360 29184 21412
rect 29236 21400 29242 21412
rect 29932 21400 29960 21440
rect 30101 21437 30113 21440
rect 30147 21437 30159 21471
rect 30101 21431 30159 21437
rect 32401 21471 32459 21477
rect 32401 21437 32413 21471
rect 32447 21468 32459 21471
rect 32490 21468 32496 21480
rect 32447 21440 32496 21468
rect 32447 21437 32459 21440
rect 32401 21431 32459 21437
rect 32490 21428 32496 21440
rect 32548 21468 32554 21480
rect 33042 21468 33048 21480
rect 32548 21440 33048 21468
rect 32548 21428 32554 21440
rect 33042 21428 33048 21440
rect 33100 21428 33106 21480
rect 33980 21468 34008 21644
rect 34238 21632 34244 21684
rect 34296 21672 34302 21684
rect 37550 21672 37556 21684
rect 34296 21644 37556 21672
rect 34296 21632 34302 21644
rect 37550 21632 37556 21644
rect 37608 21632 37614 21684
rect 37642 21632 37648 21684
rect 37700 21672 37706 21684
rect 38749 21675 38807 21681
rect 38749 21672 38761 21675
rect 37700 21644 38761 21672
rect 37700 21632 37706 21644
rect 38749 21641 38761 21644
rect 38795 21641 38807 21675
rect 38749 21635 38807 21641
rect 39669 21675 39727 21681
rect 39669 21641 39681 21675
rect 39715 21672 39727 21675
rect 39850 21672 39856 21684
rect 39715 21644 39856 21672
rect 39715 21641 39727 21644
rect 39669 21635 39727 21641
rect 39850 21632 39856 21644
rect 39908 21632 39914 21684
rect 40034 21632 40040 21684
rect 40092 21672 40098 21684
rect 41601 21675 41659 21681
rect 41601 21672 41613 21675
rect 40092 21644 41613 21672
rect 40092 21632 40098 21644
rect 41601 21641 41613 21644
rect 41647 21641 41659 21675
rect 44082 21672 44088 21684
rect 44043 21644 44088 21672
rect 41601 21635 41659 21641
rect 44082 21632 44088 21644
rect 44140 21632 44146 21684
rect 58158 21672 58164 21684
rect 58119 21644 58164 21672
rect 58158 21632 58164 21644
rect 58216 21632 58222 21684
rect 34606 21604 34612 21616
rect 34567 21576 34612 21604
rect 34606 21564 34612 21576
rect 34664 21564 34670 21616
rect 35618 21564 35624 21616
rect 35676 21564 35682 21616
rect 39945 21607 40003 21613
rect 38626 21576 39896 21604
rect 34054 21496 34060 21548
rect 34112 21536 34118 21548
rect 34333 21539 34391 21545
rect 34333 21536 34345 21539
rect 34112 21508 34345 21536
rect 34112 21496 34118 21508
rect 34333 21505 34345 21508
rect 34379 21505 34391 21539
rect 34333 21499 34391 21505
rect 36630 21496 36636 21548
rect 36688 21536 36694 21548
rect 36725 21539 36783 21545
rect 36725 21536 36737 21539
rect 36688 21508 36737 21536
rect 36688 21496 36694 21508
rect 36725 21505 36737 21508
rect 36771 21505 36783 21539
rect 36725 21499 36783 21505
rect 36906 21496 36912 21548
rect 36964 21536 36970 21548
rect 37553 21539 37611 21545
rect 37553 21536 37565 21539
rect 36964 21508 37565 21536
rect 36964 21496 36970 21508
rect 37553 21505 37565 21508
rect 37599 21536 37611 21539
rect 38626 21536 38654 21576
rect 37599 21508 38654 21536
rect 37599 21505 37611 21508
rect 37553 21499 37611 21505
rect 38838 21496 38844 21548
rect 38896 21536 38902 21548
rect 39669 21539 39727 21545
rect 39669 21536 39681 21539
rect 38896 21508 39681 21536
rect 38896 21496 38902 21508
rect 39669 21505 39681 21508
rect 39715 21505 39727 21539
rect 39868 21536 39896 21576
rect 39945 21573 39957 21607
rect 39991 21604 40003 21607
rect 40218 21604 40224 21616
rect 39991 21576 40224 21604
rect 39991 21573 40003 21576
rect 39945 21567 40003 21573
rect 40218 21564 40224 21576
rect 40276 21564 40282 21616
rect 40310 21536 40316 21548
rect 39868 21508 40316 21536
rect 39669 21499 39727 21505
rect 40310 21496 40316 21508
rect 40368 21496 40374 21548
rect 40586 21536 40592 21548
rect 40547 21508 40592 21536
rect 40586 21496 40592 21508
rect 40644 21536 40650 21548
rect 41141 21539 41199 21545
rect 41141 21536 41153 21539
rect 40644 21508 41153 21536
rect 40644 21496 40650 21508
rect 41141 21505 41153 21508
rect 41187 21505 41199 21539
rect 41141 21499 41199 21505
rect 35066 21468 35072 21480
rect 33980 21440 35072 21468
rect 35066 21428 35072 21440
rect 35124 21428 35130 21480
rect 37277 21471 37335 21477
rect 36004 21440 37228 21468
rect 31846 21400 31852 21412
rect 29236 21372 29960 21400
rect 31496 21372 31852 21400
rect 29236 21360 29242 21372
rect 27724 21304 28994 21332
rect 29365 21335 29423 21341
rect 29365 21301 29377 21335
rect 29411 21332 29423 21335
rect 31496 21332 31524 21372
rect 31846 21360 31852 21372
rect 31904 21360 31910 21412
rect 35618 21360 35624 21412
rect 35676 21400 35682 21412
rect 36004 21400 36032 21440
rect 35676 21372 36032 21400
rect 35676 21360 35682 21372
rect 36078 21360 36084 21412
rect 36136 21400 36142 21412
rect 37200 21400 37228 21440
rect 37277 21437 37289 21471
rect 37323 21468 37335 21471
rect 37458 21468 37464 21480
rect 37323 21440 37464 21468
rect 37323 21437 37335 21440
rect 37277 21431 37335 21437
rect 37458 21428 37464 21440
rect 37516 21428 37522 21480
rect 37568 21440 38976 21468
rect 37568 21400 37596 21440
rect 38838 21400 38844 21412
rect 36136 21372 37136 21400
rect 37200 21372 37596 21400
rect 38799 21372 38844 21400
rect 36136 21360 36142 21372
rect 29411 21304 31524 21332
rect 31573 21335 31631 21341
rect 29411 21301 29423 21304
rect 29365 21295 29423 21301
rect 31573 21301 31585 21335
rect 31619 21332 31631 21335
rect 33594 21332 33600 21344
rect 31619 21304 33600 21332
rect 31619 21301 31631 21304
rect 31573 21295 31631 21301
rect 33594 21292 33600 21304
rect 33652 21292 33658 21344
rect 33873 21335 33931 21341
rect 33873 21301 33885 21335
rect 33919 21332 33931 21335
rect 35802 21332 35808 21344
rect 33919 21304 35808 21332
rect 33919 21301 33931 21304
rect 33873 21295 33931 21301
rect 35802 21292 35808 21304
rect 35860 21292 35866 21344
rect 36630 21332 36636 21344
rect 36591 21304 36636 21332
rect 36630 21292 36636 21304
rect 36688 21292 36694 21344
rect 37108 21332 37136 21372
rect 38838 21360 38844 21372
rect 38896 21360 38902 21412
rect 38948 21400 38976 21440
rect 39114 21428 39120 21480
rect 39172 21468 39178 21480
rect 39209 21471 39267 21477
rect 39209 21468 39221 21471
rect 39172 21440 39221 21468
rect 39172 21428 39178 21440
rect 39209 21437 39221 21440
rect 39255 21468 39267 21471
rect 40034 21468 40040 21480
rect 39255 21440 40040 21468
rect 39255 21437 39267 21440
rect 39209 21431 39267 21437
rect 40034 21428 40040 21440
rect 40092 21428 40098 21480
rect 40494 21428 40500 21480
rect 40552 21468 40558 21480
rect 41046 21468 41052 21480
rect 40552 21440 41052 21468
rect 40552 21428 40558 21440
rect 41046 21428 41052 21440
rect 41104 21428 41110 21480
rect 41506 21428 41512 21480
rect 41564 21468 41570 21480
rect 43073 21471 43131 21477
rect 43073 21468 43085 21471
rect 41564 21440 43085 21468
rect 41564 21428 41570 21440
rect 43073 21437 43085 21440
rect 43119 21468 43131 21471
rect 43119 21440 51074 21468
rect 43119 21437 43131 21440
rect 43073 21431 43131 21437
rect 39761 21403 39819 21409
rect 39761 21400 39773 21403
rect 38948 21372 39773 21400
rect 39761 21369 39773 21372
rect 39807 21400 39819 21403
rect 39850 21400 39856 21412
rect 39807 21372 39856 21400
rect 39807 21369 39819 21372
rect 39761 21363 39819 21369
rect 39850 21360 39856 21372
rect 39908 21360 39914 21412
rect 39942 21360 39948 21412
rect 40000 21400 40006 21412
rect 43533 21403 43591 21409
rect 43533 21400 43545 21403
rect 40000 21372 43545 21400
rect 40000 21360 40006 21372
rect 43533 21369 43545 21372
rect 43579 21369 43591 21403
rect 51046 21400 51074 21440
rect 57882 21400 57888 21412
rect 51046 21372 57888 21400
rect 43533 21363 43591 21369
rect 57882 21360 57888 21372
rect 57940 21360 57946 21412
rect 39482 21332 39488 21344
rect 37108 21304 39488 21332
rect 39482 21292 39488 21304
rect 39540 21292 39546 21344
rect 40494 21332 40500 21344
rect 40455 21304 40500 21332
rect 40494 21292 40500 21304
rect 40552 21292 40558 21344
rect 42518 21332 42524 21344
rect 42479 21304 42524 21332
rect 42518 21292 42524 21304
rect 42576 21292 42582 21344
rect 44542 21292 44548 21344
rect 44600 21332 44606 21344
rect 44729 21335 44787 21341
rect 44729 21332 44741 21335
rect 44600 21304 44741 21332
rect 44600 21292 44606 21304
rect 44729 21301 44741 21304
rect 44775 21332 44787 21335
rect 44818 21332 44824 21344
rect 44775 21304 44824 21332
rect 44775 21301 44787 21304
rect 44729 21295 44787 21301
rect 44818 21292 44824 21304
rect 44876 21292 44882 21344
rect 45281 21335 45339 21341
rect 45281 21301 45293 21335
rect 45327 21332 45339 21335
rect 46198 21332 46204 21344
rect 45327 21304 46204 21332
rect 45327 21301 45339 21304
rect 45281 21295 45339 21301
rect 46198 21292 46204 21304
rect 46256 21292 46262 21344
rect 1104 21242 58880 21264
rect 1104 21190 10582 21242
rect 10634 21190 10646 21242
rect 10698 21190 10710 21242
rect 10762 21190 10774 21242
rect 10826 21190 10838 21242
rect 10890 21190 29846 21242
rect 29898 21190 29910 21242
rect 29962 21190 29974 21242
rect 30026 21190 30038 21242
rect 30090 21190 30102 21242
rect 30154 21190 49110 21242
rect 49162 21190 49174 21242
rect 49226 21190 49238 21242
rect 49290 21190 49302 21242
rect 49354 21190 49366 21242
rect 49418 21190 58880 21242
rect 1104 21168 58880 21190
rect 15746 21128 15752 21140
rect 15707 21100 15752 21128
rect 15746 21088 15752 21100
rect 15804 21088 15810 21140
rect 16758 21088 16764 21140
rect 16816 21128 16822 21140
rect 17954 21128 17960 21140
rect 16816 21100 17960 21128
rect 16816 21088 16822 21100
rect 17954 21088 17960 21100
rect 18012 21088 18018 21140
rect 21818 21128 21824 21140
rect 21779 21100 21824 21128
rect 21818 21088 21824 21100
rect 21876 21088 21882 21140
rect 23753 21131 23811 21137
rect 23753 21097 23765 21131
rect 23799 21128 23811 21131
rect 24397 21131 24455 21137
rect 23799 21100 24348 21128
rect 23799 21097 23811 21100
rect 23753 21091 23811 21097
rect 18046 21020 18052 21072
rect 18104 21060 18110 21072
rect 19334 21060 19340 21072
rect 18104 21032 19340 21060
rect 18104 21020 18110 21032
rect 19334 21020 19340 21032
rect 19392 21020 19398 21072
rect 20070 21020 20076 21072
rect 20128 21060 20134 21072
rect 22094 21060 22100 21072
rect 20128 21032 22100 21060
rect 20128 21020 20134 21032
rect 22094 21020 22100 21032
rect 22152 21020 22158 21072
rect 24320 21060 24348 21100
rect 24397 21097 24409 21131
rect 24443 21128 24455 21131
rect 24486 21128 24492 21140
rect 24443 21100 24492 21128
rect 24443 21097 24455 21100
rect 24397 21091 24455 21097
rect 24486 21088 24492 21100
rect 24544 21088 24550 21140
rect 24946 21088 24952 21140
rect 25004 21128 25010 21140
rect 25130 21128 25136 21140
rect 25004 21100 25136 21128
rect 25004 21088 25010 21100
rect 25130 21088 25136 21100
rect 25188 21088 25194 21140
rect 27246 21128 27252 21140
rect 27207 21100 27252 21128
rect 27246 21088 27252 21100
rect 27304 21088 27310 21140
rect 30558 21128 30564 21140
rect 27724 21100 30564 21128
rect 25314 21060 25320 21072
rect 23124 21032 23888 21060
rect 24320 21032 25320 21060
rect 16850 20952 16856 21004
rect 16908 20992 16914 21004
rect 17862 20992 17868 21004
rect 16908 20964 17868 20992
rect 16908 20952 16914 20964
rect 17862 20952 17868 20964
rect 17920 20992 17926 21004
rect 17957 20995 18015 21001
rect 17957 20992 17969 20995
rect 17920 20964 17969 20992
rect 17920 20952 17926 20964
rect 17957 20961 17969 20964
rect 18003 20961 18015 20995
rect 17957 20955 18015 20961
rect 18693 20995 18751 21001
rect 18693 20961 18705 20995
rect 18739 20992 18751 20995
rect 22554 20992 22560 21004
rect 18739 20964 22324 20992
rect 22515 20964 22560 20992
rect 18739 20961 18751 20964
rect 18693 20955 18751 20961
rect 17678 20884 17684 20936
rect 17736 20924 17742 20936
rect 19889 20927 19947 20933
rect 19889 20924 19901 20927
rect 17736 20896 19901 20924
rect 17736 20884 17742 20896
rect 19889 20893 19901 20896
rect 19935 20893 19947 20927
rect 19889 20887 19947 20893
rect 20162 20884 20168 20936
rect 20220 20924 20226 20936
rect 20990 20924 20996 20936
rect 20220 20896 20996 20924
rect 20220 20884 20226 20896
rect 20990 20884 20996 20896
rect 21048 20884 21054 20936
rect 21177 20927 21235 20933
rect 21177 20893 21189 20927
rect 21223 20924 21235 20927
rect 21450 20924 21456 20936
rect 21223 20896 21456 20924
rect 21223 20893 21235 20896
rect 21177 20887 21235 20893
rect 21450 20884 21456 20896
rect 21508 20884 21514 20936
rect 21634 20924 21640 20936
rect 21595 20896 21640 20924
rect 21634 20884 21640 20896
rect 21692 20884 21698 20936
rect 22296 20918 22324 20964
rect 22554 20952 22560 20964
rect 22612 20952 22618 21004
rect 23014 20992 23020 21004
rect 22756 20964 23020 20992
rect 22465 20927 22523 20933
rect 22465 20918 22477 20927
rect 22296 20893 22477 20918
rect 22511 20924 22523 20927
rect 22756 20924 22784 20964
rect 23014 20952 23020 20964
rect 23072 20952 23078 21004
rect 23124 20924 23152 21032
rect 23385 20995 23443 21001
rect 23385 20961 23397 20995
rect 23431 20992 23443 20995
rect 23750 20992 23756 21004
rect 23431 20964 23756 20992
rect 23431 20961 23443 20964
rect 23385 20955 23443 20961
rect 23750 20952 23756 20964
rect 23808 20952 23814 21004
rect 22511 20896 22784 20924
rect 22848 20896 23152 20924
rect 23477 20927 23535 20933
rect 22511 20893 22523 20896
rect 22296 20890 22523 20893
rect 22465 20887 22523 20890
rect 15102 20816 15108 20868
rect 15160 20856 15166 20868
rect 21085 20859 21143 20865
rect 21085 20856 21097 20859
rect 15160 20828 21097 20856
rect 15160 20816 15166 20828
rect 21085 20825 21097 20828
rect 21131 20856 21143 20859
rect 22848 20856 22876 20896
rect 23477 20893 23489 20927
rect 23523 20924 23535 20927
rect 23566 20924 23572 20936
rect 23523 20896 23572 20924
rect 23523 20893 23535 20896
rect 23477 20887 23535 20893
rect 23566 20884 23572 20896
rect 23624 20884 23630 20936
rect 23860 20924 23888 21032
rect 25314 21020 25320 21032
rect 25372 21020 25378 21072
rect 26970 21020 26976 21072
rect 27028 21060 27034 21072
rect 27724 21060 27752 21100
rect 30558 21088 30564 21100
rect 30616 21088 30622 21140
rect 31570 21088 31576 21140
rect 31628 21128 31634 21140
rect 31628 21100 32260 21128
rect 31628 21088 31634 21100
rect 27028 21032 27752 21060
rect 27028 21020 27034 21032
rect 29546 21020 29552 21072
rect 29604 21060 29610 21072
rect 29604 21032 30696 21060
rect 29604 21020 29610 21032
rect 24670 20952 24676 21004
rect 24728 20992 24734 21004
rect 24949 20995 25007 21001
rect 24949 20992 24961 20995
rect 24728 20964 24961 20992
rect 24728 20952 24734 20964
rect 24949 20961 24961 20964
rect 24995 20961 25007 20995
rect 24949 20955 25007 20961
rect 25406 20952 25412 21004
rect 25464 20992 25470 21004
rect 25593 20995 25651 21001
rect 25593 20992 25605 20995
rect 25464 20964 25605 20992
rect 25464 20952 25470 20964
rect 25593 20961 25605 20964
rect 25639 20961 25651 20995
rect 26602 20992 26608 21004
rect 25593 20955 25651 20961
rect 26252 20964 26608 20992
rect 24486 20924 24492 20936
rect 23860 20896 24492 20924
rect 24486 20884 24492 20896
rect 24544 20924 24550 20936
rect 24544 20896 24808 20924
rect 24544 20884 24550 20896
rect 21131 20828 22876 20856
rect 21131 20825 21143 20828
rect 21085 20819 21143 20825
rect 22922 20816 22928 20868
rect 22980 20856 22986 20868
rect 24780 20856 24808 20896
rect 24854 20884 24860 20936
rect 24912 20924 24918 20936
rect 24912 20896 24957 20924
rect 24912 20884 24918 20896
rect 25774 20884 25780 20936
rect 25832 20924 25838 20936
rect 25869 20927 25927 20933
rect 25869 20924 25881 20927
rect 25832 20896 25881 20924
rect 25832 20884 25838 20896
rect 25869 20893 25881 20896
rect 25915 20893 25927 20927
rect 25869 20887 25927 20893
rect 26252 20856 26280 20964
rect 26602 20952 26608 20964
rect 26660 20952 26666 21004
rect 28626 20952 28632 21004
rect 28684 20992 28690 21004
rect 28721 20995 28779 21001
rect 28721 20992 28733 20995
rect 28684 20964 28733 20992
rect 28684 20952 28690 20964
rect 28721 20961 28733 20964
rect 28767 20961 28779 20995
rect 28721 20955 28779 20961
rect 28997 20995 29055 21001
rect 28997 20961 29009 20995
rect 29043 20992 29055 20995
rect 29270 20992 29276 21004
rect 29043 20964 29276 20992
rect 29043 20961 29055 20964
rect 28997 20955 29055 20961
rect 29270 20952 29276 20964
rect 29328 20952 29334 21004
rect 30006 20992 30012 21004
rect 29748 20964 30012 20992
rect 26326 20884 26332 20936
rect 26384 20924 26390 20936
rect 26513 20927 26571 20933
rect 26513 20924 26525 20927
rect 26384 20896 26525 20924
rect 26384 20884 26390 20896
rect 26513 20893 26525 20896
rect 26559 20924 26571 20927
rect 26878 20924 26884 20936
rect 26559 20896 26884 20924
rect 26559 20893 26571 20896
rect 26513 20887 26571 20893
rect 26878 20884 26884 20896
rect 26936 20884 26942 20936
rect 29178 20884 29184 20936
rect 29236 20924 29242 20936
rect 29748 20933 29776 20964
rect 30006 20952 30012 20964
rect 30064 20952 30070 21004
rect 30101 20995 30159 21001
rect 30101 20961 30113 20995
rect 30147 20992 30159 20995
rect 30466 20992 30472 21004
rect 30147 20964 30472 20992
rect 30147 20961 30159 20964
rect 30101 20955 30159 20961
rect 30466 20952 30472 20964
rect 30524 20952 30530 21004
rect 29733 20927 29791 20933
rect 29733 20924 29745 20927
rect 29236 20896 29745 20924
rect 29236 20884 29242 20896
rect 29733 20893 29745 20896
rect 29779 20893 29791 20927
rect 29733 20887 29791 20893
rect 29822 20884 29828 20936
rect 29880 20924 29886 20936
rect 30668 20933 30696 21032
rect 30929 20995 30987 21001
rect 30929 20961 30941 20995
rect 30975 20992 30987 20995
rect 32122 20992 32128 21004
rect 30975 20964 32128 20992
rect 30975 20961 30987 20964
rect 30929 20955 30987 20961
rect 32122 20952 32128 20964
rect 32180 20952 32186 21004
rect 30193 20927 30251 20933
rect 30193 20924 30205 20927
rect 29880 20896 29925 20924
rect 30116 20896 30205 20924
rect 29880 20884 29886 20896
rect 22980 20828 24532 20856
rect 24780 20828 26280 20856
rect 22980 20816 22986 20828
rect 13722 20748 13728 20800
rect 13780 20788 13786 20800
rect 16209 20791 16267 20797
rect 16209 20788 16221 20791
rect 13780 20760 16221 20788
rect 13780 20748 13786 20760
rect 16209 20757 16221 20760
rect 16255 20788 16267 20791
rect 16758 20788 16764 20800
rect 16255 20760 16764 20788
rect 16255 20757 16267 20760
rect 16209 20751 16267 20757
rect 16758 20748 16764 20760
rect 16816 20748 16822 20800
rect 17402 20788 17408 20800
rect 17315 20760 17408 20788
rect 17402 20748 17408 20760
rect 17460 20788 17466 20800
rect 17770 20788 17776 20800
rect 17460 20760 17776 20788
rect 17460 20748 17466 20760
rect 17770 20748 17776 20760
rect 17828 20748 17834 20800
rect 19429 20791 19487 20797
rect 19429 20757 19441 20791
rect 19475 20788 19487 20791
rect 19702 20788 19708 20800
rect 19475 20760 19708 20788
rect 19475 20757 19487 20760
rect 19429 20751 19487 20757
rect 19702 20748 19708 20760
rect 19760 20748 19766 20800
rect 20533 20791 20591 20797
rect 20533 20757 20545 20791
rect 20579 20788 20591 20791
rect 21634 20788 21640 20800
rect 20579 20760 21640 20788
rect 20579 20757 20591 20760
rect 20533 20751 20591 20757
rect 21634 20748 21640 20760
rect 21692 20748 21698 20800
rect 22830 20788 22836 20800
rect 22791 20760 22836 20788
rect 22830 20748 22836 20760
rect 22888 20748 22894 20800
rect 24504 20788 24532 20828
rect 26786 20816 26792 20868
rect 26844 20856 26850 20868
rect 26844 20828 26937 20856
rect 28290 20828 29224 20856
rect 26844 20816 26850 20828
rect 24765 20791 24823 20797
rect 24765 20788 24777 20791
rect 24504 20760 24777 20788
rect 24765 20757 24777 20760
rect 24811 20757 24823 20791
rect 26804 20788 26832 20816
rect 28442 20788 28448 20800
rect 26804 20760 28448 20788
rect 24765 20751 24823 20757
rect 28442 20748 28448 20760
rect 28500 20748 28506 20800
rect 29196 20788 29224 20828
rect 29270 20816 29276 20868
rect 29328 20856 29334 20868
rect 29549 20859 29607 20865
rect 29549 20856 29561 20859
rect 29328 20828 29561 20856
rect 29328 20816 29334 20828
rect 29549 20825 29561 20828
rect 29595 20825 29607 20859
rect 29549 20819 29607 20825
rect 29638 20816 29644 20868
rect 29696 20856 29702 20868
rect 30116 20856 30144 20896
rect 30193 20893 30205 20896
rect 30239 20893 30251 20927
rect 30193 20887 30251 20893
rect 30653 20927 30711 20933
rect 30653 20893 30665 20927
rect 30699 20893 30711 20927
rect 32232 20924 32260 21100
rect 32398 21088 32404 21140
rect 32456 21128 32462 21140
rect 32953 21131 33011 21137
rect 32953 21128 32965 21131
rect 32456 21100 32965 21128
rect 32456 21088 32462 21100
rect 32953 21097 32965 21100
rect 32999 21097 33011 21131
rect 39114 21128 39120 21140
rect 32953 21091 33011 21097
rect 33520 21100 39120 21128
rect 33520 21060 33548 21100
rect 39114 21088 39120 21100
rect 39172 21088 39178 21140
rect 39942 21088 39948 21140
rect 40000 21128 40006 21140
rect 40037 21131 40095 21137
rect 40037 21128 40049 21131
rect 40000 21100 40049 21128
rect 40000 21088 40006 21100
rect 40037 21097 40049 21100
rect 40083 21097 40095 21131
rect 40037 21091 40095 21097
rect 40586 21088 40592 21140
rect 40644 21128 40650 21140
rect 40770 21128 40776 21140
rect 40644 21100 40776 21128
rect 40644 21088 40650 21100
rect 40770 21088 40776 21100
rect 40828 21088 40834 21140
rect 42058 21128 42064 21140
rect 42019 21100 42064 21128
rect 42058 21088 42064 21100
rect 42116 21088 42122 21140
rect 42150 21088 42156 21140
rect 42208 21128 42214 21140
rect 42208 21100 43852 21128
rect 42208 21088 42214 21100
rect 32416 21032 33548 21060
rect 32416 21001 32444 21032
rect 34330 21020 34336 21072
rect 34388 21060 34394 21072
rect 34701 21063 34759 21069
rect 34701 21060 34713 21063
rect 34388 21032 34713 21060
rect 34388 21020 34394 21032
rect 34701 21029 34713 21032
rect 34747 21029 34759 21063
rect 38010 21060 38016 21072
rect 34701 21023 34759 21029
rect 36464 21032 38016 21060
rect 32401 20995 32459 21001
rect 32401 20961 32413 20995
rect 32447 20961 32459 20995
rect 32401 20955 32459 20961
rect 34054 20952 34060 21004
rect 34112 20992 34118 21004
rect 34422 20992 34428 21004
rect 34112 20964 34428 20992
rect 34112 20952 34118 20964
rect 34422 20952 34428 20964
rect 34480 20952 34486 21004
rect 32950 20924 32956 20936
rect 32062 20896 32956 20924
rect 30653 20887 30711 20893
rect 29696 20828 30144 20856
rect 29696 20816 29702 20828
rect 29914 20788 29920 20800
rect 29196 20760 29920 20788
rect 29914 20748 29920 20760
rect 29972 20748 29978 20800
rect 30009 20791 30067 20797
rect 30009 20757 30021 20791
rect 30055 20788 30067 20791
rect 30374 20788 30380 20800
rect 30055 20760 30380 20788
rect 30055 20757 30067 20760
rect 30009 20751 30067 20757
rect 30374 20748 30380 20760
rect 30432 20748 30438 20800
rect 30668 20788 30696 20887
rect 32950 20884 32956 20896
rect 33008 20924 33014 20936
rect 33137 20927 33195 20933
rect 33137 20924 33149 20927
rect 33008 20896 33149 20924
rect 33008 20884 33014 20896
rect 33137 20893 33149 20896
rect 33183 20893 33195 20927
rect 33137 20887 33195 20893
rect 33781 20927 33839 20933
rect 33781 20893 33793 20927
rect 33827 20924 33839 20927
rect 34514 20924 34520 20936
rect 33827 20896 34520 20924
rect 33827 20893 33839 20896
rect 33781 20887 33839 20893
rect 32398 20816 32404 20868
rect 32456 20856 32462 20868
rect 33796 20856 33824 20887
rect 34514 20884 34520 20896
rect 34572 20884 34578 20936
rect 36464 20933 36492 21032
rect 38010 21020 38016 21032
rect 38068 21020 38074 21072
rect 40310 21020 40316 21072
rect 40368 21060 40374 21072
rect 42613 21063 42671 21069
rect 42613 21060 42625 21063
rect 40368 21032 42625 21060
rect 40368 21020 40374 21032
rect 42613 21029 42625 21032
rect 42659 21029 42671 21063
rect 42613 21023 42671 21029
rect 36998 20952 37004 21004
rect 37056 20992 37062 21004
rect 43714 20992 43720 21004
rect 37056 20964 40724 20992
rect 37056 20952 37062 20964
rect 36449 20927 36507 20933
rect 36449 20893 36461 20927
rect 36495 20893 36507 20927
rect 38378 20924 38384 20936
rect 36449 20887 36507 20893
rect 36740 20896 38384 20924
rect 32456 20828 33824 20856
rect 32456 20816 32462 20828
rect 35710 20816 35716 20868
rect 35768 20816 35774 20868
rect 36173 20859 36231 20865
rect 36173 20825 36185 20859
rect 36219 20856 36231 20859
rect 36740 20856 36768 20896
rect 38378 20884 38384 20896
rect 38436 20884 38442 20936
rect 38746 20884 38752 20936
rect 38804 20924 38810 20936
rect 39301 20927 39359 20933
rect 39301 20924 39313 20927
rect 38804 20896 39313 20924
rect 38804 20884 38810 20896
rect 39301 20893 39313 20896
rect 39347 20893 39359 20927
rect 39301 20887 39359 20893
rect 39482 20884 39488 20936
rect 39540 20924 39546 20936
rect 40696 20933 40724 20964
rect 40788 20964 43720 20992
rect 40681 20927 40739 20933
rect 39540 20896 40080 20924
rect 39540 20884 39546 20896
rect 36906 20856 36912 20868
rect 36219 20828 36768 20856
rect 36867 20828 36912 20856
rect 36219 20825 36231 20828
rect 36173 20819 36231 20825
rect 36906 20816 36912 20828
rect 36964 20816 36970 20868
rect 38657 20859 38715 20865
rect 38657 20825 38669 20859
rect 38703 20856 38715 20859
rect 39942 20856 39948 20868
rect 38703 20828 39948 20856
rect 38703 20825 38715 20828
rect 38657 20819 38715 20825
rect 39942 20816 39948 20828
rect 40000 20816 40006 20868
rect 40052 20856 40080 20896
rect 40681 20893 40693 20927
rect 40727 20893 40739 20927
rect 40681 20887 40739 20893
rect 40788 20856 40816 20964
rect 43714 20952 43720 20964
rect 43772 20952 43778 21004
rect 41322 20924 41328 20936
rect 41283 20896 41328 20924
rect 41322 20884 41328 20896
rect 41380 20884 41386 20936
rect 41506 20924 41512 20936
rect 41467 20896 41512 20924
rect 41506 20884 41512 20896
rect 41564 20884 41570 20936
rect 43824 20933 43852 21100
rect 44082 21088 44088 21140
rect 44140 21128 44146 21140
rect 45005 21131 45063 21137
rect 45005 21128 45017 21131
rect 44140 21100 45017 21128
rect 44140 21088 44146 21100
rect 45005 21097 45017 21100
rect 45051 21128 45063 21131
rect 46474 21128 46480 21140
rect 45051 21100 46480 21128
rect 45051 21097 45063 21100
rect 45005 21091 45063 21097
rect 46474 21088 46480 21100
rect 46532 21088 46538 21140
rect 42153 20927 42211 20933
rect 42153 20893 42165 20927
rect 42199 20924 42211 20927
rect 43809 20927 43867 20933
rect 42199 20896 43300 20924
rect 42199 20893 42211 20896
rect 42153 20887 42211 20893
rect 43272 20868 43300 20896
rect 43809 20893 43821 20927
rect 43855 20924 43867 20927
rect 47854 20924 47860 20936
rect 43855 20896 47860 20924
rect 43855 20893 43867 20896
rect 43809 20887 43867 20893
rect 47854 20884 47860 20896
rect 47912 20884 47918 20936
rect 40052 20828 40816 20856
rect 40865 20859 40923 20865
rect 40865 20825 40877 20859
rect 40911 20856 40923 20859
rect 42978 20856 42984 20868
rect 40911 20828 42984 20856
rect 40911 20825 40923 20828
rect 40865 20819 40923 20825
rect 42978 20816 42984 20828
rect 43036 20816 43042 20868
rect 43254 20816 43260 20868
rect 43312 20856 43318 20868
rect 44361 20859 44419 20865
rect 44361 20856 44373 20859
rect 43312 20828 44373 20856
rect 43312 20816 43318 20828
rect 44361 20825 44373 20828
rect 44407 20856 44419 20859
rect 44407 20828 46244 20856
rect 44407 20825 44419 20828
rect 44361 20819 44419 20825
rect 46216 20800 46244 20828
rect 34146 20788 34152 20800
rect 30668 20760 34152 20788
rect 34146 20748 34152 20760
rect 34204 20748 34210 20800
rect 36538 20748 36544 20800
rect 36596 20788 36602 20800
rect 38746 20788 38752 20800
rect 36596 20760 38752 20788
rect 36596 20748 36602 20760
rect 38746 20748 38752 20760
rect 38804 20748 38810 20800
rect 39114 20748 39120 20800
rect 39172 20788 39178 20800
rect 39209 20791 39267 20797
rect 39209 20788 39221 20791
rect 39172 20760 39221 20788
rect 39172 20748 39178 20760
rect 39209 20757 39221 20760
rect 39255 20757 39267 20791
rect 39209 20751 39267 20757
rect 41417 20791 41475 20797
rect 41417 20757 41429 20791
rect 41463 20788 41475 20791
rect 41690 20788 41696 20800
rect 41463 20760 41696 20788
rect 41463 20757 41475 20760
rect 41417 20751 41475 20757
rect 41690 20748 41696 20760
rect 41748 20748 41754 20800
rect 43070 20748 43076 20800
rect 43128 20788 43134 20800
rect 43165 20791 43223 20797
rect 43165 20788 43177 20791
rect 43128 20760 43177 20788
rect 43128 20748 43134 20760
rect 43165 20757 43177 20760
rect 43211 20757 43223 20791
rect 43165 20751 43223 20757
rect 44818 20748 44824 20800
rect 44876 20788 44882 20800
rect 45649 20791 45707 20797
rect 45649 20788 45661 20791
rect 44876 20760 45661 20788
rect 44876 20748 44882 20760
rect 45649 20757 45661 20760
rect 45695 20788 45707 20791
rect 46014 20788 46020 20800
rect 45695 20760 46020 20788
rect 45695 20757 45707 20760
rect 45649 20751 45707 20757
rect 46014 20748 46020 20760
rect 46072 20748 46078 20800
rect 46198 20788 46204 20800
rect 46159 20760 46204 20788
rect 46198 20748 46204 20760
rect 46256 20748 46262 20800
rect 1104 20698 58880 20720
rect 1104 20646 20214 20698
rect 20266 20646 20278 20698
rect 20330 20646 20342 20698
rect 20394 20646 20406 20698
rect 20458 20646 20470 20698
rect 20522 20646 39478 20698
rect 39530 20646 39542 20698
rect 39594 20646 39606 20698
rect 39658 20646 39670 20698
rect 39722 20646 39734 20698
rect 39786 20646 58880 20698
rect 1104 20624 58880 20646
rect 12710 20544 12716 20596
rect 12768 20584 12774 20596
rect 16114 20584 16120 20596
rect 12768 20556 16120 20584
rect 12768 20544 12774 20556
rect 16114 20544 16120 20556
rect 16172 20544 16178 20596
rect 17034 20584 17040 20596
rect 16995 20556 17040 20584
rect 17034 20544 17040 20556
rect 17092 20544 17098 20596
rect 18141 20587 18199 20593
rect 18141 20553 18153 20587
rect 18187 20584 18199 20587
rect 18782 20584 18788 20596
rect 18187 20556 18788 20584
rect 18187 20553 18199 20556
rect 18141 20547 18199 20553
rect 18782 20544 18788 20556
rect 18840 20584 18846 20596
rect 20622 20584 20628 20596
rect 18840 20556 20628 20584
rect 18840 20544 18846 20556
rect 20622 20544 20628 20556
rect 20680 20544 20686 20596
rect 20993 20587 21051 20593
rect 20993 20553 21005 20587
rect 21039 20584 21051 20587
rect 21358 20584 21364 20596
rect 21039 20556 21364 20584
rect 21039 20553 21051 20556
rect 20993 20547 21051 20553
rect 21358 20544 21364 20556
rect 21416 20544 21422 20596
rect 21450 20544 21456 20596
rect 21508 20584 21514 20596
rect 25222 20584 25228 20596
rect 21508 20556 25228 20584
rect 21508 20544 21514 20556
rect 25222 20544 25228 20556
rect 25280 20544 25286 20596
rect 25498 20544 25504 20596
rect 25556 20584 25562 20596
rect 25556 20556 25820 20584
rect 25556 20544 25562 20556
rect 19794 20516 19800 20528
rect 19755 20488 19800 20516
rect 19794 20476 19800 20488
rect 19852 20476 19858 20528
rect 20806 20516 20812 20528
rect 20548 20488 20812 20516
rect 17586 20408 17592 20460
rect 17644 20448 17650 20460
rect 19889 20451 19947 20457
rect 17644 20420 18920 20448
rect 17644 20408 17650 20420
rect 18892 20380 18920 20420
rect 19889 20417 19901 20451
rect 19935 20448 19947 20451
rect 20070 20448 20076 20460
rect 19935 20420 20076 20448
rect 19935 20417 19947 20420
rect 19889 20411 19947 20417
rect 20070 20408 20076 20420
rect 20128 20408 20134 20460
rect 20548 20457 20576 20488
rect 20806 20476 20812 20488
rect 20864 20476 20870 20528
rect 22278 20516 22284 20528
rect 21284 20488 22284 20516
rect 21284 20457 21312 20488
rect 22278 20476 22284 20488
rect 22336 20476 22342 20528
rect 23750 20516 23756 20528
rect 22480 20488 23756 20516
rect 20533 20451 20591 20457
rect 20533 20417 20545 20451
rect 20579 20417 20591 20451
rect 21269 20451 21327 20457
rect 20533 20411 20591 20417
rect 20640 20420 21220 20448
rect 20640 20380 20668 20420
rect 18892 20352 20668 20380
rect 20806 20340 20812 20392
rect 20864 20380 20870 20392
rect 20993 20383 21051 20389
rect 20993 20380 21005 20383
rect 20864 20352 21005 20380
rect 20864 20340 20870 20352
rect 20993 20349 21005 20352
rect 21039 20380 21051 20383
rect 21082 20380 21088 20392
rect 21039 20352 21088 20380
rect 21039 20349 21051 20352
rect 20993 20343 21051 20349
rect 21082 20340 21088 20352
rect 21140 20340 21146 20392
rect 21192 20380 21220 20420
rect 21269 20417 21281 20451
rect 21315 20417 21327 20451
rect 21269 20411 21327 20417
rect 21634 20408 21640 20460
rect 21692 20448 21698 20460
rect 21821 20451 21879 20457
rect 21821 20448 21833 20451
rect 21692 20420 21833 20448
rect 21692 20408 21698 20420
rect 21821 20417 21833 20420
rect 21867 20448 21879 20451
rect 22480 20448 22508 20488
rect 23750 20476 23756 20488
rect 23808 20476 23814 20528
rect 24026 20516 24032 20528
rect 23987 20488 24032 20516
rect 24026 20476 24032 20488
rect 24084 20476 24090 20528
rect 24121 20519 24179 20525
rect 24121 20485 24133 20519
rect 24167 20516 24179 20519
rect 24302 20516 24308 20528
rect 24167 20488 24308 20516
rect 24167 20485 24179 20488
rect 24121 20479 24179 20485
rect 24302 20476 24308 20488
rect 24360 20476 24366 20528
rect 25792 20516 25820 20556
rect 26694 20544 26700 20596
rect 26752 20584 26758 20596
rect 29178 20584 29184 20596
rect 26752 20556 29184 20584
rect 26752 20544 26758 20556
rect 29178 20544 29184 20556
rect 29236 20544 29242 20596
rect 32122 20584 32128 20596
rect 29288 20556 31984 20584
rect 32083 20556 32128 20584
rect 26878 20516 26884 20528
rect 25714 20488 26884 20516
rect 26878 20476 26884 20488
rect 26936 20476 26942 20528
rect 29288 20516 29316 20556
rect 29454 20516 29460 20528
rect 28474 20488 29316 20516
rect 29415 20488 29460 20516
rect 29454 20476 29460 20488
rect 29512 20476 29518 20528
rect 30834 20516 30840 20528
rect 30682 20488 30840 20516
rect 30834 20476 30840 20488
rect 30892 20516 30898 20528
rect 31478 20516 31484 20528
rect 30892 20488 31484 20516
rect 30892 20476 30898 20488
rect 31478 20476 31484 20488
rect 31536 20476 31542 20528
rect 21867 20420 22508 20448
rect 22649 20451 22707 20457
rect 21867 20417 21879 20420
rect 21821 20411 21879 20417
rect 22649 20417 22661 20451
rect 22695 20448 22707 20451
rect 23198 20448 23204 20460
rect 22695 20420 23204 20448
rect 22695 20417 22707 20420
rect 22649 20411 22707 20417
rect 23198 20408 23204 20420
rect 23256 20408 23262 20460
rect 26421 20451 26479 20457
rect 26421 20417 26433 20451
rect 26467 20448 26479 20451
rect 26602 20448 26608 20460
rect 26467 20420 26608 20448
rect 26467 20417 26479 20420
rect 26421 20411 26479 20417
rect 26602 20408 26608 20420
rect 26660 20408 26666 20460
rect 26970 20448 26976 20460
rect 26931 20420 26976 20448
rect 26970 20408 26976 20420
rect 27028 20408 27034 20460
rect 31573 20451 31631 20457
rect 31573 20417 31585 20451
rect 31619 20448 31631 20451
rect 31662 20448 31668 20460
rect 31619 20420 31668 20448
rect 31619 20417 31631 20420
rect 31573 20411 31631 20417
rect 31662 20408 31668 20420
rect 31720 20408 31726 20460
rect 21192 20352 22094 20380
rect 15562 20312 15568 20324
rect 15523 20284 15568 20312
rect 15562 20272 15568 20284
rect 15620 20272 15626 20324
rect 18506 20272 18512 20324
rect 18564 20312 18570 20324
rect 18564 20284 18920 20312
rect 18564 20272 18570 20284
rect 18892 20256 18920 20284
rect 20070 20272 20076 20324
rect 20128 20312 20134 20324
rect 20441 20315 20499 20321
rect 20441 20312 20453 20315
rect 20128 20284 20453 20312
rect 20128 20272 20134 20284
rect 20441 20281 20453 20284
rect 20487 20281 20499 20315
rect 22066 20312 22094 20352
rect 22278 20340 22284 20392
rect 22336 20380 22342 20392
rect 22557 20383 22615 20389
rect 22557 20380 22569 20383
rect 22336 20352 22569 20380
rect 22336 20340 22342 20352
rect 22557 20349 22569 20352
rect 22603 20349 22615 20383
rect 23658 20380 23664 20392
rect 22557 20343 22615 20349
rect 22848 20352 23520 20380
rect 23619 20352 23664 20380
rect 22848 20312 22876 20352
rect 23014 20312 23020 20324
rect 22066 20284 22876 20312
rect 22975 20284 23020 20312
rect 20441 20275 20499 20281
rect 23014 20272 23020 20284
rect 23072 20272 23078 20324
rect 23492 20312 23520 20352
rect 23658 20340 23664 20352
rect 23716 20340 23722 20392
rect 23750 20340 23756 20392
rect 23808 20380 23814 20392
rect 24026 20380 24032 20392
rect 23808 20352 24032 20380
rect 23808 20340 23814 20352
rect 24026 20340 24032 20352
rect 24084 20340 24090 20392
rect 25774 20380 25780 20392
rect 24780 20352 25780 20380
rect 24302 20312 24308 20324
rect 23492 20284 24308 20312
rect 24302 20272 24308 20284
rect 24360 20312 24366 20324
rect 24673 20315 24731 20321
rect 24673 20312 24685 20315
rect 24360 20284 24685 20312
rect 24360 20272 24366 20284
rect 24673 20281 24685 20284
rect 24719 20281 24731 20315
rect 24673 20275 24731 20281
rect 13814 20204 13820 20256
rect 13872 20244 13878 20256
rect 14921 20247 14979 20253
rect 14921 20244 14933 20247
rect 13872 20216 14933 20244
rect 13872 20204 13878 20216
rect 14921 20213 14933 20216
rect 14967 20244 14979 20247
rect 15010 20244 15016 20256
rect 14967 20216 15016 20244
rect 14967 20213 14979 20216
rect 14921 20207 14979 20213
rect 15010 20204 15016 20216
rect 15068 20204 15074 20256
rect 17402 20204 17408 20256
rect 17460 20244 17466 20256
rect 17497 20247 17555 20253
rect 17497 20244 17509 20247
rect 17460 20216 17509 20244
rect 17460 20204 17466 20216
rect 17497 20213 17509 20216
rect 17543 20213 17555 20247
rect 17497 20207 17555 20213
rect 18046 20204 18052 20256
rect 18104 20244 18110 20256
rect 18601 20247 18659 20253
rect 18601 20244 18613 20247
rect 18104 20216 18613 20244
rect 18104 20204 18110 20216
rect 18601 20213 18613 20216
rect 18647 20213 18659 20247
rect 18601 20207 18659 20213
rect 18874 20204 18880 20256
rect 18932 20244 18938 20256
rect 19153 20247 19211 20253
rect 19153 20244 19165 20247
rect 18932 20216 19165 20244
rect 18932 20204 18938 20216
rect 19153 20213 19165 20216
rect 19199 20213 19211 20247
rect 21174 20244 21180 20256
rect 21087 20216 21180 20244
rect 19153 20207 19211 20213
rect 21174 20204 21180 20216
rect 21232 20244 21238 20256
rect 21358 20244 21364 20256
rect 21232 20216 21364 20244
rect 21232 20204 21238 20216
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 21818 20204 21824 20256
rect 21876 20244 21882 20256
rect 21913 20247 21971 20253
rect 21913 20244 21925 20247
rect 21876 20216 21925 20244
rect 21876 20204 21882 20216
rect 21913 20213 21925 20216
rect 21959 20213 21971 20247
rect 21913 20207 21971 20213
rect 22002 20204 22008 20256
rect 22060 20244 22066 20256
rect 24780 20244 24808 20352
rect 25774 20340 25780 20352
rect 25832 20340 25838 20392
rect 26050 20340 26056 20392
rect 26108 20380 26114 20392
rect 26145 20383 26203 20389
rect 26145 20380 26157 20383
rect 26108 20352 26157 20380
rect 26108 20340 26114 20352
rect 26145 20349 26157 20352
rect 26191 20380 26203 20383
rect 26694 20380 26700 20392
rect 26191 20352 26700 20380
rect 26191 20349 26203 20352
rect 26145 20343 26203 20349
rect 26694 20340 26700 20352
rect 26752 20340 26758 20392
rect 27249 20383 27307 20389
rect 27249 20380 27261 20383
rect 26804 20352 27261 20380
rect 24946 20272 24952 20324
rect 25004 20312 25010 20324
rect 25130 20312 25136 20324
rect 25004 20284 25136 20312
rect 25004 20272 25010 20284
rect 25130 20272 25136 20284
rect 25188 20272 25194 20324
rect 22060 20216 24808 20244
rect 22060 20204 22066 20216
rect 25038 20204 25044 20256
rect 25096 20244 25102 20256
rect 26804 20244 26832 20352
rect 27249 20349 27261 20352
rect 27295 20349 27307 20383
rect 27249 20343 27307 20349
rect 27338 20340 27344 20392
rect 27396 20380 27402 20392
rect 29181 20383 29239 20389
rect 29181 20380 29193 20383
rect 27396 20352 29193 20380
rect 27396 20340 27402 20352
rect 29181 20349 29193 20352
rect 29227 20349 29239 20383
rect 31956 20380 31984 20556
rect 32122 20544 32128 20556
rect 32180 20544 32186 20596
rect 32950 20544 32956 20596
rect 33008 20584 33014 20596
rect 33008 20556 35480 20584
rect 33008 20544 33014 20556
rect 33244 20516 33272 20556
rect 33594 20516 33600 20528
rect 33166 20488 33272 20516
rect 33507 20488 33600 20516
rect 33594 20476 33600 20488
rect 33652 20516 33658 20528
rect 33652 20488 34560 20516
rect 33652 20476 33658 20488
rect 33873 20451 33931 20457
rect 33873 20417 33885 20451
rect 33919 20448 33931 20451
rect 34146 20448 34152 20460
rect 33919 20420 34152 20448
rect 33919 20417 33931 20420
rect 33873 20411 33931 20417
rect 34146 20408 34152 20420
rect 34204 20408 34210 20460
rect 34532 20448 34560 20488
rect 35342 20476 35348 20528
rect 35400 20516 35406 20528
rect 35452 20516 35480 20556
rect 35710 20544 35716 20596
rect 35768 20584 35774 20596
rect 36633 20587 36691 20593
rect 36633 20584 36645 20587
rect 35768 20556 36645 20584
rect 35768 20544 35774 20556
rect 36633 20553 36645 20556
rect 36679 20553 36691 20587
rect 39114 20584 39120 20596
rect 36633 20547 36691 20553
rect 37384 20556 39120 20584
rect 35400 20488 35480 20516
rect 35400 20476 35406 20488
rect 36446 20476 36452 20528
rect 36504 20516 36510 20528
rect 36998 20516 37004 20528
rect 36504 20488 37004 20516
rect 36504 20476 36510 20488
rect 36998 20476 37004 20488
rect 37056 20476 37062 20528
rect 34532 20420 34652 20448
rect 34330 20380 34336 20392
rect 31956 20352 34336 20380
rect 29181 20343 29239 20349
rect 34330 20340 34336 20352
rect 34388 20340 34394 20392
rect 34514 20380 34520 20392
rect 34440 20352 34520 20380
rect 25096 20216 26832 20244
rect 28721 20247 28779 20253
rect 25096 20204 25102 20216
rect 28721 20213 28733 20247
rect 28767 20244 28779 20247
rect 30742 20244 30748 20256
rect 28767 20216 30748 20244
rect 28767 20213 28779 20216
rect 28721 20207 28779 20213
rect 30742 20204 30748 20216
rect 30800 20204 30806 20256
rect 30926 20204 30932 20256
rect 30984 20244 30990 20256
rect 31478 20244 31484 20256
rect 30984 20216 31029 20244
rect 31439 20216 31484 20244
rect 30984 20204 30990 20216
rect 31478 20204 31484 20216
rect 31536 20204 31542 20256
rect 34333 20247 34391 20253
rect 34333 20213 34345 20247
rect 34379 20244 34391 20247
rect 34440 20244 34468 20352
rect 34514 20340 34520 20352
rect 34572 20340 34578 20392
rect 34624 20380 34652 20420
rect 36078 20408 36084 20460
rect 36136 20448 36142 20460
rect 36725 20451 36783 20457
rect 36136 20420 36181 20448
rect 36136 20408 36142 20420
rect 36725 20417 36737 20451
rect 36771 20448 36783 20451
rect 37384 20448 37412 20556
rect 39114 20544 39120 20556
rect 39172 20584 39178 20596
rect 40865 20587 40923 20593
rect 40865 20584 40877 20587
rect 39172 20556 40877 20584
rect 39172 20544 39178 20556
rect 40865 20553 40877 20556
rect 40911 20553 40923 20587
rect 43162 20584 43168 20596
rect 43123 20556 43168 20584
rect 40865 20547 40923 20553
rect 43162 20544 43168 20556
rect 43220 20544 43226 20596
rect 45370 20584 45376 20596
rect 45331 20556 45376 20584
rect 45370 20544 45376 20556
rect 45428 20544 45434 20596
rect 46474 20584 46480 20596
rect 46435 20556 46480 20584
rect 46474 20544 46480 20556
rect 46532 20544 46538 20596
rect 38194 20476 38200 20528
rect 38252 20516 38258 20528
rect 39025 20519 39083 20525
rect 39025 20516 39037 20519
rect 38252 20488 39037 20516
rect 38252 20476 38258 20488
rect 39025 20485 39037 20488
rect 39071 20485 39083 20519
rect 39025 20479 39083 20485
rect 39942 20476 39948 20528
rect 40000 20516 40006 20528
rect 40957 20519 41015 20525
rect 40957 20516 40969 20519
rect 40000 20488 40969 20516
rect 40000 20476 40006 20488
rect 40957 20485 40969 20488
rect 41003 20485 41015 20519
rect 42518 20516 42524 20528
rect 40957 20479 41015 20485
rect 42076 20488 42524 20516
rect 42076 20460 42104 20488
rect 42518 20476 42524 20488
rect 42576 20476 42582 20528
rect 44269 20519 44327 20525
rect 44269 20516 44281 20519
rect 42628 20488 44281 20516
rect 42628 20460 42656 20488
rect 44269 20485 44281 20488
rect 44315 20485 44327 20519
rect 44269 20479 44327 20485
rect 37642 20448 37648 20460
rect 36771 20420 37412 20448
rect 37603 20420 37648 20448
rect 36771 20417 36783 20420
rect 36725 20411 36783 20417
rect 37642 20408 37648 20420
rect 37700 20408 37706 20460
rect 37918 20448 37924 20460
rect 37879 20420 37924 20448
rect 37918 20408 37924 20420
rect 37976 20408 37982 20460
rect 40037 20451 40095 20457
rect 40037 20417 40049 20451
rect 40083 20417 40095 20451
rect 40310 20448 40316 20460
rect 40271 20420 40316 20448
rect 40037 20411 40095 20417
rect 35158 20380 35164 20392
rect 34624 20352 35164 20380
rect 35158 20340 35164 20352
rect 35216 20340 35222 20392
rect 35805 20383 35863 20389
rect 35805 20349 35817 20383
rect 35851 20380 35863 20383
rect 35851 20352 36032 20380
rect 35851 20349 35863 20352
rect 35805 20343 35863 20349
rect 36004 20312 36032 20352
rect 36630 20340 36636 20392
rect 36688 20380 36694 20392
rect 37369 20383 37427 20389
rect 37369 20380 37381 20383
rect 36688 20352 37381 20380
rect 36688 20340 36694 20352
rect 37369 20349 37381 20352
rect 37415 20349 37427 20383
rect 38930 20380 38936 20392
rect 38891 20352 38936 20380
rect 37369 20343 37427 20349
rect 38930 20340 38936 20352
rect 38988 20340 38994 20392
rect 39206 20380 39212 20392
rect 39167 20352 39212 20380
rect 39206 20340 39212 20352
rect 39264 20340 39270 20392
rect 37274 20312 37280 20324
rect 36004 20284 37280 20312
rect 37274 20272 37280 20284
rect 37332 20272 37338 20324
rect 38838 20312 38844 20324
rect 37384 20284 38844 20312
rect 34379 20216 34468 20244
rect 34379 20213 34391 20216
rect 34333 20207 34391 20213
rect 35158 20204 35164 20256
rect 35216 20244 35222 20256
rect 37384 20244 37412 20284
rect 38838 20272 38844 20284
rect 38896 20312 38902 20324
rect 39942 20312 39948 20324
rect 38896 20284 39948 20312
rect 38896 20272 38902 20284
rect 39942 20272 39948 20284
rect 40000 20272 40006 20324
rect 40052 20312 40080 20411
rect 40310 20408 40316 20420
rect 40368 20408 40374 20460
rect 41693 20451 41751 20457
rect 41693 20417 41705 20451
rect 41739 20448 41751 20451
rect 42058 20448 42064 20460
rect 41739 20420 42064 20448
rect 41739 20417 41751 20420
rect 41693 20411 41751 20417
rect 42058 20408 42064 20420
rect 42116 20408 42122 20460
rect 42610 20448 42616 20460
rect 42523 20420 42616 20448
rect 42610 20408 42616 20420
rect 42668 20408 42674 20460
rect 43254 20448 43260 20460
rect 43215 20420 43260 20448
rect 43254 20408 43260 20420
rect 43312 20408 43318 20460
rect 40129 20383 40187 20389
rect 40129 20349 40141 20383
rect 40175 20380 40187 20383
rect 40218 20380 40224 20392
rect 40175 20352 40224 20380
rect 40175 20349 40187 20352
rect 40129 20343 40187 20349
rect 40218 20340 40224 20352
rect 40276 20380 40282 20392
rect 40954 20380 40960 20392
rect 40276 20352 40960 20380
rect 40276 20340 40282 20352
rect 40954 20340 40960 20352
rect 41012 20380 41018 20392
rect 43717 20383 43775 20389
rect 43717 20380 43729 20383
rect 41012 20352 43729 20380
rect 41012 20340 41018 20352
rect 43717 20349 43729 20352
rect 43763 20349 43775 20383
rect 43717 20343 43775 20349
rect 40494 20312 40500 20324
rect 40052 20284 40500 20312
rect 40494 20272 40500 20284
rect 40552 20312 40558 20324
rect 41138 20312 41144 20324
rect 40552 20284 41144 20312
rect 40552 20272 40558 20284
rect 41138 20272 41144 20284
rect 41196 20272 41202 20324
rect 35216 20216 37412 20244
rect 35216 20204 35222 20216
rect 39298 20204 39304 20256
rect 39356 20244 39362 20256
rect 40126 20244 40132 20256
rect 39356 20216 40132 20244
rect 39356 20204 39362 20216
rect 40126 20204 40132 20216
rect 40184 20204 40190 20256
rect 40221 20247 40279 20253
rect 40221 20213 40233 20247
rect 40267 20244 40279 20247
rect 40678 20244 40684 20256
rect 40267 20216 40684 20244
rect 40267 20213 40279 20216
rect 40221 20207 40279 20213
rect 40678 20204 40684 20216
rect 40736 20204 40742 20256
rect 41598 20244 41604 20256
rect 41559 20216 41604 20244
rect 41598 20204 41604 20216
rect 41656 20204 41662 20256
rect 42518 20244 42524 20256
rect 42479 20216 42524 20244
rect 42518 20204 42524 20216
rect 42576 20204 42582 20256
rect 44818 20244 44824 20256
rect 44779 20216 44824 20244
rect 44818 20204 44824 20216
rect 44876 20204 44882 20256
rect 46014 20244 46020 20256
rect 45975 20216 46020 20244
rect 46014 20204 46020 20216
rect 46072 20204 46078 20256
rect 1104 20154 58880 20176
rect 1104 20102 10582 20154
rect 10634 20102 10646 20154
rect 10698 20102 10710 20154
rect 10762 20102 10774 20154
rect 10826 20102 10838 20154
rect 10890 20102 29846 20154
rect 29898 20102 29910 20154
rect 29962 20102 29974 20154
rect 30026 20102 30038 20154
rect 30090 20102 30102 20154
rect 30154 20102 49110 20154
rect 49162 20102 49174 20154
rect 49226 20102 49238 20154
rect 49290 20102 49302 20154
rect 49354 20102 49366 20154
rect 49418 20102 58880 20154
rect 1104 20080 58880 20102
rect 15381 20043 15439 20049
rect 15381 20009 15393 20043
rect 15427 20040 15439 20043
rect 16574 20040 16580 20052
rect 15427 20012 16580 20040
rect 15427 20009 15439 20012
rect 15381 20003 15439 20009
rect 16574 20000 16580 20012
rect 16632 20000 16638 20052
rect 17589 20043 17647 20049
rect 17589 20009 17601 20043
rect 17635 20040 17647 20043
rect 18966 20040 18972 20052
rect 17635 20012 18972 20040
rect 17635 20009 17647 20012
rect 17589 20003 17647 20009
rect 18966 20000 18972 20012
rect 19024 20000 19030 20052
rect 19978 20000 19984 20052
rect 20036 20040 20042 20052
rect 20073 20043 20131 20049
rect 20073 20040 20085 20043
rect 20036 20012 20085 20040
rect 20036 20000 20042 20012
rect 20073 20009 20085 20012
rect 20119 20009 20131 20043
rect 20073 20003 20131 20009
rect 22097 20043 22155 20049
rect 22097 20009 22109 20043
rect 22143 20040 22155 20043
rect 27982 20040 27988 20052
rect 22143 20012 27988 20040
rect 22143 20009 22155 20012
rect 22097 20003 22155 20009
rect 27982 20000 27988 20012
rect 28040 20000 28046 20052
rect 28994 20000 29000 20052
rect 29052 20040 29058 20052
rect 36078 20040 36084 20052
rect 29052 20012 29097 20040
rect 34716 20012 36084 20040
rect 29052 20000 29058 20012
rect 12250 19972 12256 19984
rect 12211 19944 12256 19972
rect 12250 19932 12256 19944
rect 12308 19932 12314 19984
rect 17037 19975 17095 19981
rect 17037 19941 17049 19975
rect 17083 19972 17095 19975
rect 19150 19972 19156 19984
rect 17083 19944 19156 19972
rect 17083 19941 17095 19944
rect 17037 19935 17095 19941
rect 19150 19932 19156 19944
rect 19208 19972 19214 19984
rect 21174 19972 21180 19984
rect 19208 19944 20852 19972
rect 21135 19944 21180 19972
rect 19208 19932 19214 19944
rect 19426 19864 19432 19916
rect 19484 19904 19490 19916
rect 19484 19876 20116 19904
rect 19484 19864 19490 19876
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19836 1731 19839
rect 12066 19836 12072 19848
rect 1719 19808 12072 19836
rect 1719 19805 1731 19808
rect 1673 19799 1731 19805
rect 12066 19796 12072 19808
rect 12124 19796 12130 19848
rect 12437 19839 12495 19845
rect 12437 19805 12449 19839
rect 12483 19836 12495 19839
rect 15102 19836 15108 19848
rect 12483 19808 15108 19836
rect 12483 19805 12495 19808
rect 12437 19799 12495 19805
rect 15102 19796 15108 19808
rect 15160 19796 15166 19848
rect 16390 19796 16396 19848
rect 16448 19836 16454 19848
rect 19536 19845 19564 19876
rect 18601 19839 18659 19845
rect 18601 19836 18613 19839
rect 16448 19808 18613 19836
rect 16448 19796 16454 19808
rect 18601 19805 18613 19808
rect 18647 19805 18659 19839
rect 18601 19799 18659 19805
rect 19521 19839 19579 19845
rect 19521 19805 19533 19839
rect 19567 19805 19579 19839
rect 19521 19799 19579 19805
rect 19981 19839 20039 19845
rect 19981 19805 19993 19839
rect 20027 19805 20039 19839
rect 20088 19836 20116 19876
rect 20622 19864 20628 19916
rect 20680 19904 20686 19916
rect 20717 19907 20775 19913
rect 20717 19904 20729 19907
rect 20680 19876 20729 19904
rect 20680 19864 20686 19876
rect 20717 19873 20729 19876
rect 20763 19873 20775 19907
rect 20717 19867 20775 19873
rect 20824 19845 20852 19944
rect 21174 19932 21180 19944
rect 21232 19932 21238 19984
rect 23658 19972 23664 19984
rect 23584 19944 23664 19972
rect 21913 19907 21971 19913
rect 21913 19873 21925 19907
rect 21959 19904 21971 19907
rect 22002 19904 22008 19916
rect 21959 19876 22008 19904
rect 21959 19873 21971 19876
rect 21913 19867 21971 19873
rect 22002 19864 22008 19876
rect 22060 19864 22066 19916
rect 22462 19864 22468 19916
rect 22520 19904 22526 19916
rect 22646 19904 22652 19916
rect 22520 19876 22652 19904
rect 22520 19864 22526 19876
rect 22646 19864 22652 19876
rect 22704 19864 22710 19916
rect 20809 19839 20867 19845
rect 20088 19808 20760 19836
rect 19981 19799 20039 19805
rect 15933 19771 15991 19777
rect 15933 19737 15945 19771
rect 15979 19768 15991 19771
rect 18506 19768 18512 19780
rect 15979 19740 18512 19768
rect 15979 19737 15991 19740
rect 15933 19731 15991 19737
rect 18506 19728 18512 19740
rect 18564 19728 18570 19780
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 12986 19660 12992 19712
rect 13044 19700 13050 19712
rect 13722 19700 13728 19712
rect 13044 19672 13728 19700
rect 13044 19660 13050 19672
rect 13722 19660 13728 19672
rect 13780 19700 13786 19712
rect 14185 19703 14243 19709
rect 14185 19700 14197 19703
rect 13780 19672 14197 19700
rect 13780 19660 13786 19672
rect 14185 19669 14197 19672
rect 14231 19669 14243 19703
rect 14826 19700 14832 19712
rect 14787 19672 14832 19700
rect 14185 19663 14243 19669
rect 14826 19660 14832 19672
rect 14884 19660 14890 19712
rect 16206 19660 16212 19712
rect 16264 19700 16270 19712
rect 16393 19703 16451 19709
rect 16393 19700 16405 19703
rect 16264 19672 16405 19700
rect 16264 19660 16270 19672
rect 16393 19669 16405 19672
rect 16439 19669 16451 19703
rect 16393 19663 16451 19669
rect 17862 19660 17868 19712
rect 17920 19700 17926 19712
rect 18049 19703 18107 19709
rect 18049 19700 18061 19703
rect 17920 19672 18061 19700
rect 17920 19660 17926 19672
rect 18049 19669 18061 19672
rect 18095 19669 18107 19703
rect 18616 19700 18644 19799
rect 19426 19768 19432 19780
rect 19387 19740 19432 19768
rect 19426 19728 19432 19740
rect 19484 19728 19490 19780
rect 19996 19700 20024 19799
rect 18616 19672 20024 19700
rect 20732 19700 20760 19808
rect 20809 19805 20821 19839
rect 20855 19805 20867 19839
rect 20809 19799 20867 19805
rect 21174 19796 21180 19848
rect 21232 19836 21238 19848
rect 21821 19839 21879 19845
rect 21821 19836 21833 19839
rect 21232 19808 21833 19836
rect 21232 19796 21238 19808
rect 21821 19805 21833 19808
rect 21867 19805 21879 19839
rect 22922 19836 22928 19848
rect 22883 19808 22928 19836
rect 21821 19799 21879 19805
rect 22922 19796 22928 19808
rect 22980 19796 22986 19848
rect 23584 19845 23612 19944
rect 23658 19932 23664 19944
rect 23716 19932 23722 19984
rect 24489 19975 24547 19981
rect 24489 19941 24501 19975
rect 24535 19972 24547 19975
rect 24578 19972 24584 19984
rect 24535 19944 24584 19972
rect 24535 19941 24547 19944
rect 24489 19935 24547 19941
rect 24578 19932 24584 19944
rect 24636 19932 24642 19984
rect 26789 19975 26847 19981
rect 26789 19941 26801 19975
rect 26835 19972 26847 19975
rect 27154 19972 27160 19984
rect 26835 19944 27160 19972
rect 26835 19941 26847 19944
rect 26789 19935 26847 19941
rect 27154 19932 27160 19944
rect 27212 19932 27218 19984
rect 28718 19932 28724 19984
rect 28776 19972 28782 19984
rect 29549 19975 29607 19981
rect 29549 19972 29561 19975
rect 28776 19944 29561 19972
rect 28776 19932 28782 19944
rect 29549 19941 29561 19944
rect 29595 19941 29607 19975
rect 29549 19935 29607 19941
rect 25317 19907 25375 19913
rect 25317 19904 25329 19907
rect 23676 19876 25329 19904
rect 23569 19839 23627 19845
rect 23569 19805 23581 19839
rect 23615 19805 23627 19839
rect 23569 19799 23627 19805
rect 20990 19728 20996 19780
rect 21048 19768 21054 19780
rect 23676 19768 23704 19876
rect 25317 19873 25329 19876
rect 25363 19873 25375 19907
rect 25317 19867 25375 19873
rect 25406 19864 25412 19916
rect 25464 19904 25470 19916
rect 26602 19904 26608 19916
rect 25464 19876 26608 19904
rect 25464 19864 25470 19876
rect 26602 19864 26608 19876
rect 26660 19864 26666 19916
rect 26694 19864 26700 19916
rect 26752 19904 26758 19916
rect 27249 19907 27307 19913
rect 27249 19904 27261 19907
rect 26752 19876 27261 19904
rect 26752 19864 26758 19876
rect 27249 19873 27261 19876
rect 27295 19873 27307 19907
rect 27249 19867 27307 19873
rect 27525 19907 27583 19913
rect 27525 19873 27537 19907
rect 27571 19904 27583 19907
rect 28258 19904 28264 19916
rect 27571 19876 28264 19904
rect 27571 19873 27583 19876
rect 27525 19867 27583 19873
rect 28258 19864 28264 19876
rect 28316 19864 28322 19916
rect 30193 19907 30251 19913
rect 30193 19873 30205 19907
rect 30239 19904 30251 19907
rect 30558 19904 30564 19916
rect 30239 19876 30564 19904
rect 30239 19873 30251 19876
rect 30193 19867 30251 19873
rect 30558 19864 30564 19876
rect 30616 19864 30622 19916
rect 32585 19907 32643 19913
rect 32585 19873 32597 19907
rect 32631 19904 32643 19907
rect 32674 19904 32680 19916
rect 32631 19876 32680 19904
rect 32631 19873 32643 19876
rect 32585 19867 32643 19873
rect 32674 19864 32680 19876
rect 32732 19864 32738 19916
rect 33318 19864 33324 19916
rect 33376 19904 33382 19916
rect 33376 19876 33732 19904
rect 33376 19864 33382 19876
rect 33704 19848 33732 19876
rect 33870 19864 33876 19916
rect 33928 19904 33934 19916
rect 34716 19913 34744 20012
rect 36078 20000 36084 20012
rect 36136 20000 36142 20052
rect 37550 20000 37556 20052
rect 37608 20040 37614 20052
rect 37918 20040 37924 20052
rect 37608 20012 37924 20040
rect 37608 20000 37614 20012
rect 37918 20000 37924 20012
rect 37976 20000 37982 20052
rect 38654 20040 38660 20052
rect 38615 20012 38660 20040
rect 38654 20000 38660 20012
rect 38712 20000 38718 20052
rect 39390 20000 39396 20052
rect 39448 20040 39454 20052
rect 39853 20043 39911 20049
rect 39853 20040 39865 20043
rect 39448 20012 39865 20040
rect 39448 20000 39454 20012
rect 39853 20009 39865 20012
rect 39899 20009 39911 20043
rect 40770 20040 40776 20052
rect 40731 20012 40776 20040
rect 39853 20003 39911 20009
rect 40770 20000 40776 20012
rect 40828 20000 40834 20052
rect 41782 20040 41788 20052
rect 41743 20012 41788 20040
rect 41782 20000 41788 20012
rect 41840 20000 41846 20052
rect 44269 20043 44327 20049
rect 44269 20009 44281 20043
rect 44315 20040 44327 20043
rect 44818 20040 44824 20052
rect 44315 20012 44824 20040
rect 44315 20009 44327 20012
rect 44269 20003 44327 20009
rect 39206 19972 39212 19984
rect 38212 19944 39212 19972
rect 34701 19907 34759 19913
rect 34701 19904 34713 19907
rect 33928 19876 34713 19904
rect 33928 19864 33934 19876
rect 34701 19873 34713 19876
rect 34747 19873 34759 19907
rect 34974 19904 34980 19916
rect 34935 19876 34980 19904
rect 34701 19867 34759 19873
rect 34974 19864 34980 19876
rect 35032 19864 35038 19916
rect 36909 19907 36967 19913
rect 36909 19873 36921 19907
rect 36955 19904 36967 19907
rect 38212 19904 38240 19944
rect 39206 19932 39212 19944
rect 39264 19932 39270 19984
rect 40034 19972 40040 19984
rect 39995 19944 40040 19972
rect 40034 19932 40040 19944
rect 40092 19932 40098 19984
rect 40862 19932 40868 19984
rect 40920 19972 40926 19984
rect 40920 19944 40965 19972
rect 40920 19932 40926 19944
rect 43073 19907 43131 19913
rect 43073 19904 43085 19907
rect 36955 19876 38240 19904
rect 38304 19876 43085 19904
rect 36955 19873 36967 19876
rect 36909 19867 36967 19873
rect 24118 19796 24124 19848
rect 24176 19836 24182 19848
rect 24397 19839 24455 19845
rect 24397 19836 24409 19839
rect 24176 19808 24409 19836
rect 24176 19796 24182 19808
rect 24397 19805 24409 19808
rect 24443 19836 24455 19839
rect 24762 19836 24768 19848
rect 24443 19808 24768 19836
rect 24443 19805 24455 19808
rect 24397 19799 24455 19805
rect 24762 19796 24768 19808
rect 24820 19796 24826 19848
rect 25041 19839 25099 19845
rect 25041 19805 25053 19839
rect 25087 19805 25099 19839
rect 25041 19799 25099 19805
rect 21048 19740 23704 19768
rect 23845 19771 23903 19777
rect 21048 19728 21054 19740
rect 23845 19737 23857 19771
rect 23891 19737 23903 19771
rect 25056 19768 25084 19799
rect 28626 19796 28632 19848
rect 28684 19796 28690 19848
rect 29730 19796 29736 19848
rect 29788 19836 29794 19848
rect 30745 19839 30803 19845
rect 30745 19836 30757 19839
rect 29788 19808 30757 19836
rect 29788 19796 29794 19808
rect 30745 19805 30757 19808
rect 30791 19805 30803 19839
rect 30745 19799 30803 19805
rect 25406 19768 25412 19780
rect 25056 19740 25412 19768
rect 23845 19731 23903 19737
rect 22094 19700 22100 19712
rect 20732 19672 22100 19700
rect 18049 19663 18107 19669
rect 22094 19660 22100 19672
rect 22152 19660 22158 19712
rect 23566 19660 23572 19712
rect 23624 19700 23630 19712
rect 23860 19700 23888 19731
rect 25406 19728 25412 19740
rect 25464 19728 25470 19780
rect 26878 19768 26884 19780
rect 26542 19740 26884 19768
rect 26878 19728 26884 19740
rect 26936 19768 26942 19780
rect 30760 19768 30788 19799
rect 33686 19796 33692 19848
rect 33744 19836 33750 19848
rect 34057 19839 34115 19845
rect 33744 19808 33789 19836
rect 33744 19796 33750 19808
rect 34057 19805 34069 19839
rect 34103 19805 34115 19839
rect 38304 19822 38332 19876
rect 43073 19873 43085 19876
rect 43119 19873 43131 19907
rect 43073 19867 43131 19873
rect 34057 19799 34115 19805
rect 32306 19768 32312 19780
rect 26936 19740 27108 19768
rect 26936 19728 26942 19740
rect 24210 19700 24216 19712
rect 23624 19672 24216 19700
rect 23624 19660 23630 19672
rect 24210 19660 24216 19672
rect 24268 19700 24274 19712
rect 26694 19700 26700 19712
rect 24268 19672 26700 19700
rect 24268 19660 24274 19672
rect 26694 19660 26700 19672
rect 26752 19660 26758 19712
rect 27080 19700 27108 19740
rect 28966 19740 30328 19768
rect 30760 19740 32312 19768
rect 28966 19700 28994 19740
rect 27080 19672 28994 19700
rect 29362 19660 29368 19712
rect 29420 19700 29426 19712
rect 29917 19703 29975 19709
rect 29917 19700 29929 19703
rect 29420 19672 29929 19700
rect 29420 19660 29426 19672
rect 29917 19669 29929 19672
rect 29963 19669 29975 19703
rect 29917 19663 29975 19669
rect 30009 19703 30067 19709
rect 30009 19669 30021 19703
rect 30055 19700 30067 19703
rect 30190 19700 30196 19712
rect 30055 19672 30196 19700
rect 30055 19669 30067 19672
rect 30009 19663 30067 19669
rect 30190 19660 30196 19672
rect 30248 19660 30254 19712
rect 30300 19700 30328 19740
rect 32306 19728 32312 19740
rect 32364 19728 32370 19780
rect 32401 19771 32459 19777
rect 32401 19737 32413 19771
rect 32447 19768 32459 19771
rect 33045 19771 33103 19777
rect 33045 19768 33057 19771
rect 32447 19740 33057 19768
rect 32447 19737 32459 19740
rect 32401 19731 32459 19737
rect 33045 19737 33057 19740
rect 33091 19737 33103 19771
rect 34072 19768 34100 19799
rect 38746 19796 38752 19848
rect 38804 19836 38810 19848
rect 38930 19836 38936 19848
rect 38804 19808 38936 19836
rect 38804 19796 38810 19808
rect 38930 19796 38936 19808
rect 38988 19836 38994 19848
rect 39117 19839 39175 19845
rect 39117 19836 39129 19839
rect 38988 19808 39129 19836
rect 38988 19796 38994 19808
rect 39117 19805 39129 19808
rect 39163 19805 39175 19839
rect 39117 19799 39175 19805
rect 39209 19839 39267 19845
rect 39209 19805 39221 19839
rect 39255 19805 39267 19839
rect 39209 19799 39267 19805
rect 34882 19768 34888 19780
rect 34072 19740 34888 19768
rect 33045 19731 33103 19737
rect 34882 19728 34888 19740
rect 34940 19728 34946 19780
rect 35434 19728 35440 19780
rect 35492 19728 35498 19780
rect 37090 19728 37096 19780
rect 37148 19768 37154 19780
rect 37185 19771 37243 19777
rect 37185 19768 37197 19771
rect 37148 19740 37197 19768
rect 37148 19728 37154 19740
rect 37185 19737 37197 19740
rect 37231 19737 37243 19771
rect 37185 19731 37243 19737
rect 37458 19728 37464 19780
rect 37516 19728 37522 19780
rect 38838 19728 38844 19780
rect 38896 19768 38902 19780
rect 39224 19768 39252 19799
rect 39758 19796 39764 19848
rect 39816 19836 39822 19848
rect 40034 19836 40040 19848
rect 39816 19808 40040 19836
rect 39816 19796 39822 19808
rect 40034 19796 40040 19808
rect 40092 19796 40098 19848
rect 40144 19808 40448 19836
rect 40144 19768 40172 19808
rect 38896 19740 39252 19768
rect 39868 19740 40172 19768
rect 40313 19771 40371 19777
rect 38896 19728 38902 19740
rect 30834 19700 30840 19712
rect 30300 19672 30840 19700
rect 30834 19660 30840 19672
rect 30892 19660 30898 19712
rect 31846 19660 31852 19712
rect 31904 19700 31910 19712
rect 36446 19700 36452 19712
rect 31904 19672 36452 19700
rect 31904 19660 31910 19672
rect 36446 19660 36452 19672
rect 36504 19700 36510 19712
rect 37476 19700 37504 19728
rect 36504 19672 37504 19700
rect 36504 19660 36510 19672
rect 37550 19660 37556 19712
rect 37608 19700 37614 19712
rect 39868 19700 39896 19740
rect 40313 19737 40325 19771
rect 40359 19737 40371 19771
rect 40313 19731 40371 19737
rect 37608 19672 39896 19700
rect 37608 19660 37614 19672
rect 39942 19660 39948 19712
rect 40000 19700 40006 19712
rect 40328 19700 40356 19731
rect 40000 19672 40356 19700
rect 40420 19700 40448 19808
rect 41046 19796 41052 19848
rect 41104 19836 41110 19848
rect 41877 19839 41935 19845
rect 41104 19808 41414 19836
rect 41104 19796 41110 19808
rect 41138 19728 41144 19780
rect 41196 19768 41202 19780
rect 41233 19771 41291 19777
rect 41233 19768 41245 19771
rect 41196 19740 41245 19768
rect 41196 19728 41202 19740
rect 41233 19737 41245 19740
rect 41279 19737 41291 19771
rect 41386 19768 41414 19808
rect 41877 19805 41889 19839
rect 41923 19836 41935 19839
rect 42150 19836 42156 19848
rect 41923 19808 42156 19836
rect 41923 19805 41935 19808
rect 41877 19799 41935 19805
rect 42150 19796 42156 19808
rect 42208 19796 42214 19848
rect 42521 19839 42579 19845
rect 42521 19805 42533 19839
rect 42567 19805 42579 19839
rect 42521 19799 42579 19805
rect 42536 19768 42564 19799
rect 42978 19796 42984 19848
rect 43036 19836 43042 19848
rect 43165 19839 43223 19845
rect 43165 19836 43177 19839
rect 43036 19808 43177 19836
rect 43036 19796 43042 19808
rect 43165 19805 43177 19808
rect 43211 19836 43223 19839
rect 43806 19836 43812 19848
rect 43211 19808 43812 19836
rect 43211 19805 43223 19808
rect 43165 19799 43223 19805
rect 43806 19796 43812 19808
rect 43864 19796 43870 19848
rect 44284 19768 44312 20003
rect 44818 20000 44824 20012
rect 44876 20000 44882 20052
rect 46474 20000 46480 20052
rect 46532 20040 46538 20052
rect 46658 20040 46664 20052
rect 46532 20012 46664 20040
rect 46532 20000 46538 20012
rect 46658 20000 46664 20012
rect 46716 20000 46722 20052
rect 46934 19864 46940 19916
rect 46992 19904 46998 19916
rect 46992 19876 51074 19904
rect 46992 19864 46998 19876
rect 46198 19796 46204 19848
rect 46256 19836 46262 19848
rect 47305 19839 47363 19845
rect 47305 19836 47317 19839
rect 46256 19808 47317 19836
rect 46256 19796 46262 19808
rect 47305 19805 47317 19808
rect 47351 19836 47363 19839
rect 47351 19808 47992 19836
rect 47351 19805 47363 19808
rect 47305 19799 47363 19805
rect 41386 19740 44312 19768
rect 41233 19731 41291 19737
rect 42429 19703 42487 19709
rect 42429 19700 42441 19703
rect 40420 19672 42441 19700
rect 40000 19660 40006 19672
rect 42429 19669 42441 19672
rect 42475 19669 42487 19703
rect 42429 19663 42487 19669
rect 43717 19703 43775 19709
rect 43717 19669 43729 19703
rect 43763 19700 43775 19703
rect 44082 19700 44088 19712
rect 43763 19672 44088 19700
rect 43763 19669 43775 19672
rect 43717 19663 43775 19669
rect 44082 19660 44088 19672
rect 44140 19660 44146 19712
rect 44542 19660 44548 19712
rect 44600 19700 44606 19712
rect 45005 19703 45063 19709
rect 45005 19700 45017 19703
rect 44600 19672 45017 19700
rect 44600 19660 44606 19672
rect 45005 19669 45017 19672
rect 45051 19669 45063 19703
rect 45005 19663 45063 19669
rect 45554 19660 45560 19712
rect 45612 19700 45618 19712
rect 45649 19703 45707 19709
rect 45649 19700 45661 19703
rect 45612 19672 45661 19700
rect 45612 19660 45618 19672
rect 45649 19669 45661 19672
rect 45695 19700 45707 19703
rect 46106 19700 46112 19712
rect 45695 19672 46112 19700
rect 45695 19669 45707 19672
rect 45649 19663 45707 19669
rect 46106 19660 46112 19672
rect 46164 19660 46170 19712
rect 46201 19703 46259 19709
rect 46201 19669 46213 19703
rect 46247 19700 46259 19703
rect 46290 19700 46296 19712
rect 46247 19672 46296 19700
rect 46247 19669 46259 19672
rect 46201 19663 46259 19669
rect 46290 19660 46296 19672
rect 46348 19660 46354 19712
rect 47762 19700 47768 19712
rect 47723 19672 47768 19700
rect 47762 19660 47768 19672
rect 47820 19660 47826 19712
rect 47964 19700 47992 19808
rect 51046 19768 51074 19876
rect 58158 19836 58164 19848
rect 58119 19808 58164 19836
rect 58158 19796 58164 19808
rect 58216 19796 58222 19848
rect 57885 19771 57943 19777
rect 57885 19768 57897 19771
rect 51046 19740 57897 19768
rect 57885 19737 57897 19740
rect 57931 19737 57943 19771
rect 57885 19731 57943 19737
rect 51718 19700 51724 19712
rect 47964 19672 51724 19700
rect 51718 19660 51724 19672
rect 51776 19660 51782 19712
rect 1104 19610 58880 19632
rect 1104 19558 20214 19610
rect 20266 19558 20278 19610
rect 20330 19558 20342 19610
rect 20394 19558 20406 19610
rect 20458 19558 20470 19610
rect 20522 19558 39478 19610
rect 39530 19558 39542 19610
rect 39594 19558 39606 19610
rect 39658 19558 39670 19610
rect 39722 19558 39734 19610
rect 39786 19558 58880 19610
rect 1104 19536 58880 19558
rect 12066 19496 12072 19508
rect 12027 19468 12072 19496
rect 12066 19456 12072 19468
rect 12124 19456 12130 19508
rect 16117 19499 16175 19505
rect 16117 19465 16129 19499
rect 16163 19496 16175 19499
rect 20714 19496 20720 19508
rect 16163 19468 19932 19496
rect 20675 19468 20720 19496
rect 16163 19465 16175 19468
rect 16117 19459 16175 19465
rect 17313 19431 17371 19437
rect 17313 19397 17325 19431
rect 17359 19428 17371 19431
rect 17359 19400 18184 19428
rect 17359 19397 17371 19400
rect 17313 19391 17371 19397
rect 12253 19363 12311 19369
rect 12253 19329 12265 19363
rect 12299 19329 12311 19363
rect 17770 19360 17776 19372
rect 17731 19332 17776 19360
rect 12253 19323 12311 19329
rect 12268 19292 12296 19323
rect 17770 19320 17776 19332
rect 17828 19320 17834 19372
rect 18156 19360 18184 19400
rect 18230 19388 18236 19440
rect 18288 19428 18294 19440
rect 18509 19431 18567 19437
rect 18509 19428 18521 19431
rect 18288 19400 18521 19428
rect 18288 19388 18294 19400
rect 18509 19397 18521 19400
rect 18555 19397 18567 19431
rect 19426 19428 19432 19440
rect 18509 19391 18567 19397
rect 18800 19400 19432 19428
rect 18156 19332 18276 19360
rect 12342 19292 12348 19304
rect 12268 19264 12348 19292
rect 12342 19252 12348 19264
rect 12400 19292 12406 19304
rect 12713 19295 12771 19301
rect 12713 19292 12725 19295
rect 12400 19264 12725 19292
rect 12400 19252 12406 19264
rect 12713 19261 12725 19264
rect 12759 19261 12771 19295
rect 12713 19255 12771 19261
rect 13541 19295 13599 19301
rect 13541 19261 13553 19295
rect 13587 19292 13599 19295
rect 15194 19292 15200 19304
rect 13587 19264 15200 19292
rect 13587 19261 13599 19264
rect 13541 19255 13599 19261
rect 15194 19252 15200 19264
rect 15252 19252 15258 19304
rect 15565 19295 15623 19301
rect 15565 19261 15577 19295
rect 15611 19292 15623 19295
rect 17218 19292 17224 19304
rect 15611 19264 17224 19292
rect 15611 19261 15623 19264
rect 15565 19255 15623 19261
rect 17218 19252 17224 19264
rect 17276 19252 17282 19304
rect 17954 19292 17960 19304
rect 17696 19264 17960 19292
rect 14461 19227 14519 19233
rect 14461 19193 14473 19227
rect 14507 19224 14519 19227
rect 16758 19224 16764 19236
rect 14507 19196 16620 19224
rect 16719 19196 16764 19224
rect 14507 19193 14519 19196
rect 14461 19187 14519 19193
rect 15010 19156 15016 19168
rect 14971 19128 15016 19156
rect 15010 19116 15016 19128
rect 15068 19116 15074 19168
rect 16592 19156 16620 19196
rect 16758 19184 16764 19196
rect 16816 19184 16822 19236
rect 17696 19156 17724 19264
rect 17954 19252 17960 19264
rect 18012 19252 18018 19304
rect 18248 19292 18276 19332
rect 18322 19320 18328 19372
rect 18380 19360 18386 19372
rect 18417 19363 18475 19369
rect 18417 19360 18429 19363
rect 18380 19332 18429 19360
rect 18380 19320 18386 19332
rect 18417 19329 18429 19332
rect 18463 19329 18475 19363
rect 18417 19323 18475 19329
rect 18800 19292 18828 19400
rect 19426 19388 19432 19400
rect 19484 19388 19490 19440
rect 18874 19320 18880 19372
rect 18932 19360 18938 19372
rect 19053 19363 19111 19369
rect 19053 19360 19065 19363
rect 18932 19332 19065 19360
rect 18932 19320 18938 19332
rect 19053 19329 19065 19332
rect 19099 19329 19111 19363
rect 19053 19323 19111 19329
rect 19518 19320 19524 19372
rect 19576 19360 19582 19372
rect 19904 19369 19932 19468
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 20898 19496 20904 19508
rect 20859 19468 20904 19496
rect 20898 19456 20904 19468
rect 20956 19456 20962 19508
rect 20993 19499 21051 19505
rect 20993 19465 21005 19499
rect 21039 19496 21051 19499
rect 21450 19496 21456 19508
rect 21039 19468 21456 19496
rect 21039 19465 21051 19468
rect 20993 19459 21051 19465
rect 21450 19456 21456 19468
rect 21508 19456 21514 19508
rect 22186 19456 22192 19508
rect 22244 19496 22250 19508
rect 22281 19499 22339 19505
rect 22281 19496 22293 19499
rect 22244 19468 22293 19496
rect 22244 19456 22250 19468
rect 22281 19465 22293 19468
rect 22327 19465 22339 19499
rect 22281 19459 22339 19465
rect 22557 19499 22615 19505
rect 22557 19465 22569 19499
rect 22603 19496 22615 19499
rect 23198 19496 23204 19508
rect 22603 19468 23204 19496
rect 22603 19465 22615 19468
rect 22557 19459 22615 19465
rect 23198 19456 23204 19468
rect 23256 19456 23262 19508
rect 23658 19456 23664 19508
rect 23716 19496 23722 19508
rect 25590 19496 25596 19508
rect 23716 19468 25596 19496
rect 23716 19456 23722 19468
rect 19978 19388 19984 19440
rect 20036 19428 20042 19440
rect 20438 19428 20444 19440
rect 20036 19400 20444 19428
rect 20036 19388 20042 19400
rect 20438 19388 20444 19400
rect 20496 19388 20502 19440
rect 20640 19400 23704 19428
rect 19889 19363 19947 19369
rect 19889 19360 19901 19363
rect 19576 19332 19901 19360
rect 19576 19320 19582 19332
rect 19889 19329 19901 19332
rect 19935 19329 19947 19363
rect 19889 19323 19947 19329
rect 19150 19292 19156 19304
rect 18248 19264 18828 19292
rect 19111 19264 19156 19292
rect 19150 19252 19156 19264
rect 19208 19252 19214 19304
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 19794 19292 19800 19304
rect 19392 19264 19800 19292
rect 19392 19252 19398 19264
rect 19794 19252 19800 19264
rect 19852 19252 19858 19304
rect 19981 19295 20039 19301
rect 19981 19261 19993 19295
rect 20027 19292 20039 19295
rect 20346 19292 20352 19304
rect 20027 19264 20352 19292
rect 20027 19261 20039 19264
rect 19981 19255 20039 19261
rect 20346 19252 20352 19264
rect 20404 19252 20410 19304
rect 20640 19292 20668 19400
rect 20898 19320 20904 19372
rect 20956 19360 20962 19372
rect 21085 19363 21143 19369
rect 21085 19360 21097 19363
rect 20956 19332 21097 19360
rect 20956 19320 20962 19332
rect 21085 19329 21097 19332
rect 21131 19360 21143 19363
rect 21726 19360 21732 19372
rect 21131 19332 21732 19360
rect 21131 19329 21143 19332
rect 21085 19323 21143 19329
rect 21726 19320 21732 19332
rect 21784 19320 21790 19372
rect 22186 19360 22192 19372
rect 22147 19332 22192 19360
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 22370 19320 22376 19372
rect 22428 19369 22434 19372
rect 22428 19363 22456 19369
rect 22444 19329 22456 19363
rect 22428 19323 22456 19329
rect 22428 19320 22434 19323
rect 22646 19320 22652 19372
rect 22704 19360 22710 19372
rect 22704 19332 22876 19360
rect 22704 19320 22710 19332
rect 20456 19264 20668 19292
rect 21913 19295 21971 19301
rect 17865 19227 17923 19233
rect 17865 19193 17877 19227
rect 17911 19224 17923 19227
rect 20456 19224 20484 19264
rect 21913 19261 21925 19295
rect 21959 19292 21971 19295
rect 22848 19292 22876 19332
rect 22922 19320 22928 19372
rect 22980 19360 22986 19372
rect 23293 19363 23351 19369
rect 23293 19360 23305 19363
rect 22980 19332 23305 19360
rect 22980 19320 22986 19332
rect 23293 19329 23305 19332
rect 23339 19329 23351 19363
rect 23293 19323 23351 19329
rect 23017 19295 23075 19301
rect 23017 19292 23029 19295
rect 21959 19264 22232 19292
rect 22848 19264 23029 19292
rect 21959 19261 21971 19264
rect 21913 19255 21971 19261
rect 22204 19236 22232 19264
rect 23017 19261 23029 19264
rect 23063 19261 23075 19295
rect 23676 19292 23704 19400
rect 23952 19369 23980 19468
rect 25590 19456 25596 19468
rect 25648 19456 25654 19508
rect 25958 19456 25964 19508
rect 26016 19496 26022 19508
rect 26421 19499 26479 19505
rect 26421 19496 26433 19499
rect 26016 19468 26433 19496
rect 26016 19456 26022 19468
rect 26421 19465 26433 19468
rect 26467 19465 26479 19499
rect 26421 19459 26479 19465
rect 27065 19499 27123 19505
rect 27065 19465 27077 19499
rect 27111 19496 27123 19499
rect 30190 19496 30196 19508
rect 27111 19468 30196 19496
rect 27111 19465 27123 19468
rect 27065 19459 27123 19465
rect 30190 19456 30196 19468
rect 30248 19456 30254 19508
rect 36630 19496 36636 19508
rect 31726 19468 36636 19496
rect 24044 19400 25438 19428
rect 23937 19363 23995 19369
rect 23937 19329 23949 19363
rect 23983 19329 23995 19363
rect 23937 19323 23995 19329
rect 24044 19292 24072 19400
rect 26234 19388 26240 19440
rect 26292 19428 26298 19440
rect 29730 19428 29736 19440
rect 26292 19400 28290 19428
rect 29691 19400 29736 19428
rect 26292 19388 26298 19400
rect 29730 19388 29736 19400
rect 29788 19388 29794 19440
rect 31389 19431 31447 19437
rect 31389 19397 31401 19431
rect 31435 19428 31447 19431
rect 31726 19428 31754 19468
rect 36630 19456 36636 19468
rect 36688 19456 36694 19508
rect 38286 19496 38292 19508
rect 37292 19468 38292 19496
rect 31435 19400 31754 19428
rect 33781 19431 33839 19437
rect 31435 19397 31447 19400
rect 31389 19391 31447 19397
rect 33781 19397 33793 19431
rect 33827 19428 33839 19431
rect 34606 19428 34612 19440
rect 33827 19400 34612 19428
rect 33827 19397 33839 19400
rect 33781 19391 33839 19397
rect 34606 19388 34612 19400
rect 34664 19388 34670 19440
rect 35434 19388 35440 19440
rect 35492 19388 35498 19440
rect 35894 19388 35900 19440
rect 35952 19428 35958 19440
rect 35952 19400 36216 19428
rect 35952 19388 35958 19400
rect 24210 19360 24216 19372
rect 24171 19332 24216 19360
rect 24210 19320 24216 19332
rect 24268 19320 24274 19372
rect 24486 19320 24492 19372
rect 24544 19360 24550 19372
rect 24673 19363 24731 19369
rect 24673 19360 24685 19363
rect 24544 19332 24685 19360
rect 24544 19320 24550 19332
rect 24673 19329 24685 19332
rect 24719 19329 24731 19363
rect 24673 19323 24731 19329
rect 27430 19320 27436 19372
rect 27488 19360 27494 19372
rect 27525 19363 27583 19369
rect 27525 19360 27537 19363
rect 27488 19332 27537 19360
rect 27488 19320 27494 19332
rect 27525 19329 27537 19332
rect 27571 19329 27583 19363
rect 27525 19323 27583 19329
rect 29270 19320 29276 19372
rect 29328 19360 29334 19372
rect 29454 19360 29460 19372
rect 29328 19332 29460 19360
rect 29328 19320 29334 19332
rect 29454 19320 29460 19332
rect 29512 19320 29518 19372
rect 31570 19320 31576 19372
rect 31628 19360 31634 19372
rect 33965 19363 34023 19369
rect 31628 19332 31673 19360
rect 31628 19320 31634 19332
rect 33965 19329 33977 19363
rect 34011 19360 34023 19363
rect 34514 19360 34520 19372
rect 34011 19332 34520 19360
rect 34011 19329 34023 19332
rect 33965 19323 34023 19329
rect 34514 19320 34520 19332
rect 34572 19320 34578 19372
rect 36188 19369 36216 19400
rect 37292 19369 37320 19468
rect 38286 19456 38292 19468
rect 38344 19456 38350 19508
rect 39025 19499 39083 19505
rect 39025 19465 39037 19499
rect 39071 19496 39083 19499
rect 39298 19496 39304 19508
rect 39071 19468 39304 19496
rect 39071 19465 39083 19468
rect 39025 19459 39083 19465
rect 39298 19456 39304 19468
rect 39356 19456 39362 19508
rect 46474 19496 46480 19508
rect 40052 19468 46480 19496
rect 37550 19428 37556 19440
rect 37511 19400 37556 19428
rect 37550 19388 37556 19400
rect 37608 19388 37614 19440
rect 40052 19428 40080 19468
rect 46474 19456 46480 19468
rect 46532 19456 46538 19508
rect 46658 19496 46664 19508
rect 46619 19468 46664 19496
rect 46658 19456 46664 19468
rect 46716 19456 46722 19508
rect 58158 19496 58164 19508
rect 58119 19468 58164 19496
rect 58158 19456 58164 19468
rect 58216 19456 58222 19508
rect 38778 19400 40080 19428
rect 40402 19388 40408 19440
rect 40460 19428 40466 19440
rect 40862 19428 40868 19440
rect 40460 19400 40868 19428
rect 40460 19388 40466 19400
rect 40862 19388 40868 19400
rect 40920 19388 40926 19440
rect 41230 19388 41236 19440
rect 41288 19428 41294 19440
rect 43901 19431 43959 19437
rect 43901 19428 43913 19431
rect 41288 19400 43913 19428
rect 41288 19388 41294 19400
rect 43901 19397 43913 19400
rect 43947 19397 43959 19431
rect 43901 19391 43959 19397
rect 44082 19388 44088 19440
rect 44140 19428 44146 19440
rect 48866 19428 48872 19440
rect 44140 19400 48872 19428
rect 44140 19388 44146 19400
rect 48866 19388 48872 19400
rect 48924 19388 48930 19440
rect 36173 19363 36231 19369
rect 36173 19329 36185 19363
rect 36219 19329 36231 19363
rect 36173 19323 36231 19329
rect 37277 19363 37335 19369
rect 37277 19329 37289 19363
rect 37323 19329 37335 19363
rect 37277 19323 37335 19329
rect 39298 19320 39304 19372
rect 39356 19360 39362 19372
rect 39853 19363 39911 19369
rect 39853 19360 39865 19363
rect 39356 19332 39865 19360
rect 39356 19320 39362 19332
rect 39853 19329 39865 19332
rect 39899 19329 39911 19363
rect 40126 19360 40132 19372
rect 40087 19332 40132 19360
rect 39853 19323 39911 19329
rect 40126 19320 40132 19332
rect 40184 19320 40190 19372
rect 40880 19360 40908 19388
rect 41509 19363 41567 19369
rect 41509 19360 41521 19363
rect 40880 19332 41521 19360
rect 41509 19329 41521 19332
rect 41555 19329 41567 19363
rect 42702 19360 42708 19372
rect 42663 19332 42708 19360
rect 41509 19323 41567 19329
rect 42702 19320 42708 19332
rect 42760 19320 42766 19372
rect 42794 19320 42800 19372
rect 42852 19360 42858 19372
rect 42978 19360 42984 19372
rect 42852 19332 42984 19360
rect 42852 19320 42858 19332
rect 42978 19320 42984 19332
rect 43036 19320 43042 19372
rect 43162 19360 43168 19372
rect 43123 19332 43168 19360
rect 43162 19320 43168 19332
rect 43220 19320 43226 19372
rect 43254 19320 43260 19372
rect 43312 19360 43318 19372
rect 43806 19360 43812 19372
rect 43312 19332 43357 19360
rect 43767 19332 43812 19360
rect 43312 19320 43318 19332
rect 43806 19320 43812 19332
rect 43864 19320 43870 19372
rect 44545 19363 44603 19369
rect 44545 19329 44557 19363
rect 44591 19360 44603 19363
rect 44634 19360 44640 19372
rect 44591 19332 44640 19360
rect 44591 19329 44603 19332
rect 44545 19323 44603 19329
rect 44634 19320 44640 19332
rect 44692 19320 44698 19372
rect 24949 19295 25007 19301
rect 24949 19292 24961 19295
rect 23676 19264 24072 19292
rect 24504 19264 24961 19292
rect 23017 19255 23075 19261
rect 24504 19236 24532 19264
rect 24949 19261 24961 19264
rect 24995 19261 25007 19295
rect 27801 19295 27859 19301
rect 27801 19292 27813 19295
rect 24949 19255 25007 19261
rect 25976 19264 27813 19292
rect 21266 19224 21272 19236
rect 17911 19196 20484 19224
rect 20548 19196 20852 19224
rect 21227 19196 21272 19224
rect 17911 19193 17923 19196
rect 17865 19187 17923 19193
rect 16592 19128 17724 19156
rect 18414 19116 18420 19168
rect 18472 19156 18478 19168
rect 18690 19156 18696 19168
rect 18472 19128 18696 19156
rect 18472 19116 18478 19128
rect 18690 19116 18696 19128
rect 18748 19116 18754 19168
rect 19150 19116 19156 19168
rect 19208 19156 19214 19168
rect 20165 19159 20223 19165
rect 20165 19156 20177 19159
rect 19208 19128 20177 19156
rect 19208 19116 19214 19128
rect 20165 19125 20177 19128
rect 20211 19125 20223 19159
rect 20165 19119 20223 19125
rect 20254 19116 20260 19168
rect 20312 19156 20318 19168
rect 20548 19156 20576 19196
rect 20312 19128 20576 19156
rect 20824 19156 20852 19196
rect 21266 19184 21272 19196
rect 21324 19184 21330 19236
rect 22186 19184 22192 19236
rect 22244 19184 22250 19236
rect 24486 19184 24492 19236
rect 24544 19184 24550 19236
rect 25976 19156 26004 19264
rect 27801 19261 27813 19264
rect 27847 19261 27859 19295
rect 30926 19292 30932 19304
rect 27801 19255 27859 19261
rect 28828 19264 30932 19292
rect 20824 19128 26004 19156
rect 20312 19116 20318 19128
rect 26050 19116 26056 19168
rect 26108 19156 26114 19168
rect 28828 19156 28856 19264
rect 30926 19252 30932 19264
rect 30984 19252 30990 19304
rect 32306 19252 32312 19304
rect 32364 19292 32370 19304
rect 33410 19292 33416 19304
rect 32364 19264 33416 19292
rect 32364 19252 32370 19264
rect 33410 19252 33416 19264
rect 33468 19252 33474 19304
rect 35802 19252 35808 19304
rect 35860 19292 35866 19304
rect 35897 19295 35955 19301
rect 35897 19292 35909 19295
rect 35860 19264 35909 19292
rect 35860 19252 35866 19264
rect 35897 19261 35909 19264
rect 35943 19292 35955 19295
rect 35943 19264 36124 19292
rect 35943 19261 35955 19264
rect 35897 19255 35955 19261
rect 28994 19184 29000 19236
rect 29052 19224 29058 19236
rect 36096 19224 36124 19264
rect 36538 19252 36544 19304
rect 36596 19292 36602 19304
rect 36633 19295 36691 19301
rect 36633 19292 36645 19295
rect 36596 19264 36645 19292
rect 36596 19252 36602 19264
rect 36633 19261 36645 19264
rect 36679 19261 36691 19295
rect 39482 19292 39488 19304
rect 36633 19255 36691 19261
rect 37384 19264 38608 19292
rect 39443 19264 39488 19292
rect 37384 19224 37412 19264
rect 29052 19196 34744 19224
rect 36096 19196 37412 19224
rect 38580 19224 38608 19264
rect 39482 19252 39488 19264
rect 39540 19252 39546 19304
rect 39574 19252 39580 19304
rect 39632 19292 39638 19304
rect 48133 19295 48191 19301
rect 48133 19292 48145 19295
rect 39632 19264 48145 19292
rect 39632 19252 39638 19264
rect 48133 19261 48145 19264
rect 48179 19261 48191 19295
rect 48682 19292 48688 19304
rect 48643 19264 48688 19292
rect 48133 19255 48191 19261
rect 48682 19252 48688 19264
rect 48740 19252 48746 19304
rect 41138 19224 41144 19236
rect 38580 19196 41144 19224
rect 29052 19184 29058 19196
rect 29270 19156 29276 19168
rect 26108 19128 28856 19156
rect 29231 19128 29276 19156
rect 26108 19116 26114 19128
rect 29270 19116 29276 19128
rect 29328 19116 29334 19168
rect 29454 19116 29460 19168
rect 29512 19156 29518 19168
rect 30282 19156 30288 19168
rect 29512 19128 30288 19156
rect 29512 19116 29518 19128
rect 30282 19116 30288 19128
rect 30340 19116 30346 19168
rect 30374 19116 30380 19168
rect 30432 19156 30438 19168
rect 34146 19156 34152 19168
rect 30432 19128 34152 19156
rect 30432 19116 30438 19128
rect 34146 19116 34152 19128
rect 34204 19116 34210 19168
rect 34425 19159 34483 19165
rect 34425 19125 34437 19159
rect 34471 19156 34483 19159
rect 34606 19156 34612 19168
rect 34471 19128 34612 19156
rect 34471 19125 34483 19128
rect 34425 19119 34483 19125
rect 34606 19116 34612 19128
rect 34664 19116 34670 19168
rect 34716 19156 34744 19196
rect 41138 19184 41144 19196
rect 41196 19184 41202 19236
rect 41874 19184 41880 19236
rect 41932 19224 41938 19236
rect 42521 19227 42579 19233
rect 42521 19224 42533 19227
rect 41932 19196 42533 19224
rect 41932 19184 41938 19196
rect 42521 19193 42533 19196
rect 42567 19193 42579 19227
rect 42521 19187 42579 19193
rect 42794 19184 42800 19236
rect 42852 19224 42858 19236
rect 45557 19227 45615 19233
rect 45557 19224 45569 19227
rect 42852 19196 45569 19224
rect 42852 19184 42858 19196
rect 45557 19193 45569 19196
rect 45603 19193 45615 19227
rect 45557 19187 45615 19193
rect 47673 19227 47731 19233
rect 47673 19193 47685 19227
rect 47719 19224 47731 19227
rect 49694 19224 49700 19236
rect 47719 19196 49700 19224
rect 47719 19193 47731 19196
rect 47673 19187 47731 19193
rect 49694 19184 49700 19196
rect 49752 19184 49758 19236
rect 36538 19156 36544 19168
rect 34716 19128 36544 19156
rect 36538 19116 36544 19128
rect 36596 19116 36602 19168
rect 36722 19116 36728 19168
rect 36780 19156 36786 19168
rect 39390 19156 39396 19168
rect 36780 19128 39396 19156
rect 36780 19116 36786 19128
rect 39390 19116 39396 19128
rect 39448 19116 39454 19168
rect 40954 19116 40960 19168
rect 41012 19156 41018 19168
rect 41049 19159 41107 19165
rect 41049 19156 41061 19159
rect 41012 19128 41061 19156
rect 41012 19116 41018 19128
rect 41049 19125 41061 19128
rect 41095 19125 41107 19159
rect 41049 19119 41107 19125
rect 41782 19116 41788 19168
rect 41840 19156 41846 19168
rect 42978 19156 42984 19168
rect 41840 19128 42984 19156
rect 41840 19116 41846 19128
rect 42978 19116 42984 19128
rect 43036 19116 43042 19168
rect 43622 19116 43628 19168
rect 43680 19156 43686 19168
rect 45005 19159 45063 19165
rect 45005 19156 45017 19159
rect 43680 19128 45017 19156
rect 43680 19116 43686 19128
rect 45005 19125 45017 19128
rect 45051 19125 45063 19159
rect 46198 19156 46204 19168
rect 46159 19128 46204 19156
rect 45005 19119 45063 19125
rect 46198 19116 46204 19128
rect 46256 19116 46262 19168
rect 1104 19066 58880 19088
rect 1104 19014 10582 19066
rect 10634 19014 10646 19066
rect 10698 19014 10710 19066
rect 10762 19014 10774 19066
rect 10826 19014 10838 19066
rect 10890 19014 29846 19066
rect 29898 19014 29910 19066
rect 29962 19014 29974 19066
rect 30026 19014 30038 19066
rect 30090 19014 30102 19066
rect 30154 19014 49110 19066
rect 49162 19014 49174 19066
rect 49226 19014 49238 19066
rect 49290 19014 49302 19066
rect 49354 19014 49366 19066
rect 49418 19014 58880 19066
rect 1104 18992 58880 19014
rect 12250 18912 12256 18964
rect 12308 18952 12314 18964
rect 12437 18955 12495 18961
rect 12437 18952 12449 18955
rect 12308 18924 12449 18952
rect 12308 18912 12314 18924
rect 12437 18921 12449 18924
rect 12483 18952 12495 18955
rect 12989 18955 13047 18961
rect 12989 18952 13001 18955
rect 12483 18924 13001 18952
rect 12483 18921 12495 18924
rect 12437 18915 12495 18921
rect 12989 18921 13001 18924
rect 13035 18952 13047 18955
rect 15746 18952 15752 18964
rect 13035 18924 15752 18952
rect 13035 18921 13047 18924
rect 12989 18915 13047 18921
rect 15746 18912 15752 18924
rect 15804 18912 15810 18964
rect 16114 18912 16120 18964
rect 16172 18952 16178 18964
rect 17126 18952 17132 18964
rect 16172 18924 17132 18952
rect 16172 18912 16178 18924
rect 17126 18912 17132 18924
rect 17184 18912 17190 18964
rect 17586 18912 17592 18964
rect 17644 18952 17650 18964
rect 20254 18952 20260 18964
rect 17644 18924 17689 18952
rect 18708 18924 20260 18952
rect 17644 18912 17650 18924
rect 14737 18887 14795 18893
rect 14737 18853 14749 18887
rect 14783 18884 14795 18887
rect 16482 18884 16488 18896
rect 14783 18856 16488 18884
rect 14783 18853 14795 18856
rect 14737 18847 14795 18853
rect 16482 18844 16488 18856
rect 16540 18844 16546 18896
rect 17034 18844 17040 18896
rect 17092 18884 17098 18896
rect 18046 18884 18052 18896
rect 17092 18856 18052 18884
rect 17092 18844 17098 18856
rect 18046 18844 18052 18856
rect 18104 18844 18110 18896
rect 14182 18816 14188 18828
rect 14143 18788 14188 18816
rect 14182 18776 14188 18788
rect 14240 18776 14246 18828
rect 14550 18776 14556 18828
rect 14608 18816 14614 18828
rect 15654 18816 15660 18828
rect 14608 18788 15660 18816
rect 14608 18776 14614 18788
rect 15654 18776 15660 18788
rect 15712 18776 15718 18828
rect 17310 18776 17316 18828
rect 17368 18776 17374 18828
rect 17402 18776 17408 18828
rect 17460 18816 17466 18828
rect 17586 18816 17592 18828
rect 17460 18788 17592 18816
rect 17460 18776 17466 18788
rect 17586 18776 17592 18788
rect 17644 18776 17650 18828
rect 18417 18819 18475 18825
rect 18417 18816 18429 18819
rect 17696 18788 18429 18816
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18748 13599 18751
rect 14568 18748 14596 18776
rect 13587 18720 14596 18748
rect 13587 18717 13599 18720
rect 13541 18711 13599 18717
rect 16574 18708 16580 18760
rect 16632 18748 16638 18760
rect 16853 18751 16911 18757
rect 16853 18748 16865 18751
rect 16632 18720 16865 18748
rect 16632 18708 16638 18720
rect 16853 18717 16865 18720
rect 16899 18717 16911 18751
rect 17328 18748 17356 18776
rect 17505 18751 17563 18757
rect 17505 18748 17517 18751
rect 17328 18720 17517 18748
rect 16853 18711 16911 18717
rect 17505 18717 17517 18720
rect 17551 18717 17563 18751
rect 17505 18711 17563 18717
rect 15197 18683 15255 18689
rect 15197 18649 15209 18683
rect 15243 18680 15255 18683
rect 15243 18652 17356 18680
rect 15243 18649 15255 18652
rect 15197 18643 15255 18649
rect 15470 18572 15476 18624
rect 15528 18612 15534 18624
rect 15749 18615 15807 18621
rect 15749 18612 15761 18615
rect 15528 18584 15761 18612
rect 15528 18572 15534 18584
rect 15749 18581 15761 18584
rect 15795 18581 15807 18615
rect 16298 18612 16304 18624
rect 16259 18584 16304 18612
rect 15749 18575 15807 18581
rect 16298 18572 16304 18584
rect 16356 18572 16362 18624
rect 16942 18572 16948 18624
rect 17000 18612 17006 18624
rect 17328 18612 17356 18652
rect 17402 18640 17408 18692
rect 17460 18680 17466 18692
rect 17696 18680 17724 18788
rect 18417 18785 18429 18788
rect 18463 18816 18475 18819
rect 18708 18816 18736 18924
rect 20254 18912 20260 18924
rect 20312 18912 20318 18964
rect 20438 18952 20444 18964
rect 20399 18924 20444 18952
rect 20438 18912 20444 18924
rect 20496 18912 20502 18964
rect 20530 18912 20536 18964
rect 20588 18952 20594 18964
rect 26050 18952 26056 18964
rect 20588 18924 26056 18952
rect 20588 18912 20594 18924
rect 26050 18912 26056 18924
rect 26108 18912 26114 18964
rect 26789 18955 26847 18961
rect 26789 18921 26801 18955
rect 26835 18952 26847 18955
rect 28994 18952 29000 18964
rect 26835 18924 28580 18952
rect 28955 18924 29000 18952
rect 26835 18921 26847 18924
rect 26789 18915 26847 18921
rect 19242 18844 19248 18896
rect 19300 18884 19306 18896
rect 19886 18884 19892 18896
rect 19300 18856 19892 18884
rect 19300 18844 19306 18856
rect 19886 18844 19892 18856
rect 19944 18844 19950 18896
rect 21266 18844 21272 18896
rect 21324 18884 21330 18896
rect 22002 18884 22008 18896
rect 21324 18856 22008 18884
rect 21324 18844 21330 18856
rect 22002 18844 22008 18856
rect 22060 18844 22066 18896
rect 28552 18884 28580 18924
rect 28994 18912 29000 18924
rect 29052 18912 29058 18964
rect 33686 18952 33692 18964
rect 29288 18924 33692 18952
rect 29288 18884 29316 18924
rect 33686 18912 33692 18924
rect 33744 18912 33750 18964
rect 41601 18955 41659 18961
rect 34532 18924 41414 18952
rect 28552 18856 29316 18884
rect 31202 18844 31208 18896
rect 31260 18884 31266 18896
rect 34422 18884 34428 18896
rect 31260 18856 34428 18884
rect 31260 18844 31266 18856
rect 34422 18844 34428 18856
rect 34480 18844 34486 18896
rect 18463 18788 18736 18816
rect 18463 18785 18475 18788
rect 18417 18779 18475 18785
rect 19978 18776 19984 18828
rect 20036 18816 20042 18828
rect 20073 18819 20131 18825
rect 20073 18816 20085 18819
rect 20036 18788 20085 18816
rect 20036 18776 20042 18788
rect 20073 18785 20085 18788
rect 20119 18785 20131 18819
rect 20898 18816 20904 18828
rect 20073 18779 20131 18785
rect 20364 18788 20904 18816
rect 20364 18760 20392 18788
rect 20898 18776 20904 18788
rect 20956 18776 20962 18828
rect 21082 18776 21088 18828
rect 21140 18816 21146 18828
rect 21177 18819 21235 18825
rect 21177 18816 21189 18819
rect 21140 18788 21189 18816
rect 21140 18776 21146 18788
rect 21177 18785 21189 18788
rect 21223 18785 21235 18819
rect 21177 18779 21235 18785
rect 21358 18776 21364 18828
rect 21416 18816 21422 18828
rect 21637 18819 21695 18825
rect 21637 18816 21649 18819
rect 21416 18788 21649 18816
rect 21416 18776 21422 18788
rect 21637 18785 21649 18788
rect 21683 18785 21695 18819
rect 21637 18779 21695 18785
rect 21726 18776 21732 18828
rect 21784 18816 21790 18828
rect 21910 18816 21916 18828
rect 21784 18788 21916 18816
rect 21784 18776 21790 18788
rect 21910 18776 21916 18788
rect 21968 18776 21974 18828
rect 23842 18816 23848 18828
rect 23803 18788 23848 18816
rect 23842 18776 23848 18788
rect 23900 18776 23906 18828
rect 23934 18776 23940 18828
rect 23992 18816 23998 18828
rect 24210 18816 24216 18828
rect 23992 18788 24216 18816
rect 23992 18776 23998 18788
rect 24210 18776 24216 18788
rect 24268 18776 24274 18828
rect 31754 18816 31760 18828
rect 24596 18788 31760 18816
rect 24596 18760 24624 18788
rect 31754 18776 31760 18788
rect 31812 18776 31818 18828
rect 32217 18819 32275 18825
rect 32217 18785 32229 18819
rect 32263 18816 32275 18819
rect 34532 18816 34560 18924
rect 36538 18844 36544 18896
rect 36596 18884 36602 18896
rect 38657 18887 38715 18893
rect 36596 18856 37044 18884
rect 36596 18844 36602 18856
rect 32263 18788 34560 18816
rect 32263 18785 32275 18788
rect 32217 18779 32275 18785
rect 18322 18748 18328 18760
rect 18235 18720 18328 18748
rect 18322 18708 18328 18720
rect 18380 18748 18386 18760
rect 18690 18748 18696 18760
rect 18380 18720 18696 18748
rect 18380 18708 18386 18720
rect 18690 18708 18696 18720
rect 18748 18708 18754 18760
rect 19426 18708 19432 18760
rect 19484 18748 19490 18760
rect 20165 18751 20223 18757
rect 19484 18742 20116 18748
rect 20165 18742 20177 18751
rect 19484 18720 20177 18742
rect 19484 18708 19490 18720
rect 20088 18717 20177 18720
rect 20211 18717 20223 18751
rect 20088 18714 20223 18717
rect 20165 18711 20223 18714
rect 20346 18708 20352 18760
rect 20404 18708 20410 18760
rect 20438 18708 20444 18760
rect 20496 18748 20502 18760
rect 20993 18751 21051 18757
rect 20993 18748 21005 18751
rect 20496 18720 21005 18748
rect 20496 18708 20502 18720
rect 20993 18717 21005 18720
rect 21039 18717 21051 18751
rect 20993 18711 21051 18717
rect 21266 18708 21272 18760
rect 21324 18748 21330 18760
rect 21324 18720 21369 18748
rect 21324 18708 21330 18720
rect 21450 18708 21456 18760
rect 21508 18748 21514 18760
rect 22097 18751 22155 18757
rect 22097 18748 22109 18751
rect 21508 18720 22109 18748
rect 21508 18708 21514 18720
rect 22097 18717 22109 18720
rect 22143 18717 22155 18751
rect 24578 18748 24584 18760
rect 24491 18720 24584 18748
rect 22097 18711 22155 18717
rect 24578 18708 24584 18720
rect 24636 18708 24642 18760
rect 24670 18708 24676 18760
rect 24728 18748 24734 18760
rect 25041 18751 25099 18757
rect 25041 18748 25053 18751
rect 24728 18720 25053 18748
rect 24728 18708 24734 18720
rect 25041 18717 25053 18720
rect 25087 18717 25099 18751
rect 27246 18748 27252 18760
rect 27207 18720 27252 18748
rect 25041 18711 25099 18717
rect 27246 18708 27252 18720
rect 27304 18708 27310 18760
rect 29454 18708 29460 18760
rect 29512 18748 29518 18760
rect 29917 18751 29975 18757
rect 29917 18748 29929 18751
rect 29512 18720 29929 18748
rect 29512 18708 29518 18720
rect 29917 18717 29929 18720
rect 29963 18717 29975 18751
rect 30285 18751 30343 18757
rect 30285 18748 30297 18751
rect 29917 18711 29975 18717
rect 30005 18720 30297 18748
rect 19242 18680 19248 18692
rect 17460 18652 17724 18680
rect 17926 18652 19248 18680
rect 17460 18640 17466 18652
rect 17926 18612 17954 18652
rect 19242 18640 19248 18652
rect 19300 18640 19306 18692
rect 19337 18683 19395 18689
rect 19337 18649 19349 18683
rect 19383 18680 19395 18683
rect 20714 18680 20720 18692
rect 19383 18652 20720 18680
rect 19383 18649 19395 18652
rect 19337 18643 19395 18649
rect 20714 18640 20720 18652
rect 20772 18640 20778 18692
rect 22370 18680 22376 18692
rect 22331 18652 22376 18680
rect 22370 18640 22376 18652
rect 22428 18640 22434 18692
rect 24489 18683 24547 18689
rect 24489 18680 24501 18683
rect 23598 18652 24501 18680
rect 24489 18649 24501 18652
rect 24535 18649 24547 18683
rect 24489 18643 24547 18649
rect 24946 18640 24952 18692
rect 25004 18680 25010 18692
rect 25317 18683 25375 18689
rect 25317 18680 25329 18683
rect 25004 18652 25329 18680
rect 25004 18640 25010 18652
rect 25317 18649 25329 18652
rect 25363 18649 25375 18683
rect 25317 18643 25375 18649
rect 25424 18652 25806 18680
rect 17000 18584 17045 18612
rect 17328 18584 17954 18612
rect 17000 18572 17006 18584
rect 18230 18572 18236 18624
rect 18288 18612 18294 18624
rect 18693 18615 18751 18621
rect 18693 18612 18705 18615
rect 18288 18584 18705 18612
rect 18288 18572 18294 18584
rect 18693 18581 18705 18584
rect 18739 18581 18751 18615
rect 18693 18575 18751 18581
rect 19429 18615 19487 18621
rect 19429 18581 19441 18615
rect 19475 18612 19487 18615
rect 21082 18612 21088 18624
rect 19475 18584 21088 18612
rect 19475 18581 19487 18584
rect 19429 18575 19487 18581
rect 21082 18572 21088 18584
rect 21140 18572 21146 18624
rect 21358 18612 21364 18624
rect 21319 18584 21364 18612
rect 21358 18572 21364 18584
rect 21416 18572 21422 18624
rect 21545 18615 21603 18621
rect 21545 18581 21557 18615
rect 21591 18612 21603 18615
rect 21634 18612 21640 18624
rect 21591 18584 21640 18612
rect 21591 18581 21603 18584
rect 21545 18575 21603 18581
rect 21634 18572 21640 18584
rect 21692 18572 21698 18624
rect 21818 18572 21824 18624
rect 21876 18612 21882 18624
rect 25424 18612 25452 18652
rect 26970 18640 26976 18692
rect 27028 18680 27034 18692
rect 27525 18683 27583 18689
rect 27525 18680 27537 18683
rect 27028 18652 27537 18680
rect 27028 18640 27034 18652
rect 27525 18649 27537 18652
rect 27571 18649 27583 18683
rect 27525 18643 27583 18649
rect 27816 18652 28014 18680
rect 21876 18584 25452 18612
rect 21876 18572 21882 18584
rect 25590 18572 25596 18624
rect 25648 18612 25654 18624
rect 27816 18612 27844 18652
rect 29730 18640 29736 18692
rect 29788 18680 29794 18692
rect 30005 18680 30033 18720
rect 30285 18717 30297 18720
rect 30331 18717 30343 18751
rect 30285 18711 30343 18717
rect 31202 18708 31208 18760
rect 31260 18748 31266 18760
rect 31260 18720 31432 18748
rect 31260 18708 31266 18720
rect 29788 18652 30033 18680
rect 29788 18640 29794 18652
rect 31018 18640 31024 18692
rect 31076 18640 31082 18692
rect 31404 18680 31432 18720
rect 32232 18680 32260 18779
rect 34606 18776 34612 18828
rect 34664 18816 34670 18828
rect 34977 18819 35035 18825
rect 34977 18816 34989 18819
rect 34664 18788 34989 18816
rect 34664 18776 34670 18788
rect 34977 18785 34989 18788
rect 35023 18785 35035 18819
rect 34977 18779 35035 18785
rect 36354 18776 36360 18828
rect 36412 18816 36418 18828
rect 36909 18819 36967 18825
rect 36909 18816 36921 18819
rect 36412 18788 36921 18816
rect 36412 18776 36418 18788
rect 36909 18785 36921 18788
rect 36955 18785 36967 18819
rect 37016 18816 37044 18856
rect 38657 18853 38669 18887
rect 38703 18884 38715 18887
rect 38746 18884 38752 18896
rect 38703 18856 38752 18884
rect 38703 18853 38715 18856
rect 38657 18847 38715 18853
rect 38746 18844 38752 18856
rect 38804 18844 38810 18896
rect 39574 18884 39580 18896
rect 38856 18856 39580 18884
rect 38562 18816 38568 18828
rect 37016 18788 38568 18816
rect 36909 18779 36967 18785
rect 38562 18776 38568 18788
rect 38620 18776 38626 18828
rect 34698 18748 34704 18760
rect 34659 18720 34704 18748
rect 34698 18708 34704 18720
rect 34756 18708 34762 18760
rect 38470 18708 38476 18760
rect 38528 18748 38534 18760
rect 38856 18748 38884 18856
rect 39574 18844 39580 18856
rect 39632 18844 39638 18896
rect 41386 18884 41414 18924
rect 41601 18921 41613 18955
rect 41647 18952 41659 18955
rect 41966 18952 41972 18964
rect 41647 18924 41972 18952
rect 41647 18921 41659 18924
rect 41601 18915 41659 18921
rect 41966 18912 41972 18924
rect 42024 18912 42030 18964
rect 49421 18955 49479 18961
rect 49421 18952 49433 18955
rect 42076 18924 49433 18952
rect 42076 18884 42104 18924
rect 49421 18921 49433 18924
rect 49467 18921 49479 18955
rect 49421 18915 49479 18921
rect 41386 18856 42104 18884
rect 42429 18887 42487 18893
rect 42429 18853 42441 18887
rect 42475 18884 42487 18887
rect 42518 18884 42524 18896
rect 42475 18856 42524 18884
rect 42475 18853 42487 18856
rect 42429 18847 42487 18853
rect 42518 18844 42524 18856
rect 42576 18844 42582 18896
rect 43622 18884 43628 18896
rect 42628 18856 43628 18884
rect 39206 18776 39212 18828
rect 39264 18816 39270 18828
rect 39853 18819 39911 18825
rect 39853 18816 39865 18819
rect 39264 18788 39865 18816
rect 39264 18776 39270 18788
rect 39853 18785 39865 18788
rect 39899 18785 39911 18819
rect 39853 18779 39911 18785
rect 40129 18819 40187 18825
rect 40129 18785 40141 18819
rect 40175 18816 40187 18819
rect 40586 18816 40592 18828
rect 40175 18788 40592 18816
rect 40175 18785 40187 18788
rect 40129 18779 40187 18785
rect 40586 18776 40592 18788
rect 40644 18776 40650 18828
rect 42061 18819 42119 18825
rect 42061 18785 42073 18819
rect 42107 18816 42119 18819
rect 42628 18816 42656 18856
rect 43622 18844 43628 18856
rect 43680 18844 43686 18896
rect 46658 18844 46664 18896
rect 46716 18844 46722 18896
rect 47854 18884 47860 18896
rect 47815 18856 47860 18884
rect 47854 18844 47860 18856
rect 47912 18844 47918 18896
rect 42107 18788 42656 18816
rect 42981 18819 43039 18825
rect 42107 18785 42119 18788
rect 42061 18779 42119 18785
rect 42981 18785 42993 18819
rect 43027 18816 43039 18819
rect 43070 18816 43076 18828
rect 43027 18788 43076 18816
rect 43027 18785 43039 18788
rect 42981 18779 43039 18785
rect 39114 18748 39120 18760
rect 38528 18720 38884 18748
rect 39075 18720 39120 18748
rect 38528 18708 38534 18720
rect 39114 18708 39120 18720
rect 39172 18708 39178 18760
rect 41230 18708 41236 18760
rect 41288 18708 41294 18760
rect 32398 18680 32404 18692
rect 31404 18652 32260 18680
rect 32359 18652 32404 18680
rect 32398 18640 32404 18652
rect 32456 18640 32462 18692
rect 33962 18640 33968 18692
rect 34020 18680 34026 18692
rect 34057 18683 34115 18689
rect 34057 18680 34069 18683
rect 34020 18652 34069 18680
rect 34020 18640 34026 18652
rect 34057 18649 34069 18652
rect 34103 18649 34115 18683
rect 34057 18643 34115 18649
rect 35250 18640 35256 18692
rect 35308 18680 35314 18692
rect 35434 18680 35440 18692
rect 35308 18652 35440 18680
rect 35308 18640 35314 18652
rect 35434 18640 35440 18652
rect 35492 18640 35498 18692
rect 36262 18640 36268 18692
rect 36320 18680 36326 18692
rect 37185 18683 37243 18689
rect 37185 18680 37197 18683
rect 36320 18652 37197 18680
rect 36320 18640 36326 18652
rect 37185 18649 37197 18652
rect 37231 18649 37243 18683
rect 37185 18643 37243 18649
rect 38194 18640 38200 18692
rect 38252 18640 38258 18692
rect 40402 18680 40408 18692
rect 39040 18652 40408 18680
rect 25648 18584 27844 18612
rect 25648 18572 25654 18584
rect 27890 18572 27896 18624
rect 27948 18612 27954 18624
rect 29822 18612 29828 18624
rect 27948 18584 29828 18612
rect 27948 18572 27954 18584
rect 29822 18572 29828 18584
rect 29880 18612 29886 18624
rect 30374 18612 30380 18624
rect 29880 18584 30380 18612
rect 29880 18572 29886 18584
rect 30374 18572 30380 18584
rect 30432 18572 30438 18624
rect 31711 18615 31769 18621
rect 31711 18581 31723 18615
rect 31757 18612 31769 18615
rect 32122 18612 32128 18624
rect 31757 18584 32128 18612
rect 31757 18581 31769 18584
rect 31711 18575 31769 18581
rect 32122 18572 32128 18584
rect 32180 18572 32186 18624
rect 34698 18572 34704 18624
rect 34756 18612 34762 18624
rect 35066 18612 35072 18624
rect 34756 18584 35072 18612
rect 34756 18572 34762 18584
rect 35066 18572 35072 18584
rect 35124 18612 35130 18624
rect 35802 18612 35808 18624
rect 35124 18584 35808 18612
rect 35124 18572 35130 18584
rect 35802 18572 35808 18584
rect 35860 18572 35866 18624
rect 36449 18615 36507 18621
rect 36449 18581 36461 18615
rect 36495 18612 36507 18615
rect 39040 18612 39068 18652
rect 40402 18640 40408 18652
rect 40460 18640 40466 18692
rect 39206 18612 39212 18624
rect 36495 18584 39068 18612
rect 39167 18584 39212 18612
rect 36495 18581 36507 18584
rect 36449 18575 36507 18581
rect 39206 18572 39212 18584
rect 39264 18572 39270 18624
rect 40310 18572 40316 18624
rect 40368 18612 40374 18624
rect 42076 18612 42104 18779
rect 43070 18776 43076 18788
rect 43128 18776 43134 18828
rect 43165 18819 43223 18825
rect 43165 18785 43177 18819
rect 43211 18816 43223 18819
rect 44450 18816 44456 18828
rect 43211 18788 44456 18816
rect 43211 18785 43223 18788
rect 43165 18779 43223 18785
rect 44450 18776 44456 18788
rect 44508 18816 44514 18828
rect 46109 18819 46167 18825
rect 46109 18816 46121 18819
rect 44508 18788 46121 18816
rect 44508 18776 44514 18788
rect 46109 18785 46121 18788
rect 46155 18785 46167 18819
rect 46676 18816 46704 18844
rect 48317 18819 48375 18825
rect 48317 18816 48329 18819
rect 46676 18788 48329 18816
rect 46109 18779 46167 18785
rect 48317 18785 48329 18788
rect 48363 18816 48375 18819
rect 48682 18816 48688 18828
rect 48363 18788 48688 18816
rect 48363 18785 48375 18788
rect 48317 18779 48375 18785
rect 48682 18776 48688 18788
rect 48740 18816 48746 18828
rect 48869 18819 48927 18825
rect 48869 18816 48881 18819
rect 48740 18788 48881 18816
rect 48740 18776 48746 18788
rect 48869 18785 48881 18788
rect 48915 18785 48927 18819
rect 48869 18779 48927 18785
rect 43254 18748 43260 18760
rect 42812 18720 43260 18748
rect 40368 18584 42104 18612
rect 42521 18615 42579 18621
rect 40368 18572 40374 18584
rect 42521 18581 42533 18615
rect 42567 18612 42579 18615
rect 42812 18612 42840 18720
rect 43254 18708 43260 18720
rect 43312 18708 43318 18760
rect 43714 18748 43720 18760
rect 43675 18720 43720 18748
rect 43714 18708 43720 18720
rect 43772 18708 43778 18760
rect 46661 18751 46719 18757
rect 46661 18748 46673 18751
rect 44100 18720 46673 18748
rect 42886 18640 42892 18692
rect 42944 18680 42950 18692
rect 44100 18680 44128 18720
rect 46661 18717 46673 18720
rect 46707 18717 46719 18751
rect 58158 18748 58164 18760
rect 58119 18720 58164 18748
rect 46661 18711 46719 18717
rect 58158 18708 58164 18720
rect 58216 18708 58222 18760
rect 42944 18652 44128 18680
rect 42944 18640 42950 18652
rect 46290 18640 46296 18692
rect 46348 18680 46354 18692
rect 47213 18683 47271 18689
rect 47213 18680 47225 18683
rect 46348 18652 47225 18680
rect 46348 18640 46354 18652
rect 47213 18649 47225 18652
rect 47259 18649 47271 18683
rect 57882 18680 57888 18692
rect 57843 18652 57888 18680
rect 47213 18643 47271 18649
rect 57882 18640 57888 18652
rect 57940 18640 57946 18692
rect 42978 18612 42984 18624
rect 42567 18584 42840 18612
rect 42939 18584 42984 18612
rect 42567 18581 42579 18584
rect 42521 18575 42579 18581
rect 42978 18572 42984 18584
rect 43036 18572 43042 18624
rect 43070 18572 43076 18624
rect 43128 18612 43134 18624
rect 43622 18612 43628 18624
rect 43128 18584 43628 18612
rect 43128 18572 43134 18584
rect 43622 18572 43628 18584
rect 43680 18572 43686 18624
rect 43806 18612 43812 18624
rect 43767 18584 43812 18612
rect 43806 18572 43812 18584
rect 43864 18572 43870 18624
rect 44453 18615 44511 18621
rect 44453 18581 44465 18615
rect 44499 18612 44511 18615
rect 44542 18612 44548 18624
rect 44499 18584 44548 18612
rect 44499 18581 44511 18584
rect 44453 18575 44511 18581
rect 44542 18572 44548 18584
rect 44600 18572 44606 18624
rect 45097 18615 45155 18621
rect 45097 18581 45109 18615
rect 45143 18612 45155 18615
rect 45186 18612 45192 18624
rect 45143 18584 45192 18612
rect 45143 18581 45155 18584
rect 45097 18575 45155 18581
rect 45186 18572 45192 18584
rect 45244 18572 45250 18624
rect 45646 18612 45652 18624
rect 45607 18584 45652 18612
rect 45646 18572 45652 18584
rect 45704 18572 45710 18624
rect 1104 18522 58880 18544
rect 1104 18470 20214 18522
rect 20266 18470 20278 18522
rect 20330 18470 20342 18522
rect 20394 18470 20406 18522
rect 20458 18470 20470 18522
rect 20522 18470 39478 18522
rect 39530 18470 39542 18522
rect 39594 18470 39606 18522
rect 39658 18470 39670 18522
rect 39722 18470 39734 18522
rect 39786 18470 58880 18522
rect 1104 18448 58880 18470
rect 13173 18411 13231 18417
rect 13173 18408 13185 18411
rect 2746 18380 13185 18408
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18272 1731 18275
rect 2746 18272 2774 18380
rect 13173 18377 13185 18380
rect 13219 18377 13231 18411
rect 17589 18411 17647 18417
rect 17589 18408 17601 18411
rect 13173 18371 13231 18377
rect 17236 18380 17601 18408
rect 12710 18340 12716 18352
rect 12671 18312 12716 18340
rect 12710 18300 12716 18312
rect 12768 18300 12774 18352
rect 13909 18343 13967 18349
rect 13909 18309 13921 18343
rect 13955 18340 13967 18343
rect 13955 18312 16712 18340
rect 13955 18309 13967 18312
rect 13909 18303 13967 18309
rect 16684 18284 16712 18312
rect 1719 18244 2774 18272
rect 13357 18275 13415 18281
rect 1719 18241 1731 18244
rect 1673 18235 1731 18241
rect 13357 18241 13369 18275
rect 13403 18272 13415 18275
rect 15194 18272 15200 18284
rect 13403 18244 15200 18272
rect 13403 18241 13415 18244
rect 13357 18235 13415 18241
rect 15194 18232 15200 18244
rect 15252 18232 15258 18284
rect 16666 18272 16672 18284
rect 16627 18244 16672 18272
rect 16666 18232 16672 18244
rect 16724 18232 16730 18284
rect 17236 18204 17264 18380
rect 17589 18377 17601 18380
rect 17635 18377 17647 18411
rect 17589 18371 17647 18377
rect 19613 18411 19671 18417
rect 19613 18377 19625 18411
rect 19659 18408 19671 18411
rect 20990 18408 20996 18420
rect 19659 18380 20996 18408
rect 19659 18377 19671 18380
rect 19613 18371 19671 18377
rect 20990 18368 20996 18380
rect 21048 18368 21054 18420
rect 21266 18368 21272 18420
rect 21324 18408 21330 18420
rect 23014 18408 23020 18420
rect 21324 18380 23020 18408
rect 21324 18368 21330 18380
rect 23014 18368 23020 18380
rect 23072 18368 23078 18420
rect 23658 18368 23664 18420
rect 23716 18408 23722 18420
rect 25590 18408 25596 18420
rect 23716 18380 25596 18408
rect 23716 18368 23722 18380
rect 25590 18368 25596 18380
rect 25648 18368 25654 18420
rect 25866 18368 25872 18420
rect 25924 18408 25930 18420
rect 25924 18380 29500 18408
rect 25924 18368 25930 18380
rect 17310 18300 17316 18352
rect 17368 18340 17374 18352
rect 17368 18312 17413 18340
rect 17368 18300 17374 18312
rect 18414 18300 18420 18352
rect 18472 18340 18478 18352
rect 21726 18340 21732 18352
rect 18472 18312 20760 18340
rect 18472 18300 18478 18312
rect 17402 18232 17408 18284
rect 17460 18270 17466 18284
rect 17497 18275 17555 18281
rect 17497 18270 17509 18275
rect 17460 18242 17509 18270
rect 17460 18232 17466 18242
rect 17497 18241 17509 18242
rect 17543 18241 17555 18275
rect 17497 18235 17555 18241
rect 17589 18275 17647 18281
rect 17589 18241 17601 18275
rect 17635 18272 17647 18275
rect 18046 18272 18052 18284
rect 17635 18244 18052 18272
rect 17635 18241 17647 18244
rect 17589 18235 17647 18241
rect 18046 18232 18052 18244
rect 18104 18232 18110 18284
rect 18233 18275 18291 18281
rect 18233 18241 18245 18275
rect 18279 18272 18291 18275
rect 18506 18272 18512 18284
rect 18279 18244 18512 18272
rect 18279 18241 18291 18244
rect 18233 18235 18291 18241
rect 18506 18232 18512 18244
rect 18564 18232 18570 18284
rect 18966 18232 18972 18284
rect 19024 18272 19030 18284
rect 19245 18275 19303 18281
rect 19245 18272 19257 18275
rect 19024 18244 19257 18272
rect 19024 18232 19030 18244
rect 19245 18241 19257 18244
rect 19291 18241 19303 18275
rect 19245 18235 19303 18241
rect 19610 18232 19616 18284
rect 19668 18272 19674 18284
rect 20346 18272 20352 18284
rect 19668 18244 20352 18272
rect 19668 18232 19674 18244
rect 20346 18232 20352 18244
rect 20404 18232 20410 18284
rect 17310 18204 17316 18216
rect 17236 18176 17316 18204
rect 17310 18164 17316 18176
rect 17368 18164 17374 18216
rect 17770 18164 17776 18216
rect 17828 18204 17834 18216
rect 18141 18207 18199 18213
rect 18141 18204 18153 18207
rect 17828 18176 18153 18204
rect 17828 18164 17834 18176
rect 18141 18173 18153 18176
rect 18187 18173 18199 18207
rect 18141 18167 18199 18173
rect 18874 18164 18880 18216
rect 18932 18204 18938 18216
rect 19153 18207 19211 18213
rect 19153 18204 19165 18207
rect 18932 18176 19165 18204
rect 18932 18164 18938 18176
rect 19153 18173 19165 18176
rect 19199 18173 19211 18207
rect 19153 18167 19211 18173
rect 20073 18207 20131 18213
rect 20073 18173 20085 18207
rect 20119 18173 20131 18207
rect 20732 18204 20760 18312
rect 21284 18312 21732 18340
rect 20898 18232 20904 18284
rect 20956 18272 20962 18284
rect 21284 18281 21312 18312
rect 21726 18300 21732 18312
rect 21784 18300 21790 18352
rect 22741 18343 22799 18349
rect 22741 18340 22753 18343
rect 22066 18312 22753 18340
rect 20993 18275 21051 18281
rect 20993 18272 21005 18275
rect 20956 18244 21005 18272
rect 20956 18232 20962 18244
rect 20993 18241 21005 18244
rect 21039 18241 21051 18275
rect 20993 18235 21051 18241
rect 21269 18275 21327 18281
rect 21269 18241 21281 18275
rect 21315 18241 21327 18275
rect 21269 18235 21327 18241
rect 21450 18232 21456 18284
rect 21508 18272 21514 18284
rect 21821 18275 21879 18281
rect 21821 18272 21833 18275
rect 21508 18244 21833 18272
rect 21508 18232 21514 18244
rect 21821 18241 21833 18244
rect 21867 18241 21879 18275
rect 21821 18235 21879 18241
rect 22066 18204 22094 18312
rect 22741 18309 22753 18312
rect 22787 18309 22799 18343
rect 24946 18340 24952 18352
rect 24907 18312 24952 18340
rect 22741 18303 22799 18309
rect 24946 18300 24952 18312
rect 25004 18300 25010 18352
rect 25406 18300 25412 18352
rect 25464 18300 25470 18352
rect 29086 18340 29092 18352
rect 29047 18312 29092 18340
rect 29086 18300 29092 18312
rect 29144 18300 29150 18352
rect 29472 18340 29500 18380
rect 30374 18368 30380 18420
rect 30432 18408 30438 18420
rect 30432 18380 31340 18408
rect 30432 18368 30438 18380
rect 30009 18343 30067 18349
rect 30009 18340 30021 18343
rect 29472 18312 30021 18340
rect 30009 18309 30021 18312
rect 30055 18309 30067 18343
rect 31312 18340 31340 18380
rect 33778 18368 33784 18420
rect 33836 18408 33842 18420
rect 38838 18408 38844 18420
rect 33836 18380 38844 18408
rect 33836 18368 33842 18380
rect 38838 18368 38844 18380
rect 38896 18368 38902 18420
rect 39022 18408 39028 18420
rect 38983 18380 39028 18408
rect 39022 18368 39028 18380
rect 39080 18368 39086 18420
rect 39298 18368 39304 18420
rect 39356 18408 39362 18420
rect 40126 18408 40132 18420
rect 39356 18380 40132 18408
rect 39356 18368 39362 18380
rect 40126 18368 40132 18380
rect 40184 18368 40190 18420
rect 40972 18380 41552 18408
rect 37458 18340 37464 18352
rect 31312 18312 36400 18340
rect 30009 18303 30067 18309
rect 22462 18272 22468 18284
rect 22423 18244 22468 18272
rect 22462 18232 22468 18244
rect 22520 18232 22526 18284
rect 23842 18232 23848 18284
rect 23900 18232 23906 18284
rect 31018 18232 31024 18284
rect 31076 18272 31082 18284
rect 31386 18272 31392 18284
rect 31076 18244 31392 18272
rect 31076 18232 31082 18244
rect 31386 18232 31392 18244
rect 31444 18232 31450 18284
rect 33965 18275 34023 18281
rect 33965 18241 33977 18275
rect 34011 18272 34023 18275
rect 34011 18244 34836 18272
rect 34011 18241 34023 18244
rect 33965 18235 34023 18241
rect 20732 18176 22094 18204
rect 20073 18167 20131 18173
rect 15565 18139 15623 18145
rect 15565 18105 15577 18139
rect 15611 18136 15623 18139
rect 16758 18136 16764 18148
rect 15611 18108 16620 18136
rect 16719 18108 16764 18136
rect 15611 18105 15623 18108
rect 15565 18099 15623 18105
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 11609 18071 11667 18077
rect 11609 18037 11621 18071
rect 11655 18068 11667 18071
rect 12158 18068 12164 18080
rect 11655 18040 12164 18068
rect 11655 18037 11667 18040
rect 11609 18031 11667 18037
rect 12158 18028 12164 18040
rect 12216 18068 12222 18080
rect 13814 18068 13820 18080
rect 12216 18040 13820 18068
rect 12216 18028 12222 18040
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 14366 18068 14372 18080
rect 14327 18040 14372 18068
rect 14366 18028 14372 18040
rect 14424 18028 14430 18080
rect 15010 18068 15016 18080
rect 14971 18040 15016 18068
rect 15010 18028 15016 18040
rect 15068 18028 15074 18080
rect 16117 18071 16175 18077
rect 16117 18037 16129 18071
rect 16163 18068 16175 18071
rect 16482 18068 16488 18080
rect 16163 18040 16488 18068
rect 16163 18037 16175 18040
rect 16117 18031 16175 18037
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 16592 18068 16620 18108
rect 16758 18096 16764 18108
rect 16816 18096 16822 18148
rect 17586 18096 17592 18148
rect 17644 18136 17650 18148
rect 17644 18108 19334 18136
rect 17644 18096 17650 18108
rect 18340 18080 18368 18108
rect 18138 18068 18144 18080
rect 16592 18040 18144 18068
rect 18138 18028 18144 18040
rect 18196 18028 18202 18080
rect 18322 18028 18328 18080
rect 18380 18028 18386 18080
rect 18506 18068 18512 18080
rect 18467 18040 18512 18068
rect 18506 18028 18512 18040
rect 18564 18028 18570 18080
rect 19306 18068 19334 18108
rect 19610 18096 19616 18148
rect 19668 18136 19674 18148
rect 19794 18136 19800 18148
rect 19668 18108 19800 18136
rect 19668 18096 19674 18108
rect 19794 18096 19800 18108
rect 19852 18136 19858 18148
rect 20088 18136 20116 18167
rect 24210 18164 24216 18216
rect 24268 18204 24274 18216
rect 24673 18207 24731 18213
rect 24673 18204 24685 18207
rect 24268 18176 24685 18204
rect 24268 18164 24274 18176
rect 24673 18173 24685 18176
rect 24719 18173 24731 18207
rect 24673 18167 24731 18173
rect 27154 18164 27160 18216
rect 27212 18204 27218 18216
rect 28813 18207 28871 18213
rect 28813 18204 28825 18207
rect 27212 18176 28825 18204
rect 27212 18164 27218 18176
rect 28813 18173 28825 18176
rect 28859 18173 28871 18207
rect 28813 18167 28871 18173
rect 29273 18207 29331 18213
rect 29273 18173 29285 18207
rect 29319 18204 29331 18207
rect 29362 18204 29368 18216
rect 29319 18176 29368 18204
rect 29319 18173 29331 18176
rect 29273 18167 29331 18173
rect 19852 18108 20116 18136
rect 19852 18096 19858 18108
rect 20714 18096 20720 18148
rect 20772 18136 20778 18148
rect 28828 18136 28856 18167
rect 29362 18164 29368 18176
rect 29420 18164 29426 18216
rect 29454 18164 29460 18216
rect 29512 18204 29518 18216
rect 29733 18207 29791 18213
rect 29733 18204 29745 18207
rect 29512 18176 29745 18204
rect 29512 18164 29518 18176
rect 29733 18173 29745 18176
rect 29779 18173 29791 18207
rect 30374 18204 30380 18216
rect 29733 18167 29791 18173
rect 29840 18176 30380 18204
rect 29840 18136 29868 18176
rect 30374 18164 30380 18176
rect 30432 18164 30438 18216
rect 31202 18164 31208 18216
rect 31260 18204 31266 18216
rect 31481 18207 31539 18213
rect 31481 18204 31493 18207
rect 31260 18176 31493 18204
rect 31260 18164 31266 18176
rect 31481 18173 31493 18176
rect 31527 18173 31539 18207
rect 31481 18167 31539 18173
rect 32306 18164 32312 18216
rect 32364 18204 32370 18216
rect 32766 18204 32772 18216
rect 32364 18176 32772 18204
rect 32364 18164 32370 18176
rect 32766 18164 32772 18176
rect 32824 18164 32830 18216
rect 33410 18204 33416 18216
rect 33371 18176 33416 18204
rect 33410 18164 33416 18176
rect 33468 18164 33474 18216
rect 33778 18204 33784 18216
rect 33739 18176 33784 18204
rect 33778 18164 33784 18176
rect 33836 18164 33842 18216
rect 20772 18108 22094 18136
rect 20772 18096 20778 18108
rect 21634 18068 21640 18080
rect 19306 18040 21640 18068
rect 21634 18028 21640 18040
rect 21692 18028 21698 18080
rect 21910 18068 21916 18080
rect 21871 18040 21916 18068
rect 21910 18028 21916 18040
rect 21968 18028 21974 18080
rect 22066 18068 22094 18108
rect 26344 18108 28028 18136
rect 28828 18108 29868 18136
rect 31404 18108 31754 18136
rect 23474 18068 23480 18080
rect 22066 18040 23480 18068
rect 23474 18028 23480 18040
rect 23532 18028 23538 18080
rect 24213 18071 24271 18077
rect 24213 18037 24225 18071
rect 24259 18068 24271 18071
rect 26344 18068 26372 18108
rect 24259 18040 26372 18068
rect 26421 18071 26479 18077
rect 24259 18037 24271 18040
rect 24213 18031 24271 18037
rect 26421 18037 26433 18071
rect 26467 18068 26479 18071
rect 27890 18068 27896 18080
rect 26467 18040 27896 18068
rect 26467 18037 26479 18040
rect 26421 18031 26479 18037
rect 27890 18028 27896 18040
rect 27948 18028 27954 18080
rect 28000 18068 28028 18108
rect 31404 18068 31432 18108
rect 28000 18040 31432 18068
rect 31726 18068 31754 18108
rect 32030 18096 32036 18148
rect 32088 18136 32094 18148
rect 32490 18136 32496 18148
rect 32088 18108 32496 18136
rect 32088 18096 32094 18108
rect 32490 18096 32496 18108
rect 32548 18096 32554 18148
rect 32674 18096 32680 18148
rect 32732 18136 32738 18148
rect 33980 18136 34008 18235
rect 34698 18204 34704 18216
rect 34659 18176 34704 18204
rect 34698 18164 34704 18176
rect 34756 18164 34762 18216
rect 34808 18204 34836 18244
rect 35066 18204 35072 18216
rect 34808 18176 35072 18204
rect 35066 18164 35072 18176
rect 35124 18164 35130 18216
rect 36081 18207 36139 18213
rect 36081 18173 36093 18207
rect 36127 18173 36139 18207
rect 36262 18204 36268 18216
rect 36223 18176 36268 18204
rect 36081 18167 36139 18173
rect 32732 18108 34008 18136
rect 32732 18096 32738 18108
rect 33042 18068 33048 18080
rect 31726 18040 33048 18068
rect 33042 18028 33048 18040
rect 33100 18028 33106 18080
rect 33410 18028 33416 18080
rect 33468 18068 33474 18080
rect 33962 18068 33968 18080
rect 33468 18040 33968 18068
rect 33468 18028 33474 18040
rect 33962 18028 33968 18040
rect 34020 18028 34026 18080
rect 36096 18068 36124 18167
rect 36262 18164 36268 18176
rect 36320 18164 36326 18216
rect 36372 18204 36400 18312
rect 37292 18312 37464 18340
rect 37292 18281 37320 18312
rect 37458 18300 37464 18312
rect 37516 18300 37522 18352
rect 37553 18343 37611 18349
rect 37553 18309 37565 18343
rect 37599 18340 37611 18343
rect 37642 18340 37648 18352
rect 37599 18312 37648 18340
rect 37599 18309 37611 18312
rect 37553 18303 37611 18309
rect 37642 18300 37648 18312
rect 37700 18300 37706 18352
rect 39206 18300 39212 18352
rect 39264 18340 39270 18352
rect 40972 18349 41000 18380
rect 40957 18343 41015 18349
rect 39264 18312 39790 18340
rect 39264 18300 39270 18312
rect 40957 18309 40969 18343
rect 41003 18309 41015 18343
rect 41524 18340 41552 18380
rect 41598 18368 41604 18420
rect 41656 18408 41662 18420
rect 41785 18411 41843 18417
rect 41785 18408 41797 18411
rect 41656 18380 41797 18408
rect 41656 18368 41662 18380
rect 41785 18377 41797 18380
rect 41831 18377 41843 18411
rect 41785 18371 41843 18377
rect 42426 18368 42432 18420
rect 42484 18408 42490 18420
rect 43533 18411 43591 18417
rect 43533 18408 43545 18411
rect 42484 18380 43545 18408
rect 42484 18368 42490 18380
rect 43533 18377 43545 18380
rect 43579 18377 43591 18411
rect 43533 18371 43591 18377
rect 44174 18368 44180 18420
rect 44232 18408 44238 18420
rect 44450 18408 44456 18420
rect 44232 18380 44456 18408
rect 44232 18368 44238 18380
rect 44450 18368 44456 18380
rect 44508 18368 44514 18420
rect 45002 18408 45008 18420
rect 44963 18380 45008 18408
rect 45002 18368 45008 18380
rect 45060 18368 45066 18420
rect 45094 18368 45100 18420
rect 45152 18408 45158 18420
rect 45554 18408 45560 18420
rect 45152 18380 45560 18408
rect 45152 18368 45158 18380
rect 45554 18368 45560 18380
rect 45612 18368 45618 18420
rect 46106 18408 46112 18420
rect 46067 18380 46112 18408
rect 46106 18368 46112 18380
rect 46164 18368 46170 18420
rect 46934 18368 46940 18420
rect 46992 18408 46998 18420
rect 48133 18411 48191 18417
rect 48133 18408 48145 18411
rect 46992 18380 48145 18408
rect 46992 18368 46998 18380
rect 48133 18377 48145 18380
rect 48179 18377 48191 18411
rect 48682 18408 48688 18420
rect 48643 18380 48688 18408
rect 48133 18371 48191 18377
rect 48682 18368 48688 18380
rect 48740 18368 48746 18420
rect 58158 18408 58164 18420
rect 58119 18380 58164 18408
rect 58158 18368 58164 18380
rect 58216 18368 58222 18420
rect 43806 18340 43812 18352
rect 41524 18312 43812 18340
rect 40957 18303 41015 18309
rect 43806 18300 43812 18312
rect 43864 18300 43870 18352
rect 44376 18312 44588 18340
rect 37277 18275 37335 18281
rect 37277 18241 37289 18275
rect 37323 18241 37335 18275
rect 37277 18235 37335 18241
rect 38654 18232 38660 18284
rect 38712 18232 38718 18284
rect 41233 18275 41291 18281
rect 41233 18241 41245 18275
rect 41279 18272 41291 18275
rect 41322 18272 41328 18284
rect 41279 18244 41328 18272
rect 41279 18241 41291 18244
rect 41233 18235 41291 18241
rect 41322 18232 41328 18244
rect 41380 18232 41386 18284
rect 41874 18272 41880 18284
rect 41835 18244 41880 18272
rect 41874 18232 41880 18244
rect 41932 18232 41938 18284
rect 42794 18272 42800 18284
rect 42755 18244 42800 18272
rect 42794 18232 42800 18244
rect 42852 18232 42858 18284
rect 43162 18232 43168 18284
rect 43220 18272 43226 18284
rect 43533 18275 43591 18281
rect 43533 18272 43545 18275
rect 43220 18244 43545 18272
rect 43220 18232 43226 18244
rect 43533 18241 43545 18244
rect 43579 18272 43591 18275
rect 44376 18272 44404 18312
rect 43579 18244 44404 18272
rect 44453 18275 44511 18281
rect 43579 18241 43591 18244
rect 43533 18235 43591 18241
rect 44453 18241 44465 18275
rect 44499 18241 44511 18275
rect 44560 18272 44588 18312
rect 44910 18300 44916 18352
rect 44968 18340 44974 18352
rect 46661 18343 46719 18349
rect 46661 18340 46673 18343
rect 44968 18312 46673 18340
rect 44968 18300 44974 18312
rect 46661 18309 46673 18312
rect 46707 18309 46719 18343
rect 46661 18303 46719 18309
rect 45002 18272 45008 18284
rect 44560 18244 45008 18272
rect 44453 18235 44511 18241
rect 36372 18176 41460 18204
rect 38562 18096 38568 18148
rect 38620 18136 38626 18148
rect 41432 18136 41460 18176
rect 42058 18164 42064 18216
rect 42116 18204 42122 18216
rect 42702 18204 42708 18216
rect 42116 18176 42708 18204
rect 42116 18164 42122 18176
rect 42702 18164 42708 18176
rect 42760 18164 42766 18216
rect 42886 18204 42892 18216
rect 42847 18176 42892 18204
rect 42886 18164 42892 18176
rect 42944 18164 42950 18216
rect 43898 18164 43904 18216
rect 43956 18204 43962 18216
rect 44177 18207 44235 18213
rect 44177 18204 44189 18207
rect 43956 18176 44189 18204
rect 43956 18164 43962 18176
rect 44177 18173 44189 18176
rect 44223 18173 44235 18207
rect 44177 18167 44235 18173
rect 44468 18136 44496 18235
rect 45002 18232 45008 18244
rect 45060 18232 45066 18284
rect 45097 18275 45155 18281
rect 45097 18241 45109 18275
rect 45143 18272 45155 18275
rect 46198 18272 46204 18284
rect 45143 18244 46204 18272
rect 45143 18241 45155 18244
rect 45097 18235 45155 18241
rect 46198 18232 46204 18244
rect 46256 18272 46262 18284
rect 46566 18272 46572 18284
rect 46256 18244 46572 18272
rect 46256 18232 46262 18244
rect 46566 18232 46572 18244
rect 46624 18232 46630 18284
rect 48314 18232 48320 18284
rect 48372 18272 48378 18284
rect 49789 18275 49847 18281
rect 49789 18272 49801 18275
rect 48372 18244 49801 18272
rect 48372 18232 48378 18244
rect 49789 18241 49801 18244
rect 49835 18241 49847 18275
rect 49789 18235 49847 18241
rect 51046 18244 55214 18272
rect 47581 18207 47639 18213
rect 47581 18204 47593 18207
rect 45112 18176 47593 18204
rect 45112 18136 45140 18176
rect 47581 18173 47593 18176
rect 47627 18173 47639 18207
rect 51046 18204 51074 18244
rect 47581 18167 47639 18173
rect 47688 18176 51074 18204
rect 55186 18204 55214 18244
rect 57882 18204 57888 18216
rect 55186 18176 57888 18204
rect 38620 18108 39712 18136
rect 41432 18108 45140 18136
rect 38620 18096 38626 18108
rect 39390 18068 39396 18080
rect 36096 18040 39396 18068
rect 39390 18028 39396 18040
rect 39448 18028 39454 18080
rect 39482 18028 39488 18080
rect 39540 18068 39546 18080
rect 39684 18068 39712 18108
rect 45554 18096 45560 18148
rect 45612 18136 45618 18148
rect 47688 18136 47716 18176
rect 57882 18164 57888 18176
rect 57940 18164 57946 18216
rect 50433 18139 50491 18145
rect 50433 18136 50445 18139
rect 45612 18108 47716 18136
rect 47780 18108 50445 18136
rect 45612 18096 45618 18108
rect 41322 18068 41328 18080
rect 39540 18040 39585 18068
rect 39684 18040 41328 18068
rect 39540 18028 39546 18040
rect 41322 18028 41328 18040
rect 41380 18028 41386 18080
rect 41414 18028 41420 18080
rect 41472 18068 41478 18080
rect 42429 18071 42487 18077
rect 42429 18068 42441 18071
rect 41472 18040 42441 18068
rect 41472 18028 41478 18040
rect 42429 18037 42441 18040
rect 42475 18037 42487 18071
rect 42429 18031 42487 18037
rect 42702 18028 42708 18080
rect 42760 18068 42766 18080
rect 47780 18068 47808 18108
rect 50433 18105 50445 18108
rect 50479 18105 50491 18139
rect 50433 18099 50491 18105
rect 42760 18040 47808 18068
rect 49329 18071 49387 18077
rect 42760 18028 42766 18040
rect 49329 18037 49341 18071
rect 49375 18068 49387 18071
rect 49602 18068 49608 18080
rect 49375 18040 49608 18068
rect 49375 18037 49387 18040
rect 49329 18031 49387 18037
rect 49602 18028 49608 18040
rect 49660 18028 49666 18080
rect 1104 17978 58880 18000
rect 1104 17926 10582 17978
rect 10634 17926 10646 17978
rect 10698 17926 10710 17978
rect 10762 17926 10774 17978
rect 10826 17926 10838 17978
rect 10890 17926 29846 17978
rect 29898 17926 29910 17978
rect 29962 17926 29974 17978
rect 30026 17926 30038 17978
rect 30090 17926 30102 17978
rect 30154 17926 49110 17978
rect 49162 17926 49174 17978
rect 49226 17926 49238 17978
rect 49290 17926 49302 17978
rect 49354 17926 49366 17978
rect 49418 17926 58880 17978
rect 1104 17904 58880 17926
rect 12989 17867 13047 17873
rect 12989 17833 13001 17867
rect 13035 17864 13047 17867
rect 13906 17864 13912 17876
rect 13035 17836 13912 17864
rect 13035 17833 13047 17836
rect 12989 17827 13047 17833
rect 13906 17824 13912 17836
rect 13964 17864 13970 17876
rect 14550 17864 14556 17876
rect 13964 17836 14556 17864
rect 13964 17824 13970 17836
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 15930 17864 15936 17876
rect 15891 17836 15936 17864
rect 15930 17824 15936 17836
rect 15988 17824 15994 17876
rect 16114 17824 16120 17876
rect 16172 17864 16178 17876
rect 16577 17867 16635 17873
rect 16577 17864 16589 17867
rect 16172 17836 16589 17864
rect 16172 17824 16178 17836
rect 16577 17833 16589 17836
rect 16623 17833 16635 17867
rect 18046 17864 18052 17876
rect 16577 17827 16635 17833
rect 17236 17836 18052 17864
rect 14829 17799 14887 17805
rect 14829 17765 14841 17799
rect 14875 17796 14887 17799
rect 14875 17768 16804 17796
rect 14875 17765 14887 17768
rect 14829 17759 14887 17765
rect 13541 17731 13599 17737
rect 13541 17697 13553 17731
rect 13587 17728 13599 17731
rect 16776 17728 16804 17768
rect 17236 17728 17264 17836
rect 18046 17824 18052 17836
rect 18104 17864 18110 17876
rect 18104 17836 18552 17864
rect 18104 17824 18110 17836
rect 18138 17756 18144 17808
rect 18196 17796 18202 17808
rect 18524 17796 18552 17836
rect 18598 17824 18604 17876
rect 18656 17864 18662 17876
rect 18693 17867 18751 17873
rect 18693 17864 18705 17867
rect 18656 17836 18705 17864
rect 18656 17824 18662 17836
rect 18693 17833 18705 17836
rect 18739 17833 18751 17867
rect 18693 17827 18751 17833
rect 19981 17867 20039 17873
rect 19981 17833 19993 17867
rect 20027 17864 20039 17867
rect 20714 17864 20720 17876
rect 20027 17836 20720 17864
rect 20027 17833 20039 17836
rect 19981 17827 20039 17833
rect 20714 17824 20720 17836
rect 20772 17824 20778 17876
rect 21542 17824 21548 17876
rect 21600 17864 21606 17876
rect 21726 17864 21732 17876
rect 21600 17836 21732 17864
rect 21600 17824 21606 17836
rect 21726 17824 21732 17836
rect 21784 17824 21790 17876
rect 22094 17824 22100 17876
rect 22152 17864 22158 17876
rect 24489 17867 24547 17873
rect 22152 17836 23428 17864
rect 22152 17824 22158 17836
rect 19426 17796 19432 17808
rect 18196 17768 18368 17796
rect 18524 17768 19432 17796
rect 18196 17756 18202 17768
rect 17402 17728 17408 17740
rect 13587 17700 16712 17728
rect 16776 17700 17264 17728
rect 17363 17700 17408 17728
rect 13587 17697 13599 17700
rect 13541 17691 13599 17697
rect 16684 17672 16712 17700
rect 17402 17688 17408 17700
rect 17460 17688 17466 17740
rect 18340 17737 18368 17768
rect 19426 17756 19432 17768
rect 19484 17756 19490 17808
rect 23400 17796 23428 17836
rect 24489 17833 24501 17867
rect 24535 17864 24547 17867
rect 24578 17864 24584 17876
rect 24535 17836 24584 17864
rect 24535 17833 24547 17836
rect 24489 17827 24547 17833
rect 24578 17824 24584 17836
rect 24636 17824 24642 17876
rect 25682 17864 25688 17876
rect 25056 17836 25688 17864
rect 24949 17799 25007 17805
rect 24949 17796 24961 17799
rect 23400 17768 24961 17796
rect 24949 17765 24961 17768
rect 24995 17765 25007 17799
rect 24949 17759 25007 17765
rect 18233 17731 18291 17737
rect 18233 17728 18245 17731
rect 17512 17700 18245 17728
rect 16025 17663 16083 17669
rect 16025 17629 16037 17663
rect 16071 17660 16083 17663
rect 16390 17660 16396 17672
rect 16071 17632 16396 17660
rect 16071 17629 16083 17632
rect 16025 17623 16083 17629
rect 16390 17620 16396 17632
rect 16448 17620 16454 17672
rect 16482 17620 16488 17672
rect 16540 17660 16546 17672
rect 16540 17632 16585 17660
rect 16540 17620 16546 17632
rect 16666 17620 16672 17672
rect 16724 17660 16730 17672
rect 17313 17663 17371 17669
rect 17313 17660 17325 17663
rect 16724 17632 17325 17660
rect 16724 17620 16730 17632
rect 17313 17629 17325 17632
rect 17359 17629 17371 17663
rect 17512 17660 17540 17700
rect 18233 17697 18245 17700
rect 18279 17697 18291 17731
rect 18233 17691 18291 17697
rect 18325 17731 18383 17737
rect 18325 17697 18337 17731
rect 18371 17697 18383 17731
rect 18325 17691 18383 17697
rect 18417 17731 18475 17737
rect 18417 17697 18429 17731
rect 18463 17728 18475 17731
rect 19058 17728 19064 17740
rect 18463 17700 19064 17728
rect 18463 17697 18475 17700
rect 18417 17691 18475 17697
rect 19058 17688 19064 17700
rect 19116 17688 19122 17740
rect 19260 17700 19564 17728
rect 17313 17623 17371 17629
rect 17420 17632 17540 17660
rect 14277 17595 14335 17601
rect 14277 17561 14289 17595
rect 14323 17592 14335 17595
rect 16850 17592 16856 17604
rect 14323 17564 16856 17592
rect 14323 17561 14335 17564
rect 14277 17555 14335 17561
rect 16850 17552 16856 17564
rect 16908 17552 16914 17604
rect 16942 17552 16948 17604
rect 17000 17592 17006 17604
rect 17420 17592 17448 17632
rect 17586 17620 17592 17672
rect 17644 17660 17650 17672
rect 18509 17663 18567 17669
rect 18509 17660 18521 17663
rect 17644 17632 18521 17660
rect 17644 17620 17650 17632
rect 18509 17629 18521 17632
rect 18555 17660 18567 17663
rect 18782 17660 18788 17672
rect 18555 17632 18788 17660
rect 18555 17629 18567 17632
rect 18509 17623 18567 17629
rect 18782 17620 18788 17632
rect 18840 17620 18846 17672
rect 19260 17660 19288 17700
rect 19426 17660 19432 17672
rect 18984 17632 19288 17660
rect 19387 17632 19432 17660
rect 18984 17592 19012 17632
rect 19426 17620 19432 17632
rect 19484 17620 19490 17672
rect 19536 17669 19564 17700
rect 19610 17688 19616 17740
rect 19668 17728 19674 17740
rect 20441 17731 20499 17737
rect 20441 17728 20453 17731
rect 19668 17700 20453 17728
rect 19668 17688 19674 17700
rect 20441 17697 20453 17700
rect 20487 17697 20499 17731
rect 20441 17691 20499 17697
rect 21174 17688 21180 17740
rect 21232 17728 21238 17740
rect 22373 17731 22431 17737
rect 22373 17728 22385 17731
rect 21232 17700 22385 17728
rect 21232 17688 21238 17700
rect 22373 17697 22385 17700
rect 22419 17697 22431 17731
rect 22373 17691 22431 17697
rect 22462 17688 22468 17740
rect 22520 17728 22526 17740
rect 22922 17728 22928 17740
rect 22520 17700 22928 17728
rect 22520 17688 22526 17700
rect 22922 17688 22928 17700
rect 22980 17728 22986 17740
rect 25056 17728 25084 17836
rect 25682 17824 25688 17836
rect 25740 17864 25746 17876
rect 25740 17836 27200 17864
rect 25740 17824 25746 17836
rect 22980 17700 25084 17728
rect 22980 17688 22986 17700
rect 26050 17688 26056 17740
rect 26108 17728 26114 17740
rect 27172 17737 27200 17836
rect 28534 17824 28540 17876
rect 28592 17864 28598 17876
rect 28902 17864 28908 17876
rect 28592 17836 28908 17864
rect 28592 17824 28598 17836
rect 28902 17824 28908 17836
rect 28960 17864 28966 17876
rect 30650 17864 30656 17876
rect 28960 17836 30656 17864
rect 28960 17824 28966 17836
rect 30650 17824 30656 17836
rect 30708 17824 30714 17876
rect 31481 17867 31539 17873
rect 31481 17833 31493 17867
rect 31527 17864 31539 17867
rect 31570 17864 31576 17876
rect 31527 17836 31576 17864
rect 31527 17833 31539 17836
rect 31481 17827 31539 17833
rect 31570 17824 31576 17836
rect 31628 17824 31634 17876
rect 31754 17824 31760 17876
rect 31812 17864 31818 17876
rect 39758 17864 39764 17876
rect 31812 17836 39764 17864
rect 31812 17824 31818 17836
rect 39758 17824 39764 17836
rect 39816 17824 39822 17876
rect 44174 17864 44180 17876
rect 39960 17836 44180 17864
rect 33686 17756 33692 17808
rect 33744 17796 33750 17808
rect 33781 17799 33839 17805
rect 33781 17796 33793 17799
rect 33744 17768 33793 17796
rect 33744 17756 33750 17768
rect 33781 17765 33793 17768
rect 33827 17796 33839 17799
rect 35894 17796 35900 17808
rect 33827 17768 35900 17796
rect 33827 17765 33839 17768
rect 33781 17759 33839 17765
rect 35894 17756 35900 17768
rect 35952 17796 35958 17808
rect 36722 17796 36728 17808
rect 35952 17768 36728 17796
rect 35952 17756 35958 17768
rect 36722 17756 36728 17768
rect 36780 17756 36786 17808
rect 38930 17756 38936 17808
rect 38988 17796 38994 17808
rect 39209 17799 39267 17805
rect 39209 17796 39221 17799
rect 38988 17768 39221 17796
rect 38988 17756 38994 17768
rect 39209 17765 39221 17768
rect 39255 17765 39267 17799
rect 39209 17759 39267 17765
rect 39298 17756 39304 17808
rect 39356 17796 39362 17808
rect 39960 17796 39988 17836
rect 44174 17824 44180 17836
rect 44232 17824 44238 17876
rect 44266 17824 44272 17876
rect 44324 17864 44330 17876
rect 44361 17867 44419 17873
rect 44361 17864 44373 17867
rect 44324 17836 44373 17864
rect 44324 17824 44330 17836
rect 44361 17833 44373 17836
rect 44407 17833 44419 17867
rect 45094 17864 45100 17876
rect 45055 17836 45100 17864
rect 44361 17827 44419 17833
rect 45094 17824 45100 17836
rect 45152 17824 45158 17876
rect 46474 17864 46480 17876
rect 46435 17836 46480 17864
rect 46474 17824 46480 17836
rect 46532 17824 46538 17876
rect 48682 17824 48688 17876
rect 48740 17864 48746 17876
rect 49237 17867 49295 17873
rect 49237 17864 49249 17867
rect 48740 17836 49249 17864
rect 48740 17824 48746 17836
rect 49237 17833 49249 17836
rect 49283 17833 49295 17867
rect 49237 17827 49295 17833
rect 39356 17768 39988 17796
rect 39356 17756 39362 17768
rect 42242 17756 42248 17808
rect 42300 17796 42306 17808
rect 43254 17796 43260 17808
rect 42300 17768 42564 17796
rect 43215 17768 43260 17796
rect 42300 17756 42306 17768
rect 26697 17731 26755 17737
rect 26697 17728 26709 17731
rect 26108 17700 26709 17728
rect 26108 17688 26114 17700
rect 26697 17697 26709 17700
rect 26743 17697 26755 17731
rect 26697 17691 26755 17697
rect 27157 17731 27215 17737
rect 27157 17697 27169 17731
rect 27203 17697 27215 17731
rect 27157 17691 27215 17697
rect 19521 17663 19579 17669
rect 19521 17629 19533 17663
rect 19567 17629 19579 17663
rect 19521 17623 19579 17629
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17629 19763 17663
rect 19705 17623 19763 17629
rect 19797 17663 19855 17669
rect 19797 17629 19809 17663
rect 19843 17629 19855 17663
rect 19797 17623 19855 17629
rect 17000 17564 17448 17592
rect 17604 17564 19012 17592
rect 17000 17552 17006 17564
rect 11333 17527 11391 17533
rect 11333 17493 11345 17527
rect 11379 17524 11391 17527
rect 11793 17527 11851 17533
rect 11793 17524 11805 17527
rect 11379 17496 11805 17524
rect 11379 17493 11391 17496
rect 11333 17487 11391 17493
rect 11793 17493 11805 17496
rect 11839 17524 11851 17527
rect 12437 17527 12495 17533
rect 12437 17524 12449 17527
rect 11839 17496 12449 17524
rect 11839 17493 11851 17496
rect 11793 17487 11851 17493
rect 12437 17493 12449 17496
rect 12483 17524 12495 17527
rect 12986 17524 12992 17536
rect 12483 17496 12992 17524
rect 12483 17493 12495 17496
rect 12437 17487 12495 17493
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 15381 17527 15439 17533
rect 15381 17493 15393 17527
rect 15427 17524 15439 17527
rect 17604 17524 17632 17564
rect 15427 17496 17632 17524
rect 17681 17527 17739 17533
rect 15427 17493 15439 17496
rect 15381 17487 15439 17493
rect 17681 17493 17693 17527
rect 17727 17524 17739 17527
rect 18598 17524 18604 17536
rect 17727 17496 18604 17524
rect 17727 17493 17739 17496
rect 17681 17487 17739 17493
rect 18598 17484 18604 17496
rect 18656 17484 18662 17536
rect 18984 17524 19012 17564
rect 19242 17552 19248 17604
rect 19300 17592 19306 17604
rect 19720 17592 19748 17623
rect 19300 17564 19748 17592
rect 19812 17592 19840 17623
rect 20346 17620 20352 17672
rect 20404 17660 20410 17672
rect 20714 17660 20720 17672
rect 20404 17632 20720 17660
rect 20404 17620 20410 17632
rect 20714 17620 20720 17632
rect 20772 17620 20778 17672
rect 20898 17620 20904 17672
rect 20956 17660 20962 17672
rect 21361 17663 21419 17669
rect 20956 17632 21128 17660
rect 20956 17620 20962 17632
rect 20990 17592 20996 17604
rect 19812 17564 20996 17592
rect 19300 17552 19306 17564
rect 20990 17552 20996 17564
rect 21048 17552 21054 17604
rect 21100 17592 21128 17632
rect 21361 17629 21373 17663
rect 21407 17629 21419 17663
rect 21361 17623 21419 17629
rect 22097 17663 22155 17669
rect 22097 17629 22109 17663
rect 22143 17629 22155 17663
rect 22097 17623 22155 17629
rect 21376 17592 21404 17623
rect 22112 17592 22140 17623
rect 23658 17620 23664 17672
rect 23716 17660 23722 17672
rect 24394 17660 24400 17672
rect 23716 17632 24400 17660
rect 23716 17620 23722 17632
rect 24394 17620 24400 17632
rect 24452 17620 24458 17672
rect 26712 17660 26740 17691
rect 27982 17688 27988 17740
rect 28040 17728 28046 17740
rect 28813 17731 28871 17737
rect 28813 17728 28825 17731
rect 28040 17700 28825 17728
rect 28040 17688 28046 17700
rect 28813 17697 28825 17700
rect 28859 17697 28871 17731
rect 28813 17691 28871 17697
rect 28997 17731 29055 17737
rect 28997 17697 29009 17731
rect 29043 17728 29055 17731
rect 29043 17700 31340 17728
rect 29043 17697 29055 17700
rect 28997 17691 29055 17697
rect 26712 17632 27660 17660
rect 22370 17592 22376 17604
rect 21100 17564 21441 17592
rect 22112 17564 22376 17592
rect 21266 17524 21272 17536
rect 18984 17496 21272 17524
rect 21266 17484 21272 17496
rect 21324 17484 21330 17536
rect 21376 17524 21404 17564
rect 22370 17552 22376 17564
rect 22428 17552 22434 17604
rect 22830 17552 22836 17604
rect 22888 17552 22894 17604
rect 24302 17552 24308 17604
rect 24360 17592 24366 17604
rect 24360 17564 25084 17592
rect 24360 17552 24366 17564
rect 23014 17524 23020 17536
rect 21376 17496 23020 17524
rect 23014 17484 23020 17496
rect 23072 17484 23078 17536
rect 23845 17527 23903 17533
rect 23845 17493 23857 17527
rect 23891 17524 23903 17527
rect 24762 17524 24768 17536
rect 23891 17496 24768 17524
rect 23891 17493 23903 17496
rect 23845 17487 23903 17493
rect 24762 17484 24768 17496
rect 24820 17484 24826 17536
rect 25056 17524 25084 17564
rect 25130 17552 25136 17604
rect 25188 17592 25194 17604
rect 26421 17595 26479 17601
rect 25188 17564 25254 17592
rect 25188 17552 25194 17564
rect 26421 17561 26433 17595
rect 26467 17592 26479 17595
rect 27062 17592 27068 17604
rect 26467 17564 27068 17592
rect 26467 17561 26479 17564
rect 26421 17555 26479 17561
rect 27062 17552 27068 17564
rect 27120 17552 27126 17604
rect 27522 17524 27528 17536
rect 25056 17496 27528 17524
rect 27522 17484 27528 17496
rect 27580 17484 27586 17536
rect 27632 17524 27660 17632
rect 29454 17620 29460 17672
rect 29512 17660 29518 17672
rect 29733 17663 29791 17669
rect 29733 17660 29745 17663
rect 29512 17632 29745 17660
rect 29512 17620 29518 17632
rect 29733 17629 29745 17632
rect 29779 17629 29791 17663
rect 29733 17623 29791 17629
rect 29546 17552 29552 17604
rect 29604 17592 29610 17604
rect 30009 17595 30067 17601
rect 30009 17592 30021 17595
rect 29604 17564 30021 17592
rect 29604 17552 29610 17564
rect 30009 17561 30021 17564
rect 30055 17561 30067 17595
rect 30009 17555 30067 17561
rect 30834 17524 30840 17536
rect 27632 17496 30840 17524
rect 30834 17484 30840 17496
rect 30892 17484 30898 17536
rect 30926 17484 30932 17536
rect 30984 17524 30990 17536
rect 31128 17524 31156 17646
rect 31312 17592 31340 17700
rect 35986 17688 35992 17740
rect 36044 17728 36050 17740
rect 36541 17731 36599 17737
rect 36541 17728 36553 17731
rect 36044 17700 36553 17728
rect 36044 17688 36050 17700
rect 36541 17697 36553 17700
rect 36587 17728 36599 17731
rect 36814 17728 36820 17740
rect 36587 17700 36820 17728
rect 36587 17697 36599 17700
rect 36541 17691 36599 17697
rect 36814 17688 36820 17700
rect 36872 17688 36878 17740
rect 36998 17728 37004 17740
rect 36959 17700 37004 17728
rect 36998 17688 37004 17700
rect 37056 17688 37062 17740
rect 37274 17728 37280 17740
rect 37235 17700 37280 17728
rect 37274 17688 37280 17700
rect 37332 17688 37338 17740
rect 37366 17688 37372 17740
rect 37424 17728 37430 17740
rect 40954 17728 40960 17740
rect 37424 17700 40960 17728
rect 37424 17688 37430 17700
rect 40954 17688 40960 17700
rect 41012 17688 41018 17740
rect 42536 17737 42564 17768
rect 43254 17756 43260 17768
rect 43312 17756 43318 17808
rect 47581 17799 47639 17805
rect 47581 17796 47593 17799
rect 43456 17768 47593 17796
rect 42521 17731 42579 17737
rect 42521 17697 42533 17731
rect 42567 17697 42579 17731
rect 42521 17691 42579 17697
rect 42610 17688 42616 17740
rect 42668 17728 42674 17740
rect 42705 17731 42763 17737
rect 42705 17728 42717 17731
rect 42668 17700 42717 17728
rect 42668 17688 42674 17700
rect 42705 17697 42717 17700
rect 42751 17728 42763 17731
rect 43456 17728 43484 17768
rect 47581 17765 47593 17768
rect 47627 17765 47639 17799
rect 47581 17759 47639 17765
rect 42751 17700 43484 17728
rect 43717 17731 43775 17737
rect 42751 17697 42763 17700
rect 42705 17691 42763 17697
rect 43717 17697 43729 17731
rect 43763 17728 43775 17731
rect 44634 17728 44640 17740
rect 43763 17700 44640 17728
rect 43763 17697 43775 17700
rect 43717 17691 43775 17697
rect 44634 17688 44640 17700
rect 44692 17728 44698 17740
rect 44818 17728 44824 17740
rect 44692 17700 44824 17728
rect 44692 17688 44698 17700
rect 44818 17688 44824 17700
rect 44876 17688 44882 17740
rect 48222 17728 48228 17740
rect 45296 17700 48228 17728
rect 31662 17620 31668 17672
rect 31720 17660 31726 17672
rect 32033 17663 32091 17669
rect 32033 17660 32045 17663
rect 31720 17632 32045 17660
rect 31720 17620 31726 17632
rect 32033 17629 32045 17632
rect 32079 17629 32091 17663
rect 32033 17623 32091 17629
rect 41594 17663 41652 17669
rect 41594 17629 41606 17663
rect 41640 17660 41652 17663
rect 41782 17660 41788 17672
rect 41640 17632 41788 17660
rect 41640 17629 41652 17632
rect 41594 17623 41652 17629
rect 41782 17620 41788 17632
rect 41840 17620 41846 17672
rect 43625 17663 43683 17669
rect 43625 17629 43637 17663
rect 43671 17660 43683 17663
rect 44082 17660 44088 17672
rect 43671 17632 44088 17660
rect 43671 17629 43683 17632
rect 43625 17623 43683 17629
rect 44082 17620 44088 17632
rect 44140 17620 44146 17672
rect 44269 17663 44327 17669
rect 44269 17629 44281 17663
rect 44315 17660 44327 17663
rect 44542 17660 44548 17672
rect 44315 17632 44548 17660
rect 44315 17629 44327 17632
rect 44269 17623 44327 17629
rect 31846 17592 31852 17604
rect 31312 17564 31852 17592
rect 31846 17552 31852 17564
rect 31904 17552 31910 17604
rect 32309 17595 32367 17601
rect 32309 17561 32321 17595
rect 32355 17592 32367 17595
rect 32355 17564 32536 17592
rect 32355 17561 32367 17564
rect 32309 17555 32367 17561
rect 32508 17536 32536 17564
rect 33042 17552 33048 17604
rect 33100 17552 33106 17604
rect 34698 17552 34704 17604
rect 34756 17592 34762 17604
rect 35066 17592 35072 17604
rect 34756 17564 35072 17592
rect 34756 17552 34762 17564
rect 35066 17552 35072 17564
rect 35124 17552 35130 17604
rect 36357 17595 36415 17601
rect 36357 17561 36369 17595
rect 36403 17592 36415 17595
rect 37366 17592 37372 17604
rect 36403 17564 37372 17592
rect 36403 17561 36415 17564
rect 36357 17555 36415 17561
rect 37366 17552 37372 17564
rect 37424 17552 37430 17604
rect 38502 17564 40080 17592
rect 31386 17524 31392 17536
rect 30984 17496 31392 17524
rect 30984 17484 30990 17496
rect 31386 17484 31392 17496
rect 31444 17484 31450 17536
rect 32490 17484 32496 17536
rect 32548 17484 32554 17536
rect 34882 17484 34888 17536
rect 34940 17524 34946 17536
rect 38749 17527 38807 17533
rect 38749 17524 38761 17527
rect 34940 17496 38761 17524
rect 34940 17484 34946 17496
rect 38749 17493 38761 17496
rect 38795 17493 38807 17527
rect 38749 17487 38807 17493
rect 39022 17484 39028 17536
rect 39080 17524 39086 17536
rect 39853 17527 39911 17533
rect 39853 17524 39865 17527
rect 39080 17496 39865 17524
rect 39080 17484 39086 17496
rect 39853 17493 39865 17496
rect 39899 17493 39911 17527
rect 40052 17524 40080 17564
rect 40586 17552 40592 17604
rect 40644 17552 40650 17604
rect 41322 17592 41328 17604
rect 41283 17564 41328 17592
rect 41322 17552 41328 17564
rect 41380 17552 41386 17604
rect 41874 17552 41880 17604
rect 41932 17592 41938 17604
rect 44284 17592 44312 17623
rect 44542 17620 44548 17632
rect 44600 17620 44606 17672
rect 45296 17669 45324 17700
rect 48222 17688 48228 17700
rect 48280 17688 48286 17740
rect 45281 17663 45339 17669
rect 45281 17629 45293 17663
rect 45327 17629 45339 17663
rect 45281 17623 45339 17629
rect 45925 17663 45983 17669
rect 45925 17629 45937 17663
rect 45971 17660 45983 17663
rect 46474 17660 46480 17672
rect 45971 17632 46480 17660
rect 45971 17629 45983 17632
rect 45925 17623 45983 17629
rect 46474 17620 46480 17632
rect 46532 17620 46538 17672
rect 46569 17663 46627 17669
rect 46569 17629 46581 17663
rect 46615 17660 46627 17663
rect 46658 17660 46664 17672
rect 46615 17632 46664 17660
rect 46615 17629 46627 17632
rect 46569 17623 46627 17629
rect 46658 17620 46664 17632
rect 46716 17660 46722 17672
rect 48685 17663 48743 17669
rect 48685 17660 48697 17663
rect 46716 17632 48697 17660
rect 46716 17620 46722 17632
rect 48685 17629 48697 17632
rect 48731 17629 48743 17663
rect 48685 17623 48743 17629
rect 41932 17564 44312 17592
rect 41932 17552 41938 17564
rect 41690 17524 41696 17536
rect 40052 17496 41696 17524
rect 39853 17487 39911 17493
rect 41690 17484 41696 17496
rect 41748 17484 41754 17536
rect 42058 17524 42064 17536
rect 42019 17496 42064 17524
rect 42058 17484 42064 17496
rect 42116 17484 42122 17536
rect 42426 17524 42432 17536
rect 42387 17496 42432 17524
rect 42426 17484 42432 17496
rect 42484 17484 42490 17536
rect 42794 17484 42800 17536
rect 42852 17524 42858 17536
rect 45833 17527 45891 17533
rect 45833 17524 45845 17527
rect 42852 17496 45845 17524
rect 42852 17484 42858 17496
rect 45833 17493 45845 17496
rect 45879 17493 45891 17527
rect 47026 17524 47032 17536
rect 46987 17496 47032 17524
rect 45833 17487 45891 17493
rect 47026 17484 47032 17496
rect 47084 17484 47090 17536
rect 48222 17524 48228 17536
rect 48183 17496 48228 17524
rect 48222 17484 48228 17496
rect 48280 17484 48286 17536
rect 50154 17524 50160 17536
rect 50115 17496 50160 17524
rect 50154 17484 50160 17496
rect 50212 17484 50218 17536
rect 1104 17434 58880 17456
rect 1104 17382 20214 17434
rect 20266 17382 20278 17434
rect 20330 17382 20342 17434
rect 20394 17382 20406 17434
rect 20458 17382 20470 17434
rect 20522 17382 39478 17434
rect 39530 17382 39542 17434
rect 39594 17382 39606 17434
rect 39658 17382 39670 17434
rect 39722 17382 39734 17434
rect 39786 17382 58880 17434
rect 1104 17360 58880 17382
rect 12069 17323 12127 17329
rect 12069 17289 12081 17323
rect 12115 17320 12127 17323
rect 12710 17320 12716 17332
rect 12115 17292 12716 17320
rect 12115 17289 12127 17292
rect 12069 17283 12127 17289
rect 12710 17280 12716 17292
rect 12768 17280 12774 17332
rect 16022 17280 16028 17332
rect 16080 17320 16086 17332
rect 21174 17320 21180 17332
rect 16080 17292 21180 17320
rect 16080 17280 16086 17292
rect 21174 17280 21180 17292
rect 21232 17280 21238 17332
rect 21910 17280 21916 17332
rect 21968 17320 21974 17332
rect 22830 17320 22836 17332
rect 21968 17292 22836 17320
rect 21968 17280 21974 17292
rect 22830 17280 22836 17292
rect 22888 17280 22894 17332
rect 27706 17320 27712 17332
rect 22940 17292 27712 17320
rect 18966 17252 18972 17264
rect 16132 17224 18972 17252
rect 10965 17187 11023 17193
rect 10965 17153 10977 17187
rect 11011 17184 11023 17187
rect 13265 17187 13323 17193
rect 13265 17184 13277 17187
rect 11011 17156 13277 17184
rect 11011 17153 11023 17156
rect 10965 17147 11023 17153
rect 13265 17153 13277 17156
rect 13311 17184 13323 17187
rect 14274 17184 14280 17196
rect 13311 17156 14280 17184
rect 13311 17153 13323 17156
rect 13265 17147 13323 17153
rect 14274 17144 14280 17156
rect 14332 17144 14338 17196
rect 16132 17193 16160 17224
rect 18966 17212 18972 17224
rect 19024 17212 19030 17264
rect 19334 17252 19340 17264
rect 19295 17224 19340 17252
rect 19334 17212 19340 17224
rect 19392 17212 19398 17264
rect 19426 17212 19432 17264
rect 19484 17252 19490 17264
rect 19484 17224 19840 17252
rect 19484 17212 19490 17224
rect 15197 17187 15255 17193
rect 15197 17184 15209 17187
rect 14752 17156 15209 17184
rect 12618 17076 12624 17128
rect 12676 17116 12682 17128
rect 14752 17116 14780 17156
rect 15197 17153 15209 17156
rect 15243 17153 15255 17187
rect 15197 17147 15255 17153
rect 16117 17187 16175 17193
rect 16117 17153 16129 17187
rect 16163 17153 16175 17187
rect 16117 17147 16175 17153
rect 16850 17144 16856 17196
rect 16908 17184 16914 17196
rect 17207 17187 17265 17193
rect 17207 17184 17219 17187
rect 16908 17156 17219 17184
rect 16908 17144 16914 17156
rect 17207 17153 17219 17156
rect 17253 17153 17265 17187
rect 17207 17147 17265 17153
rect 18141 17187 18199 17193
rect 18141 17153 18153 17187
rect 18187 17184 18199 17187
rect 19058 17184 19064 17196
rect 18187 17156 19064 17184
rect 18187 17153 18199 17156
rect 18141 17147 18199 17153
rect 19058 17144 19064 17156
rect 19116 17144 19122 17196
rect 19812 17184 19840 17224
rect 19978 17212 19984 17264
rect 20036 17252 20042 17264
rect 22094 17252 22100 17264
rect 20036 17224 22100 17252
rect 20036 17212 20042 17224
rect 22094 17212 22100 17224
rect 22152 17212 22158 17264
rect 22741 17255 22799 17261
rect 22741 17221 22753 17255
rect 22787 17252 22799 17255
rect 22940 17252 22968 17292
rect 27706 17280 27712 17292
rect 27764 17280 27770 17332
rect 28626 17280 28632 17332
rect 28684 17320 28690 17332
rect 28813 17323 28871 17329
rect 28813 17320 28825 17323
rect 28684 17292 28825 17320
rect 28684 17280 28690 17292
rect 28813 17289 28825 17292
rect 28859 17320 28871 17323
rect 28902 17320 28908 17332
rect 28859 17292 28908 17320
rect 28859 17289 28871 17292
rect 28813 17283 28871 17289
rect 28902 17280 28908 17292
rect 28960 17280 28966 17332
rect 29546 17280 29552 17332
rect 29604 17320 29610 17332
rect 31662 17320 31668 17332
rect 29604 17292 31668 17320
rect 29604 17280 29610 17292
rect 31662 17280 31668 17292
rect 31720 17320 31726 17332
rect 31720 17292 31800 17320
rect 31720 17280 31726 17292
rect 22787 17224 22968 17252
rect 22787 17221 22799 17224
rect 22741 17215 22799 17221
rect 23014 17212 23020 17264
rect 23072 17252 23078 17264
rect 24949 17255 25007 17261
rect 23072 17224 23230 17252
rect 23072 17212 23078 17224
rect 24949 17221 24961 17255
rect 24995 17252 25007 17255
rect 25038 17252 25044 17264
rect 24995 17224 25044 17252
rect 24995 17221 25007 17224
rect 24949 17215 25007 17221
rect 25038 17212 25044 17224
rect 25096 17212 25102 17264
rect 27338 17252 27344 17264
rect 27299 17224 27344 17252
rect 27338 17212 27344 17224
rect 27396 17212 27402 17264
rect 27798 17212 27804 17264
rect 27856 17212 27862 17264
rect 30650 17252 30656 17264
rect 30498 17224 30656 17252
rect 30650 17212 30656 17224
rect 30708 17212 30714 17264
rect 31478 17212 31484 17264
rect 31536 17212 31542 17264
rect 20254 17184 20260 17196
rect 19812 17156 20260 17184
rect 20254 17144 20260 17156
rect 20312 17144 20318 17196
rect 20349 17187 20407 17193
rect 20349 17153 20361 17187
rect 20395 17184 20407 17187
rect 20438 17184 20444 17196
rect 20395 17156 20444 17184
rect 20395 17153 20407 17156
rect 20349 17147 20407 17153
rect 20438 17144 20444 17156
rect 20496 17144 20502 17196
rect 20622 17144 20628 17196
rect 20680 17184 20686 17196
rect 20993 17187 21051 17193
rect 20993 17184 21005 17187
rect 20680 17156 21005 17184
rect 20680 17144 20686 17156
rect 20993 17153 21005 17156
rect 21039 17153 21051 17187
rect 20993 17147 21051 17153
rect 21082 17144 21088 17196
rect 21140 17184 21146 17196
rect 21818 17184 21824 17196
rect 21140 17156 21824 17184
rect 21140 17144 21146 17156
rect 21818 17144 21824 17156
rect 21876 17144 21882 17196
rect 24670 17184 24676 17196
rect 24631 17156 24676 17184
rect 24670 17144 24676 17156
rect 24728 17144 24734 17196
rect 26050 17144 26056 17196
rect 26108 17144 26114 17196
rect 26602 17144 26608 17196
rect 26660 17184 26666 17196
rect 26786 17184 26792 17196
rect 26660 17156 26792 17184
rect 26660 17144 26666 17156
rect 26786 17144 26792 17156
rect 26844 17184 26850 17196
rect 27065 17187 27123 17193
rect 27065 17184 27077 17187
rect 26844 17156 27077 17184
rect 26844 17144 26850 17156
rect 27065 17153 27077 17156
rect 27111 17153 27123 17187
rect 27065 17147 27123 17153
rect 31205 17187 31263 17193
rect 31205 17153 31217 17187
rect 31251 17184 31263 17187
rect 31496 17184 31524 17212
rect 31251 17156 31524 17184
rect 31251 17153 31263 17156
rect 31205 17147 31263 17153
rect 31772 17128 31800 17292
rect 31846 17280 31852 17332
rect 31904 17320 31910 17332
rect 33226 17320 33232 17332
rect 31904 17292 33232 17320
rect 31904 17280 31910 17292
rect 33226 17280 33232 17292
rect 33284 17280 33290 17332
rect 36722 17280 36728 17332
rect 36780 17320 36786 17332
rect 37826 17320 37832 17332
rect 36780 17292 37832 17320
rect 36780 17280 36786 17292
rect 37826 17280 37832 17292
rect 37884 17280 37890 17332
rect 39592 17292 41184 17320
rect 33042 17212 33048 17264
rect 33100 17212 33106 17264
rect 37461 17255 37519 17261
rect 37461 17221 37473 17255
rect 37507 17252 37519 17255
rect 37550 17252 37556 17264
rect 37507 17224 37556 17252
rect 37507 17221 37519 17224
rect 37461 17215 37519 17221
rect 37550 17212 37556 17224
rect 37608 17212 37614 17264
rect 37642 17212 37648 17264
rect 37700 17252 37706 17264
rect 39592 17252 39620 17292
rect 37700 17224 39620 17252
rect 37700 17212 37706 17224
rect 39592 17193 39620 17224
rect 39853 17255 39911 17261
rect 39853 17221 39865 17255
rect 39899 17252 39911 17255
rect 39942 17252 39948 17264
rect 39899 17224 39948 17252
rect 39899 17221 39911 17224
rect 39853 17215 39911 17221
rect 39942 17212 39948 17224
rect 40000 17212 40006 17264
rect 40586 17212 40592 17264
rect 40644 17212 40650 17264
rect 41156 17252 41184 17292
rect 41230 17280 41236 17332
rect 41288 17320 41294 17332
rect 41325 17323 41383 17329
rect 41325 17320 41337 17323
rect 41288 17292 41337 17320
rect 41288 17280 41294 17292
rect 41325 17289 41337 17292
rect 41371 17289 41383 17323
rect 41325 17283 41383 17289
rect 42702 17280 42708 17332
rect 42760 17320 42766 17332
rect 43717 17323 43775 17329
rect 43717 17320 43729 17323
rect 42760 17292 43729 17320
rect 42760 17280 42766 17292
rect 43717 17289 43729 17292
rect 43763 17289 43775 17323
rect 47026 17320 47032 17332
rect 43717 17283 43775 17289
rect 44100 17292 47032 17320
rect 41782 17252 41788 17264
rect 41156 17224 41788 17252
rect 41782 17212 41788 17224
rect 41840 17212 41846 17264
rect 44100 17252 44128 17292
rect 42720 17224 44128 17252
rect 39577 17187 39635 17193
rect 39577 17153 39589 17187
rect 39623 17153 39635 17187
rect 39577 17147 39635 17153
rect 42150 17144 42156 17196
rect 42208 17184 42214 17196
rect 42720 17193 42748 17224
rect 44174 17212 44180 17264
rect 44232 17252 44238 17264
rect 44232 17224 45784 17252
rect 44232 17212 44238 17224
rect 42705 17187 42763 17193
rect 42705 17184 42717 17187
rect 42208 17156 42717 17184
rect 42208 17144 42214 17156
rect 42705 17153 42717 17156
rect 42751 17153 42763 17187
rect 42705 17147 42763 17153
rect 44085 17187 44143 17193
rect 44085 17153 44097 17187
rect 44131 17184 44143 17187
rect 45005 17187 45063 17193
rect 44131 17156 44864 17184
rect 44131 17153 44143 17156
rect 44085 17147 44143 17153
rect 12676 17088 14780 17116
rect 12676 17076 12682 17088
rect 14826 17076 14832 17128
rect 14884 17116 14890 17128
rect 15841 17119 15899 17125
rect 15841 17116 15853 17119
rect 14884 17088 15853 17116
rect 14884 17076 14890 17088
rect 15841 17085 15853 17088
rect 15887 17085 15899 17119
rect 15841 17079 15899 17085
rect 17129 17119 17187 17125
rect 17129 17085 17141 17119
rect 17175 17085 17187 17119
rect 17129 17079 17187 17085
rect 18233 17119 18291 17125
rect 18233 17085 18245 17119
rect 18279 17116 18291 17119
rect 18782 17116 18788 17128
rect 18279 17088 18788 17116
rect 18279 17085 18291 17088
rect 18233 17079 18291 17085
rect 11882 17008 11888 17060
rect 11940 17048 11946 17060
rect 13998 17048 14004 17060
rect 11940 17020 14004 17048
rect 11940 17008 11946 17020
rect 13998 17008 14004 17020
rect 14056 17008 14062 17060
rect 14366 17008 14372 17060
rect 14424 17048 14430 17060
rect 14424 17020 16896 17048
rect 14424 17008 14430 17020
rect 12618 16980 12624 16992
rect 12579 16952 12624 16980
rect 12618 16940 12624 16952
rect 12676 16940 12682 16992
rect 13078 16980 13084 16992
rect 13039 16952 13084 16980
rect 13078 16940 13084 16952
rect 13136 16940 13142 16992
rect 14090 16980 14096 16992
rect 14051 16952 14096 16980
rect 14090 16940 14096 16952
rect 14148 16940 14154 16992
rect 14642 16980 14648 16992
rect 14603 16952 14648 16980
rect 14642 16940 14648 16952
rect 14700 16940 14706 16992
rect 15286 16980 15292 16992
rect 15247 16952 15292 16980
rect 15286 16940 15292 16952
rect 15344 16940 15350 16992
rect 15930 16980 15936 16992
rect 15891 16952 15936 16980
rect 15930 16940 15936 16952
rect 15988 16940 15994 16992
rect 16025 16983 16083 16989
rect 16025 16949 16037 16983
rect 16071 16980 16083 16983
rect 16390 16980 16396 16992
rect 16071 16952 16396 16980
rect 16071 16949 16083 16952
rect 16025 16943 16083 16949
rect 16390 16940 16396 16952
rect 16448 16940 16454 16992
rect 16868 16980 16896 17020
rect 17144 16980 17172 17079
rect 18782 17076 18788 17088
rect 18840 17076 18846 17128
rect 18874 17076 18880 17128
rect 18932 17116 18938 17128
rect 18969 17119 19027 17125
rect 18969 17116 18981 17119
rect 18932 17088 18981 17116
rect 18932 17076 18938 17088
rect 18969 17085 18981 17088
rect 19015 17085 19027 17119
rect 18969 17079 19027 17085
rect 19150 17076 19156 17128
rect 19208 17116 19214 17128
rect 19245 17119 19303 17125
rect 19245 17116 19257 17119
rect 19208 17088 19257 17116
rect 19208 17076 19214 17088
rect 19245 17085 19257 17088
rect 19291 17085 19303 17119
rect 19245 17079 19303 17085
rect 17494 17048 17500 17060
rect 17455 17020 17500 17048
rect 17494 17008 17500 17020
rect 17552 17008 17558 17060
rect 18509 17051 18567 17057
rect 18509 17017 18521 17051
rect 18555 17017 18567 17051
rect 19260 17048 19288 17079
rect 19426 17076 19432 17128
rect 19484 17125 19490 17128
rect 19484 17119 19512 17125
rect 19500 17085 19512 17119
rect 19484 17079 19512 17085
rect 19484 17076 19490 17079
rect 19610 17076 19616 17128
rect 19668 17116 19674 17128
rect 21269 17119 21327 17125
rect 19668 17088 20484 17116
rect 19668 17076 19674 17088
rect 19794 17048 19800 17060
rect 19260 17020 19800 17048
rect 18509 17011 18567 17017
rect 16868 16952 17172 16980
rect 18524 16980 18552 17011
rect 19794 17008 19800 17020
rect 19852 17008 19858 17060
rect 18690 16980 18696 16992
rect 18524 16952 18696 16980
rect 18690 16940 18696 16952
rect 18748 16940 18754 16992
rect 19610 16980 19616 16992
rect 19571 16952 19616 16980
rect 19610 16940 19616 16952
rect 19668 16940 19674 16992
rect 20165 16983 20223 16989
rect 20165 16949 20177 16983
rect 20211 16980 20223 16983
rect 20346 16980 20352 16992
rect 20211 16952 20352 16980
rect 20211 16949 20223 16952
rect 20165 16943 20223 16949
rect 20346 16940 20352 16952
rect 20404 16940 20410 16992
rect 20456 16980 20484 17088
rect 21269 17085 21281 17119
rect 21315 17116 21327 17119
rect 22370 17116 22376 17128
rect 21315 17088 22376 17116
rect 21315 17085 21327 17088
rect 21269 17079 21327 17085
rect 21284 16980 21312 17079
rect 22370 17076 22376 17088
rect 22428 17076 22434 17128
rect 22465 17119 22523 17125
rect 22465 17085 22477 17119
rect 22511 17116 22523 17119
rect 23290 17116 23296 17128
rect 22511 17088 23296 17116
rect 22511 17085 22523 17088
rect 22465 17079 22523 17085
rect 23290 17076 23296 17088
rect 23348 17076 23354 17128
rect 24213 17119 24271 17125
rect 24213 17085 24225 17119
rect 24259 17116 24271 17119
rect 28534 17116 28540 17128
rect 24259 17088 28540 17116
rect 24259 17085 24271 17088
rect 24213 17079 24271 17085
rect 28534 17076 28540 17088
rect 28592 17076 28598 17128
rect 30929 17119 30987 17125
rect 30929 17085 30941 17119
rect 30975 17116 30987 17119
rect 31662 17116 31668 17128
rect 30975 17088 31668 17116
rect 30975 17085 30987 17088
rect 30929 17079 30987 17085
rect 31662 17076 31668 17088
rect 31720 17076 31726 17128
rect 31754 17076 31760 17128
rect 31812 17116 31818 17128
rect 32125 17119 32183 17125
rect 32125 17116 32137 17119
rect 31812 17088 32137 17116
rect 31812 17076 31818 17088
rect 32125 17085 32137 17088
rect 32171 17085 32183 17119
rect 32401 17119 32459 17125
rect 32401 17116 32413 17119
rect 32125 17079 32183 17085
rect 32232 17088 32413 17116
rect 21910 17048 21916 17060
rect 21871 17020 21916 17048
rect 21910 17008 21916 17020
rect 21968 17008 21974 17060
rect 28902 17008 28908 17060
rect 28960 17048 28966 17060
rect 28960 17020 29592 17048
rect 28960 17008 28966 17020
rect 20456 16952 21312 16980
rect 21634 16940 21640 16992
rect 21692 16980 21698 16992
rect 26234 16980 26240 16992
rect 21692 16952 26240 16980
rect 21692 16940 21698 16952
rect 26234 16940 26240 16952
rect 26292 16940 26298 16992
rect 26421 16983 26479 16989
rect 26421 16949 26433 16983
rect 26467 16980 26479 16983
rect 29270 16980 29276 16992
rect 26467 16952 29276 16980
rect 26467 16949 26479 16952
rect 26421 16943 26479 16949
rect 29270 16940 29276 16952
rect 29328 16940 29334 16992
rect 29454 16980 29460 16992
rect 29415 16952 29460 16980
rect 29454 16940 29460 16952
rect 29512 16940 29518 16992
rect 29564 16980 29592 17020
rect 31386 17008 31392 17060
rect 31444 17048 31450 17060
rect 31444 17020 31984 17048
rect 31444 17008 31450 17020
rect 31846 16980 31852 16992
rect 29564 16952 31852 16980
rect 31846 16940 31852 16952
rect 31904 16940 31910 16992
rect 31956 16980 31984 17020
rect 32232 16980 32260 17088
rect 32401 17085 32413 17088
rect 32447 17085 32459 17119
rect 32401 17079 32459 17085
rect 34330 17076 34336 17128
rect 34388 17116 34394 17128
rect 34425 17119 34483 17125
rect 34425 17116 34437 17119
rect 34388 17088 34437 17116
rect 34388 17076 34394 17088
rect 34425 17085 34437 17088
rect 34471 17085 34483 17119
rect 34425 17079 34483 17085
rect 34609 17119 34667 17125
rect 34609 17085 34621 17119
rect 34655 17116 34667 17119
rect 34882 17116 34888 17128
rect 34655 17088 34888 17116
rect 34655 17085 34667 17088
rect 34609 17079 34667 17085
rect 34882 17076 34888 17088
rect 34940 17076 34946 17128
rect 34977 17119 35035 17125
rect 34977 17085 34989 17119
rect 35023 17085 35035 17119
rect 34977 17079 35035 17085
rect 37277 17119 37335 17125
rect 37277 17085 37289 17119
rect 37323 17116 37335 17119
rect 37550 17116 37556 17128
rect 37323 17088 37556 17116
rect 37323 17085 37335 17088
rect 37277 17079 37335 17085
rect 33962 17008 33968 17060
rect 34020 17048 34026 17060
rect 34992 17048 35020 17079
rect 37550 17076 37556 17088
rect 37608 17116 37614 17128
rect 39022 17116 39028 17128
rect 37608 17088 39028 17116
rect 37608 17076 37614 17088
rect 39022 17076 39028 17088
rect 39080 17076 39086 17128
rect 39117 17119 39175 17125
rect 39117 17085 39129 17119
rect 39163 17116 39175 17119
rect 39298 17116 39304 17128
rect 39163 17088 39304 17116
rect 39163 17085 39175 17088
rect 39117 17079 39175 17085
rect 39298 17076 39304 17088
rect 39356 17076 39362 17128
rect 42429 17119 42487 17125
rect 42429 17116 42441 17119
rect 39684 17088 42441 17116
rect 34020 17020 35020 17048
rect 34020 17008 34026 17020
rect 35802 17008 35808 17060
rect 35860 17048 35866 17060
rect 38102 17048 38108 17060
rect 35860 17020 38108 17048
rect 35860 17008 35866 17020
rect 38102 17008 38108 17020
rect 38160 17008 38166 17060
rect 39040 17048 39068 17076
rect 39684 17048 39712 17088
rect 42429 17085 42441 17088
rect 42475 17085 42487 17119
rect 43990 17116 43996 17128
rect 43951 17088 43996 17116
rect 42429 17079 42487 17085
rect 43990 17076 43996 17088
rect 44048 17076 44054 17128
rect 44174 17076 44180 17128
rect 44232 17116 44238 17128
rect 44729 17119 44787 17125
rect 44729 17116 44741 17119
rect 44232 17088 44741 17116
rect 44232 17076 44238 17088
rect 44729 17085 44741 17088
rect 44775 17085 44787 17119
rect 44836 17116 44864 17156
rect 45005 17153 45017 17187
rect 45051 17184 45063 17187
rect 45278 17184 45284 17196
rect 45051 17156 45284 17184
rect 45051 17153 45063 17156
rect 45005 17147 45063 17153
rect 45278 17144 45284 17156
rect 45336 17144 45342 17196
rect 45756 17193 45784 17224
rect 45940 17193 45968 17292
rect 47026 17280 47032 17292
rect 47084 17280 47090 17332
rect 48130 17280 48136 17332
rect 48188 17320 48194 17332
rect 50341 17323 50399 17329
rect 50341 17320 50353 17323
rect 48188 17292 50353 17320
rect 48188 17280 48194 17292
rect 50341 17289 50353 17292
rect 50387 17289 50399 17323
rect 50341 17283 50399 17289
rect 46014 17212 46020 17264
rect 46072 17252 46078 17264
rect 48590 17252 48596 17264
rect 46072 17224 48596 17252
rect 46072 17212 46078 17224
rect 48590 17212 48596 17224
rect 48648 17252 48654 17264
rect 49237 17255 49295 17261
rect 49237 17252 49249 17255
rect 48648 17224 49249 17252
rect 48648 17212 48654 17224
rect 49237 17221 49249 17224
rect 49283 17252 49295 17255
rect 49602 17252 49608 17264
rect 49283 17224 49608 17252
rect 49283 17221 49295 17224
rect 49237 17215 49295 17221
rect 49602 17212 49608 17224
rect 49660 17252 49666 17264
rect 49789 17255 49847 17261
rect 49789 17252 49801 17255
rect 49660 17224 49801 17252
rect 49660 17212 49666 17224
rect 49789 17221 49801 17224
rect 49835 17221 49847 17255
rect 49789 17215 49847 17221
rect 45649 17187 45707 17193
rect 45649 17153 45661 17187
rect 45695 17153 45707 17187
rect 45649 17147 45707 17153
rect 45741 17187 45799 17193
rect 45741 17153 45753 17187
rect 45787 17153 45799 17187
rect 45741 17147 45799 17153
rect 45925 17187 45983 17193
rect 45925 17153 45937 17187
rect 45971 17153 45983 17187
rect 45925 17147 45983 17153
rect 45094 17116 45100 17128
rect 44836 17088 45100 17116
rect 44729 17079 44787 17085
rect 45094 17076 45100 17088
rect 45152 17076 45158 17128
rect 42610 17048 42616 17060
rect 39040 17020 39712 17048
rect 41386 17020 42616 17048
rect 31956 16952 32260 16980
rect 32766 16940 32772 16992
rect 32824 16980 32830 16992
rect 32950 16980 32956 16992
rect 32824 16952 32956 16980
rect 32824 16940 32830 16952
rect 32950 16940 32956 16952
rect 33008 16980 33014 16992
rect 33873 16983 33931 16989
rect 33873 16980 33885 16983
rect 33008 16952 33885 16980
rect 33008 16940 33014 16952
rect 33873 16949 33885 16952
rect 33919 16949 33931 16983
rect 33873 16943 33931 16949
rect 34146 16940 34152 16992
rect 34204 16980 34210 16992
rect 38286 16980 38292 16992
rect 34204 16952 38292 16980
rect 34204 16940 34210 16952
rect 38286 16940 38292 16952
rect 38344 16940 38350 16992
rect 38654 16940 38660 16992
rect 38712 16980 38718 16992
rect 41386 16980 41414 17020
rect 42610 17008 42616 17020
rect 42668 17008 42674 17060
rect 43254 17008 43260 17060
rect 43312 17048 43318 17060
rect 45664 17048 45692 17147
rect 45756 17116 45784 17147
rect 46198 17144 46204 17196
rect 46256 17184 46262 17196
rect 46569 17187 46627 17193
rect 46569 17184 46581 17187
rect 46256 17156 46581 17184
rect 46256 17144 46262 17156
rect 46569 17153 46581 17156
rect 46615 17184 46627 17187
rect 46615 17156 48820 17184
rect 46615 17153 46627 17156
rect 46569 17147 46627 17153
rect 47581 17119 47639 17125
rect 47581 17116 47593 17119
rect 45756 17088 47593 17116
rect 47581 17085 47593 17088
rect 47627 17085 47639 17119
rect 47581 17079 47639 17085
rect 48133 17051 48191 17057
rect 48133 17048 48145 17051
rect 43312 17020 48145 17048
rect 43312 17008 43318 17020
rect 48133 17017 48145 17020
rect 48179 17017 48191 17051
rect 48133 17011 48191 17017
rect 38712 16952 41414 16980
rect 38712 16940 38718 16952
rect 41506 16940 41512 16992
rect 41564 16980 41570 16992
rect 41785 16983 41843 16989
rect 41785 16980 41797 16983
rect 41564 16952 41797 16980
rect 41564 16940 41570 16952
rect 41785 16949 41797 16952
rect 41831 16980 41843 16983
rect 41874 16980 41880 16992
rect 41831 16952 41880 16980
rect 41831 16949 41843 16952
rect 41785 16943 41843 16949
rect 41874 16940 41880 16952
rect 41932 16940 41938 16992
rect 44821 16983 44879 16989
rect 44821 16949 44833 16983
rect 44867 16980 44879 16983
rect 44910 16980 44916 16992
rect 44867 16952 44916 16980
rect 44867 16949 44879 16952
rect 44821 16943 44879 16949
rect 44910 16940 44916 16952
rect 44968 16940 44974 16992
rect 45186 16980 45192 16992
rect 45147 16952 45192 16980
rect 45186 16940 45192 16952
rect 45244 16940 45250 16992
rect 45646 16980 45652 16992
rect 45607 16952 45652 16980
rect 45646 16940 45652 16952
rect 45704 16940 45710 16992
rect 46474 16980 46480 16992
rect 46435 16952 46480 16980
rect 46474 16940 46480 16952
rect 46532 16940 46538 16992
rect 48792 16989 48820 17156
rect 48777 16983 48835 16989
rect 48777 16949 48789 16983
rect 48823 16980 48835 16983
rect 48958 16980 48964 16992
rect 48823 16952 48964 16980
rect 48823 16949 48835 16952
rect 48777 16943 48835 16949
rect 48958 16940 48964 16952
rect 49016 16940 49022 16992
rect 1104 16890 58880 16912
rect 1104 16838 10582 16890
rect 10634 16838 10646 16890
rect 10698 16838 10710 16890
rect 10762 16838 10774 16890
rect 10826 16838 10838 16890
rect 10890 16838 29846 16890
rect 29898 16838 29910 16890
rect 29962 16838 29974 16890
rect 30026 16838 30038 16890
rect 30090 16838 30102 16890
rect 30154 16838 49110 16890
rect 49162 16838 49174 16890
rect 49226 16838 49238 16890
rect 49290 16838 49302 16890
rect 49354 16838 49366 16890
rect 49418 16838 58880 16890
rect 1104 16816 58880 16838
rect 11882 16776 11888 16788
rect 11843 16748 11888 16776
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 12437 16779 12495 16785
rect 12437 16745 12449 16779
rect 12483 16776 12495 16779
rect 14090 16776 14096 16788
rect 12483 16748 14096 16776
rect 12483 16745 12495 16748
rect 12437 16739 12495 16745
rect 14090 16736 14096 16748
rect 14148 16736 14154 16788
rect 14642 16776 14648 16788
rect 14200 16748 14648 16776
rect 12989 16711 13047 16717
rect 12989 16677 13001 16711
rect 13035 16708 13047 16711
rect 14200 16708 14228 16748
rect 14642 16736 14648 16748
rect 14700 16736 14706 16788
rect 14829 16779 14887 16785
rect 14829 16745 14841 16779
rect 14875 16776 14887 16779
rect 14918 16776 14924 16788
rect 14875 16748 14924 16776
rect 14875 16745 14887 16748
rect 14829 16739 14887 16745
rect 14918 16736 14924 16748
rect 14976 16736 14982 16788
rect 15378 16776 15384 16788
rect 15339 16748 15384 16776
rect 15378 16736 15384 16748
rect 15436 16736 15442 16788
rect 16577 16779 16635 16785
rect 16577 16745 16589 16779
rect 16623 16776 16635 16779
rect 16666 16776 16672 16788
rect 16623 16748 16672 16776
rect 16623 16745 16635 16748
rect 16577 16739 16635 16745
rect 16666 16736 16672 16748
rect 16724 16736 16730 16788
rect 19426 16776 19432 16788
rect 16776 16748 19432 16776
rect 16776 16720 16804 16748
rect 19426 16736 19432 16748
rect 19484 16736 19490 16788
rect 20438 16736 20444 16788
rect 20496 16776 20502 16788
rect 20898 16776 20904 16788
rect 20496 16748 20904 16776
rect 20496 16736 20502 16748
rect 20898 16736 20904 16748
rect 20956 16736 20962 16788
rect 22186 16736 22192 16788
rect 22244 16776 22250 16788
rect 22244 16748 24900 16776
rect 22244 16736 22250 16748
rect 13035 16680 14228 16708
rect 14277 16711 14335 16717
rect 13035 16677 13047 16680
rect 12989 16671 13047 16677
rect 14277 16677 14289 16711
rect 14323 16708 14335 16711
rect 16758 16708 16764 16720
rect 14323 16680 16764 16708
rect 14323 16677 14335 16680
rect 14277 16671 14335 16677
rect 16758 16668 16764 16680
rect 16816 16668 16822 16720
rect 16942 16668 16948 16720
rect 17000 16708 17006 16720
rect 17681 16711 17739 16717
rect 17681 16708 17693 16711
rect 17000 16680 17693 16708
rect 17000 16668 17006 16680
rect 17681 16677 17693 16680
rect 17727 16677 17739 16711
rect 18690 16708 18696 16720
rect 18651 16680 18696 16708
rect 17681 16671 17739 16677
rect 18690 16668 18696 16680
rect 18748 16668 18754 16720
rect 18874 16668 18880 16720
rect 18932 16708 18938 16720
rect 20530 16708 20536 16720
rect 18932 16680 20536 16708
rect 18932 16668 18938 16680
rect 13541 16643 13599 16649
rect 13541 16609 13553 16643
rect 13587 16640 13599 16643
rect 14826 16640 14832 16652
rect 13587 16612 14832 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 14826 16600 14832 16612
rect 14884 16600 14890 16652
rect 16666 16600 16672 16652
rect 16724 16640 16730 16652
rect 17221 16643 17279 16649
rect 17221 16640 17233 16643
rect 16724 16612 17233 16640
rect 16724 16600 16730 16612
rect 17221 16609 17233 16612
rect 17267 16609 17279 16643
rect 17221 16603 17279 16609
rect 18417 16643 18475 16649
rect 18417 16609 18429 16643
rect 18463 16640 18475 16643
rect 18463 16612 19196 16640
rect 18463 16609 18475 16612
rect 18417 16603 18475 16609
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16572 1731 16575
rect 13078 16572 13084 16584
rect 1719 16544 13084 16572
rect 1719 16541 1731 16544
rect 1673 16535 1731 16541
rect 13078 16532 13084 16544
rect 13136 16532 13142 16584
rect 15838 16572 15844 16584
rect 15799 16544 15844 16572
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 15933 16575 15991 16581
rect 15933 16541 15945 16575
rect 15979 16572 15991 16575
rect 16022 16572 16028 16584
rect 15979 16544 16028 16572
rect 15979 16541 15991 16544
rect 15933 16535 15991 16541
rect 16022 16532 16028 16544
rect 16080 16532 16086 16584
rect 16298 16532 16304 16584
rect 16356 16572 16362 16584
rect 16482 16572 16488 16584
rect 16356 16544 16488 16572
rect 16356 16532 16362 16544
rect 16482 16532 16488 16544
rect 16540 16532 16546 16584
rect 17310 16572 17316 16584
rect 17271 16544 17316 16572
rect 17310 16532 17316 16544
rect 17368 16532 17374 16584
rect 18325 16575 18383 16581
rect 18325 16541 18337 16575
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 15194 16464 15200 16516
rect 15252 16504 15258 16516
rect 15746 16504 15752 16516
rect 15252 16476 15752 16504
rect 15252 16464 15258 16476
rect 15746 16464 15752 16476
rect 15804 16504 15810 16516
rect 18340 16504 18368 16535
rect 15804 16476 18368 16504
rect 19168 16504 19196 16612
rect 19260 16572 19288 16680
rect 20530 16668 20536 16680
rect 20588 16668 20594 16720
rect 20714 16668 20720 16720
rect 20772 16708 20778 16720
rect 22204 16708 22232 16736
rect 20772 16680 22232 16708
rect 24872 16708 24900 16748
rect 24946 16736 24952 16788
rect 25004 16776 25010 16788
rect 29086 16776 29092 16788
rect 25004 16748 29092 16776
rect 25004 16736 25010 16748
rect 29086 16736 29092 16748
rect 29144 16736 29150 16788
rect 29270 16736 29276 16788
rect 29328 16776 29334 16788
rect 31386 16776 31392 16788
rect 29328 16748 31392 16776
rect 29328 16736 29334 16748
rect 31386 16736 31392 16748
rect 31444 16736 31450 16788
rect 33134 16736 33140 16788
rect 33192 16776 33198 16788
rect 33778 16776 33784 16788
rect 33192 16748 33784 16776
rect 33192 16736 33198 16748
rect 33778 16736 33784 16748
rect 33836 16776 33842 16788
rect 33965 16779 34023 16785
rect 33965 16776 33977 16779
rect 33836 16748 33977 16776
rect 33836 16736 33842 16748
rect 33965 16745 33977 16748
rect 34011 16745 34023 16779
rect 37642 16776 37648 16788
rect 33965 16739 34023 16745
rect 37016 16748 37648 16776
rect 24872 16680 25084 16708
rect 20772 16668 20778 16680
rect 19334 16600 19340 16652
rect 19392 16640 19398 16652
rect 19914 16643 19972 16649
rect 19914 16640 19926 16643
rect 19392 16612 19926 16640
rect 19392 16600 19398 16612
rect 19914 16609 19926 16612
rect 19960 16609 19972 16643
rect 21634 16640 21640 16652
rect 19914 16603 19972 16609
rect 20180 16612 20668 16640
rect 21595 16612 21640 16640
rect 19429 16575 19487 16581
rect 19429 16572 19441 16575
rect 19260 16544 19441 16572
rect 19429 16541 19441 16544
rect 19475 16541 19487 16575
rect 19429 16535 19487 16541
rect 19705 16575 19763 16581
rect 19705 16541 19717 16575
rect 19751 16572 19763 16575
rect 19794 16572 19800 16584
rect 19751 16544 19800 16572
rect 19751 16541 19763 16544
rect 19705 16535 19763 16541
rect 19794 16532 19800 16544
rect 19852 16532 19858 16584
rect 19334 16504 19340 16516
rect 19168 16476 19340 16504
rect 15804 16464 15810 16476
rect 19334 16464 19340 16476
rect 19392 16464 19398 16516
rect 20180 16504 20208 16612
rect 20640 16572 20668 16612
rect 21634 16600 21640 16612
rect 21692 16600 21698 16652
rect 21726 16600 21732 16652
rect 21784 16640 21790 16652
rect 23934 16640 23940 16652
rect 21784 16612 23940 16640
rect 21784 16600 21790 16612
rect 23934 16600 23940 16612
rect 23992 16600 23998 16652
rect 24946 16640 24952 16652
rect 24907 16612 24952 16640
rect 24946 16600 24952 16612
rect 25004 16600 25010 16652
rect 25056 16640 25084 16680
rect 27522 16668 27528 16720
rect 27580 16708 27586 16720
rect 28994 16708 29000 16720
rect 27580 16680 29000 16708
rect 27580 16668 27586 16680
rect 28994 16668 29000 16680
rect 29052 16668 29058 16720
rect 29178 16668 29184 16720
rect 29236 16708 29242 16720
rect 29914 16708 29920 16720
rect 29236 16680 29920 16708
rect 29236 16668 29242 16680
rect 29914 16668 29920 16680
rect 29972 16668 29978 16720
rect 31754 16668 31760 16720
rect 31812 16708 31818 16720
rect 31812 16680 32260 16708
rect 31812 16668 31818 16680
rect 25590 16640 25596 16652
rect 25056 16612 25596 16640
rect 25590 16600 25596 16612
rect 25648 16600 25654 16652
rect 25958 16600 25964 16652
rect 26016 16640 26022 16652
rect 27798 16640 27804 16652
rect 26016 16612 27804 16640
rect 26016 16600 26022 16612
rect 27798 16600 27804 16612
rect 27856 16600 27862 16652
rect 20809 16575 20867 16581
rect 20809 16572 20821 16575
rect 20640 16544 20821 16572
rect 20809 16541 20821 16544
rect 20855 16541 20867 16575
rect 21174 16572 21180 16584
rect 21135 16544 21180 16572
rect 20809 16535 20867 16541
rect 21174 16532 21180 16544
rect 21232 16532 21238 16584
rect 21266 16532 21272 16584
rect 21324 16572 21330 16584
rect 22002 16572 22008 16584
rect 21324 16544 22008 16572
rect 21324 16532 21330 16544
rect 22002 16532 22008 16544
rect 22060 16532 22066 16584
rect 22097 16575 22155 16581
rect 22097 16541 22109 16575
rect 22143 16541 22155 16575
rect 22097 16535 22155 16541
rect 19720 16476 20208 16504
rect 19720 16448 19748 16476
rect 20254 16464 20260 16516
rect 20312 16464 20318 16516
rect 20346 16464 20352 16516
rect 20404 16504 20410 16516
rect 21542 16504 21548 16516
rect 20404 16476 21548 16504
rect 20404 16464 20410 16476
rect 21542 16464 21548 16476
rect 21600 16464 21606 16516
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 14642 16396 14648 16448
rect 14700 16436 14706 16448
rect 18874 16436 18880 16448
rect 14700 16408 18880 16436
rect 14700 16396 14706 16408
rect 18874 16396 18880 16408
rect 18932 16396 18938 16448
rect 19702 16396 19708 16448
rect 19760 16396 19766 16448
rect 19794 16396 19800 16448
rect 19852 16436 19858 16448
rect 20070 16436 20076 16448
rect 19852 16408 19897 16436
rect 20031 16408 20076 16436
rect 19852 16396 19858 16408
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 20272 16436 20300 16464
rect 21266 16436 21272 16448
rect 20272 16408 21272 16436
rect 21266 16396 21272 16408
rect 21324 16396 21330 16448
rect 22112 16436 22140 16535
rect 23750 16532 23756 16584
rect 23808 16572 23814 16584
rect 24489 16575 24547 16581
rect 24489 16572 24501 16575
rect 23808 16544 24501 16572
rect 23808 16532 23814 16544
rect 24489 16541 24501 16544
rect 24535 16572 24547 16575
rect 24670 16572 24676 16584
rect 24535 16544 24676 16572
rect 24535 16541 24547 16544
rect 24489 16535 24547 16541
rect 24670 16532 24676 16544
rect 24728 16532 24734 16584
rect 27154 16572 27160 16584
rect 27115 16544 27160 16572
rect 27154 16532 27160 16544
rect 27212 16532 27218 16584
rect 29012 16581 29040 16668
rect 29086 16600 29092 16652
rect 29144 16640 29150 16652
rect 31846 16640 31852 16652
rect 29144 16612 31852 16640
rect 29144 16600 29150 16612
rect 31846 16600 31852 16612
rect 31904 16600 31910 16652
rect 32232 16649 32260 16680
rect 33870 16668 33876 16720
rect 33928 16708 33934 16720
rect 35434 16708 35440 16720
rect 33928 16680 35440 16708
rect 33928 16668 33934 16680
rect 35434 16668 35440 16680
rect 35492 16668 35498 16720
rect 32217 16643 32275 16649
rect 32217 16609 32229 16643
rect 32263 16609 32275 16643
rect 32217 16603 32275 16609
rect 34698 16600 34704 16652
rect 34756 16640 34762 16652
rect 34756 16612 34801 16640
rect 34756 16600 34762 16612
rect 35066 16600 35072 16652
rect 35124 16640 35130 16652
rect 35161 16643 35219 16649
rect 35161 16640 35173 16643
rect 35124 16612 35173 16640
rect 35124 16600 35130 16612
rect 35161 16609 35173 16612
rect 35207 16609 35219 16643
rect 35161 16603 35219 16609
rect 28997 16575 29055 16581
rect 28997 16541 29009 16575
rect 29043 16541 29055 16575
rect 28997 16535 29055 16541
rect 29546 16532 29552 16584
rect 29604 16572 29610 16584
rect 29917 16575 29975 16581
rect 29917 16572 29929 16575
rect 29604 16544 29929 16572
rect 29604 16532 29610 16544
rect 29917 16541 29929 16544
rect 29963 16541 29975 16575
rect 30285 16575 30343 16581
rect 30285 16572 30297 16575
rect 29917 16535 29975 16541
rect 30005 16544 30297 16572
rect 22278 16464 22284 16516
rect 22336 16504 22342 16516
rect 22373 16507 22431 16513
rect 22373 16504 22385 16507
rect 22336 16476 22385 16504
rect 22336 16464 22342 16476
rect 22373 16473 22385 16476
rect 22419 16473 22431 16507
rect 25130 16504 25136 16516
rect 23598 16476 25136 16504
rect 22373 16467 22431 16473
rect 25130 16464 25136 16476
rect 25188 16464 25194 16516
rect 25225 16507 25283 16513
rect 25225 16473 25237 16507
rect 25271 16473 25283 16507
rect 26450 16476 27108 16504
rect 25225 16467 25283 16473
rect 22554 16436 22560 16448
rect 22112 16408 22560 16436
rect 22554 16396 22560 16408
rect 22612 16396 22618 16448
rect 23842 16436 23848 16448
rect 23803 16408 23848 16436
rect 23842 16396 23848 16408
rect 23900 16396 23906 16448
rect 23934 16396 23940 16448
rect 23992 16436 23998 16448
rect 25240 16436 25268 16467
rect 26694 16436 26700 16448
rect 23992 16408 25268 16436
rect 26655 16408 26700 16436
rect 23992 16396 23998 16408
rect 26694 16396 26700 16408
rect 26752 16396 26758 16448
rect 27080 16436 27108 16476
rect 28718 16464 28724 16516
rect 28776 16504 28782 16516
rect 28813 16507 28871 16513
rect 28813 16504 28825 16507
rect 28776 16476 28825 16504
rect 28776 16464 28782 16476
rect 28813 16473 28825 16476
rect 28859 16473 28871 16507
rect 28813 16467 28871 16473
rect 29270 16464 29276 16516
rect 29328 16504 29334 16516
rect 30005 16504 30033 16544
rect 30285 16541 30297 16544
rect 30331 16541 30343 16575
rect 30285 16535 30343 16541
rect 31202 16532 31208 16584
rect 31260 16572 31266 16584
rect 31711 16575 31769 16581
rect 31711 16572 31723 16575
rect 31260 16544 31723 16572
rect 31260 16532 31266 16544
rect 31711 16541 31723 16544
rect 31757 16541 31769 16575
rect 31711 16535 31769 16541
rect 36446 16532 36452 16584
rect 36504 16572 36510 16584
rect 37016 16581 37044 16748
rect 37642 16736 37648 16748
rect 37700 16736 37706 16788
rect 38838 16736 38844 16788
rect 38896 16776 38902 16788
rect 42153 16779 42211 16785
rect 42153 16776 42165 16779
rect 38896 16748 42165 16776
rect 38896 16736 38902 16748
rect 42153 16745 42165 16748
rect 42199 16745 42211 16779
rect 44266 16776 44272 16788
rect 44227 16748 44272 16776
rect 42153 16739 42211 16745
rect 44266 16736 44272 16748
rect 44324 16736 44330 16788
rect 45278 16736 45284 16788
rect 45336 16776 45342 16788
rect 45738 16776 45744 16788
rect 45336 16748 45744 16776
rect 45336 16736 45342 16748
rect 45738 16736 45744 16748
rect 45796 16776 45802 16788
rect 47489 16779 47547 16785
rect 47489 16776 47501 16779
rect 45796 16748 47501 16776
rect 45796 16736 45802 16748
rect 47489 16745 47501 16748
rect 47535 16745 47547 16779
rect 48682 16776 48688 16788
rect 48643 16748 48688 16776
rect 47489 16739 47547 16745
rect 48682 16736 48688 16748
rect 48740 16736 48746 16788
rect 49602 16736 49608 16788
rect 49660 16776 49666 16788
rect 50157 16779 50215 16785
rect 50157 16776 50169 16779
rect 49660 16748 50169 16776
rect 49660 16736 49666 16748
rect 50157 16745 50169 16748
rect 50203 16745 50215 16779
rect 50157 16739 50215 16745
rect 38930 16668 38936 16720
rect 38988 16708 38994 16720
rect 39209 16711 39267 16717
rect 39209 16708 39221 16711
rect 38988 16680 39221 16708
rect 38988 16668 38994 16680
rect 39209 16677 39221 16680
rect 39255 16677 39267 16711
rect 39209 16671 39267 16677
rect 39853 16711 39911 16717
rect 39853 16677 39865 16711
rect 39899 16677 39911 16711
rect 39853 16671 39911 16677
rect 37274 16640 37280 16652
rect 37235 16612 37280 16640
rect 37274 16600 37280 16612
rect 37332 16600 37338 16652
rect 37642 16600 37648 16652
rect 37700 16640 37706 16652
rect 39868 16640 39896 16671
rect 41598 16668 41604 16720
rect 41656 16708 41662 16720
rect 43070 16708 43076 16720
rect 41656 16680 42472 16708
rect 43031 16680 43076 16708
rect 41656 16668 41662 16680
rect 37700 16612 39252 16640
rect 37700 16600 37706 16612
rect 39224 16584 39252 16612
rect 39684 16612 39896 16640
rect 41325 16643 41383 16649
rect 37001 16575 37059 16581
rect 37001 16572 37013 16575
rect 36504 16544 37013 16572
rect 36504 16532 36510 16544
rect 37001 16541 37013 16544
rect 37047 16541 37059 16575
rect 37001 16535 37059 16541
rect 39206 16532 39212 16584
rect 39264 16532 39270 16584
rect 31478 16504 31484 16516
rect 29328 16476 30033 16504
rect 31326 16476 31484 16504
rect 29328 16464 29334 16476
rect 31478 16464 31484 16476
rect 31536 16464 31542 16516
rect 32490 16504 32496 16516
rect 32451 16476 32496 16504
rect 32490 16464 32496 16476
rect 32548 16464 32554 16516
rect 32950 16464 32956 16516
rect 33008 16464 33014 16516
rect 34514 16464 34520 16516
rect 34572 16504 34578 16516
rect 34885 16507 34943 16513
rect 34885 16504 34897 16507
rect 34572 16476 34897 16504
rect 34572 16464 34578 16476
rect 34885 16473 34897 16476
rect 34931 16473 34943 16507
rect 34885 16467 34943 16473
rect 35250 16464 35256 16516
rect 35308 16504 35314 16516
rect 39684 16504 39712 16612
rect 41325 16609 41337 16643
rect 41371 16640 41383 16643
rect 41966 16640 41972 16652
rect 41371 16612 41972 16640
rect 41371 16609 41383 16612
rect 41325 16603 41383 16609
rect 41966 16600 41972 16612
rect 42024 16600 42030 16652
rect 42242 16600 42248 16652
rect 42300 16640 42306 16652
rect 42337 16643 42395 16649
rect 42337 16640 42349 16643
rect 42300 16612 42349 16640
rect 42300 16600 42306 16612
rect 42337 16609 42349 16612
rect 42383 16609 42395 16643
rect 42444 16640 42472 16680
rect 43070 16668 43076 16680
rect 43128 16668 43134 16720
rect 44634 16708 44640 16720
rect 44376 16680 44640 16708
rect 44376 16649 44404 16680
rect 44634 16668 44640 16680
rect 44692 16708 44698 16720
rect 46937 16711 46995 16717
rect 46937 16708 46949 16711
rect 44692 16680 46949 16708
rect 44692 16668 44698 16680
rect 46937 16677 46949 16680
rect 46983 16677 46995 16711
rect 46937 16671 46995 16677
rect 43349 16643 43407 16649
rect 43349 16640 43361 16643
rect 42444 16612 43361 16640
rect 42337 16603 42395 16609
rect 43349 16609 43361 16612
rect 43395 16609 43407 16643
rect 43349 16603 43407 16609
rect 44361 16643 44419 16649
rect 44361 16609 44373 16643
rect 44407 16609 44419 16643
rect 45002 16640 45008 16652
rect 44963 16612 45008 16640
rect 44361 16603 44419 16609
rect 45002 16600 45008 16612
rect 45060 16600 45066 16652
rect 46385 16643 46443 16649
rect 46385 16640 46397 16643
rect 45572 16612 46397 16640
rect 41601 16575 41659 16581
rect 41601 16541 41613 16575
rect 41647 16572 41659 16575
rect 41782 16572 41788 16584
rect 41647 16544 41788 16572
rect 41647 16541 41659 16544
rect 41601 16535 41659 16541
rect 41782 16532 41788 16544
rect 41840 16532 41846 16584
rect 42429 16575 42487 16581
rect 42429 16541 42441 16575
rect 42475 16541 42487 16575
rect 42429 16535 42487 16541
rect 35308 16476 37766 16504
rect 38580 16476 39712 16504
rect 35308 16464 35314 16476
rect 33870 16436 33876 16448
rect 27080 16408 33876 16436
rect 33870 16396 33876 16408
rect 33928 16396 33934 16448
rect 34330 16396 34336 16448
rect 34388 16436 34394 16448
rect 38580 16436 38608 16476
rect 40586 16464 40592 16516
rect 40644 16464 40650 16516
rect 41414 16464 41420 16516
rect 41472 16504 41478 16516
rect 42444 16504 42472 16535
rect 42702 16532 42708 16584
rect 42760 16572 42766 16584
rect 43441 16575 43499 16581
rect 43441 16572 43453 16575
rect 42760 16544 43453 16572
rect 42760 16532 42766 16544
rect 43441 16541 43453 16544
rect 43487 16541 43499 16575
rect 43441 16535 43499 16541
rect 44453 16575 44511 16581
rect 44453 16541 44465 16575
rect 44499 16572 44511 16575
rect 44542 16572 44548 16584
rect 44499 16544 44548 16572
rect 44499 16541 44511 16544
rect 44453 16535 44511 16541
rect 44542 16532 44548 16544
rect 44600 16532 44606 16584
rect 45097 16575 45155 16581
rect 45097 16541 45109 16575
rect 45143 16572 45155 16575
rect 45572 16572 45600 16612
rect 46385 16609 46397 16612
rect 46431 16640 46443 16643
rect 48041 16643 48099 16649
rect 48041 16640 48053 16643
rect 46431 16612 48053 16640
rect 46431 16609 46443 16612
rect 46385 16603 46443 16609
rect 48041 16609 48053 16612
rect 48087 16609 48099 16643
rect 48041 16603 48099 16609
rect 45143 16544 45600 16572
rect 45925 16575 45983 16581
rect 45143 16541 45155 16544
rect 45097 16535 45155 16541
rect 45925 16541 45937 16575
rect 45971 16572 45983 16575
rect 47578 16572 47584 16584
rect 45971 16544 47584 16572
rect 45971 16541 45983 16544
rect 45925 16535 45983 16541
rect 45112 16504 45140 16535
rect 45940 16504 45968 16535
rect 47578 16532 47584 16544
rect 47636 16532 47642 16584
rect 58158 16572 58164 16584
rect 58119 16544 58164 16572
rect 58158 16532 58164 16544
rect 58216 16532 58222 16584
rect 41472 16476 45140 16504
rect 45204 16476 45968 16504
rect 41472 16464 41478 16476
rect 34388 16408 38608 16436
rect 38749 16439 38807 16445
rect 34388 16396 34394 16408
rect 38749 16405 38761 16439
rect 38795 16436 38807 16439
rect 39850 16436 39856 16448
rect 38795 16408 39856 16436
rect 38795 16405 38807 16408
rect 38749 16399 38807 16405
rect 39850 16396 39856 16408
rect 39908 16396 39914 16448
rect 43898 16396 43904 16448
rect 43956 16436 43962 16448
rect 44085 16439 44143 16445
rect 44085 16436 44097 16439
rect 43956 16408 44097 16436
rect 43956 16396 43962 16408
rect 44085 16405 44097 16408
rect 44131 16405 44143 16439
rect 44085 16399 44143 16405
rect 45002 16396 45008 16448
rect 45060 16436 45066 16448
rect 45204 16436 45232 16476
rect 48958 16464 48964 16516
rect 49016 16504 49022 16516
rect 57885 16507 57943 16513
rect 57885 16504 57897 16507
rect 49016 16476 57897 16504
rect 49016 16464 49022 16476
rect 57885 16473 57897 16476
rect 57931 16473 57943 16507
rect 57885 16467 57943 16473
rect 45830 16436 45836 16448
rect 45060 16408 45232 16436
rect 45791 16408 45836 16436
rect 45060 16396 45066 16408
rect 45830 16396 45836 16408
rect 45888 16396 45894 16448
rect 48590 16396 48596 16448
rect 48648 16436 48654 16448
rect 49145 16439 49203 16445
rect 49145 16436 49157 16439
rect 48648 16408 49157 16436
rect 48648 16396 48654 16408
rect 49145 16405 49157 16408
rect 49191 16405 49203 16439
rect 49145 16399 49203 16405
rect 1104 16346 58880 16368
rect 1104 16294 20214 16346
rect 20266 16294 20278 16346
rect 20330 16294 20342 16346
rect 20394 16294 20406 16346
rect 20458 16294 20470 16346
rect 20522 16294 39478 16346
rect 39530 16294 39542 16346
rect 39594 16294 39606 16346
rect 39658 16294 39670 16346
rect 39722 16294 39734 16346
rect 39786 16294 58880 16346
rect 1104 16272 58880 16294
rect 12250 16232 12256 16244
rect 12211 16204 12256 16232
rect 12250 16192 12256 16204
rect 12308 16192 12314 16244
rect 14461 16235 14519 16241
rect 14461 16201 14473 16235
rect 14507 16232 14519 16235
rect 15194 16232 15200 16244
rect 14507 16204 15200 16232
rect 14507 16201 14519 16204
rect 14461 16195 14519 16201
rect 15194 16192 15200 16204
rect 15252 16192 15258 16244
rect 15396 16204 17264 16232
rect 13357 16167 13415 16173
rect 13357 16133 13369 16167
rect 13403 16164 13415 16167
rect 15396 16164 15424 16204
rect 15562 16164 15568 16176
rect 13403 16136 15424 16164
rect 15523 16136 15568 16164
rect 13403 16133 13415 16136
rect 13357 16127 13415 16133
rect 15562 16124 15568 16136
rect 15620 16124 15626 16176
rect 17236 16164 17264 16204
rect 17310 16192 17316 16244
rect 17368 16232 17374 16244
rect 17368 16204 24808 16232
rect 17368 16192 17374 16204
rect 17770 16164 17776 16176
rect 17236 16136 17776 16164
rect 17770 16124 17776 16136
rect 17828 16164 17834 16176
rect 18049 16167 18107 16173
rect 18049 16164 18061 16167
rect 17828 16136 18061 16164
rect 17828 16124 17834 16136
rect 18049 16133 18061 16136
rect 18095 16164 18107 16167
rect 18095 16136 18828 16164
rect 18095 16133 18107 16136
rect 18049 16127 18107 16133
rect 13909 16099 13967 16105
rect 13909 16065 13921 16099
rect 13955 16096 13967 16099
rect 17034 16096 17040 16108
rect 13955 16068 17040 16096
rect 13955 16065 13967 16068
rect 13909 16059 13967 16065
rect 17034 16056 17040 16068
rect 17092 16096 17098 16108
rect 17221 16099 17279 16105
rect 17221 16096 17233 16099
rect 17092 16068 17233 16096
rect 17092 16056 17098 16068
rect 17221 16065 17233 16068
rect 17267 16065 17279 16099
rect 17221 16059 17279 16065
rect 17405 16099 17463 16105
rect 17405 16065 17417 16099
rect 17451 16096 17463 16099
rect 17451 16068 17816 16096
rect 17451 16065 17463 16068
rect 17405 16059 17463 16065
rect 12805 16031 12863 16037
rect 12805 15997 12817 16031
rect 12851 16028 12863 16031
rect 12894 16028 12900 16040
rect 12851 16000 12900 16028
rect 12851 15997 12863 16000
rect 12805 15991 12863 15997
rect 12894 15988 12900 16000
rect 12952 16028 12958 16040
rect 16114 16028 16120 16040
rect 12952 16000 16120 16028
rect 12952 15988 12958 16000
rect 16114 15988 16120 16000
rect 16172 15988 16178 16040
rect 17313 16031 17371 16037
rect 17313 15997 17325 16031
rect 17359 16028 17371 16031
rect 17678 16028 17684 16040
rect 17359 16000 17684 16028
rect 17359 15997 17371 16000
rect 17313 15991 17371 15997
rect 17678 15988 17684 16000
rect 17736 15988 17742 16040
rect 15194 15920 15200 15972
rect 15252 15960 15258 15972
rect 17788 15960 17816 16068
rect 17862 16056 17868 16108
rect 17920 16096 17926 16108
rect 18141 16099 18199 16105
rect 17920 16068 17965 16096
rect 17920 16056 17926 16068
rect 18141 16065 18153 16099
rect 18187 16096 18199 16099
rect 18414 16096 18420 16108
rect 18187 16068 18420 16096
rect 18187 16065 18199 16068
rect 18141 16059 18199 16065
rect 18414 16056 18420 16068
rect 18472 16056 18478 16108
rect 18800 16105 18828 16136
rect 18874 16124 18880 16176
rect 18932 16164 18938 16176
rect 19058 16164 19064 16176
rect 18932 16136 19064 16164
rect 18932 16124 18938 16136
rect 19058 16124 19064 16136
rect 19116 16164 19122 16176
rect 20530 16164 20536 16176
rect 19116 16136 20536 16164
rect 19116 16124 19122 16136
rect 20530 16124 20536 16136
rect 20588 16124 20594 16176
rect 20901 16167 20959 16173
rect 20901 16133 20913 16167
rect 20947 16164 20959 16167
rect 24486 16164 24492 16176
rect 20947 16136 21036 16164
rect 23966 16136 24492 16164
rect 20947 16133 20959 16136
rect 20901 16127 20959 16133
rect 18785 16099 18843 16105
rect 18785 16065 18797 16099
rect 18831 16096 18843 16099
rect 19797 16099 19855 16105
rect 18831 16068 19380 16096
rect 18831 16065 18843 16068
rect 18785 16059 18843 16065
rect 18690 16028 18696 16040
rect 18651 16000 18696 16028
rect 18690 15988 18696 16000
rect 18748 15988 18754 16040
rect 19150 15988 19156 16040
rect 19208 16028 19214 16040
rect 19208 16000 19253 16028
rect 19208 15988 19214 16000
rect 19352 15960 19380 16068
rect 19797 16065 19809 16099
rect 19843 16096 19855 16099
rect 19886 16096 19892 16108
rect 19843 16068 19892 16096
rect 19843 16065 19855 16068
rect 19797 16059 19855 16065
rect 19886 16056 19892 16068
rect 19944 16096 19950 16108
rect 20070 16096 20076 16108
rect 19944 16068 20076 16096
rect 19944 16056 19950 16068
rect 20070 16056 20076 16068
rect 20128 16056 20134 16108
rect 20625 16099 20683 16105
rect 20625 16065 20637 16099
rect 20671 16096 20683 16099
rect 20714 16096 20720 16108
rect 20671 16068 20720 16096
rect 20671 16065 20683 16068
rect 20625 16059 20683 16065
rect 20714 16056 20720 16068
rect 20772 16056 20778 16108
rect 19702 16028 19708 16040
rect 19663 16000 19708 16028
rect 19702 15988 19708 16000
rect 19760 15988 19766 16040
rect 20162 15988 20168 16040
rect 20220 16028 20226 16040
rect 20916 16028 20944 16127
rect 21008 16096 21036 16136
rect 24486 16124 24492 16136
rect 24544 16124 24550 16176
rect 21100 16096 21220 16102
rect 21634 16096 21640 16108
rect 21008 16074 21640 16096
rect 21008 16068 21128 16074
rect 21192 16068 21640 16074
rect 21634 16056 21640 16068
rect 21692 16056 21698 16108
rect 21726 16056 21732 16108
rect 21784 16096 21790 16108
rect 21821 16099 21879 16105
rect 21821 16096 21833 16099
rect 21784 16068 21833 16096
rect 21784 16056 21790 16068
rect 21821 16065 21833 16068
rect 21867 16065 21879 16099
rect 21821 16059 21879 16065
rect 20220 16000 20944 16028
rect 20993 16031 21051 16037
rect 20220 15988 20226 16000
rect 20993 15997 21005 16031
rect 21039 15997 21051 16031
rect 20993 15991 21051 15997
rect 20714 15960 20720 15972
rect 15252 15932 16804 15960
rect 17788 15932 19196 15960
rect 19352 15932 20720 15960
rect 15252 15920 15258 15932
rect 15013 15895 15071 15901
rect 15013 15861 15025 15895
rect 15059 15892 15071 15895
rect 15102 15892 15108 15904
rect 15059 15864 15108 15892
rect 15059 15861 15071 15864
rect 15013 15855 15071 15861
rect 15102 15852 15108 15864
rect 15160 15852 15166 15904
rect 16114 15892 16120 15904
rect 16075 15864 16120 15892
rect 16114 15852 16120 15864
rect 16172 15852 16178 15904
rect 16298 15852 16304 15904
rect 16356 15892 16362 15904
rect 16669 15895 16727 15901
rect 16669 15892 16681 15895
rect 16356 15864 16681 15892
rect 16356 15852 16362 15864
rect 16669 15861 16681 15864
rect 16715 15861 16727 15895
rect 16776 15892 16804 15932
rect 19168 15904 19196 15932
rect 20714 15920 20720 15932
rect 20772 15920 20778 15972
rect 17862 15892 17868 15904
rect 16776 15864 17868 15892
rect 16669 15855 16727 15861
rect 17862 15852 17868 15864
rect 17920 15852 17926 15904
rect 18138 15892 18144 15904
rect 18099 15864 18144 15892
rect 18138 15852 18144 15864
rect 18196 15852 18202 15904
rect 19150 15852 19156 15904
rect 19208 15852 19214 15904
rect 19886 15852 19892 15904
rect 19944 15892 19950 15904
rect 20073 15895 20131 15901
rect 20073 15892 20085 15895
rect 19944 15864 20085 15892
rect 19944 15852 19950 15864
rect 20073 15861 20085 15864
rect 20119 15861 20131 15895
rect 21008 15892 21036 15991
rect 21082 15988 21088 16040
rect 21140 16037 21146 16040
rect 21140 16031 21168 16037
rect 21156 15997 21168 16031
rect 22462 16028 22468 16040
rect 22423 16000 22468 16028
rect 21140 15991 21168 15997
rect 21140 15988 21146 15991
rect 22462 15988 22468 16000
rect 22520 15988 22526 16040
rect 22738 16028 22744 16040
rect 22699 16000 22744 16028
rect 22738 15988 22744 16000
rect 22796 15988 22802 16040
rect 23106 15988 23112 16040
rect 23164 16028 23170 16040
rect 24673 16031 24731 16037
rect 24673 16028 24685 16031
rect 23164 16000 24685 16028
rect 23164 15988 23170 16000
rect 24673 15997 24685 16000
rect 24719 15997 24731 16031
rect 24780 16028 24808 16204
rect 25222 16192 25228 16244
rect 25280 16232 25286 16244
rect 25498 16232 25504 16244
rect 25280 16204 25504 16232
rect 25280 16192 25286 16204
rect 25498 16192 25504 16204
rect 25556 16192 25562 16244
rect 27522 16232 27528 16244
rect 25976 16204 27528 16232
rect 25976 16164 26004 16204
rect 27522 16192 27528 16204
rect 27580 16192 27586 16244
rect 31570 16192 31576 16244
rect 31628 16232 31634 16244
rect 32950 16232 32956 16244
rect 31628 16204 32956 16232
rect 31628 16192 31634 16204
rect 32950 16192 32956 16204
rect 33008 16232 33014 16244
rect 34606 16232 34612 16244
rect 33008 16204 34612 16232
rect 33008 16192 33014 16204
rect 34606 16192 34612 16204
rect 34664 16232 34670 16244
rect 35250 16232 35256 16244
rect 34664 16204 35256 16232
rect 34664 16192 34670 16204
rect 35250 16192 35256 16204
rect 35308 16192 35314 16244
rect 35342 16192 35348 16244
rect 35400 16232 35406 16244
rect 38654 16232 38660 16244
rect 35400 16204 38660 16232
rect 35400 16192 35406 16204
rect 38654 16192 38660 16204
rect 38712 16192 38718 16244
rect 39390 16192 39396 16244
rect 39448 16232 39454 16244
rect 39485 16235 39543 16241
rect 39485 16232 39497 16235
rect 39448 16204 39497 16232
rect 39448 16192 39454 16204
rect 39485 16201 39497 16204
rect 39531 16201 39543 16235
rect 39485 16195 39543 16201
rect 41046 16192 41052 16244
rect 41104 16232 41110 16244
rect 41279 16235 41337 16241
rect 41279 16232 41291 16235
rect 41104 16204 41291 16232
rect 41104 16192 41110 16204
rect 41279 16201 41291 16204
rect 41325 16201 41337 16235
rect 41279 16195 41337 16201
rect 44542 16192 44548 16244
rect 44600 16232 44606 16244
rect 44726 16232 44732 16244
rect 44600 16204 44732 16232
rect 44600 16192 44606 16204
rect 44726 16192 44732 16204
rect 44784 16232 44790 16244
rect 46569 16235 46627 16241
rect 46569 16232 46581 16235
rect 44784 16204 46581 16232
rect 44784 16192 44790 16204
rect 46569 16201 46581 16204
rect 46615 16201 46627 16235
rect 47578 16232 47584 16244
rect 47539 16204 47584 16232
rect 46569 16195 46627 16201
rect 47578 16192 47584 16204
rect 47636 16192 47642 16244
rect 48225 16235 48283 16241
rect 48225 16201 48237 16235
rect 48271 16232 48283 16235
rect 48682 16232 48688 16244
rect 48271 16204 48688 16232
rect 48271 16201 48283 16204
rect 48225 16195 48283 16201
rect 48682 16192 48688 16204
rect 48740 16192 48746 16244
rect 58158 16232 58164 16244
rect 58119 16204 58164 16232
rect 58158 16192 58164 16204
rect 58216 16192 58222 16244
rect 26142 16164 26148 16176
rect 25714 16136 26004 16164
rect 26103 16136 26148 16164
rect 26142 16124 26148 16136
rect 26200 16124 26206 16176
rect 29454 16164 29460 16176
rect 26620 16136 29460 16164
rect 26418 16056 26424 16108
rect 26476 16096 26482 16108
rect 26476 16068 26521 16096
rect 26476 16056 26482 16068
rect 26620 16028 26648 16136
rect 29454 16124 29460 16136
rect 29512 16164 29518 16176
rect 29512 16136 29684 16164
rect 29512 16124 29518 16136
rect 27154 16056 27160 16108
rect 27212 16096 27218 16108
rect 29656 16105 29684 16136
rect 29914 16124 29920 16176
rect 29972 16164 29978 16176
rect 30742 16164 30748 16176
rect 29972 16136 30748 16164
rect 29972 16124 29978 16136
rect 30742 16124 30748 16136
rect 30800 16124 30806 16176
rect 34146 16124 34152 16176
rect 34204 16164 34210 16176
rect 37458 16164 37464 16176
rect 34204 16136 37464 16164
rect 34204 16124 34210 16136
rect 37458 16124 37464 16136
rect 37516 16124 37522 16176
rect 45830 16164 45836 16176
rect 38318 16136 45836 16164
rect 45830 16124 45836 16136
rect 45888 16124 45894 16176
rect 48130 16124 48136 16176
rect 48188 16164 48194 16176
rect 49237 16167 49295 16173
rect 49237 16164 49249 16167
rect 48188 16136 49249 16164
rect 48188 16124 48194 16136
rect 49237 16133 49249 16136
rect 49283 16133 49295 16167
rect 49237 16127 49295 16133
rect 27249 16099 27307 16105
rect 27249 16096 27261 16099
rect 27212 16068 27261 16096
rect 27212 16056 27218 16068
rect 27249 16065 27261 16068
rect 27295 16065 27307 16099
rect 27249 16059 27307 16065
rect 29641 16099 29699 16105
rect 29641 16065 29653 16099
rect 29687 16065 29699 16099
rect 30190 16096 30196 16108
rect 30151 16068 30196 16096
rect 29641 16059 29699 16065
rect 30190 16056 30196 16068
rect 30248 16056 30254 16108
rect 31202 16056 31208 16108
rect 31260 16096 31266 16108
rect 32125 16099 32183 16105
rect 32125 16096 32137 16099
rect 31260 16068 32137 16096
rect 31260 16056 31266 16068
rect 32125 16065 32137 16068
rect 32171 16065 32183 16099
rect 32125 16059 32183 16065
rect 33502 16056 33508 16108
rect 33560 16096 33566 16108
rect 33778 16096 33784 16108
rect 33560 16068 33784 16096
rect 33560 16056 33566 16068
rect 33778 16056 33784 16068
rect 33836 16096 33842 16108
rect 34425 16099 34483 16105
rect 34425 16096 34437 16099
rect 33836 16068 34437 16096
rect 33836 16056 33842 16068
rect 34425 16065 34437 16068
rect 34471 16065 34483 16099
rect 34425 16059 34483 16065
rect 39022 16056 39028 16108
rect 39080 16096 39086 16108
rect 39850 16096 39856 16108
rect 39080 16068 39125 16096
rect 39811 16068 39856 16096
rect 39080 16056 39086 16068
rect 39850 16056 39856 16068
rect 39908 16056 39914 16108
rect 40126 16096 40132 16108
rect 40087 16068 40132 16096
rect 40126 16056 40132 16068
rect 40184 16056 40190 16108
rect 42242 16096 42248 16108
rect 40236 16068 42248 16096
rect 24780 16000 26648 16028
rect 28905 16031 28963 16037
rect 24673 15991 24731 15997
rect 28905 15997 28917 16031
rect 28951 15997 28963 16031
rect 28905 15991 28963 15997
rect 29089 16031 29147 16037
rect 29089 15997 29101 16031
rect 29135 15997 29147 16031
rect 29089 15991 29147 15997
rect 21269 15963 21327 15969
rect 21269 15929 21281 15963
rect 21315 15960 21327 15963
rect 22370 15960 22376 15972
rect 21315 15932 22376 15960
rect 21315 15929 21327 15932
rect 21269 15923 21327 15929
rect 22370 15920 22376 15932
rect 22428 15920 22434 15972
rect 24210 15960 24216 15972
rect 24171 15932 24216 15960
rect 24210 15920 24216 15932
rect 24268 15920 24274 15972
rect 24854 15960 24860 15972
rect 24320 15932 24860 15960
rect 21634 15892 21640 15904
rect 21008 15864 21640 15892
rect 20073 15855 20131 15861
rect 21634 15852 21640 15864
rect 21692 15852 21698 15904
rect 21913 15895 21971 15901
rect 21913 15861 21925 15895
rect 21959 15892 21971 15895
rect 24320 15892 24348 15932
rect 24854 15920 24860 15932
rect 24912 15920 24918 15972
rect 21959 15864 24348 15892
rect 21959 15861 21971 15864
rect 21913 15855 21971 15861
rect 24762 15852 24768 15904
rect 24820 15892 24826 15904
rect 28718 15892 28724 15904
rect 24820 15864 28724 15892
rect 24820 15852 24826 15864
rect 28718 15852 28724 15864
rect 28776 15852 28782 15904
rect 28920 15892 28948 15991
rect 29104 15960 29132 15991
rect 30834 15988 30840 16040
rect 30892 16028 30898 16040
rect 31570 16028 31576 16040
rect 30892 16000 31576 16028
rect 30892 15988 30898 16000
rect 31570 15988 31576 16000
rect 31628 15988 31634 16040
rect 32309 16031 32367 16037
rect 32309 15997 32321 16031
rect 32355 16028 32367 16031
rect 33870 16028 33876 16040
rect 32355 16000 33876 16028
rect 32355 15997 32367 16000
rect 32309 15991 32367 15997
rect 33870 15988 33876 16000
rect 33928 15988 33934 16040
rect 33962 15988 33968 16040
rect 34020 16028 34026 16040
rect 34609 16031 34667 16037
rect 34020 16000 34065 16028
rect 34020 15988 34026 16000
rect 34609 15997 34621 16031
rect 34655 16028 34667 16031
rect 34790 16028 34796 16040
rect 34655 16000 34796 16028
rect 34655 15997 34667 16000
rect 34609 15991 34667 15997
rect 34790 15988 34796 16000
rect 34848 15988 34854 16040
rect 34885 16031 34943 16037
rect 34885 15997 34897 16031
rect 34931 16028 34943 16031
rect 35066 16028 35072 16040
rect 34931 16000 35072 16028
rect 34931 15997 34943 16000
rect 34885 15991 34943 15997
rect 33686 15960 33692 15972
rect 29104 15932 33692 15960
rect 33686 15920 33692 15932
rect 33744 15920 33750 15972
rect 34146 15920 34152 15972
rect 34204 15960 34210 15972
rect 34900 15960 34928 15991
rect 35066 15988 35072 16000
rect 35124 15988 35130 16040
rect 38746 16028 38752 16040
rect 38707 16000 38752 16028
rect 38746 15988 38752 16000
rect 38804 15988 38810 16040
rect 39868 16028 39896 16056
rect 40236 16028 40264 16068
rect 42242 16056 42248 16068
rect 42300 16056 42306 16108
rect 42613 16099 42671 16105
rect 42613 16096 42625 16099
rect 42444 16068 42625 16096
rect 39868 16000 40264 16028
rect 40954 15988 40960 16040
rect 41012 16028 41018 16040
rect 41049 16031 41107 16037
rect 41049 16028 41061 16031
rect 41012 16000 41061 16028
rect 41012 15988 41018 16000
rect 41049 15997 41061 16000
rect 41095 15997 41107 16031
rect 41049 15991 41107 15997
rect 34204 15932 34928 15960
rect 34204 15920 34210 15932
rect 40218 15920 40224 15972
rect 40276 15960 40282 15972
rect 42444 15960 42472 16068
rect 42613 16065 42625 16068
rect 42659 16065 42671 16099
rect 42794 16096 42800 16108
rect 42755 16068 42800 16096
rect 42613 16059 42671 16065
rect 42794 16056 42800 16068
rect 42852 16056 42858 16108
rect 42886 16056 42892 16108
rect 42944 16096 42950 16108
rect 43349 16099 43407 16105
rect 42944 16068 42989 16096
rect 42944 16056 42950 16068
rect 43349 16065 43361 16099
rect 43395 16065 43407 16099
rect 43349 16059 43407 16065
rect 42518 15988 42524 16040
rect 42576 16028 42582 16040
rect 43364 16028 43392 16059
rect 43438 16056 43444 16108
rect 43496 16096 43502 16108
rect 44358 16096 44364 16108
rect 43496 16068 43541 16096
rect 44319 16068 44364 16096
rect 43496 16056 43502 16068
rect 44358 16056 44364 16068
rect 44416 16056 44422 16108
rect 45005 16099 45063 16105
rect 45005 16065 45017 16099
rect 45051 16065 45063 16099
rect 45005 16059 45063 16065
rect 43622 16028 43628 16040
rect 42576 16000 43392 16028
rect 43583 16000 43628 16028
rect 42576 15988 42582 16000
rect 43622 15988 43628 16000
rect 43680 15988 43686 16040
rect 43806 15988 43812 16040
rect 43864 16028 43870 16040
rect 44085 16031 44143 16037
rect 44085 16028 44097 16031
rect 43864 16000 44097 16028
rect 43864 15988 43870 16000
rect 44085 15997 44097 16000
rect 44131 15997 44143 16031
rect 44085 15991 44143 15997
rect 45020 16028 45048 16059
rect 48314 16056 48320 16108
rect 48372 16096 48378 16108
rect 48685 16099 48743 16105
rect 48685 16096 48697 16099
rect 48372 16068 48697 16096
rect 48372 16056 48378 16068
rect 48685 16065 48697 16068
rect 48731 16065 48743 16099
rect 49786 16096 49792 16108
rect 49747 16068 49792 16096
rect 48685 16059 48743 16065
rect 49786 16056 49792 16068
rect 49844 16056 49850 16108
rect 46382 16028 46388 16040
rect 45020 16000 46388 16028
rect 43162 15960 43168 15972
rect 40276 15932 43168 15960
rect 40276 15920 40282 15932
rect 43162 15920 43168 15932
rect 43220 15960 43226 15972
rect 43438 15960 43444 15972
rect 43220 15932 43444 15960
rect 43220 15920 43226 15932
rect 43438 15920 43444 15932
rect 43496 15920 43502 15972
rect 43714 15920 43720 15972
rect 43772 15960 43778 15972
rect 45020 15960 45048 16000
rect 46382 15988 46388 16000
rect 46440 15988 46446 16040
rect 43772 15932 45048 15960
rect 43772 15920 43778 15932
rect 30282 15892 30288 15904
rect 28920 15864 30288 15892
rect 30282 15852 30288 15864
rect 30340 15852 30346 15904
rect 30834 15852 30840 15904
rect 30892 15892 30898 15904
rect 31481 15895 31539 15901
rect 31481 15892 31493 15895
rect 30892 15864 31493 15892
rect 30892 15852 30898 15864
rect 31481 15861 31493 15864
rect 31527 15892 31539 15895
rect 35342 15892 35348 15904
rect 31527 15864 35348 15892
rect 31527 15861 31539 15864
rect 31481 15855 31539 15861
rect 35342 15852 35348 15864
rect 35400 15852 35406 15904
rect 37277 15895 37335 15901
rect 37277 15861 37289 15895
rect 37323 15892 37335 15895
rect 39022 15892 39028 15904
rect 37323 15864 39028 15892
rect 37323 15861 37335 15864
rect 37277 15855 37335 15861
rect 39022 15852 39028 15864
rect 39080 15852 39086 15904
rect 40954 15852 40960 15904
rect 41012 15892 41018 15904
rect 41874 15892 41880 15904
rect 41012 15864 41880 15892
rect 41012 15852 41018 15864
rect 41874 15852 41880 15864
rect 41932 15852 41938 15904
rect 42426 15892 42432 15904
rect 42387 15864 42432 15892
rect 42426 15852 42432 15864
rect 42484 15852 42490 15904
rect 43533 15895 43591 15901
rect 43533 15861 43545 15895
rect 43579 15892 43591 15895
rect 43990 15892 43996 15904
rect 43579 15864 43996 15892
rect 43579 15861 43591 15864
rect 43533 15855 43591 15861
rect 43990 15852 43996 15864
rect 44048 15852 44054 15904
rect 44174 15892 44180 15904
rect 44135 15864 44180 15892
rect 44174 15852 44180 15864
rect 44232 15852 44238 15904
rect 44269 15895 44327 15901
rect 44269 15861 44281 15895
rect 44315 15892 44327 15895
rect 44542 15892 44548 15904
rect 44315 15864 44548 15892
rect 44315 15861 44327 15864
rect 44269 15855 44327 15861
rect 44542 15852 44548 15864
rect 44600 15852 44606 15904
rect 44910 15892 44916 15904
rect 44871 15864 44916 15892
rect 44910 15852 44916 15864
rect 44968 15852 44974 15904
rect 45557 15895 45615 15901
rect 45557 15861 45569 15895
rect 45603 15892 45615 15895
rect 45738 15892 45744 15904
rect 45603 15864 45744 15892
rect 45603 15861 45615 15864
rect 45557 15855 45615 15861
rect 45738 15852 45744 15864
rect 45796 15852 45802 15904
rect 46014 15892 46020 15904
rect 45975 15864 46020 15892
rect 46014 15852 46020 15864
rect 46072 15852 46078 15904
rect 1104 15802 58880 15824
rect 1104 15750 10582 15802
rect 10634 15750 10646 15802
rect 10698 15750 10710 15802
rect 10762 15750 10774 15802
rect 10826 15750 10838 15802
rect 10890 15750 29846 15802
rect 29898 15750 29910 15802
rect 29962 15750 29974 15802
rect 30026 15750 30038 15802
rect 30090 15750 30102 15802
rect 30154 15750 49110 15802
rect 49162 15750 49174 15802
rect 49226 15750 49238 15802
rect 49290 15750 49302 15802
rect 49354 15750 49366 15802
rect 49418 15750 58880 15802
rect 1104 15728 58880 15750
rect 14274 15648 14280 15700
rect 14332 15688 14338 15700
rect 15105 15691 15163 15697
rect 15105 15688 15117 15691
rect 14332 15660 15117 15688
rect 14332 15648 14338 15660
rect 15105 15657 15117 15660
rect 15151 15688 15163 15691
rect 15194 15688 15200 15700
rect 15151 15660 15200 15688
rect 15151 15657 15163 15660
rect 15105 15651 15163 15657
rect 15194 15648 15200 15660
rect 15252 15648 15258 15700
rect 15654 15688 15660 15700
rect 15615 15660 15660 15688
rect 15654 15648 15660 15660
rect 15712 15648 15718 15700
rect 16209 15691 16267 15697
rect 16209 15657 16221 15691
rect 16255 15688 16267 15691
rect 20070 15688 20076 15700
rect 16255 15660 20076 15688
rect 16255 15657 16267 15660
rect 16209 15651 16267 15657
rect 20070 15648 20076 15660
rect 20128 15688 20134 15700
rect 21082 15688 21088 15700
rect 20128 15660 21088 15688
rect 20128 15648 20134 15660
rect 21082 15648 21088 15660
rect 21140 15648 21146 15700
rect 21266 15648 21272 15700
rect 21324 15688 21330 15700
rect 21913 15691 21971 15697
rect 21324 15660 21680 15688
rect 21324 15648 21330 15660
rect 13541 15623 13599 15629
rect 13541 15589 13553 15623
rect 13587 15620 13599 15623
rect 15838 15620 15844 15632
rect 13587 15592 15844 15620
rect 13587 15589 13599 15592
rect 13541 15583 13599 15589
rect 15838 15580 15844 15592
rect 15896 15580 15902 15632
rect 16761 15623 16819 15629
rect 16761 15589 16773 15623
rect 16807 15620 16819 15623
rect 20349 15623 20407 15629
rect 20349 15620 20361 15623
rect 16807 15592 20361 15620
rect 16807 15589 16819 15592
rect 16761 15583 16819 15589
rect 20349 15589 20361 15592
rect 20395 15620 20407 15623
rect 21174 15620 21180 15632
rect 20395 15592 21180 15620
rect 20395 15589 20407 15592
rect 20349 15583 20407 15589
rect 21174 15580 21180 15592
rect 21232 15580 21238 15632
rect 15654 15512 15660 15564
rect 15712 15552 15718 15564
rect 16206 15552 16212 15564
rect 15712 15524 16212 15552
rect 15712 15512 15718 15524
rect 16206 15512 16212 15524
rect 16264 15512 16270 15564
rect 18322 15552 18328 15564
rect 17604 15524 18328 15552
rect 11425 15487 11483 15493
rect 11425 15453 11437 15487
rect 11471 15453 11483 15487
rect 11425 15447 11483 15453
rect 14553 15487 14611 15493
rect 14553 15453 14565 15487
rect 14599 15484 14611 15487
rect 17604 15484 17632 15524
rect 18322 15512 18328 15524
rect 18380 15552 18386 15564
rect 19613 15555 19671 15561
rect 18380 15524 19564 15552
rect 18380 15512 18386 15524
rect 14599 15456 17632 15484
rect 14599 15453 14611 15456
rect 14553 15447 14611 15453
rect 11440 15416 11468 15447
rect 17678 15444 17684 15496
rect 17736 15484 17742 15496
rect 19536 15493 19564 15524
rect 19613 15521 19625 15555
rect 19659 15552 19671 15555
rect 20898 15552 20904 15564
rect 19659 15524 19932 15552
rect 20859 15524 20904 15552
rect 19659 15521 19671 15524
rect 19613 15515 19671 15521
rect 17773 15487 17831 15493
rect 17773 15484 17785 15487
rect 17736 15456 17785 15484
rect 17736 15444 17742 15456
rect 17773 15453 17785 15456
rect 17819 15453 17831 15487
rect 17773 15447 17831 15453
rect 19521 15487 19579 15493
rect 19521 15453 19533 15487
rect 19567 15484 19579 15487
rect 19702 15484 19708 15496
rect 19567 15456 19708 15484
rect 19567 15453 19579 15456
rect 19521 15447 19579 15453
rect 19702 15444 19708 15456
rect 19760 15444 19766 15496
rect 19904 15484 19932 15524
rect 20898 15512 20904 15524
rect 20956 15512 20962 15564
rect 21542 15552 21548 15564
rect 21008 15524 21548 15552
rect 20162 15484 20168 15496
rect 19904 15456 20168 15484
rect 20162 15444 20168 15456
rect 20220 15444 20226 15496
rect 20530 15444 20536 15496
rect 20588 15484 20594 15496
rect 20625 15487 20683 15493
rect 20625 15484 20637 15487
rect 20588 15456 20637 15484
rect 20588 15444 20594 15456
rect 20625 15453 20637 15456
rect 20671 15453 20683 15487
rect 20625 15447 20683 15453
rect 20714 15444 20720 15496
rect 20772 15484 20778 15496
rect 21008 15484 21036 15524
rect 21542 15512 21548 15524
rect 21600 15512 21606 15564
rect 21358 15484 21364 15496
rect 20772 15456 21036 15484
rect 21319 15456 21364 15484
rect 20772 15444 20778 15456
rect 21358 15444 21364 15456
rect 21416 15444 21422 15496
rect 21652 15493 21680 15660
rect 21913 15657 21925 15691
rect 21959 15688 21971 15691
rect 22646 15688 22652 15700
rect 21959 15660 22652 15688
rect 21959 15657 21971 15660
rect 21913 15651 21971 15657
rect 22646 15648 22652 15660
rect 22704 15648 22710 15700
rect 23474 15648 23480 15700
rect 23532 15688 23538 15700
rect 24026 15688 24032 15700
rect 23532 15660 24032 15688
rect 23532 15648 23538 15660
rect 24026 15648 24032 15660
rect 24084 15688 24090 15700
rect 24397 15691 24455 15697
rect 24397 15688 24409 15691
rect 24084 15660 24409 15688
rect 24084 15648 24090 15660
rect 24397 15657 24409 15660
rect 24443 15657 24455 15691
rect 24397 15651 24455 15657
rect 25041 15691 25099 15697
rect 25041 15657 25053 15691
rect 25087 15688 25099 15691
rect 25406 15688 25412 15700
rect 25087 15660 25412 15688
rect 25087 15657 25099 15660
rect 25041 15651 25099 15657
rect 25406 15648 25412 15660
rect 25464 15648 25470 15700
rect 39209 15691 39267 15697
rect 39209 15688 39221 15691
rect 25516 15660 39221 15688
rect 21726 15580 21732 15632
rect 21784 15620 21790 15632
rect 24118 15620 24124 15632
rect 21784 15592 24124 15620
rect 21784 15580 21790 15592
rect 24118 15580 24124 15592
rect 24176 15620 24182 15632
rect 24578 15620 24584 15632
rect 24176 15592 24584 15620
rect 24176 15580 24182 15592
rect 24578 15580 24584 15592
rect 24636 15580 24642 15632
rect 25130 15580 25136 15632
rect 25188 15620 25194 15632
rect 25516 15620 25544 15660
rect 39209 15657 39221 15660
rect 39255 15657 39267 15691
rect 41046 15688 41052 15700
rect 39209 15651 39267 15657
rect 39960 15660 41052 15688
rect 25188 15592 25544 15620
rect 28997 15623 29055 15629
rect 25188 15580 25194 15592
rect 28997 15589 29009 15623
rect 29043 15620 29055 15623
rect 29546 15620 29552 15632
rect 29043 15592 29552 15620
rect 29043 15589 29055 15592
rect 28997 15583 29055 15589
rect 29546 15580 29552 15592
rect 29604 15580 29610 15632
rect 32306 15580 32312 15632
rect 32364 15620 32370 15632
rect 32766 15620 32772 15632
rect 32364 15592 32772 15620
rect 32364 15580 32370 15592
rect 32766 15580 32772 15592
rect 32824 15580 32830 15632
rect 38657 15623 38715 15629
rect 38657 15589 38669 15623
rect 38703 15620 38715 15623
rect 39850 15620 39856 15632
rect 38703 15592 39856 15620
rect 38703 15589 38715 15592
rect 38657 15583 38715 15589
rect 39850 15580 39856 15592
rect 39908 15580 39914 15632
rect 26418 15552 26424 15564
rect 22848 15524 26424 15552
rect 21637 15487 21695 15493
rect 21637 15453 21649 15487
rect 21683 15453 21695 15487
rect 21637 15447 21695 15453
rect 21781 15487 21839 15493
rect 21781 15453 21793 15487
rect 21827 15484 21839 15487
rect 22186 15484 22192 15496
rect 21827 15456 22192 15484
rect 21827 15453 21839 15456
rect 21781 15447 21839 15453
rect 22186 15444 22192 15456
rect 22244 15444 22250 15496
rect 11977 15419 12035 15425
rect 11977 15416 11989 15419
rect 11440 15388 11989 15416
rect 11977 15385 11989 15388
rect 12023 15416 12035 15419
rect 15102 15416 15108 15428
rect 12023 15388 15108 15416
rect 12023 15385 12035 15388
rect 11977 15379 12035 15385
rect 15102 15376 15108 15388
rect 15160 15376 15166 15428
rect 18506 15416 18512 15428
rect 18419 15388 18512 15416
rect 18506 15376 18512 15388
rect 18564 15416 18570 15428
rect 21545 15419 21603 15425
rect 18564 15388 21496 15416
rect 18564 15376 18570 15388
rect 11238 15348 11244 15360
rect 11199 15320 11244 15348
rect 11238 15308 11244 15320
rect 11296 15308 11302 15360
rect 12986 15348 12992 15360
rect 12947 15320 12992 15348
rect 12986 15308 12992 15320
rect 13044 15308 13050 15360
rect 17310 15348 17316 15360
rect 17271 15320 17316 15348
rect 17310 15308 17316 15320
rect 17368 15308 17374 15360
rect 17862 15348 17868 15360
rect 17823 15320 17868 15348
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 18414 15308 18420 15360
rect 18472 15348 18478 15360
rect 18601 15351 18659 15357
rect 18601 15348 18613 15351
rect 18472 15320 18613 15348
rect 18472 15308 18478 15320
rect 18601 15317 18613 15320
rect 18647 15317 18659 15351
rect 18601 15311 18659 15317
rect 19889 15351 19947 15357
rect 19889 15317 19901 15351
rect 19935 15348 19947 15351
rect 20070 15348 20076 15360
rect 19935 15320 20076 15348
rect 19935 15317 19947 15320
rect 19889 15311 19947 15317
rect 20070 15308 20076 15320
rect 20128 15308 20134 15360
rect 20533 15351 20591 15357
rect 20533 15317 20545 15351
rect 20579 15348 20591 15351
rect 20898 15348 20904 15360
rect 20579 15320 20904 15348
rect 20579 15317 20591 15320
rect 20533 15311 20591 15317
rect 20898 15308 20904 15320
rect 20956 15308 20962 15360
rect 21468 15348 21496 15388
rect 21545 15385 21557 15419
rect 21591 15416 21603 15419
rect 22094 15416 22100 15428
rect 21591 15388 22100 15416
rect 21591 15385 21603 15388
rect 21545 15379 21603 15385
rect 22094 15376 22100 15388
rect 22152 15376 22158 15428
rect 22848 15348 22876 15524
rect 26418 15512 26424 15524
rect 26476 15512 26482 15564
rect 26786 15552 26792 15564
rect 26747 15524 26792 15552
rect 26786 15512 26792 15524
rect 26844 15512 26850 15564
rect 27525 15555 27583 15561
rect 27525 15521 27537 15555
rect 27571 15552 27583 15555
rect 28534 15552 28540 15564
rect 27571 15524 28540 15552
rect 27571 15521 27583 15524
rect 27525 15515 27583 15521
rect 28534 15512 28540 15524
rect 28592 15512 28598 15564
rect 31849 15555 31907 15561
rect 31849 15521 31861 15555
rect 31895 15552 31907 15555
rect 36538 15552 36544 15564
rect 31895 15524 36544 15552
rect 31895 15521 31907 15524
rect 31849 15515 31907 15521
rect 36538 15512 36544 15524
rect 36596 15512 36602 15564
rect 36814 15512 36820 15564
rect 36872 15552 36878 15564
rect 36909 15555 36967 15561
rect 36909 15552 36921 15555
rect 36872 15524 36921 15552
rect 36872 15512 36878 15524
rect 36909 15521 36921 15524
rect 36955 15521 36967 15555
rect 36909 15515 36967 15521
rect 38378 15512 38384 15564
rect 38436 15552 38442 15564
rect 39960 15552 39988 15660
rect 41046 15648 41052 15660
rect 41104 15648 41110 15700
rect 41506 15648 41512 15700
rect 41564 15688 41570 15700
rect 41693 15691 41751 15697
rect 41693 15688 41705 15691
rect 41564 15660 41705 15688
rect 41564 15648 41570 15660
rect 41693 15657 41705 15660
rect 41739 15657 41751 15691
rect 42518 15688 42524 15700
rect 42479 15660 42524 15688
rect 41693 15651 41751 15657
rect 42518 15648 42524 15660
rect 42576 15648 42582 15700
rect 43346 15688 43352 15700
rect 43307 15660 43352 15688
rect 43346 15648 43352 15660
rect 43404 15648 43410 15700
rect 43438 15648 43444 15700
rect 43496 15688 43502 15700
rect 45005 15691 45063 15697
rect 45005 15688 45017 15691
rect 43496 15660 45017 15688
rect 43496 15648 43502 15660
rect 45005 15657 45017 15660
rect 45051 15688 45063 15691
rect 45186 15688 45192 15700
rect 45051 15660 45192 15688
rect 45051 15657 45063 15660
rect 45005 15651 45063 15657
rect 45186 15648 45192 15660
rect 45244 15648 45250 15700
rect 45554 15688 45560 15700
rect 45515 15660 45560 15688
rect 45554 15648 45560 15660
rect 45612 15648 45618 15700
rect 47305 15691 47363 15697
rect 47305 15657 47317 15691
rect 47351 15688 47363 15691
rect 47578 15688 47584 15700
rect 47351 15660 47584 15688
rect 47351 15657 47363 15660
rect 47305 15651 47363 15657
rect 47578 15648 47584 15660
rect 47636 15688 47642 15700
rect 47765 15691 47823 15697
rect 47765 15688 47777 15691
rect 47636 15660 47777 15688
rect 47636 15648 47642 15660
rect 47765 15657 47777 15660
rect 47811 15688 47823 15691
rect 48682 15688 48688 15700
rect 47811 15660 48688 15688
rect 47811 15657 47823 15660
rect 47765 15651 47823 15657
rect 48682 15648 48688 15660
rect 48740 15688 48746 15700
rect 48869 15691 48927 15697
rect 48869 15688 48881 15691
rect 48740 15660 48881 15688
rect 48740 15648 48746 15660
rect 48869 15657 48881 15660
rect 48915 15688 48927 15691
rect 49421 15691 49479 15697
rect 49421 15688 49433 15691
rect 48915 15660 49433 15688
rect 48915 15657 48927 15660
rect 48869 15651 48927 15657
rect 49421 15657 49433 15660
rect 49467 15657 49479 15691
rect 49421 15651 49479 15657
rect 42334 15580 42340 15632
rect 42392 15620 42398 15632
rect 42610 15620 42616 15632
rect 42392 15592 42616 15620
rect 42392 15580 42398 15592
rect 42610 15580 42616 15592
rect 42668 15580 42674 15632
rect 43257 15623 43315 15629
rect 43257 15589 43269 15623
rect 43303 15620 43315 15623
rect 44450 15620 44456 15632
rect 43303 15592 44456 15620
rect 43303 15589 43315 15592
rect 43257 15583 43315 15589
rect 44450 15580 44456 15592
rect 44508 15580 44514 15632
rect 38436 15524 39988 15552
rect 41049 15555 41107 15561
rect 38436 15512 38442 15524
rect 41049 15521 41061 15555
rect 41095 15552 41107 15555
rect 41690 15552 41696 15564
rect 41095 15524 41696 15552
rect 41095 15521 41107 15524
rect 41049 15515 41107 15521
rect 41690 15512 41696 15524
rect 41748 15512 41754 15564
rect 46109 15555 46167 15561
rect 46109 15552 46121 15555
rect 42720 15524 46121 15552
rect 23109 15487 23167 15493
rect 23109 15453 23121 15487
rect 23155 15453 23167 15487
rect 23109 15447 23167 15453
rect 23753 15487 23811 15493
rect 23753 15453 23765 15487
rect 23799 15453 23811 15487
rect 23753 15447 23811 15453
rect 24581 15487 24639 15493
rect 24581 15453 24593 15487
rect 24627 15484 24639 15487
rect 24670 15484 24676 15496
rect 24627 15456 24676 15484
rect 24627 15453 24639 15456
rect 24581 15447 24639 15453
rect 23124 15416 23152 15447
rect 23566 15416 23572 15428
rect 23124 15388 23572 15416
rect 23566 15376 23572 15388
rect 23624 15376 23630 15428
rect 21468 15320 22876 15348
rect 22925 15351 22983 15357
rect 22925 15317 22937 15351
rect 22971 15348 22983 15351
rect 23290 15348 23296 15360
rect 22971 15320 23296 15348
rect 22971 15317 22983 15320
rect 22925 15311 22983 15317
rect 23290 15308 23296 15320
rect 23348 15308 23354 15360
rect 23768 15348 23796 15447
rect 24670 15444 24676 15456
rect 24728 15444 24734 15496
rect 27246 15484 27252 15496
rect 27207 15456 27252 15484
rect 27246 15444 27252 15456
rect 27304 15444 27310 15496
rect 32306 15484 32312 15496
rect 32267 15456 32312 15484
rect 32306 15444 32312 15456
rect 32364 15444 32370 15496
rect 34606 15444 34612 15496
rect 34664 15484 34670 15496
rect 34664 15456 35098 15484
rect 34664 15444 34670 15456
rect 36446 15444 36452 15496
rect 36504 15484 36510 15496
rect 36504 15456 36549 15484
rect 36504 15444 36510 15456
rect 38930 15444 38936 15496
rect 38988 15484 38994 15496
rect 39117 15487 39175 15493
rect 39117 15484 39129 15487
rect 38988 15456 39129 15484
rect 38988 15444 38994 15456
rect 39117 15453 39129 15456
rect 39163 15453 39175 15487
rect 39117 15447 39175 15453
rect 39390 15444 39396 15496
rect 39448 15484 39454 15496
rect 40129 15487 40187 15493
rect 39448 15456 40080 15484
rect 39448 15444 39454 15456
rect 25958 15376 25964 15428
rect 26016 15376 26022 15428
rect 26513 15419 26571 15425
rect 26513 15385 26525 15419
rect 26559 15385 26571 15419
rect 26513 15379 26571 15385
rect 26142 15348 26148 15360
rect 23768 15320 26148 15348
rect 26142 15308 26148 15320
rect 26200 15308 26206 15360
rect 26528 15348 26556 15379
rect 27982 15376 27988 15428
rect 28040 15376 28046 15428
rect 29546 15376 29552 15428
rect 29604 15416 29610 15428
rect 30282 15416 30288 15428
rect 29604 15388 30288 15416
rect 29604 15376 29610 15388
rect 30282 15376 30288 15388
rect 30340 15376 30346 15428
rect 31570 15416 31576 15428
rect 31142 15388 31432 15416
rect 31531 15388 31576 15416
rect 28442 15348 28448 15360
rect 26528 15320 28448 15348
rect 28442 15308 28448 15320
rect 28500 15308 28506 15360
rect 29638 15308 29644 15360
rect 29696 15348 29702 15360
rect 30101 15351 30159 15357
rect 30101 15348 30113 15351
rect 29696 15320 30113 15348
rect 29696 15308 29702 15320
rect 30101 15317 30113 15320
rect 30147 15348 30159 15351
rect 30190 15348 30196 15360
rect 30147 15320 30196 15348
rect 30147 15317 30159 15320
rect 30101 15311 30159 15317
rect 30190 15308 30196 15320
rect 30248 15308 30254 15360
rect 30650 15308 30656 15360
rect 30708 15348 30714 15360
rect 30834 15348 30840 15360
rect 30708 15320 30840 15348
rect 30708 15308 30714 15320
rect 30834 15308 30840 15320
rect 30892 15308 30898 15360
rect 31404 15348 31432 15388
rect 31570 15376 31576 15388
rect 31628 15376 31634 15428
rect 31938 15376 31944 15428
rect 31996 15416 32002 15428
rect 32493 15419 32551 15425
rect 32493 15416 32505 15419
rect 31996 15388 32505 15416
rect 31996 15376 32002 15388
rect 32493 15385 32505 15388
rect 32539 15385 32551 15419
rect 32493 15379 32551 15385
rect 32582 15376 32588 15428
rect 32640 15416 32646 15428
rect 33042 15416 33048 15428
rect 32640 15388 33048 15416
rect 32640 15376 32646 15388
rect 33042 15376 33048 15388
rect 33100 15376 33106 15428
rect 33134 15376 33140 15428
rect 33192 15416 33198 15428
rect 33962 15416 33968 15428
rect 33192 15388 33968 15416
rect 33192 15376 33198 15388
rect 33962 15376 33968 15388
rect 34020 15416 34026 15428
rect 34149 15419 34207 15425
rect 34149 15416 34161 15419
rect 34020 15388 34161 15416
rect 34020 15376 34026 15388
rect 34149 15385 34161 15388
rect 34195 15385 34207 15419
rect 36170 15416 36176 15428
rect 34149 15379 34207 15385
rect 34256 15388 34836 15416
rect 36131 15388 36176 15416
rect 31478 15348 31484 15360
rect 31404 15320 31484 15348
rect 31478 15308 31484 15320
rect 31536 15308 31542 15360
rect 32306 15308 32312 15360
rect 32364 15348 32370 15360
rect 34256 15348 34284 15388
rect 32364 15320 34284 15348
rect 32364 15308 32370 15320
rect 34606 15308 34612 15360
rect 34664 15348 34670 15360
rect 34701 15351 34759 15357
rect 34701 15348 34713 15351
rect 34664 15320 34713 15348
rect 34664 15308 34670 15320
rect 34701 15317 34713 15320
rect 34747 15317 34759 15351
rect 34808 15348 34836 15388
rect 36170 15376 36176 15388
rect 36228 15376 36234 15428
rect 37185 15419 37243 15425
rect 37185 15416 37197 15419
rect 36280 15388 37197 15416
rect 36280 15348 36308 15388
rect 37185 15385 37197 15388
rect 37231 15385 37243 15419
rect 37185 15379 37243 15385
rect 37274 15376 37280 15428
rect 37332 15416 37338 15428
rect 37332 15388 37674 15416
rect 37332 15376 37338 15388
rect 38838 15376 38844 15428
rect 38896 15416 38902 15428
rect 39853 15419 39911 15425
rect 39853 15416 39865 15419
rect 38896 15388 39865 15416
rect 38896 15376 38902 15388
rect 39853 15385 39865 15388
rect 39899 15416 39911 15419
rect 39942 15416 39948 15428
rect 39899 15388 39948 15416
rect 39899 15385 39911 15388
rect 39853 15379 39911 15385
rect 39942 15376 39948 15388
rect 40000 15376 40006 15428
rect 40052 15416 40080 15456
rect 40129 15453 40141 15487
rect 40175 15484 40187 15487
rect 40586 15484 40592 15496
rect 40175 15456 40592 15484
rect 40175 15453 40187 15456
rect 40129 15447 40187 15453
rect 40586 15444 40592 15456
rect 40644 15444 40650 15496
rect 40773 15487 40831 15493
rect 40773 15453 40785 15487
rect 40819 15453 40831 15487
rect 41966 15484 41972 15496
rect 41927 15456 41972 15484
rect 40773 15447 40831 15453
rect 40788 15416 40816 15447
rect 41966 15444 41972 15456
rect 42024 15444 42030 15496
rect 42720 15493 42748 15524
rect 46109 15521 46121 15524
rect 46155 15521 46167 15555
rect 46109 15515 46167 15521
rect 42705 15487 42763 15493
rect 42705 15484 42717 15487
rect 42076 15456 42717 15484
rect 40052 15388 40816 15416
rect 41138 15376 41144 15428
rect 41196 15416 41202 15428
rect 42076 15416 42104 15456
rect 42705 15453 42717 15456
rect 42751 15453 42763 15487
rect 43162 15484 43168 15496
rect 43123 15456 43168 15484
rect 42705 15447 42763 15453
rect 43162 15444 43168 15456
rect 43220 15444 43226 15496
rect 43714 15444 43720 15496
rect 43772 15484 43778 15496
rect 44085 15487 44143 15493
rect 44085 15484 44097 15487
rect 43772 15456 44097 15484
rect 43772 15444 43778 15456
rect 44085 15453 44097 15456
rect 44131 15453 44143 15487
rect 58158 15484 58164 15496
rect 58119 15456 58164 15484
rect 44085 15447 44143 15453
rect 58158 15444 58164 15456
rect 58216 15444 58222 15496
rect 41196 15388 42104 15416
rect 42429 15419 42487 15425
rect 41196 15376 41202 15388
rect 42429 15385 42441 15419
rect 42475 15416 42487 15419
rect 42518 15416 42524 15428
rect 42475 15388 42524 15416
rect 42475 15385 42487 15388
rect 42429 15379 42487 15385
rect 42518 15376 42524 15388
rect 42576 15376 42582 15428
rect 43346 15376 43352 15428
rect 43404 15416 43410 15428
rect 43441 15419 43499 15425
rect 43441 15416 43453 15419
rect 43404 15388 43453 15416
rect 43404 15376 43410 15388
rect 43441 15385 43453 15388
rect 43487 15385 43499 15419
rect 57882 15416 57888 15428
rect 57843 15388 57888 15416
rect 43441 15379 43499 15385
rect 57882 15376 57888 15388
rect 57940 15376 57946 15428
rect 34808 15320 36308 15348
rect 34701 15311 34759 15317
rect 39298 15308 39304 15360
rect 39356 15348 39362 15360
rect 41509 15351 41567 15357
rect 41509 15348 41521 15351
rect 39356 15320 41521 15348
rect 39356 15308 39362 15320
rect 41509 15317 41521 15320
rect 41555 15317 41567 15351
rect 41509 15311 41567 15317
rect 41874 15308 41880 15360
rect 41932 15348 41938 15360
rect 42334 15348 42340 15360
rect 41932 15320 42340 15348
rect 41932 15308 41938 15320
rect 42334 15308 42340 15320
rect 42392 15308 42398 15360
rect 42978 15308 42984 15360
rect 43036 15348 43042 15360
rect 43622 15348 43628 15360
rect 43036 15320 43628 15348
rect 43036 15308 43042 15320
rect 43622 15308 43628 15320
rect 43680 15308 43686 15360
rect 43990 15348 43996 15360
rect 43951 15320 43996 15348
rect 43990 15308 43996 15320
rect 44048 15308 44054 15360
rect 46382 15308 46388 15360
rect 46440 15348 46446 15360
rect 46661 15351 46719 15357
rect 46661 15348 46673 15351
rect 46440 15320 46673 15348
rect 46440 15308 46446 15320
rect 46661 15317 46673 15320
rect 46707 15317 46719 15351
rect 48314 15348 48320 15360
rect 48275 15320 48320 15348
rect 46661 15311 46719 15317
rect 48314 15308 48320 15320
rect 48372 15348 48378 15360
rect 48590 15348 48596 15360
rect 48372 15320 48596 15348
rect 48372 15308 48378 15320
rect 48590 15308 48596 15320
rect 48648 15308 48654 15360
rect 1104 15258 58880 15280
rect 1104 15206 20214 15258
rect 20266 15206 20278 15258
rect 20330 15206 20342 15258
rect 20394 15206 20406 15258
rect 20458 15206 20470 15258
rect 20522 15206 39478 15258
rect 39530 15206 39542 15258
rect 39594 15206 39606 15258
rect 39658 15206 39670 15258
rect 39722 15206 39734 15258
rect 39786 15206 58880 15258
rect 1104 15184 58880 15206
rect 12710 15104 12716 15156
rect 12768 15144 12774 15156
rect 13630 15144 13636 15156
rect 12768 15116 13636 15144
rect 12768 15104 12774 15116
rect 13630 15104 13636 15116
rect 13688 15144 13694 15156
rect 13817 15147 13875 15153
rect 13817 15144 13829 15147
rect 13688 15116 13829 15144
rect 13688 15104 13694 15116
rect 13817 15113 13829 15116
rect 13863 15113 13875 15147
rect 13817 15107 13875 15113
rect 15013 15147 15071 15153
rect 15013 15113 15025 15147
rect 15059 15144 15071 15147
rect 15194 15144 15200 15156
rect 15059 15116 15200 15144
rect 15059 15113 15071 15116
rect 15013 15107 15071 15113
rect 15194 15104 15200 15116
rect 15252 15104 15258 15156
rect 16117 15147 16175 15153
rect 16117 15113 16129 15147
rect 16163 15144 16175 15147
rect 18506 15144 18512 15156
rect 16163 15116 18512 15144
rect 16163 15113 16175 15116
rect 16117 15107 16175 15113
rect 18506 15104 18512 15116
rect 18564 15104 18570 15156
rect 19242 15104 19248 15156
rect 19300 15104 19306 15156
rect 20898 15144 20904 15156
rect 20732 15116 20904 15144
rect 14461 15079 14519 15085
rect 14461 15045 14473 15079
rect 14507 15076 14519 15079
rect 17678 15076 17684 15088
rect 14507 15048 17684 15076
rect 14507 15045 14519 15048
rect 14461 15039 14519 15045
rect 17678 15036 17684 15048
rect 17736 15036 17742 15088
rect 17957 15079 18015 15085
rect 17957 15045 17969 15079
rect 18003 15076 18015 15079
rect 18046 15076 18052 15088
rect 18003 15048 18052 15076
rect 18003 15045 18015 15048
rect 17957 15039 18015 15045
rect 18046 15036 18052 15048
rect 18104 15036 18110 15088
rect 19153 15079 19211 15085
rect 19153 15045 19165 15079
rect 19199 15076 19211 15079
rect 19260 15076 19288 15104
rect 20732 15076 20760 15116
rect 20898 15104 20904 15116
rect 20956 15104 20962 15156
rect 21269 15147 21327 15153
rect 21269 15113 21281 15147
rect 21315 15113 21327 15147
rect 21726 15144 21732 15156
rect 21269 15107 21327 15113
rect 21468 15116 21732 15144
rect 21284 15076 21312 15107
rect 21468 15076 21496 15116
rect 21726 15104 21732 15116
rect 21784 15104 21790 15156
rect 21818 15104 21824 15156
rect 21876 15144 21882 15156
rect 22278 15144 22284 15156
rect 21876 15116 22284 15144
rect 21876 15104 21882 15116
rect 22278 15104 22284 15116
rect 22336 15104 22342 15156
rect 22465 15147 22523 15153
rect 22465 15113 22477 15147
rect 22511 15144 22523 15147
rect 23106 15144 23112 15156
rect 22511 15116 23112 15144
rect 22511 15113 22523 15116
rect 22465 15107 22523 15113
rect 23106 15104 23112 15116
rect 23164 15104 23170 15156
rect 23842 15104 23848 15156
rect 23900 15144 23906 15156
rect 25682 15144 25688 15156
rect 23900 15116 25688 15144
rect 23900 15104 23906 15116
rect 25682 15104 25688 15116
rect 25740 15104 25746 15156
rect 27065 15147 27123 15153
rect 27065 15113 27077 15147
rect 27111 15144 27123 15147
rect 30558 15144 30564 15156
rect 27111 15116 30564 15144
rect 27111 15113 27123 15116
rect 27065 15107 27123 15113
rect 30558 15104 30564 15116
rect 30616 15104 30622 15156
rect 31018 15104 31024 15156
rect 31076 15144 31082 15156
rect 31570 15144 31576 15156
rect 31076 15116 31576 15144
rect 31076 15104 31082 15116
rect 31570 15104 31576 15116
rect 31628 15104 31634 15156
rect 31846 15104 31852 15156
rect 31904 15144 31910 15156
rect 34422 15144 34428 15156
rect 31904 15116 34428 15144
rect 31904 15104 31910 15116
rect 34422 15104 34428 15116
rect 34480 15104 34486 15156
rect 35710 15104 35716 15156
rect 35768 15144 35774 15156
rect 37366 15144 37372 15156
rect 35768 15116 37372 15144
rect 35768 15104 35774 15116
rect 37366 15104 37372 15116
rect 37424 15104 37430 15156
rect 38194 15104 38200 15156
rect 38252 15144 38258 15156
rect 40586 15144 40592 15156
rect 38252 15116 40592 15144
rect 38252 15104 38258 15116
rect 40586 15104 40592 15116
rect 40644 15104 40650 15156
rect 43530 15144 43536 15156
rect 43491 15116 43536 15144
rect 43530 15104 43536 15116
rect 43588 15104 43594 15156
rect 43622 15104 43628 15156
rect 43680 15144 43686 15156
rect 44174 15144 44180 15156
rect 43680 15116 43852 15144
rect 44135 15116 44180 15144
rect 43680 15104 43686 15116
rect 19199 15048 20760 15076
rect 20824 15048 21220 15076
rect 21284 15048 21496 15076
rect 19199 15045 19211 15048
rect 19153 15039 19211 15045
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 11238 15008 11244 15020
rect 1719 14980 11244 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 11238 14968 11244 14980
rect 11296 14968 11302 15020
rect 17310 15008 17316 15020
rect 17271 14980 17316 15008
rect 17310 14968 17316 14980
rect 17368 14968 17374 15020
rect 18138 14968 18144 15020
rect 18196 15008 18202 15020
rect 18417 15011 18475 15017
rect 18417 15008 18429 15011
rect 18196 14980 18429 15008
rect 18196 14968 18202 14980
rect 18417 14977 18429 14980
rect 18463 14977 18475 15011
rect 19058 15008 19064 15020
rect 19019 14980 19064 15008
rect 18417 14971 18475 14977
rect 19058 14968 19064 14980
rect 19116 14968 19122 15020
rect 19242 15008 19248 15020
rect 19203 14980 19248 15008
rect 19242 14968 19248 14980
rect 19300 14968 19306 15020
rect 19889 15011 19947 15017
rect 19889 14977 19901 15011
rect 19935 15008 19947 15011
rect 20070 15008 20076 15020
rect 19935 14980 20076 15008
rect 19935 14977 19947 14980
rect 19889 14971 19947 14977
rect 20070 14968 20076 14980
rect 20128 14968 20134 15020
rect 16114 14900 16120 14952
rect 16172 14940 16178 14952
rect 16853 14943 16911 14949
rect 16853 14940 16865 14943
rect 16172 14912 16865 14940
rect 16172 14900 16178 14912
rect 16853 14909 16865 14912
rect 16899 14940 16911 14943
rect 18509 14943 18567 14949
rect 16899 14912 17954 14940
rect 16899 14909 16911 14912
rect 16853 14903 16911 14909
rect 1486 14872 1492 14884
rect 1447 14844 1492 14872
rect 1486 14832 1492 14844
rect 1544 14832 1550 14884
rect 15565 14875 15623 14881
rect 15565 14841 15577 14875
rect 15611 14872 15623 14875
rect 17218 14872 17224 14884
rect 15611 14844 17224 14872
rect 15611 14841 15623 14844
rect 15565 14835 15623 14841
rect 17218 14832 17224 14844
rect 17276 14832 17282 14884
rect 17926 14872 17954 14912
rect 18509 14909 18521 14943
rect 18555 14940 18567 14943
rect 19981 14943 20039 14949
rect 18555 14912 19932 14940
rect 18555 14909 18567 14912
rect 18509 14903 18567 14909
rect 18874 14872 18880 14884
rect 17926 14844 18880 14872
rect 18874 14832 18880 14844
rect 18932 14832 18938 14884
rect 18966 14832 18972 14884
rect 19024 14872 19030 14884
rect 19334 14872 19340 14884
rect 19024 14844 19340 14872
rect 19024 14832 19030 14844
rect 19334 14832 19340 14844
rect 19392 14832 19398 14884
rect 19904 14872 19932 14912
rect 19981 14909 19993 14943
rect 20027 14940 20039 14943
rect 20254 14940 20260 14952
rect 20027 14912 20260 14940
rect 20027 14909 20039 14912
rect 19981 14903 20039 14909
rect 20254 14900 20260 14912
rect 20312 14900 20318 14952
rect 20824 14949 20852 15048
rect 20979 15011 21037 15017
rect 20979 14977 20991 15011
rect 21025 15008 21037 15011
rect 21192 15008 21220 15048
rect 21542 15036 21548 15088
rect 21600 15076 21606 15088
rect 23934 15076 23940 15088
rect 21600 15048 23940 15076
rect 21600 15036 21606 15048
rect 23934 15036 23940 15048
rect 23992 15036 23998 15088
rect 24854 15036 24860 15088
rect 24912 15076 24918 15088
rect 24912 15048 25438 15076
rect 24912 15036 24918 15048
rect 28534 15036 28540 15088
rect 28592 15036 28598 15088
rect 28994 15076 29000 15088
rect 28955 15048 29000 15076
rect 28994 15036 29000 15048
rect 29052 15036 29058 15088
rect 29546 15076 29552 15088
rect 29288 15048 29552 15076
rect 21726 15008 21732 15020
rect 21025 14980 21128 15008
rect 21192 14980 21732 15008
rect 21025 14977 21037 14980
rect 20979 14971 21037 14977
rect 20809 14943 20867 14949
rect 20809 14909 20821 14943
rect 20855 14909 20867 14943
rect 21100 14940 21128 14980
rect 21726 14968 21732 14980
rect 21784 14968 21790 15020
rect 22094 14968 22100 15020
rect 22152 15008 22158 15020
rect 22557 15011 22615 15017
rect 22557 15008 22569 15011
rect 22152 14980 22569 15008
rect 22152 14968 22158 14980
rect 22557 14977 22569 14980
rect 22603 15008 22615 15011
rect 22646 15008 22652 15020
rect 22603 14980 22652 15008
rect 22603 14977 22615 14980
rect 22557 14971 22615 14977
rect 22646 14968 22652 14980
rect 22704 14968 22710 15020
rect 22922 14968 22928 15020
rect 22980 15008 22986 15020
rect 23198 15008 23204 15020
rect 22980 14980 23204 15008
rect 22980 14968 22986 14980
rect 23198 14968 23204 14980
rect 23256 14968 23262 15020
rect 23474 15008 23480 15020
rect 23308 14980 23480 15008
rect 22373 14943 22431 14949
rect 21100 14912 22324 14940
rect 20809 14903 20867 14909
rect 22296 14884 22324 14912
rect 22373 14909 22385 14943
rect 22419 14940 22431 14943
rect 23308 14940 23336 14980
rect 23474 14968 23480 14980
rect 23532 14968 23538 15020
rect 23661 15011 23719 15017
rect 23661 14977 23673 15011
rect 23707 15008 23719 15011
rect 23750 15008 23756 15020
rect 23707 14980 23756 15008
rect 23707 14977 23719 14980
rect 23661 14971 23719 14977
rect 23750 14968 23756 14980
rect 23808 15008 23814 15020
rect 24394 15008 24400 15020
rect 23808 14980 24400 15008
rect 23808 14968 23814 14980
rect 24394 14968 24400 14980
rect 24452 14968 24458 15020
rect 26786 15008 26792 15020
rect 26160 14980 26792 15008
rect 22419 14912 23336 14940
rect 22419 14909 22431 14912
rect 22373 14903 22431 14909
rect 23382 14900 23388 14952
rect 23440 14940 23446 14952
rect 24670 14940 24676 14952
rect 23440 14912 23485 14940
rect 24631 14912 24676 14940
rect 23440 14900 23446 14912
rect 24670 14900 24676 14912
rect 24728 14900 24734 14952
rect 24946 14940 24952 14952
rect 24907 14912 24952 14940
rect 24946 14900 24952 14912
rect 25004 14900 25010 14952
rect 25314 14900 25320 14952
rect 25372 14940 25378 14952
rect 26160 14940 26188 14980
rect 26786 14968 26792 14980
rect 26844 14968 26850 15020
rect 29288 15017 29316 15048
rect 29546 15036 29552 15048
rect 29604 15036 29610 15088
rect 29917 15079 29975 15085
rect 29917 15076 29929 15079
rect 29748 15048 29929 15076
rect 29273 15011 29331 15017
rect 29273 14977 29285 15011
rect 29319 14977 29331 15011
rect 29748 15008 29776 15048
rect 29917 15045 29929 15048
rect 29963 15045 29975 15079
rect 29917 15039 29975 15045
rect 30834 15036 30840 15088
rect 30892 15076 30898 15088
rect 31662 15076 31668 15088
rect 30892 15048 31668 15076
rect 30892 15036 30898 15048
rect 31662 15036 31668 15048
rect 31720 15036 31726 15088
rect 32309 15079 32367 15085
rect 32309 15045 32321 15079
rect 32355 15076 32367 15079
rect 32858 15076 32864 15088
rect 32355 15048 32864 15076
rect 32355 15045 32367 15048
rect 32309 15039 32367 15045
rect 32858 15036 32864 15048
rect 32916 15036 32922 15088
rect 32122 15008 32128 15020
rect 29273 14971 29331 14977
rect 29472 14980 29776 15008
rect 32083 14980 32128 15008
rect 25372 14912 26188 14940
rect 25372 14900 25378 14912
rect 26234 14900 26240 14952
rect 26292 14940 26298 14952
rect 29472 14940 29500 14980
rect 32122 14968 32128 14980
rect 32180 14968 32186 15020
rect 34440 15017 34468 15104
rect 35250 15036 35256 15088
rect 35308 15036 35314 15088
rect 36538 15036 36544 15088
rect 36596 15076 36602 15088
rect 36596 15048 41736 15076
rect 36596 15036 36602 15048
rect 34425 15011 34483 15017
rect 34425 14977 34437 15011
rect 34471 14977 34483 15011
rect 34425 14971 34483 14977
rect 37553 15011 37611 15017
rect 37553 14977 37565 15011
rect 37599 15008 37611 15011
rect 37642 15008 37648 15020
rect 37599 14980 37648 15008
rect 37599 14977 37611 14980
rect 37553 14971 37611 14977
rect 37642 14968 37648 14980
rect 37700 15008 37706 15020
rect 38194 15008 38200 15020
rect 37700 14980 37964 15008
rect 38155 14980 38200 15008
rect 37700 14968 37706 14980
rect 26292 14912 29500 14940
rect 29733 14943 29791 14949
rect 26292 14900 26298 14912
rect 29733 14909 29745 14943
rect 29779 14909 29791 14943
rect 30374 14940 30380 14952
rect 30335 14912 30380 14940
rect 29733 14903 29791 14909
rect 21818 14872 21824 14884
rect 19904 14844 21824 14872
rect 21818 14832 21824 14844
rect 21876 14832 21882 14884
rect 21910 14832 21916 14884
rect 21968 14872 21974 14884
rect 21968 14844 22232 14872
rect 21968 14832 21974 14844
rect 20162 14804 20168 14816
rect 20123 14776 20168 14804
rect 20162 14764 20168 14776
rect 20220 14764 20226 14816
rect 20346 14764 20352 14816
rect 20404 14804 20410 14816
rect 20622 14804 20628 14816
rect 20404 14776 20628 14804
rect 20404 14764 20410 14776
rect 20622 14764 20628 14776
rect 20680 14764 20686 14816
rect 21542 14764 21548 14816
rect 21600 14804 21606 14816
rect 22094 14804 22100 14816
rect 21600 14776 22100 14804
rect 21600 14764 21606 14776
rect 22094 14764 22100 14776
rect 22152 14764 22158 14816
rect 22204 14804 22232 14844
rect 22278 14832 22284 14884
rect 22336 14872 22342 14884
rect 22336 14844 23060 14872
rect 22336 14832 22342 14844
rect 22738 14804 22744 14816
rect 22204 14776 22744 14804
rect 22738 14764 22744 14776
rect 22796 14764 22802 14816
rect 22922 14804 22928 14816
rect 22883 14776 22928 14804
rect 22922 14764 22928 14776
rect 22980 14764 22986 14816
rect 23032 14804 23060 14844
rect 25976 14844 27660 14872
rect 25976 14804 26004 14844
rect 23032 14776 26004 14804
rect 26421 14807 26479 14813
rect 26421 14773 26433 14807
rect 26467 14804 26479 14807
rect 26694 14804 26700 14816
rect 26467 14776 26700 14804
rect 26467 14773 26479 14776
rect 26421 14767 26479 14773
rect 26694 14764 26700 14776
rect 26752 14764 26758 14816
rect 27522 14804 27528 14816
rect 27483 14776 27528 14804
rect 27522 14764 27528 14776
rect 27580 14764 27586 14816
rect 27632 14804 27660 14844
rect 29546 14832 29552 14884
rect 29604 14872 29610 14884
rect 29748 14872 29776 14903
rect 30374 14900 30380 14912
rect 30432 14940 30438 14952
rect 32585 14943 32643 14949
rect 32585 14940 32597 14943
rect 30432 14912 32597 14940
rect 30432 14900 30438 14912
rect 32585 14909 32597 14912
rect 32631 14940 32643 14943
rect 32674 14940 32680 14952
rect 32631 14912 32680 14940
rect 32631 14909 32643 14912
rect 32585 14903 32643 14909
rect 32674 14900 32680 14912
rect 32732 14940 32738 14952
rect 34146 14940 34152 14952
rect 32732 14912 34152 14940
rect 32732 14900 32738 14912
rect 34146 14900 34152 14912
rect 34204 14900 34210 14952
rect 34698 14940 34704 14952
rect 34659 14912 34704 14940
rect 34698 14900 34704 14912
rect 34756 14900 34762 14952
rect 36814 14900 36820 14952
rect 36872 14940 36878 14952
rect 37277 14943 37335 14949
rect 37277 14940 37289 14943
rect 36872 14912 37289 14940
rect 36872 14900 36878 14912
rect 37277 14909 37289 14912
rect 37323 14909 37335 14943
rect 37936 14940 37964 14980
rect 38194 14968 38200 14980
rect 38252 14968 38258 15020
rect 39209 15011 39267 15017
rect 39209 15008 39221 15011
rect 38856 14980 39221 15008
rect 38856 14940 38884 14980
rect 39209 14977 39221 14980
rect 39255 15008 39267 15011
rect 39390 15008 39396 15020
rect 39255 14980 39396 15008
rect 39255 14977 39267 14980
rect 39209 14971 39267 14977
rect 39390 14968 39396 14980
rect 39448 14968 39454 15020
rect 39853 15011 39911 15017
rect 39853 14977 39865 15011
rect 39899 14977 39911 15011
rect 39853 14971 39911 14977
rect 37936 14912 38884 14940
rect 38933 14943 38991 14949
rect 37277 14903 37335 14909
rect 38933 14909 38945 14943
rect 38979 14909 38991 14943
rect 39868 14940 39896 14971
rect 39942 14968 39948 15020
rect 40000 15008 40006 15020
rect 40129 15011 40187 15017
rect 40129 15008 40141 15011
rect 40000 14980 40141 15008
rect 40000 14968 40006 14980
rect 40129 14977 40141 14980
rect 40175 14977 40187 15011
rect 40129 14971 40187 14977
rect 40218 14968 40224 15020
rect 40276 15008 40282 15020
rect 40957 15011 41015 15017
rect 40957 15008 40969 15011
rect 40276 14980 40969 15008
rect 40276 14968 40282 14980
rect 40957 14977 40969 14980
rect 41003 14977 41015 15011
rect 40957 14971 41015 14977
rect 41046 14968 41052 15020
rect 41104 15008 41110 15020
rect 41601 15011 41659 15017
rect 41601 15008 41613 15011
rect 41104 14980 41613 15008
rect 41104 14968 41110 14980
rect 41601 14977 41613 14980
rect 41647 14977 41659 15011
rect 41708 15008 41736 15048
rect 41782 15036 41788 15088
rect 41840 15076 41846 15088
rect 42853 15079 42911 15085
rect 42853 15076 42865 15079
rect 41840 15048 42865 15076
rect 41840 15036 41846 15048
rect 42853 15045 42865 15048
rect 42899 15045 42911 15079
rect 42853 15039 42911 15045
rect 42996 15048 43760 15076
rect 41708 14998 42840 15008
rect 42996 14998 43024 15048
rect 43732 15017 43760 15048
rect 41708 14980 43024 14998
rect 41601 14971 41659 14977
rect 42812 14970 43024 14980
rect 43717 15011 43775 15017
rect 43717 14977 43729 15011
rect 43763 14977 43775 15011
rect 43824 15008 43852 15116
rect 44174 15104 44180 15116
rect 44232 15104 44238 15156
rect 46382 15144 46388 15156
rect 46343 15116 46388 15144
rect 46382 15104 46388 15116
rect 46440 15104 46446 15156
rect 46474 15104 46480 15156
rect 46532 15144 46538 15156
rect 47578 15144 47584 15156
rect 46532 15116 47584 15144
rect 46532 15104 46538 15116
rect 47578 15104 47584 15116
rect 47636 15104 47642 15156
rect 44082 15036 44088 15088
rect 44140 15076 44146 15088
rect 46658 15076 46664 15088
rect 44140 15048 46664 15076
rect 44140 15036 44146 15048
rect 46658 15036 46664 15048
rect 46716 15036 46722 15088
rect 46934 15076 46940 15088
rect 46895 15048 46940 15076
rect 46934 15036 46940 15048
rect 46992 15036 46998 15088
rect 58158 15076 58164 15088
rect 58119 15048 58164 15076
rect 58158 15036 58164 15048
rect 58216 15036 58222 15088
rect 44729 15011 44787 15017
rect 44729 15008 44741 15011
rect 43824 14980 44741 15008
rect 43717 14971 43775 14977
rect 44729 14977 44741 14980
rect 44775 15008 44787 15011
rect 45833 15011 45891 15017
rect 45833 15008 45845 15011
rect 44775 14980 45845 15008
rect 44775 14977 44787 14980
rect 44729 14971 44787 14977
rect 45833 14977 45845 14980
rect 45879 14977 45891 15011
rect 45833 14971 45891 14977
rect 40586 14940 40592 14952
rect 39868 14912 40592 14940
rect 38933 14903 38991 14909
rect 32030 14872 32036 14884
rect 29604 14844 32036 14872
rect 29604 14832 29610 14844
rect 32030 14832 32036 14844
rect 32088 14872 32094 14884
rect 33686 14872 33692 14884
rect 32088 14844 33692 14872
rect 32088 14832 32094 14844
rect 33686 14832 33692 14844
rect 33744 14832 33750 14884
rect 38948 14872 38976 14903
rect 40586 14900 40592 14912
rect 40644 14900 40650 14952
rect 40862 14940 40868 14952
rect 40823 14912 40868 14940
rect 40862 14900 40868 14912
rect 40920 14900 40926 14952
rect 41693 14943 41751 14949
rect 41693 14909 41705 14943
rect 41739 14940 41751 14943
rect 41782 14940 41788 14952
rect 41739 14912 41788 14940
rect 41739 14909 41751 14912
rect 41693 14903 41751 14909
rect 41782 14900 41788 14912
rect 41840 14900 41846 14952
rect 41877 14943 41935 14949
rect 41877 14909 41889 14943
rect 41923 14940 41935 14943
rect 41923 14912 42104 14940
rect 41923 14909 41935 14912
rect 41877 14903 41935 14909
rect 40770 14872 40776 14884
rect 35728 14844 36768 14872
rect 38948 14844 39068 14872
rect 33410 14804 33416 14816
rect 27632 14776 33416 14804
rect 33410 14764 33416 14776
rect 33468 14804 33474 14816
rect 35728 14804 35756 14844
rect 36170 14804 36176 14816
rect 33468 14776 35756 14804
rect 36131 14776 36176 14804
rect 33468 14764 33474 14776
rect 36170 14764 36176 14776
rect 36228 14764 36234 14816
rect 36630 14804 36636 14816
rect 36591 14776 36636 14804
rect 36630 14764 36636 14776
rect 36688 14764 36694 14816
rect 36740 14804 36768 14844
rect 37918 14804 37924 14816
rect 36740 14776 37924 14804
rect 37918 14764 37924 14776
rect 37976 14764 37982 14816
rect 38102 14764 38108 14816
rect 38160 14804 38166 14816
rect 38381 14807 38439 14813
rect 38381 14804 38393 14807
rect 38160 14776 38393 14804
rect 38160 14764 38166 14776
rect 38381 14773 38393 14776
rect 38427 14804 38439 14807
rect 38838 14804 38844 14816
rect 38427 14776 38844 14804
rect 38427 14773 38439 14776
rect 38381 14767 38439 14773
rect 38838 14764 38844 14776
rect 38896 14764 38902 14816
rect 39040 14804 39068 14844
rect 39500 14844 40776 14872
rect 39500 14804 39528 14844
rect 40770 14832 40776 14844
rect 40828 14832 40834 14884
rect 39040 14776 39528 14804
rect 40034 14764 40040 14816
rect 40092 14804 40098 14816
rect 40402 14804 40408 14816
rect 40092 14776 40408 14804
rect 40092 14764 40098 14776
rect 40402 14764 40408 14776
rect 40460 14764 40466 14816
rect 40678 14804 40684 14816
rect 40639 14776 40684 14804
rect 40678 14764 40684 14776
rect 40736 14764 40742 14816
rect 41782 14764 41788 14816
rect 41840 14804 41846 14816
rect 42076 14804 42104 14912
rect 42150 14900 42156 14952
rect 42208 14940 42214 14952
rect 42518 14940 42524 14952
rect 42208 14912 42524 14940
rect 42208 14900 42214 14912
rect 42518 14900 42524 14912
rect 42576 14940 42582 14952
rect 44174 14940 44180 14952
rect 42576 14912 44180 14940
rect 42576 14900 42582 14912
rect 44174 14900 44180 14912
rect 44232 14940 44238 14952
rect 44634 14940 44640 14952
rect 44232 14912 44640 14940
rect 44232 14900 44238 14912
rect 44634 14900 44640 14912
rect 44692 14900 44698 14952
rect 45278 14872 45284 14884
rect 45239 14844 45284 14872
rect 45278 14832 45284 14844
rect 45336 14832 45342 14884
rect 42886 14804 42892 14816
rect 41840 14776 41885 14804
rect 42076 14776 42892 14804
rect 41840 14764 41846 14776
rect 42886 14764 42892 14776
rect 42944 14764 42950 14816
rect 42981 14807 43039 14813
rect 42981 14773 42993 14807
rect 43027 14804 43039 14807
rect 43070 14804 43076 14816
rect 43027 14776 43076 14804
rect 43027 14773 43039 14776
rect 42981 14767 43039 14773
rect 43070 14764 43076 14776
rect 43128 14804 43134 14816
rect 44082 14804 44088 14816
rect 43128 14776 44088 14804
rect 43128 14764 43134 14776
rect 44082 14764 44088 14776
rect 44140 14764 44146 14816
rect 48130 14804 48136 14816
rect 48091 14776 48136 14804
rect 48130 14764 48136 14776
rect 48188 14764 48194 14816
rect 1104 14714 58880 14736
rect 1104 14662 10582 14714
rect 10634 14662 10646 14714
rect 10698 14662 10710 14714
rect 10762 14662 10774 14714
rect 10826 14662 10838 14714
rect 10890 14662 29846 14714
rect 29898 14662 29910 14714
rect 29962 14662 29974 14714
rect 30026 14662 30038 14714
rect 30090 14662 30102 14714
rect 30154 14662 49110 14714
rect 49162 14662 49174 14714
rect 49226 14662 49238 14714
rect 49290 14662 49302 14714
rect 49354 14662 49366 14714
rect 49418 14662 58880 14714
rect 1104 14640 58880 14662
rect 14274 14600 14280 14612
rect 14235 14572 14280 14600
rect 14274 14560 14280 14572
rect 14332 14560 14338 14612
rect 15378 14600 15384 14612
rect 15339 14572 15384 14600
rect 15378 14560 15384 14572
rect 15436 14560 15442 14612
rect 15470 14560 15476 14612
rect 15528 14600 15534 14612
rect 15841 14603 15899 14609
rect 15841 14600 15853 14603
rect 15528 14572 15853 14600
rect 15528 14560 15534 14572
rect 15841 14569 15853 14572
rect 15887 14569 15899 14603
rect 15841 14563 15899 14569
rect 17589 14603 17647 14609
rect 17589 14569 17601 14603
rect 17635 14600 17647 14603
rect 19518 14600 19524 14612
rect 17635 14572 19524 14600
rect 17635 14569 17647 14572
rect 17589 14563 17647 14569
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 19705 14603 19763 14609
rect 19705 14569 19717 14603
rect 19751 14600 19763 14603
rect 24486 14600 24492 14612
rect 19751 14572 23520 14600
rect 24447 14572 24492 14600
rect 19751 14569 19763 14572
rect 19705 14563 19763 14569
rect 18693 14535 18751 14541
rect 18693 14501 18705 14535
rect 18739 14532 18751 14535
rect 19058 14532 19064 14544
rect 18739 14504 19064 14532
rect 18739 14501 18751 14504
rect 18693 14495 18751 14501
rect 19058 14492 19064 14504
rect 19116 14492 19122 14544
rect 19242 14492 19248 14544
rect 19300 14532 19306 14544
rect 19610 14532 19616 14544
rect 19300 14504 19616 14532
rect 19300 14492 19306 14504
rect 19610 14492 19616 14504
rect 19668 14492 19674 14544
rect 20346 14532 20352 14544
rect 20307 14504 20352 14532
rect 20346 14492 20352 14504
rect 20404 14492 20410 14544
rect 20438 14492 20444 14544
rect 20496 14532 20502 14544
rect 20622 14532 20628 14544
rect 20496 14504 20628 14532
rect 20496 14492 20502 14504
rect 20622 14492 20628 14504
rect 20680 14492 20686 14544
rect 20714 14492 20720 14544
rect 20772 14532 20778 14544
rect 20772 14504 21220 14532
rect 20772 14492 20778 14504
rect 20070 14424 20076 14476
rect 20128 14464 20134 14476
rect 20257 14467 20315 14473
rect 20257 14464 20269 14467
rect 20128 14436 20269 14464
rect 20128 14424 20134 14436
rect 20257 14433 20269 14436
rect 20303 14464 20315 14467
rect 20806 14464 20812 14476
rect 20303 14436 20812 14464
rect 20303 14433 20315 14436
rect 20257 14427 20315 14433
rect 20806 14424 20812 14436
rect 20864 14424 20870 14476
rect 21085 14467 21143 14473
rect 21085 14433 21097 14467
rect 21131 14433 21143 14467
rect 21192 14464 21220 14504
rect 21266 14492 21272 14544
rect 21324 14532 21330 14544
rect 22830 14532 22836 14544
rect 21324 14504 22836 14532
rect 21324 14492 21330 14504
rect 22830 14492 22836 14504
rect 22888 14532 22894 14544
rect 23247 14535 23305 14541
rect 23247 14532 23259 14535
rect 22888 14504 23259 14532
rect 22888 14492 22894 14504
rect 23247 14501 23259 14504
rect 23293 14501 23305 14535
rect 23492 14532 23520 14572
rect 24486 14560 24492 14572
rect 24544 14560 24550 14612
rect 25130 14560 25136 14612
rect 25188 14600 25194 14612
rect 29638 14600 29644 14612
rect 25188 14572 29644 14600
rect 25188 14560 25194 14572
rect 29638 14560 29644 14572
rect 29696 14560 29702 14612
rect 32582 14600 32588 14612
rect 29840 14572 32588 14600
rect 29840 14544 29868 14572
rect 32582 14560 32588 14572
rect 32640 14560 32646 14612
rect 33870 14560 33876 14612
rect 33928 14600 33934 14612
rect 38657 14603 38715 14609
rect 38657 14600 38669 14603
rect 33928 14572 38669 14600
rect 33928 14560 33934 14572
rect 38657 14569 38669 14572
rect 38703 14569 38715 14603
rect 40218 14600 40224 14612
rect 38657 14563 38715 14569
rect 38764 14572 40224 14600
rect 25038 14532 25044 14544
rect 23492 14504 25044 14532
rect 23247 14495 23305 14501
rect 25038 14492 25044 14504
rect 25096 14492 25102 14544
rect 26418 14492 26424 14544
rect 26476 14532 26482 14544
rect 26789 14535 26847 14541
rect 26789 14532 26801 14535
rect 26476 14504 26801 14532
rect 26476 14492 26482 14504
rect 26789 14501 26801 14504
rect 26835 14532 26847 14535
rect 26878 14532 26884 14544
rect 26835 14504 26884 14532
rect 26835 14501 26847 14504
rect 26789 14495 26847 14501
rect 26878 14492 26884 14504
rect 26936 14492 26942 14544
rect 27249 14535 27307 14541
rect 27249 14501 27261 14535
rect 27295 14532 27307 14535
rect 27338 14532 27344 14544
rect 27295 14504 27344 14532
rect 27295 14501 27307 14504
rect 27249 14495 27307 14501
rect 27338 14492 27344 14504
rect 27396 14492 27402 14544
rect 29822 14492 29828 14544
rect 29880 14492 29886 14544
rect 30668 14504 31708 14532
rect 21542 14464 21548 14476
rect 21192 14436 21548 14464
rect 21085 14427 21143 14433
rect 10781 14399 10839 14405
rect 10781 14365 10793 14399
rect 10827 14396 10839 14399
rect 10827 14368 11376 14396
rect 10827 14365 10839 14368
rect 10781 14359 10839 14365
rect 10594 14260 10600 14272
rect 10555 14232 10600 14260
rect 10594 14220 10600 14232
rect 10652 14220 10658 14272
rect 11348 14269 11376 14368
rect 19518 14356 19524 14408
rect 19576 14396 19582 14408
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 19576 14368 19625 14396
rect 19576 14356 19582 14368
rect 19613 14365 19625 14368
rect 19659 14396 19671 14399
rect 19978 14396 19984 14408
rect 19659 14368 19984 14396
rect 19659 14365 19671 14368
rect 19613 14359 19671 14365
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 20162 14356 20168 14408
rect 20220 14396 20226 14408
rect 20220 14368 20484 14396
rect 20220 14356 20226 14368
rect 18141 14331 18199 14337
rect 18141 14297 18153 14331
rect 18187 14328 18199 14331
rect 18322 14328 18328 14340
rect 18187 14300 18328 14328
rect 18187 14297 18199 14300
rect 18141 14291 18199 14297
rect 18322 14288 18328 14300
rect 18380 14328 18386 14340
rect 20346 14328 20352 14340
rect 18380 14300 20352 14328
rect 18380 14288 18386 14300
rect 20346 14288 20352 14300
rect 20404 14288 20410 14340
rect 20456 14328 20484 14368
rect 20530 14356 20536 14408
rect 20588 14396 20594 14408
rect 20588 14368 20632 14396
rect 20588 14356 20594 14368
rect 20898 14356 20904 14408
rect 20956 14396 20962 14408
rect 21100 14396 21128 14427
rect 21542 14424 21548 14436
rect 21600 14424 21606 14476
rect 21818 14424 21824 14476
rect 21876 14464 21882 14476
rect 22278 14464 22284 14476
rect 21876 14436 22284 14464
rect 21876 14424 21882 14436
rect 22278 14424 22284 14436
rect 22336 14424 22342 14476
rect 22557 14467 22615 14473
rect 22557 14433 22569 14467
rect 22603 14464 22615 14467
rect 25317 14467 25375 14473
rect 25317 14464 25329 14467
rect 22603 14436 25329 14464
rect 22603 14433 22615 14436
rect 22557 14427 22615 14433
rect 25317 14433 25329 14436
rect 25363 14433 25375 14467
rect 28997 14467 29055 14473
rect 28997 14464 29009 14467
rect 25317 14427 25375 14433
rect 26620 14436 29009 14464
rect 21266 14405 21272 14408
rect 20956 14368 21128 14396
rect 21255 14399 21272 14405
rect 20956 14356 20962 14368
rect 21255 14365 21267 14399
rect 21255 14359 21272 14365
rect 21266 14356 21272 14359
rect 21324 14356 21330 14408
rect 21358 14356 21364 14408
rect 21416 14396 21422 14408
rect 21416 14368 22048 14396
rect 21416 14356 21422 14368
rect 21910 14328 21916 14340
rect 20456 14300 21916 14328
rect 21910 14288 21916 14300
rect 21968 14288 21974 14340
rect 22020 14328 22048 14368
rect 22094 14356 22100 14408
rect 22152 14398 22158 14408
rect 22189 14399 22247 14405
rect 22189 14398 22201 14399
rect 22152 14370 22201 14398
rect 22152 14356 22158 14370
rect 22189 14365 22201 14370
rect 22235 14365 22247 14399
rect 22189 14359 22247 14365
rect 23017 14399 23075 14405
rect 23017 14365 23029 14399
rect 23063 14396 23075 14399
rect 23198 14396 23204 14408
rect 23063 14368 23204 14396
rect 23063 14365 23075 14368
rect 23017 14359 23075 14365
rect 23198 14356 23204 14368
rect 23256 14396 23262 14408
rect 23382 14396 23388 14408
rect 23256 14368 23388 14396
rect 23256 14356 23262 14368
rect 23382 14356 23388 14368
rect 23440 14356 23446 14408
rect 24578 14396 24584 14408
rect 24539 14368 24584 14396
rect 24578 14356 24584 14368
rect 24636 14356 24642 14408
rect 25041 14399 25099 14405
rect 25041 14365 25053 14399
rect 25087 14365 25099 14399
rect 25041 14359 25099 14365
rect 22462 14328 22468 14340
rect 22020 14300 22468 14328
rect 22462 14288 22468 14300
rect 22520 14288 22526 14340
rect 23290 14288 23296 14340
rect 23348 14328 23354 14340
rect 25056 14328 25084 14359
rect 25314 14328 25320 14340
rect 23348 14300 25320 14328
rect 23348 14288 23354 14300
rect 25314 14288 25320 14300
rect 25372 14288 25378 14340
rect 25958 14288 25964 14340
rect 26016 14288 26022 14340
rect 11333 14263 11391 14269
rect 11333 14229 11345 14263
rect 11379 14260 11391 14263
rect 12618 14260 12624 14272
rect 11379 14232 12624 14260
rect 11379 14229 11391 14232
rect 11333 14223 11391 14229
rect 12618 14220 12624 14232
rect 12676 14260 12682 14272
rect 13722 14260 13728 14272
rect 12676 14232 13728 14260
rect 12676 14220 12682 14232
rect 13722 14220 13728 14232
rect 13780 14220 13786 14272
rect 14829 14263 14887 14269
rect 14829 14229 14841 14263
rect 14875 14260 14887 14263
rect 14918 14260 14924 14272
rect 14875 14232 14924 14260
rect 14875 14229 14887 14232
rect 14829 14223 14887 14229
rect 14918 14220 14924 14232
rect 14976 14220 14982 14272
rect 16390 14260 16396 14272
rect 16351 14232 16396 14260
rect 16390 14220 16396 14232
rect 16448 14220 16454 14272
rect 17037 14263 17095 14269
rect 17037 14229 17049 14263
rect 17083 14260 17095 14263
rect 19058 14260 19064 14272
rect 17083 14232 19064 14260
rect 17083 14229 17095 14232
rect 17037 14223 17095 14229
rect 19058 14220 19064 14232
rect 19116 14220 19122 14272
rect 19334 14220 19340 14272
rect 19392 14260 19398 14272
rect 20714 14260 20720 14272
rect 19392 14232 20720 14260
rect 19392 14220 19398 14232
rect 20714 14220 20720 14232
rect 20772 14220 20778 14272
rect 21542 14260 21548 14272
rect 21503 14232 21548 14260
rect 21542 14220 21548 14232
rect 21600 14220 21606 14272
rect 22094 14220 22100 14272
rect 22152 14260 22158 14272
rect 24210 14260 24216 14272
rect 22152 14232 24216 14260
rect 22152 14220 22158 14232
rect 24210 14220 24216 14232
rect 24268 14220 24274 14272
rect 24486 14220 24492 14272
rect 24544 14260 24550 14272
rect 26620 14260 26648 14436
rect 28997 14433 29009 14436
rect 29043 14464 29055 14467
rect 30668 14464 30696 14504
rect 29043 14436 29224 14464
rect 29043 14433 29055 14436
rect 28997 14427 29055 14433
rect 28258 14288 28264 14340
rect 28316 14288 28322 14340
rect 28626 14288 28632 14340
rect 28684 14328 28690 14340
rect 28721 14331 28779 14337
rect 28721 14328 28733 14331
rect 28684 14300 28733 14328
rect 28684 14288 28690 14300
rect 28721 14297 28733 14300
rect 28767 14297 28779 14331
rect 29196 14328 29224 14436
rect 29564 14436 30696 14464
rect 29564 14408 29592 14436
rect 30742 14424 30748 14476
rect 30800 14464 30806 14476
rect 30837 14467 30895 14473
rect 30837 14464 30849 14467
rect 30800 14436 30849 14464
rect 30800 14424 30806 14436
rect 30837 14433 30849 14436
rect 30883 14433 30895 14467
rect 30837 14427 30895 14433
rect 31021 14467 31079 14473
rect 31021 14433 31033 14467
rect 31067 14464 31079 14467
rect 31110 14464 31116 14476
rect 31067 14436 31116 14464
rect 31067 14433 31079 14436
rect 31021 14427 31079 14433
rect 31110 14424 31116 14436
rect 31168 14424 31174 14476
rect 31680 14464 31708 14504
rect 31754 14492 31760 14544
rect 31812 14532 31818 14544
rect 34514 14532 34520 14544
rect 31812 14504 34520 14532
rect 31812 14492 31818 14504
rect 34514 14492 34520 14504
rect 34572 14492 34578 14544
rect 36446 14532 36452 14544
rect 36407 14504 36452 14532
rect 36446 14492 36452 14504
rect 36504 14492 36510 14544
rect 37918 14492 37924 14544
rect 37976 14532 37982 14544
rect 38764 14532 38792 14572
rect 40218 14560 40224 14572
rect 40276 14560 40282 14612
rect 40586 14560 40592 14612
rect 40644 14600 40650 14612
rect 40862 14600 40868 14612
rect 40644 14572 40868 14600
rect 40644 14560 40650 14572
rect 40862 14560 40868 14572
rect 40920 14560 40926 14612
rect 41046 14600 41052 14612
rect 41007 14572 41052 14600
rect 41046 14560 41052 14572
rect 41104 14560 41110 14612
rect 41322 14560 41328 14612
rect 41380 14600 41386 14612
rect 41506 14600 41512 14612
rect 41380 14572 41512 14600
rect 41380 14560 41386 14572
rect 41506 14560 41512 14572
rect 41564 14600 41570 14612
rect 42889 14603 42947 14609
rect 42889 14600 42901 14603
rect 41564 14572 42901 14600
rect 41564 14560 41570 14572
rect 42889 14569 42901 14572
rect 42935 14600 42947 14603
rect 42935 14572 43576 14600
rect 42935 14569 42947 14572
rect 42889 14563 42947 14569
rect 39853 14535 39911 14541
rect 39853 14532 39865 14535
rect 37976 14504 38792 14532
rect 38856 14504 39865 14532
rect 37976 14492 37982 14504
rect 33689 14467 33747 14473
rect 33689 14464 33701 14467
rect 31680 14436 33701 14464
rect 33689 14433 33701 14436
rect 33735 14464 33747 14467
rect 36354 14464 36360 14476
rect 33735 14436 36360 14464
rect 33735 14433 33747 14436
rect 33689 14427 33747 14433
rect 36354 14424 36360 14436
rect 36412 14424 36418 14476
rect 38562 14424 38568 14476
rect 38620 14464 38626 14476
rect 38856 14464 38884 14504
rect 39853 14501 39865 14504
rect 39899 14501 39911 14535
rect 40126 14532 40132 14544
rect 39853 14495 39911 14501
rect 40052 14504 40132 14532
rect 38620 14436 38884 14464
rect 39025 14467 39083 14473
rect 38620 14424 38626 14436
rect 39025 14433 39037 14467
rect 39071 14464 39083 14467
rect 39390 14464 39396 14476
rect 39071 14436 39396 14464
rect 39071 14433 39083 14436
rect 39025 14427 39083 14433
rect 39390 14424 39396 14436
rect 39448 14424 39454 14476
rect 40052 14464 40080 14504
rect 40126 14492 40132 14504
rect 40184 14492 40190 14544
rect 40954 14532 40960 14544
rect 40788 14504 40960 14532
rect 40788 14473 40816 14504
rect 40954 14492 40960 14504
rect 41012 14532 41018 14544
rect 42978 14532 42984 14544
rect 41012 14504 42984 14532
rect 41012 14492 41018 14504
rect 42978 14492 42984 14504
rect 43036 14492 43042 14544
rect 43548 14541 43576 14572
rect 44358 14560 44364 14612
rect 44416 14600 44422 14612
rect 45005 14603 45063 14609
rect 45005 14600 45017 14603
rect 44416 14572 45017 14600
rect 44416 14560 44422 14572
rect 45005 14569 45017 14572
rect 45051 14569 45063 14603
rect 45005 14563 45063 14569
rect 45186 14560 45192 14612
rect 45244 14600 45250 14612
rect 46661 14603 46719 14609
rect 46661 14600 46673 14603
rect 45244 14572 46673 14600
rect 45244 14560 45250 14572
rect 46661 14569 46673 14572
rect 46707 14569 46719 14603
rect 46661 14563 46719 14569
rect 43533 14535 43591 14541
rect 43533 14501 43545 14535
rect 43579 14532 43591 14535
rect 46198 14532 46204 14544
rect 43579 14504 46204 14532
rect 43579 14501 43591 14504
rect 43533 14495 43591 14501
rect 46198 14492 46204 14504
rect 46256 14492 46262 14544
rect 40773 14467 40831 14473
rect 40052 14436 40172 14464
rect 29546 14396 29552 14408
rect 29507 14368 29552 14396
rect 29546 14356 29552 14368
rect 29604 14356 29610 14408
rect 29825 14399 29883 14405
rect 29825 14365 29837 14399
rect 29871 14396 29883 14399
rect 29914 14396 29920 14408
rect 29871 14368 29920 14396
rect 29871 14365 29883 14368
rect 29825 14359 29883 14365
rect 29914 14356 29920 14368
rect 29972 14396 29978 14408
rect 30650 14396 30656 14408
rect 29972 14368 30656 14396
rect 29972 14356 29978 14368
rect 30650 14356 30656 14368
rect 30708 14356 30714 14408
rect 32677 14399 32735 14405
rect 32677 14365 32689 14399
rect 32723 14396 32735 14399
rect 33134 14396 33140 14408
rect 32723 14368 33140 14396
rect 32723 14365 32735 14368
rect 32677 14359 32735 14365
rect 33134 14356 33140 14368
rect 33192 14356 33198 14408
rect 33962 14396 33968 14408
rect 33923 14368 33968 14396
rect 33962 14356 33968 14368
rect 34020 14356 34026 14408
rect 34514 14356 34520 14408
rect 34572 14396 34578 14408
rect 34701 14399 34759 14405
rect 34701 14396 34713 14399
rect 34572 14368 34713 14396
rect 34572 14356 34578 14368
rect 34701 14365 34713 14368
rect 34747 14365 34759 14399
rect 34701 14359 34759 14365
rect 36078 14356 36084 14408
rect 36136 14356 36142 14408
rect 36814 14356 36820 14408
rect 36872 14396 36878 14408
rect 36909 14399 36967 14405
rect 36909 14396 36921 14399
rect 36872 14368 36921 14396
rect 36872 14356 36878 14368
rect 36909 14365 36921 14368
rect 36955 14365 36967 14399
rect 36909 14359 36967 14365
rect 37090 14356 37096 14408
rect 37148 14396 37154 14408
rect 37185 14399 37243 14405
rect 37185 14396 37197 14399
rect 37148 14368 37197 14396
rect 37148 14356 37154 14368
rect 37185 14365 37197 14368
rect 37231 14396 37243 14399
rect 37642 14396 37648 14408
rect 37231 14368 37648 14396
rect 37231 14365 37243 14368
rect 37185 14359 37243 14365
rect 37642 14356 37648 14368
rect 37700 14356 37706 14408
rect 37829 14399 37887 14405
rect 37829 14365 37841 14399
rect 37875 14396 37887 14399
rect 38194 14396 38200 14408
rect 37875 14368 38200 14396
rect 37875 14365 37887 14368
rect 37829 14359 37887 14365
rect 34146 14328 34152 14340
rect 29196 14300 34152 14328
rect 28721 14291 28779 14297
rect 34146 14288 34152 14300
rect 34204 14288 34210 14340
rect 34974 14288 34980 14340
rect 35032 14328 35038 14340
rect 35032 14300 35077 14328
rect 36280 14300 36584 14328
rect 35032 14288 35038 14300
rect 24544 14232 26648 14260
rect 24544 14220 24550 14232
rect 27154 14220 27160 14272
rect 27212 14260 27218 14272
rect 30374 14260 30380 14272
rect 27212 14232 30380 14260
rect 27212 14220 27218 14232
rect 30374 14220 30380 14232
rect 30432 14220 30438 14272
rect 30650 14220 30656 14272
rect 30708 14260 30714 14272
rect 32398 14260 32404 14272
rect 30708 14232 32404 14260
rect 30708 14220 30714 14232
rect 32398 14220 32404 14232
rect 32456 14220 32462 14272
rect 33778 14220 33784 14272
rect 33836 14260 33842 14272
rect 36280 14260 36308 14300
rect 33836 14232 36308 14260
rect 36556 14260 36584 14300
rect 37366 14288 37372 14340
rect 37424 14328 37430 14340
rect 37844 14328 37872 14359
rect 38194 14356 38200 14368
rect 38252 14356 38258 14408
rect 38855 14399 38913 14405
rect 38855 14365 38867 14399
rect 38901 14365 38913 14399
rect 38855 14359 38913 14365
rect 37918 14328 37924 14340
rect 37424 14300 37924 14328
rect 37424 14288 37430 14300
rect 37918 14288 37924 14300
rect 37976 14288 37982 14340
rect 38102 14328 38108 14340
rect 38063 14300 38108 14328
rect 38102 14288 38108 14300
rect 38160 14288 38166 14340
rect 38746 14288 38752 14340
rect 38804 14328 38810 14340
rect 38856 14328 38884 14359
rect 39758 14356 39764 14408
rect 39816 14396 39822 14408
rect 40144 14405 40172 14436
rect 40773 14433 40785 14467
rect 40819 14433 40831 14467
rect 40773 14427 40831 14433
rect 40862 14424 40868 14476
rect 40920 14464 40926 14476
rect 43993 14467 44051 14473
rect 43993 14464 44005 14467
rect 40920 14436 44005 14464
rect 40920 14424 40926 14436
rect 40037 14399 40095 14405
rect 40037 14398 40049 14399
rect 39960 14396 40049 14398
rect 39816 14370 40049 14396
rect 39816 14368 39988 14370
rect 39816 14356 39822 14368
rect 40037 14365 40049 14370
rect 40083 14365 40095 14399
rect 40037 14359 40095 14365
rect 40129 14399 40187 14405
rect 40129 14365 40141 14399
rect 40175 14365 40187 14399
rect 40129 14359 40187 14365
rect 40221 14399 40279 14405
rect 40221 14365 40233 14399
rect 40267 14396 40279 14399
rect 40402 14396 40408 14408
rect 40267 14368 40408 14396
rect 40267 14365 40279 14368
rect 40221 14359 40279 14365
rect 40402 14356 40408 14368
rect 40460 14356 40466 14408
rect 40954 14396 40960 14408
rect 40915 14368 40960 14396
rect 40954 14356 40960 14368
rect 41012 14356 41018 14408
rect 41064 14405 41092 14436
rect 43993 14433 44005 14436
rect 44039 14433 44051 14467
rect 48314 14464 48320 14476
rect 43993 14427 44051 14433
rect 48240 14436 48320 14464
rect 41049 14399 41107 14405
rect 41049 14365 41061 14399
rect 41095 14365 41107 14399
rect 41690 14396 41696 14408
rect 41651 14368 41696 14396
rect 41049 14359 41107 14365
rect 41690 14356 41696 14368
rect 41748 14356 41754 14408
rect 42242 14396 42248 14408
rect 42203 14368 42248 14396
rect 42242 14356 42248 14368
rect 42300 14356 42306 14408
rect 46566 14396 46572 14408
rect 44560 14368 46572 14396
rect 38804 14300 38884 14328
rect 38804 14288 38810 14300
rect 40770 14288 40776 14340
rect 40828 14328 40834 14340
rect 41708 14328 41736 14356
rect 44560 14328 44588 14368
rect 46566 14356 46572 14368
rect 46624 14356 46630 14408
rect 40828 14300 41736 14328
rect 42168 14300 44588 14328
rect 40828 14288 40834 14300
rect 41506 14260 41512 14272
rect 36556 14232 41512 14260
rect 33836 14220 33842 14232
rect 41506 14220 41512 14232
rect 41564 14220 41570 14272
rect 41601 14263 41659 14269
rect 41601 14229 41613 14263
rect 41647 14260 41659 14263
rect 42168 14260 42196 14300
rect 44634 14288 44640 14340
rect 44692 14328 44698 14340
rect 47213 14331 47271 14337
rect 47213 14328 47225 14331
rect 44692 14300 47225 14328
rect 44692 14288 44698 14300
rect 47213 14297 47225 14300
rect 47259 14328 47271 14331
rect 47765 14331 47823 14337
rect 47765 14328 47777 14331
rect 47259 14300 47777 14328
rect 47259 14297 47271 14300
rect 47213 14291 47271 14297
rect 47765 14297 47777 14300
rect 47811 14328 47823 14331
rect 48130 14328 48136 14340
rect 47811 14300 48136 14328
rect 47811 14297 47823 14300
rect 47765 14291 47823 14297
rect 48130 14288 48136 14300
rect 48188 14288 48194 14340
rect 42334 14260 42340 14272
rect 41647 14232 42196 14260
rect 42295 14232 42340 14260
rect 41647 14229 41659 14232
rect 41601 14223 41659 14229
rect 42334 14220 42340 14232
rect 42392 14220 42398 14272
rect 45554 14260 45560 14272
rect 45515 14232 45560 14260
rect 45554 14220 45560 14232
rect 45612 14220 45618 14272
rect 45922 14220 45928 14272
rect 45980 14260 45986 14272
rect 46109 14263 46167 14269
rect 46109 14260 46121 14263
rect 45980 14232 46121 14260
rect 45980 14220 45986 14232
rect 46109 14229 46121 14232
rect 46155 14260 46167 14263
rect 48240 14260 48268 14436
rect 48314 14424 48320 14436
rect 48372 14424 48378 14476
rect 46155 14232 48268 14260
rect 46155 14229 46167 14232
rect 46109 14223 46167 14229
rect 1104 14170 58880 14192
rect 1104 14118 20214 14170
rect 20266 14118 20278 14170
rect 20330 14118 20342 14170
rect 20394 14118 20406 14170
rect 20458 14118 20470 14170
rect 20522 14118 39478 14170
rect 39530 14118 39542 14170
rect 39594 14118 39606 14170
rect 39658 14118 39670 14170
rect 39722 14118 39734 14170
rect 39786 14118 58880 14170
rect 1104 14096 58880 14118
rect 14458 14016 14464 14068
rect 14516 14056 14522 14068
rect 15102 14056 15108 14068
rect 14516 14028 15108 14056
rect 14516 14016 14522 14028
rect 15102 14016 15108 14028
rect 15160 14016 15166 14068
rect 16117 14059 16175 14065
rect 16117 14025 16129 14059
rect 16163 14056 16175 14059
rect 16482 14056 16488 14068
rect 16163 14028 16488 14056
rect 16163 14025 16175 14028
rect 16117 14019 16175 14025
rect 16482 14016 16488 14028
rect 16540 14056 16546 14068
rect 16666 14056 16672 14068
rect 16540 14028 16672 14056
rect 16540 14016 16546 14028
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 17770 14056 17776 14068
rect 17731 14028 17776 14056
rect 17770 14016 17776 14028
rect 17828 14016 17834 14068
rect 18322 14056 18328 14068
rect 18283 14028 18328 14056
rect 18322 14016 18328 14028
rect 18380 14016 18386 14068
rect 19429 14059 19487 14065
rect 19429 14025 19441 14059
rect 19475 14056 19487 14059
rect 19610 14056 19616 14068
rect 19475 14028 19616 14056
rect 19475 14025 19487 14028
rect 19429 14019 19487 14025
rect 19610 14016 19616 14028
rect 19668 14016 19674 14068
rect 20990 14016 20996 14068
rect 21048 14056 21054 14068
rect 21821 14059 21879 14065
rect 21821 14056 21833 14059
rect 21048 14028 21833 14056
rect 21048 14016 21054 14028
rect 21821 14025 21833 14028
rect 21867 14025 21879 14059
rect 24486 14056 24492 14068
rect 21821 14019 21879 14025
rect 22020 14028 24492 14056
rect 16390 13948 16396 14000
rect 16448 13988 16454 14000
rect 17221 13991 17279 13997
rect 17221 13988 17233 13991
rect 16448 13960 17233 13988
rect 16448 13948 16454 13960
rect 17221 13957 17233 13960
rect 17267 13988 17279 13991
rect 17954 13988 17960 14000
rect 17267 13960 17960 13988
rect 17267 13957 17279 13960
rect 17221 13951 17279 13957
rect 17954 13948 17960 13960
rect 18012 13948 18018 14000
rect 18877 13991 18935 13997
rect 18877 13957 18889 13991
rect 18923 13988 18935 13991
rect 18923 13960 21036 13988
rect 18923 13957 18935 13960
rect 18877 13951 18935 13957
rect 21008 13932 21036 13960
rect 21174 13948 21180 14000
rect 21232 13988 21238 14000
rect 21269 13991 21327 13997
rect 21269 13988 21281 13991
rect 21232 13960 21281 13988
rect 21232 13948 21238 13960
rect 21269 13957 21281 13960
rect 21315 13957 21327 13991
rect 21269 13951 21327 13957
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 10594 13920 10600 13932
rect 1719 13892 10600 13920
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 10594 13880 10600 13892
rect 10652 13880 10658 13932
rect 13722 13880 13728 13932
rect 13780 13920 13786 13932
rect 15565 13923 15623 13929
rect 15565 13920 15577 13923
rect 13780 13892 15577 13920
rect 13780 13880 13786 13892
rect 15565 13889 15577 13892
rect 15611 13920 15623 13923
rect 15611 13892 19334 13920
rect 15611 13889 15623 13892
rect 15565 13883 15623 13889
rect 13630 13812 13636 13864
rect 13688 13852 13694 13864
rect 14734 13852 14740 13864
rect 13688 13824 14740 13852
rect 13688 13812 13694 13824
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 19306 13784 19334 13892
rect 19978 13880 19984 13932
rect 20036 13920 20042 13932
rect 20530 13920 20536 13932
rect 20036 13892 20536 13920
rect 20036 13880 20042 13892
rect 20530 13880 20536 13892
rect 20588 13880 20594 13932
rect 20990 13920 20996 13932
rect 20951 13892 20996 13920
rect 20990 13880 20996 13892
rect 21048 13880 21054 13932
rect 20438 13852 20444 13864
rect 20399 13824 20444 13852
rect 20438 13812 20444 13824
rect 20496 13812 20502 13864
rect 20806 13812 20812 13864
rect 20864 13852 20870 13864
rect 21269 13855 21327 13861
rect 21269 13852 21281 13855
rect 20864 13824 21281 13852
rect 20864 13812 20870 13824
rect 21269 13821 21281 13824
rect 21315 13821 21327 13855
rect 22020 13852 22048 14028
rect 24486 14016 24492 14028
rect 24544 14016 24550 14068
rect 24578 14016 24584 14068
rect 24636 14056 24642 14068
rect 25958 14056 25964 14068
rect 24636 14028 25964 14056
rect 24636 14016 24642 14028
rect 25222 13988 25228 14000
rect 22848 13960 24532 13988
rect 22848 13932 22876 13960
rect 22186 13880 22192 13932
rect 22244 13920 22250 13932
rect 22830 13920 22836 13932
rect 22244 13892 22289 13920
rect 22743 13892 22836 13920
rect 22244 13880 22250 13892
rect 22830 13880 22836 13892
rect 22888 13880 22894 13932
rect 23014 13880 23020 13932
rect 23072 13920 23078 13932
rect 23842 13920 23848 13932
rect 23072 13892 23704 13920
rect 23803 13892 23848 13920
rect 23072 13880 23078 13892
rect 21269 13815 21327 13821
rect 21376 13824 22048 13852
rect 22097 13855 22155 13861
rect 21376 13784 21404 13824
rect 22097 13821 22109 13855
rect 22143 13821 22155 13855
rect 22097 13815 22155 13821
rect 19306 13756 21404 13784
rect 21542 13744 21548 13796
rect 21600 13784 21606 13796
rect 22002 13784 22008 13796
rect 21600 13756 22008 13784
rect 21600 13744 21606 13756
rect 22002 13744 22008 13756
rect 22060 13784 22066 13796
rect 22101 13784 22129 13815
rect 22370 13812 22376 13864
rect 22428 13852 22434 13864
rect 22741 13855 22799 13861
rect 22741 13852 22753 13855
rect 22428 13824 22753 13852
rect 22428 13812 22434 13824
rect 22741 13821 22753 13824
rect 22787 13821 22799 13855
rect 23198 13852 23204 13864
rect 23159 13824 23204 13852
rect 22741 13815 22799 13821
rect 23198 13812 23204 13824
rect 23256 13812 23262 13864
rect 23676 13852 23704 13892
rect 23842 13880 23848 13892
rect 23900 13880 23906 13932
rect 23934 13880 23940 13932
rect 23992 13920 23998 13932
rect 24118 13920 24124 13932
rect 23992 13892 24037 13920
rect 24079 13892 24124 13920
rect 23992 13880 23998 13892
rect 24118 13880 24124 13892
rect 24176 13880 24182 13932
rect 24210 13880 24216 13932
rect 24268 13920 24274 13932
rect 24268 13892 24313 13920
rect 24268 13880 24274 13892
rect 24504 13852 24532 13960
rect 24688 13960 25228 13988
rect 24688 13929 24716 13960
rect 25222 13948 25228 13960
rect 25280 13948 25286 14000
rect 25332 13988 25360 14028
rect 25958 14016 25964 14028
rect 26016 14056 26022 14068
rect 27890 14056 27896 14068
rect 26016 14028 27896 14056
rect 26016 14016 26022 14028
rect 27890 14016 27896 14028
rect 27948 14016 27954 14068
rect 28534 14016 28540 14068
rect 28592 14056 28598 14068
rect 29638 14056 29644 14068
rect 28592 14028 29132 14056
rect 29599 14028 29644 14056
rect 28592 14016 28598 14028
rect 25332 13960 25438 13988
rect 27338 13948 27344 14000
rect 27396 13988 27402 14000
rect 27709 13991 27767 13997
rect 27709 13988 27721 13991
rect 27396 13960 27721 13988
rect 27396 13948 27402 13960
rect 27709 13957 27721 13960
rect 27755 13957 27767 13991
rect 27908 13988 27936 14016
rect 27908 13960 28198 13988
rect 27709 13951 27767 13957
rect 24673 13923 24731 13929
rect 24673 13889 24685 13923
rect 24719 13889 24731 13923
rect 24673 13883 24731 13889
rect 26786 13880 26792 13932
rect 26844 13920 26850 13932
rect 27154 13920 27160 13932
rect 26844 13892 27160 13920
rect 26844 13880 26850 13892
rect 27154 13880 27160 13892
rect 27212 13920 27218 13932
rect 27433 13923 27491 13929
rect 27433 13920 27445 13923
rect 27212 13892 27445 13920
rect 27212 13880 27218 13892
rect 27433 13889 27445 13892
rect 27479 13889 27491 13923
rect 29104 13920 29132 14028
rect 29638 14016 29644 14028
rect 29696 14056 29702 14068
rect 36630 14056 36636 14068
rect 29696 14028 36636 14056
rect 29696 14016 29702 14028
rect 36630 14016 36636 14028
rect 36688 14016 36694 14068
rect 36725 14059 36783 14065
rect 36725 14025 36737 14059
rect 36771 14056 36783 14059
rect 36906 14056 36912 14068
rect 36771 14028 36912 14056
rect 36771 14025 36783 14028
rect 36725 14019 36783 14025
rect 36906 14016 36912 14028
rect 36964 14016 36970 14068
rect 39206 14016 39212 14068
rect 39264 14016 39270 14068
rect 39945 14059 40003 14065
rect 39945 14025 39957 14059
rect 39991 14056 40003 14059
rect 40126 14056 40132 14068
rect 39991 14028 40132 14056
rect 39991 14025 40003 14028
rect 39945 14019 40003 14025
rect 40126 14016 40132 14028
rect 40184 14016 40190 14068
rect 42978 14056 42984 14068
rect 42939 14028 42984 14056
rect 42978 14016 42984 14028
rect 43036 14016 43042 14068
rect 44177 14059 44235 14065
rect 44177 14025 44189 14059
rect 44223 14056 44235 14059
rect 44266 14056 44272 14068
rect 44223 14028 44272 14056
rect 44223 14025 44235 14028
rect 44177 14019 44235 14025
rect 44266 14016 44272 14028
rect 44324 14056 44330 14068
rect 44450 14056 44456 14068
rect 44324 14028 44456 14056
rect 44324 14016 44330 14028
rect 44450 14016 44456 14028
rect 44508 14016 44514 14068
rect 45278 14016 45284 14068
rect 45336 14056 45342 14068
rect 46293 14059 46351 14065
rect 46293 14056 46305 14059
rect 45336 14028 46305 14056
rect 45336 14016 45342 14028
rect 46293 14025 46305 14028
rect 46339 14025 46351 14059
rect 46293 14019 46351 14025
rect 29178 13948 29184 14000
rect 29236 13988 29242 14000
rect 29236 13960 29946 13988
rect 29236 13948 29242 13960
rect 31478 13948 31484 14000
rect 31536 13988 31542 14000
rect 32858 13988 32864 14000
rect 31536 13960 32864 13988
rect 31536 13948 31542 13960
rect 32858 13948 32864 13960
rect 32916 13948 32922 14000
rect 34609 13991 34667 13997
rect 34609 13988 34621 13991
rect 34072 13960 34621 13988
rect 31662 13920 31668 13932
rect 29104 13892 29960 13920
rect 27433 13883 27491 13889
rect 29932 13864 29960 13892
rect 31404 13892 31668 13920
rect 26418 13852 26424 13864
rect 23676 13824 24440 13852
rect 24504 13824 26004 13852
rect 26379 13824 26424 13852
rect 22060 13756 22129 13784
rect 22060 13744 22066 13756
rect 22462 13744 22468 13796
rect 22520 13784 22526 13796
rect 23661 13787 23719 13793
rect 23661 13784 23673 13787
rect 22520 13756 23673 13784
rect 22520 13744 22526 13756
rect 23661 13753 23673 13756
rect 23707 13753 23719 13787
rect 24412 13784 24440 13824
rect 24578 13784 24584 13796
rect 24412 13756 24584 13784
rect 23661 13747 23719 13753
rect 24578 13744 24584 13756
rect 24636 13744 24642 13796
rect 25976 13784 26004 13824
rect 26418 13812 26424 13824
rect 26476 13812 26482 13864
rect 29181 13855 29239 13861
rect 29181 13852 29193 13855
rect 26528 13824 29193 13852
rect 26528 13784 26556 13824
rect 29181 13821 29193 13824
rect 29227 13852 29239 13855
rect 29638 13852 29644 13864
rect 29227 13824 29644 13852
rect 29227 13821 29239 13824
rect 29181 13815 29239 13821
rect 29638 13812 29644 13824
rect 29696 13852 29702 13864
rect 29822 13852 29828 13864
rect 29696 13824 29828 13852
rect 29696 13812 29702 13824
rect 29822 13812 29828 13824
rect 29880 13812 29886 13864
rect 29914 13812 29920 13864
rect 29972 13812 29978 13864
rect 30558 13812 30564 13864
rect 30616 13852 30622 13864
rect 31404 13861 31432 13892
rect 31662 13880 31668 13892
rect 31720 13880 31726 13932
rect 31389 13855 31447 13861
rect 31389 13852 31401 13855
rect 30616 13824 31401 13852
rect 30616 13812 30622 13824
rect 31389 13821 31401 13824
rect 31435 13821 31447 13855
rect 31389 13815 31447 13821
rect 31846 13812 31852 13864
rect 31904 13852 31910 13864
rect 32125 13855 32183 13861
rect 32125 13852 32137 13855
rect 31904 13824 32137 13852
rect 31904 13812 31910 13824
rect 32125 13821 32137 13824
rect 32171 13821 32183 13855
rect 32125 13815 32183 13821
rect 33594 13812 33600 13864
rect 33652 13852 33658 13864
rect 33873 13855 33931 13861
rect 33873 13852 33885 13855
rect 33652 13824 33885 13852
rect 33652 13812 33658 13824
rect 33873 13821 33885 13824
rect 33919 13821 33931 13855
rect 33873 13815 33931 13821
rect 25976 13756 26556 13784
rect 1486 13716 1492 13728
rect 1447 13688 1492 13716
rect 1486 13676 1492 13688
rect 1544 13676 1550 13728
rect 17586 13676 17592 13728
rect 17644 13716 17650 13728
rect 20898 13716 20904 13728
rect 17644 13688 20904 13716
rect 17644 13676 17650 13688
rect 20898 13676 20904 13688
rect 20956 13716 20962 13728
rect 21085 13719 21143 13725
rect 21085 13716 21097 13719
rect 20956 13688 21097 13716
rect 20956 13676 20962 13688
rect 21085 13685 21097 13688
rect 21131 13685 21143 13719
rect 21085 13679 21143 13685
rect 21266 13676 21272 13728
rect 21324 13716 21330 13728
rect 22097 13719 22155 13725
rect 22097 13716 22109 13719
rect 21324 13688 22109 13716
rect 21324 13676 21330 13688
rect 22097 13685 22109 13688
rect 22143 13716 22155 13719
rect 22370 13716 22376 13728
rect 22143 13688 22376 13716
rect 22143 13685 22155 13688
rect 22097 13679 22155 13685
rect 22370 13676 22376 13688
rect 22428 13676 22434 13728
rect 22738 13676 22744 13728
rect 22796 13716 22802 13728
rect 24930 13719 24988 13725
rect 24930 13716 24942 13719
rect 22796 13688 24942 13716
rect 22796 13676 22802 13688
rect 24930 13685 24942 13688
rect 24976 13685 24988 13719
rect 24930 13679 24988 13685
rect 26050 13676 26056 13728
rect 26108 13716 26114 13728
rect 30742 13716 30748 13728
rect 26108 13688 30748 13716
rect 26108 13676 26114 13688
rect 30742 13676 30748 13688
rect 30800 13716 30806 13728
rect 30926 13716 30932 13728
rect 30800 13688 30932 13716
rect 30800 13676 30806 13688
rect 30926 13676 30932 13688
rect 30984 13676 30990 13728
rect 31131 13719 31189 13725
rect 31131 13685 31143 13719
rect 31177 13716 31189 13719
rect 31938 13716 31944 13728
rect 31177 13688 31944 13716
rect 31177 13685 31189 13688
rect 31131 13679 31189 13685
rect 31938 13676 31944 13688
rect 31996 13676 32002 13728
rect 32030 13676 32036 13728
rect 32088 13716 32094 13728
rect 32382 13719 32440 13725
rect 32382 13716 32394 13719
rect 32088 13688 32394 13716
rect 32088 13676 32094 13688
rect 32382 13685 32394 13688
rect 32428 13685 32440 13719
rect 32382 13679 32440 13685
rect 32950 13676 32956 13728
rect 33008 13716 33014 13728
rect 34072 13716 34100 13960
rect 34609 13957 34621 13960
rect 34655 13957 34667 13991
rect 34609 13951 34667 13957
rect 35066 13948 35072 14000
rect 35124 13948 35130 14000
rect 38654 13988 38660 14000
rect 36188 13960 38660 13988
rect 34146 13880 34152 13932
rect 34204 13920 34210 13932
rect 34333 13923 34391 13929
rect 34333 13920 34345 13923
rect 34204 13892 34345 13920
rect 34204 13880 34210 13892
rect 34333 13889 34345 13892
rect 34379 13889 34391 13923
rect 34333 13883 34391 13889
rect 34348 13852 34376 13883
rect 35342 13852 35348 13864
rect 34348 13824 35348 13852
rect 35342 13812 35348 13824
rect 35400 13852 35406 13864
rect 36188 13852 36216 13960
rect 38654 13948 38660 13960
rect 38712 13948 38718 14000
rect 36538 13920 36544 13932
rect 36499 13892 36544 13920
rect 36538 13880 36544 13892
rect 36596 13880 36602 13932
rect 37090 13880 37096 13932
rect 37148 13920 37154 13932
rect 37553 13923 37611 13929
rect 37553 13920 37565 13923
rect 37148 13892 37565 13920
rect 37148 13880 37154 13892
rect 37553 13889 37565 13892
rect 37599 13889 37611 13923
rect 37553 13883 37611 13889
rect 37918 13880 37924 13932
rect 37976 13920 37982 13932
rect 38197 13923 38255 13929
rect 38197 13920 38209 13923
rect 37976 13892 38209 13920
rect 37976 13880 37982 13892
rect 38197 13889 38209 13892
rect 38243 13889 38255 13923
rect 39114 13920 39120 13932
rect 38197 13883 38255 13889
rect 38948 13892 39120 13920
rect 35400 13824 36216 13852
rect 35400 13812 35406 13824
rect 36262 13812 36268 13864
rect 36320 13852 36326 13864
rect 36814 13852 36820 13864
rect 36320 13824 36820 13852
rect 36320 13812 36326 13824
rect 36814 13812 36820 13824
rect 36872 13852 36878 13864
rect 38948 13861 38976 13892
rect 39114 13880 39120 13892
rect 39172 13880 39178 13932
rect 39224 13920 39252 14016
rect 41414 13988 41420 14000
rect 39868 13960 41420 13988
rect 39301 13923 39359 13929
rect 39301 13920 39313 13923
rect 39224 13892 39313 13920
rect 39301 13889 39313 13892
rect 39347 13920 39359 13923
rect 39482 13920 39488 13932
rect 39347 13892 39488 13920
rect 39347 13889 39359 13892
rect 39301 13883 39359 13889
rect 39482 13880 39488 13892
rect 39540 13880 39546 13932
rect 37277 13855 37335 13861
rect 37277 13852 37289 13855
rect 36872 13824 37289 13852
rect 36872 13812 36878 13824
rect 37277 13821 37289 13824
rect 37323 13821 37335 13855
rect 37277 13815 37335 13821
rect 38933 13855 38991 13861
rect 38933 13821 38945 13855
rect 38979 13821 38991 13855
rect 39206 13852 39212 13864
rect 39167 13824 39212 13852
rect 38933 13815 38991 13821
rect 39206 13812 39212 13824
rect 39264 13812 39270 13864
rect 39390 13812 39396 13864
rect 39448 13852 39454 13864
rect 39868 13852 39896 13960
rect 41414 13948 41420 13960
rect 41472 13948 41478 14000
rect 41506 13948 41512 14000
rect 41564 13988 41570 14000
rect 41564 13960 41644 13988
rect 41564 13948 41570 13960
rect 40126 13880 40132 13932
rect 40184 13920 40190 13932
rect 40221 13923 40279 13929
rect 40221 13920 40233 13923
rect 40184 13892 40233 13920
rect 40184 13880 40190 13892
rect 40221 13889 40233 13892
rect 40267 13889 40279 13923
rect 40770 13920 40776 13932
rect 40731 13892 40776 13920
rect 40221 13883 40279 13889
rect 40770 13880 40776 13892
rect 40828 13880 40834 13932
rect 40957 13923 41015 13929
rect 40957 13889 40969 13923
rect 41003 13920 41015 13923
rect 41138 13920 41144 13932
rect 41003 13892 41144 13920
rect 41003 13889 41015 13892
rect 40957 13883 41015 13889
rect 41138 13880 41144 13892
rect 41196 13920 41202 13932
rect 41616 13929 41644 13960
rect 42794 13948 42800 14000
rect 42852 13988 42858 14000
rect 45189 13991 45247 13997
rect 45189 13988 45201 13991
rect 42852 13960 45201 13988
rect 42852 13948 42858 13960
rect 45189 13957 45201 13960
rect 45235 13988 45247 13991
rect 45738 13988 45744 14000
rect 45235 13960 45744 13988
rect 45235 13957 45247 13960
rect 45189 13951 45247 13957
rect 45738 13948 45744 13960
rect 45796 13948 45802 14000
rect 45833 13991 45891 13997
rect 45833 13957 45845 13991
rect 45879 13988 45891 13991
rect 46474 13988 46480 14000
rect 45879 13960 46480 13988
rect 45879 13957 45891 13960
rect 45833 13951 45891 13957
rect 46474 13948 46480 13960
rect 46532 13948 46538 14000
rect 41601 13923 41659 13929
rect 41196 13892 41414 13920
rect 41196 13880 41202 13892
rect 39448 13824 39896 13852
rect 39945 13855 40003 13861
rect 39448 13812 39454 13824
rect 39945 13821 39957 13855
rect 39991 13852 40003 13855
rect 39991 13824 41322 13852
rect 39991 13821 40003 13824
rect 39945 13815 40003 13821
rect 35986 13744 35992 13796
rect 36044 13784 36050 13796
rect 36081 13787 36139 13793
rect 36081 13784 36093 13787
rect 36044 13756 36093 13784
rect 36044 13744 36050 13756
rect 36081 13753 36093 13756
rect 36127 13753 36139 13787
rect 36081 13747 36139 13753
rect 36446 13744 36452 13796
rect 36504 13784 36510 13796
rect 36722 13784 36728 13796
rect 36504 13756 36728 13784
rect 36504 13744 36510 13756
rect 36722 13744 36728 13756
rect 36780 13744 36786 13796
rect 40218 13744 40224 13796
rect 40276 13784 40282 13796
rect 40770 13784 40776 13796
rect 40276 13756 40776 13784
rect 40276 13744 40282 13756
rect 40770 13744 40776 13756
rect 40828 13744 40834 13796
rect 33008 13688 34100 13716
rect 33008 13676 33014 13688
rect 37642 13676 37648 13728
rect 37700 13716 37706 13728
rect 38102 13716 38108 13728
rect 37700 13688 38108 13716
rect 37700 13676 37706 13688
rect 38102 13676 38108 13688
rect 38160 13716 38166 13728
rect 38381 13719 38439 13725
rect 38381 13716 38393 13719
rect 38160 13688 38393 13716
rect 38160 13676 38166 13688
rect 38381 13685 38393 13688
rect 38427 13685 38439 13719
rect 38381 13679 38439 13685
rect 39206 13676 39212 13728
rect 39264 13716 39270 13728
rect 39574 13716 39580 13728
rect 39264 13688 39580 13716
rect 39264 13676 39270 13688
rect 39574 13676 39580 13688
rect 39632 13676 39638 13728
rect 40126 13676 40132 13728
rect 40184 13716 40190 13728
rect 41294 13716 41322 13824
rect 41386 13784 41414 13892
rect 41601 13889 41613 13923
rect 41647 13920 41659 13923
rect 42702 13920 42708 13932
rect 41647 13892 42708 13920
rect 41647 13889 41659 13892
rect 41601 13883 41659 13889
rect 42702 13880 42708 13892
rect 42760 13880 42766 13932
rect 43625 13923 43683 13929
rect 43625 13889 43637 13923
rect 43671 13920 43683 13923
rect 44174 13920 44180 13932
rect 43671 13892 44180 13920
rect 43671 13889 43683 13892
rect 43625 13883 43683 13889
rect 44174 13880 44180 13892
rect 44232 13880 44238 13932
rect 41506 13852 41512 13864
rect 41467 13824 41512 13852
rect 41506 13812 41512 13824
rect 41564 13812 41570 13864
rect 41690 13812 41696 13864
rect 41748 13852 41754 13864
rect 43530 13852 43536 13864
rect 41748 13824 43536 13852
rect 41748 13812 41754 13824
rect 43530 13812 43536 13824
rect 43588 13812 43594 13864
rect 43806 13812 43812 13864
rect 43864 13852 43870 13864
rect 44637 13855 44695 13861
rect 44637 13852 44649 13855
rect 43864 13824 44649 13852
rect 43864 13812 43870 13824
rect 44637 13821 44649 13824
rect 44683 13821 44695 13855
rect 44637 13815 44695 13821
rect 45002 13784 45008 13796
rect 41386 13756 45008 13784
rect 45002 13744 45008 13756
rect 45060 13744 45066 13796
rect 41690 13716 41696 13728
rect 40184 13688 40229 13716
rect 41294 13688 41696 13716
rect 40184 13676 40190 13688
rect 41690 13676 41696 13688
rect 41748 13676 41754 13728
rect 41966 13676 41972 13728
rect 42024 13716 42030 13728
rect 42518 13716 42524 13728
rect 42024 13688 42524 13716
rect 42024 13676 42030 13688
rect 42518 13676 42524 13688
rect 42576 13676 42582 13728
rect 45554 13676 45560 13728
rect 45612 13716 45618 13728
rect 46845 13719 46903 13725
rect 46845 13716 46857 13719
rect 45612 13688 46857 13716
rect 45612 13676 45618 13688
rect 46845 13685 46857 13688
rect 46891 13685 46903 13719
rect 46845 13679 46903 13685
rect 1104 13626 58880 13648
rect 1104 13574 10582 13626
rect 10634 13574 10646 13626
rect 10698 13574 10710 13626
rect 10762 13574 10774 13626
rect 10826 13574 10838 13626
rect 10890 13574 29846 13626
rect 29898 13574 29910 13626
rect 29962 13574 29974 13626
rect 30026 13574 30038 13626
rect 30090 13574 30102 13626
rect 30154 13574 49110 13626
rect 49162 13574 49174 13626
rect 49226 13574 49238 13626
rect 49290 13574 49302 13626
rect 49354 13574 49366 13626
rect 49418 13574 58880 13626
rect 1104 13552 58880 13574
rect 12069 13515 12127 13521
rect 12069 13481 12081 13515
rect 12115 13512 12127 13515
rect 14182 13512 14188 13524
rect 12115 13484 14188 13512
rect 12115 13481 12127 13484
rect 12069 13475 12127 13481
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13308 11575 13311
rect 12084 13308 12112 13475
rect 14182 13472 14188 13484
rect 14240 13472 14246 13524
rect 16669 13515 16727 13521
rect 16669 13481 16681 13515
rect 16715 13512 16727 13515
rect 16758 13512 16764 13524
rect 16715 13484 16764 13512
rect 16715 13481 16727 13484
rect 16669 13475 16727 13481
rect 16758 13472 16764 13484
rect 16816 13512 16822 13524
rect 19334 13512 19340 13524
rect 16816 13484 19340 13512
rect 16816 13472 16822 13484
rect 19334 13472 19340 13484
rect 19392 13472 19398 13524
rect 19613 13515 19671 13521
rect 19613 13481 19625 13515
rect 19659 13512 19671 13515
rect 20070 13512 20076 13524
rect 19659 13484 20076 13512
rect 19659 13481 19671 13484
rect 19613 13475 19671 13481
rect 20070 13472 20076 13484
rect 20128 13472 20134 13524
rect 21269 13515 21327 13521
rect 21269 13481 21281 13515
rect 21315 13512 21327 13515
rect 22002 13512 22008 13524
rect 21315 13484 22008 13512
rect 21315 13481 21327 13484
rect 21269 13475 21327 13481
rect 22002 13472 22008 13484
rect 22060 13472 22066 13524
rect 22186 13472 22192 13524
rect 22244 13512 22250 13524
rect 24765 13515 24823 13521
rect 24765 13512 24777 13515
rect 22244 13484 24777 13512
rect 22244 13472 22250 13484
rect 24765 13481 24777 13484
rect 24811 13481 24823 13515
rect 24765 13475 24823 13481
rect 25590 13472 25596 13524
rect 25648 13512 25654 13524
rect 27338 13512 27344 13524
rect 25648 13484 27344 13512
rect 25648 13472 25654 13484
rect 27338 13472 27344 13484
rect 27396 13472 27402 13524
rect 28074 13512 28080 13524
rect 27586 13484 28080 13512
rect 12158 13404 12164 13456
rect 12216 13444 12222 13456
rect 16025 13447 16083 13453
rect 16025 13444 16037 13447
rect 12216 13416 16037 13444
rect 12216 13404 12222 13416
rect 16025 13413 16037 13416
rect 16071 13413 16083 13447
rect 17126 13444 17132 13456
rect 17087 13416 17132 13444
rect 16025 13407 16083 13413
rect 17126 13404 17132 13416
rect 17184 13404 17190 13456
rect 17773 13447 17831 13453
rect 17773 13413 17785 13447
rect 17819 13444 17831 13447
rect 21726 13444 21732 13456
rect 17819 13416 21732 13444
rect 17819 13413 17831 13416
rect 17773 13407 17831 13413
rect 21726 13404 21732 13416
rect 21784 13404 21790 13456
rect 24670 13404 24676 13456
rect 24728 13444 24734 13456
rect 27249 13447 27307 13453
rect 27249 13444 27261 13447
rect 24728 13416 27261 13444
rect 24728 13404 24734 13416
rect 27249 13413 27261 13416
rect 27295 13413 27307 13447
rect 27586 13444 27614 13484
rect 28074 13472 28080 13484
rect 28132 13512 28138 13524
rect 28350 13512 28356 13524
rect 28132 13484 28356 13512
rect 28132 13472 28138 13484
rect 28350 13472 28356 13484
rect 28408 13472 28414 13524
rect 30190 13472 30196 13524
rect 30248 13512 30254 13524
rect 31202 13512 31208 13524
rect 30248 13484 31208 13512
rect 30248 13472 30254 13484
rect 31202 13472 31208 13484
rect 31260 13472 31266 13524
rect 32030 13512 32036 13524
rect 31726 13484 32036 13512
rect 27249 13407 27307 13413
rect 27448 13416 27614 13444
rect 19150 13336 19156 13388
rect 19208 13376 19214 13388
rect 19208 13348 21956 13376
rect 19208 13336 19214 13348
rect 11563 13280 12112 13308
rect 11563 13277 11575 13280
rect 11517 13271 11575 13277
rect 18046 13268 18052 13320
rect 18104 13308 18110 13320
rect 20165 13311 20223 13317
rect 20165 13308 20177 13311
rect 18104 13280 20177 13308
rect 18104 13268 18110 13280
rect 18340 13252 18368 13280
rect 20165 13277 20177 13280
rect 20211 13308 20223 13311
rect 20806 13308 20812 13320
rect 20211 13280 20812 13308
rect 20211 13277 20223 13280
rect 20165 13271 20223 13277
rect 20806 13268 20812 13280
rect 20864 13268 20870 13320
rect 21358 13308 21364 13320
rect 21319 13280 21364 13308
rect 21358 13268 21364 13280
rect 21416 13268 21422 13320
rect 21928 13308 21956 13348
rect 22002 13336 22008 13388
rect 22060 13376 22066 13388
rect 23566 13376 23572 13388
rect 22060 13348 23572 13376
rect 22060 13336 22066 13348
rect 23566 13336 23572 13348
rect 23624 13336 23630 13388
rect 25409 13379 25467 13385
rect 25409 13345 25421 13379
rect 25455 13376 25467 13379
rect 25774 13376 25780 13388
rect 25455 13348 25780 13376
rect 25455 13345 25467 13348
rect 25409 13339 25467 13345
rect 25774 13336 25780 13348
rect 25832 13336 25838 13388
rect 26237 13379 26295 13385
rect 26237 13345 26249 13379
rect 26283 13376 26295 13379
rect 27448 13376 27476 13416
rect 29270 13404 29276 13456
rect 29328 13444 29334 13456
rect 29546 13444 29552 13456
rect 29328 13416 29552 13444
rect 29328 13404 29334 13416
rect 29546 13404 29552 13416
rect 29604 13404 29610 13456
rect 31110 13404 31116 13456
rect 31168 13444 31174 13456
rect 31726 13444 31754 13484
rect 32030 13472 32036 13484
rect 32088 13472 32094 13524
rect 33502 13512 33508 13524
rect 32140 13484 33508 13512
rect 31168 13416 31754 13444
rect 31168 13404 31174 13416
rect 26283 13348 27476 13376
rect 26283 13345 26295 13348
rect 26237 13339 26295 13345
rect 28258 13336 28264 13388
rect 28316 13376 28322 13388
rect 30101 13379 30159 13385
rect 30101 13376 30113 13379
rect 28316 13348 30113 13376
rect 28316 13336 28322 13348
rect 30101 13345 30113 13348
rect 30147 13345 30159 13379
rect 32140 13376 32168 13484
rect 33502 13472 33508 13484
rect 33560 13472 33566 13524
rect 33778 13512 33784 13524
rect 33739 13484 33784 13512
rect 33778 13472 33784 13484
rect 33836 13472 33842 13524
rect 40589 13515 40647 13521
rect 40589 13512 40601 13515
rect 34716 13484 40601 13512
rect 30101 13339 30159 13345
rect 31726 13348 32168 13376
rect 32309 13379 32367 13385
rect 22186 13308 22192 13320
rect 21928 13280 22192 13308
rect 22186 13268 22192 13280
rect 22244 13268 22250 13320
rect 23842 13268 23848 13320
rect 23900 13308 23906 13320
rect 23900 13280 23945 13308
rect 23900 13268 23906 13280
rect 24762 13268 24768 13320
rect 24820 13308 24826 13320
rect 25961 13311 26019 13317
rect 25961 13308 25973 13311
rect 24820 13280 25973 13308
rect 24820 13268 24826 13280
rect 25961 13277 25973 13280
rect 26007 13277 26019 13311
rect 25961 13271 26019 13277
rect 18322 13200 18328 13252
rect 18380 13200 18386 13252
rect 19610 13200 19616 13252
rect 19668 13240 19674 13252
rect 20625 13243 20683 13249
rect 20625 13240 20637 13243
rect 19668 13212 20637 13240
rect 19668 13200 19674 13212
rect 20625 13209 20637 13212
rect 20671 13209 20683 13243
rect 20625 13203 20683 13209
rect 11330 13172 11336 13184
rect 11291 13144 11336 13172
rect 11330 13132 11336 13144
rect 11388 13132 11394 13184
rect 18233 13175 18291 13181
rect 18233 13141 18245 13175
rect 18279 13172 18291 13175
rect 18414 13172 18420 13184
rect 18279 13144 18420 13172
rect 18279 13141 18291 13144
rect 18233 13135 18291 13141
rect 18414 13132 18420 13144
rect 18472 13132 18478 13184
rect 20640 13172 20668 13203
rect 20990 13200 20996 13252
rect 21048 13240 21054 13252
rect 21821 13243 21879 13249
rect 21821 13240 21833 13243
rect 21048 13212 21833 13240
rect 21048 13200 21054 13212
rect 21821 13209 21833 13212
rect 21867 13209 21879 13243
rect 21821 13203 21879 13209
rect 23014 13200 23020 13252
rect 23072 13200 23078 13252
rect 24946 13200 24952 13252
rect 25004 13240 25010 13252
rect 25225 13243 25283 13249
rect 25225 13240 25237 13243
rect 25004 13212 25237 13240
rect 25004 13200 25010 13212
rect 25225 13209 25237 13212
rect 25271 13209 25283 13243
rect 25976 13240 26004 13271
rect 26142 13268 26148 13320
rect 26200 13308 26206 13320
rect 26970 13308 26976 13320
rect 26200 13280 26976 13308
rect 26200 13268 26206 13280
rect 26970 13268 26976 13280
rect 27028 13268 27034 13320
rect 28994 13268 29000 13320
rect 29052 13308 29058 13320
rect 29822 13308 29828 13320
rect 29052 13280 29097 13308
rect 29783 13280 29828 13308
rect 29052 13268 29058 13280
rect 29822 13268 29828 13280
rect 29880 13268 29886 13320
rect 31202 13268 31208 13320
rect 31260 13268 31266 13320
rect 26234 13240 26240 13252
rect 25976 13212 26240 13240
rect 25225 13203 25283 13209
rect 26234 13200 26240 13212
rect 26292 13200 26298 13252
rect 28166 13200 28172 13252
rect 28224 13200 28230 13252
rect 28718 13240 28724 13252
rect 28679 13212 28724 13240
rect 28718 13200 28724 13212
rect 28776 13200 28782 13252
rect 31726 13240 31754 13348
rect 32309 13345 32321 13379
rect 32355 13376 32367 13379
rect 34716 13376 34744 13484
rect 40589 13481 40601 13484
rect 40635 13481 40647 13515
rect 41230 13512 41236 13524
rect 41191 13484 41236 13512
rect 40589 13475 40647 13481
rect 41230 13472 41236 13484
rect 41288 13472 41294 13524
rect 42610 13472 42616 13524
rect 42668 13512 42674 13524
rect 42797 13515 42855 13521
rect 42797 13512 42809 13515
rect 42668 13484 42809 13512
rect 42668 13472 42674 13484
rect 42797 13481 42809 13484
rect 42843 13481 42855 13515
rect 42797 13475 42855 13481
rect 43530 13472 43536 13524
rect 43588 13512 43594 13524
rect 43901 13515 43959 13521
rect 43901 13512 43913 13515
rect 43588 13484 43913 13512
rect 43588 13472 43594 13484
rect 43901 13481 43913 13484
rect 43947 13481 43959 13515
rect 43901 13475 43959 13481
rect 38010 13444 38016 13456
rect 37971 13416 38016 13444
rect 38010 13404 38016 13416
rect 38068 13404 38074 13456
rect 38470 13404 38476 13456
rect 38528 13444 38534 13456
rect 39945 13447 40003 13453
rect 39945 13444 39957 13447
rect 38528 13416 39957 13444
rect 38528 13404 38534 13416
rect 39945 13413 39957 13416
rect 39991 13444 40003 13447
rect 43916 13444 43944 13475
rect 46106 13472 46112 13524
rect 46164 13512 46170 13524
rect 46201 13515 46259 13521
rect 46201 13512 46213 13515
rect 46164 13484 46213 13512
rect 46164 13472 46170 13484
rect 46201 13481 46213 13484
rect 46247 13512 46259 13515
rect 46474 13512 46480 13524
rect 46247 13484 46480 13512
rect 46247 13481 46259 13484
rect 46201 13475 46259 13481
rect 46474 13472 46480 13484
rect 46532 13472 46538 13524
rect 45554 13444 45560 13456
rect 39991 13416 41414 13444
rect 43916 13416 45560 13444
rect 39991 13413 40003 13416
rect 39945 13407 40003 13413
rect 36262 13376 36268 13388
rect 32355 13348 34744 13376
rect 35360 13348 36268 13376
rect 32355 13345 32367 13348
rect 32309 13339 32367 13345
rect 31846 13268 31852 13320
rect 31904 13308 31910 13320
rect 32033 13311 32091 13317
rect 32033 13308 32045 13311
rect 31904 13280 32045 13308
rect 31904 13268 31910 13280
rect 32033 13277 32045 13280
rect 32079 13277 32091 13311
rect 32033 13271 32091 13277
rect 34054 13268 34060 13320
rect 34112 13308 34118 13320
rect 34701 13311 34759 13317
rect 34701 13308 34713 13311
rect 34112 13280 34713 13308
rect 34112 13268 34118 13280
rect 34701 13277 34713 13280
rect 34747 13277 34759 13311
rect 34701 13271 34759 13277
rect 34977 13311 35035 13317
rect 34977 13277 34989 13311
rect 35023 13308 35035 13311
rect 35158 13308 35164 13320
rect 35023 13280 35164 13308
rect 35023 13277 35035 13280
rect 34977 13271 35035 13277
rect 34238 13240 34244 13252
rect 31404 13212 31754 13240
rect 33534 13212 34244 13240
rect 21266 13172 21272 13184
rect 20640 13144 21272 13172
rect 21266 13132 21272 13144
rect 21324 13132 21330 13184
rect 21910 13132 21916 13184
rect 21968 13172 21974 13184
rect 24118 13172 24124 13184
rect 21968 13144 24124 13172
rect 21968 13132 21974 13144
rect 24118 13132 24124 13144
rect 24176 13132 24182 13184
rect 25130 13172 25136 13184
rect 25091 13144 25136 13172
rect 25130 13132 25136 13144
rect 25188 13132 25194 13184
rect 25958 13132 25964 13184
rect 26016 13172 26022 13184
rect 31404 13172 31432 13212
rect 34238 13200 34244 13212
rect 34296 13200 34302 13252
rect 34716 13240 34744 13271
rect 35158 13268 35164 13280
rect 35216 13268 35222 13320
rect 35360 13240 35388 13348
rect 36262 13336 36268 13348
rect 36320 13376 36326 13388
rect 36357 13379 36415 13385
rect 36357 13376 36369 13379
rect 36320 13348 36369 13376
rect 36320 13336 36326 13348
rect 36357 13345 36369 13348
rect 36403 13345 36415 13379
rect 38102 13376 38108 13388
rect 36357 13339 36415 13345
rect 37108 13348 38108 13376
rect 37108 13320 37136 13348
rect 38102 13336 38108 13348
rect 38160 13336 38166 13388
rect 38286 13376 38292 13388
rect 38247 13348 38292 13376
rect 38286 13336 38292 13348
rect 38344 13336 38350 13388
rect 38654 13336 38660 13388
rect 38712 13376 38718 13388
rect 41386 13376 41414 13416
rect 45554 13404 45560 13416
rect 45612 13404 45618 13456
rect 42794 13376 42800 13388
rect 38712 13348 40724 13376
rect 41386 13348 42800 13376
rect 38712 13336 38718 13348
rect 35621 13311 35679 13317
rect 35621 13277 35633 13311
rect 35667 13308 35679 13311
rect 35710 13308 35716 13320
rect 35667 13280 35716 13308
rect 35667 13277 35679 13280
rect 35621 13271 35679 13277
rect 35710 13268 35716 13280
rect 35768 13268 35774 13320
rect 35802 13268 35808 13320
rect 35860 13308 35866 13320
rect 36633 13311 36691 13317
rect 36633 13308 36645 13311
rect 35860 13280 36645 13308
rect 35860 13268 35866 13280
rect 36633 13277 36645 13280
rect 36679 13308 36691 13311
rect 37090 13308 37096 13320
rect 36679 13280 37096 13308
rect 36679 13277 36691 13280
rect 36633 13271 36691 13277
rect 37090 13268 37096 13280
rect 37148 13268 37154 13320
rect 37277 13311 37335 13317
rect 37277 13277 37289 13311
rect 37323 13308 37335 13311
rect 37366 13308 37372 13320
rect 37323 13280 37372 13308
rect 37323 13277 37335 13280
rect 37277 13271 37335 13277
rect 37366 13268 37372 13280
rect 37424 13268 37430 13320
rect 37918 13268 37924 13320
rect 37976 13308 37982 13320
rect 38378 13308 38384 13320
rect 37976 13280 38384 13308
rect 37976 13268 37982 13280
rect 38378 13268 38384 13280
rect 38436 13268 38442 13320
rect 40034 13308 40040 13320
rect 39995 13280 40040 13308
rect 40034 13268 40040 13280
rect 40092 13268 40098 13320
rect 40696 13317 40724 13348
rect 42794 13336 42800 13348
rect 42852 13336 42858 13388
rect 45097 13379 45155 13385
rect 45097 13345 45109 13379
rect 45143 13376 45155 13379
rect 46198 13376 46204 13388
rect 45143 13348 46204 13376
rect 45143 13345 45155 13348
rect 45097 13339 45155 13345
rect 46198 13336 46204 13348
rect 46256 13336 46262 13388
rect 40681 13311 40739 13317
rect 40681 13277 40693 13311
rect 40727 13308 40739 13311
rect 41598 13308 41604 13320
rect 40727 13280 41604 13308
rect 40727 13277 40739 13280
rect 40681 13271 40739 13277
rect 41598 13268 41604 13280
rect 41656 13268 41662 13320
rect 43346 13308 43352 13320
rect 43307 13280 43352 13308
rect 43346 13268 43352 13280
rect 43404 13268 43410 13320
rect 58158 13308 58164 13320
rect 58119 13280 58164 13308
rect 58158 13268 58164 13280
rect 58216 13268 58222 13320
rect 34716 13212 35388 13240
rect 35434 13200 35440 13252
rect 35492 13240 35498 13252
rect 35897 13243 35955 13249
rect 35897 13240 35909 13243
rect 35492 13212 35909 13240
rect 35492 13200 35498 13212
rect 35897 13209 35909 13212
rect 35943 13240 35955 13243
rect 37553 13243 37611 13249
rect 37553 13240 37565 13243
rect 35943 13212 37565 13240
rect 35943 13209 35955 13212
rect 35897 13203 35955 13209
rect 37553 13209 37565 13212
rect 37599 13240 37611 13243
rect 37642 13240 37648 13252
rect 37599 13212 37648 13240
rect 37599 13209 37611 13212
rect 37553 13203 37611 13209
rect 37642 13200 37648 13212
rect 37700 13200 37706 13252
rect 38838 13200 38844 13252
rect 38896 13240 38902 13252
rect 39209 13243 39267 13249
rect 39209 13240 39221 13243
rect 38896 13212 39221 13240
rect 38896 13200 38902 13212
rect 39209 13209 39221 13212
rect 39255 13209 39267 13243
rect 39209 13203 39267 13209
rect 26016 13144 31432 13172
rect 31573 13175 31631 13181
rect 26016 13132 26022 13144
rect 31573 13141 31585 13175
rect 31619 13172 31631 13175
rect 38930 13172 38936 13184
rect 31619 13144 38936 13172
rect 31619 13141 31631 13144
rect 31573 13135 31631 13141
rect 38930 13132 38936 13144
rect 38988 13132 38994 13184
rect 39114 13172 39120 13184
rect 39075 13144 39120 13172
rect 39114 13132 39120 13144
rect 39172 13132 39178 13184
rect 39224 13172 39252 13203
rect 39482 13200 39488 13252
rect 39540 13240 39546 13252
rect 41230 13240 41236 13252
rect 39540 13212 41236 13240
rect 39540 13200 39546 13212
rect 41230 13200 41236 13212
rect 41288 13200 41294 13252
rect 41322 13200 41328 13252
rect 41380 13240 41386 13252
rect 41693 13243 41751 13249
rect 41693 13240 41705 13243
rect 41380 13212 41705 13240
rect 41380 13200 41386 13212
rect 41693 13209 41705 13212
rect 41739 13209 41751 13243
rect 57882 13240 57888 13252
rect 57843 13212 57888 13240
rect 41693 13203 41751 13209
rect 57882 13200 57888 13212
rect 57940 13200 57946 13252
rect 40218 13172 40224 13184
rect 39224 13144 40224 13172
rect 40218 13132 40224 13144
rect 40276 13172 40282 13184
rect 41414 13172 41420 13184
rect 40276 13144 41420 13172
rect 40276 13132 40282 13144
rect 41414 13132 41420 13144
rect 41472 13132 41478 13184
rect 41598 13132 41604 13184
rect 41656 13172 41662 13184
rect 42245 13175 42303 13181
rect 42245 13172 42257 13175
rect 41656 13144 42257 13172
rect 41656 13132 41662 13144
rect 42245 13141 42257 13144
rect 42291 13172 42303 13175
rect 42886 13172 42892 13184
rect 42291 13144 42892 13172
rect 42291 13141 42303 13144
rect 42245 13135 42303 13141
rect 42886 13132 42892 13144
rect 42944 13132 42950 13184
rect 1104 13082 58880 13104
rect 1104 13030 20214 13082
rect 20266 13030 20278 13082
rect 20330 13030 20342 13082
rect 20394 13030 20406 13082
rect 20458 13030 20470 13082
rect 20522 13030 39478 13082
rect 39530 13030 39542 13082
rect 39594 13030 39606 13082
rect 39658 13030 39670 13082
rect 39722 13030 39734 13082
rect 39786 13030 58880 13082
rect 1104 13008 58880 13030
rect 18506 12968 18512 12980
rect 18467 12940 18512 12968
rect 18506 12928 18512 12940
rect 18564 12928 18570 12980
rect 20070 12968 20076 12980
rect 20031 12940 20076 12968
rect 20070 12928 20076 12940
rect 20128 12928 20134 12980
rect 21269 12971 21327 12977
rect 21269 12937 21281 12971
rect 21315 12968 21327 12971
rect 21910 12968 21916 12980
rect 21315 12940 21916 12968
rect 21315 12937 21327 12940
rect 21269 12931 21327 12937
rect 21910 12928 21916 12940
rect 21968 12928 21974 12980
rect 22373 12971 22431 12977
rect 22373 12937 22385 12971
rect 22419 12968 22431 12971
rect 22646 12968 22652 12980
rect 22419 12940 22652 12968
rect 22419 12937 22431 12940
rect 22373 12931 22431 12937
rect 22646 12928 22652 12940
rect 22704 12928 22710 12980
rect 24578 12968 24584 12980
rect 23032 12940 24584 12968
rect 17954 12900 17960 12912
rect 17867 12872 17960 12900
rect 17954 12860 17960 12872
rect 18012 12900 18018 12912
rect 19242 12900 19248 12912
rect 18012 12872 19248 12900
rect 18012 12860 18018 12872
rect 19242 12860 19248 12872
rect 19300 12860 19306 12912
rect 19613 12903 19671 12909
rect 19613 12869 19625 12903
rect 19659 12900 19671 12903
rect 19702 12900 19708 12912
rect 19659 12872 19708 12900
rect 19659 12869 19671 12872
rect 19613 12863 19671 12869
rect 18414 12792 18420 12844
rect 18472 12832 18478 12844
rect 19628 12832 19656 12863
rect 19702 12860 19708 12872
rect 19760 12900 19766 12912
rect 21818 12900 21824 12912
rect 19760 12872 21824 12900
rect 19760 12860 19766 12872
rect 21818 12860 21824 12872
rect 21876 12860 21882 12912
rect 22186 12860 22192 12912
rect 22244 12900 22250 12912
rect 23032 12900 23060 12940
rect 24578 12928 24584 12940
rect 24636 12928 24642 12980
rect 24762 12928 24768 12980
rect 24820 12968 24826 12980
rect 26418 12968 26424 12980
rect 24820 12940 26004 12968
rect 26379 12940 26424 12968
rect 24820 12928 24826 12940
rect 22244 12872 23060 12900
rect 22244 12860 22250 12872
rect 20714 12832 20720 12844
rect 18472 12804 19656 12832
rect 20627 12804 20720 12832
rect 18472 12792 18478 12804
rect 20714 12792 20720 12804
rect 20772 12832 20778 12844
rect 22204 12832 22232 12860
rect 20772 12804 22232 12832
rect 20772 12792 20778 12804
rect 22278 12792 22284 12844
rect 22336 12832 22342 12844
rect 22465 12835 22523 12841
rect 22465 12832 22477 12835
rect 22336 12804 22477 12832
rect 22336 12792 22342 12804
rect 22465 12801 22477 12804
rect 22511 12801 22523 12835
rect 22465 12795 22523 12801
rect 22830 12792 22836 12844
rect 22888 12832 22894 12844
rect 22925 12835 22983 12841
rect 22925 12832 22937 12835
rect 22888 12804 22937 12832
rect 22888 12792 22894 12804
rect 22925 12801 22937 12804
rect 22971 12801 22983 12835
rect 23032 12832 23060 12872
rect 23109 12903 23167 12909
rect 23109 12869 23121 12903
rect 23155 12900 23167 12903
rect 23155 12872 24992 12900
rect 23155 12869 23167 12872
rect 23109 12863 23167 12869
rect 23201 12835 23259 12841
rect 23201 12832 23213 12835
rect 23032 12804 23213 12832
rect 22925 12795 22983 12801
rect 23201 12801 23213 12804
rect 23247 12801 23259 12835
rect 23201 12795 23259 12801
rect 23474 12792 23480 12844
rect 23532 12832 23538 12844
rect 23845 12835 23903 12841
rect 23845 12832 23857 12835
rect 23532 12804 23857 12832
rect 23532 12792 23538 12804
rect 23845 12801 23857 12804
rect 23891 12832 23903 12835
rect 24118 12832 24124 12844
rect 23891 12804 24124 12832
rect 23891 12801 23903 12804
rect 23845 12795 23903 12801
rect 24118 12792 24124 12804
rect 24176 12792 24182 12844
rect 24964 12776 24992 12872
rect 25041 12835 25099 12841
rect 25041 12801 25053 12835
rect 25087 12801 25099 12835
rect 25041 12795 25099 12801
rect 15470 12724 15476 12776
rect 15528 12764 15534 12776
rect 18969 12767 19027 12773
rect 18969 12764 18981 12767
rect 15528 12736 18981 12764
rect 15528 12724 15534 12736
rect 18969 12733 18981 12736
rect 19015 12764 19027 12767
rect 23382 12764 23388 12776
rect 19015 12736 23388 12764
rect 19015 12733 19027 12736
rect 18969 12727 19027 12733
rect 23382 12724 23388 12736
rect 23440 12724 23446 12776
rect 23750 12764 23756 12776
rect 23711 12736 23756 12764
rect 23750 12724 23756 12736
rect 23808 12724 23814 12776
rect 24946 12764 24952 12776
rect 24907 12736 24952 12764
rect 24946 12724 24952 12736
rect 25004 12724 25010 12776
rect 21634 12656 21640 12708
rect 21692 12696 21698 12708
rect 24673 12699 24731 12705
rect 24673 12696 24685 12699
rect 21692 12668 24685 12696
rect 21692 12656 21698 12668
rect 24673 12665 24685 12668
rect 24719 12665 24731 12699
rect 25056 12696 25084 12795
rect 24673 12659 24731 12665
rect 24780 12668 25084 12696
rect 25148 12696 25176 12940
rect 25406 12860 25412 12912
rect 25464 12900 25470 12912
rect 25464 12872 25912 12900
rect 25464 12860 25470 12872
rect 25222 12792 25228 12844
rect 25280 12832 25286 12844
rect 25884 12841 25912 12872
rect 25685 12835 25743 12841
rect 25685 12832 25697 12835
rect 25280 12804 25697 12832
rect 25280 12792 25286 12804
rect 25685 12801 25697 12804
rect 25731 12801 25743 12835
rect 25685 12795 25743 12801
rect 25869 12835 25927 12841
rect 25869 12801 25881 12835
rect 25915 12801 25927 12835
rect 25976 12832 26004 12940
rect 26418 12928 26424 12940
rect 26476 12928 26482 12980
rect 26970 12928 26976 12980
rect 27028 12928 27034 12980
rect 27338 12928 27344 12980
rect 27396 12968 27402 12980
rect 27798 12968 27804 12980
rect 27396 12940 27804 12968
rect 27396 12928 27402 12940
rect 27798 12928 27804 12940
rect 27856 12928 27862 12980
rect 29086 12968 29092 12980
rect 28000 12940 28994 12968
rect 29047 12940 29092 12968
rect 26988 12900 27016 12928
rect 28000 12900 28028 12940
rect 28966 12900 28994 12940
rect 29086 12928 29092 12940
rect 29144 12928 29150 12980
rect 31110 12968 31116 12980
rect 29656 12940 31116 12968
rect 29656 12900 29684 12940
rect 31110 12928 31116 12940
rect 31168 12928 31174 12980
rect 31294 12968 31300 12980
rect 31255 12940 31300 12968
rect 31294 12928 31300 12940
rect 31352 12928 31358 12980
rect 36170 12968 36176 12980
rect 31726 12940 36176 12968
rect 31726 12900 31754 12940
rect 36170 12928 36176 12940
rect 36228 12928 36234 12980
rect 36906 12968 36912 12980
rect 36556 12940 36912 12968
rect 32398 12900 32404 12912
rect 26988 12872 28106 12900
rect 28966 12872 29684 12900
rect 31050 12872 31754 12900
rect 32359 12872 32404 12900
rect 32398 12860 32404 12872
rect 32456 12860 32462 12912
rect 34422 12900 34428 12912
rect 33626 12872 34428 12900
rect 34422 12860 34428 12872
rect 34480 12860 34486 12912
rect 26170 12835 26228 12841
rect 26170 12832 26182 12835
rect 25976 12804 26182 12832
rect 25869 12795 25927 12801
rect 26170 12801 26182 12804
rect 26216 12801 26228 12835
rect 26170 12795 26228 12801
rect 25884 12764 25912 12795
rect 31202 12792 31208 12844
rect 31260 12832 31266 12844
rect 31662 12832 31668 12844
rect 31260 12804 31668 12832
rect 31260 12792 31266 12804
rect 31662 12792 31668 12804
rect 31720 12792 31726 12844
rect 34146 12832 34152 12844
rect 33888 12804 34152 12832
rect 27338 12764 27344 12776
rect 25884 12736 26188 12764
rect 27299 12736 27344 12764
rect 25406 12696 25412 12708
rect 25148 12668 25412 12696
rect 12986 12588 12992 12640
rect 13044 12628 13050 12640
rect 16853 12631 16911 12637
rect 16853 12628 16865 12631
rect 13044 12600 16865 12628
rect 13044 12588 13050 12600
rect 16853 12597 16865 12600
rect 16899 12628 16911 12631
rect 17405 12631 17463 12637
rect 17405 12628 17417 12631
rect 16899 12600 17417 12628
rect 16899 12597 16911 12600
rect 16853 12591 16911 12597
rect 17405 12597 17417 12600
rect 17451 12628 17463 12631
rect 20070 12628 20076 12640
rect 17451 12600 20076 12628
rect 17451 12597 17463 12600
rect 17405 12591 17463 12597
rect 20070 12588 20076 12600
rect 20128 12628 20134 12640
rect 23014 12628 23020 12640
rect 20128 12600 23020 12628
rect 20128 12588 20134 12600
rect 23014 12588 23020 12600
rect 23072 12588 23078 12640
rect 23198 12628 23204 12640
rect 23159 12600 23204 12628
rect 23198 12588 23204 12600
rect 23256 12588 23262 12640
rect 23658 12588 23664 12640
rect 23716 12628 23722 12640
rect 24026 12628 24032 12640
rect 23716 12600 24032 12628
rect 23716 12588 23722 12600
rect 24026 12588 24032 12600
rect 24084 12588 24090 12640
rect 24121 12631 24179 12637
rect 24121 12597 24133 12631
rect 24167 12628 24179 12631
rect 24302 12628 24308 12640
rect 24167 12600 24308 12628
rect 24167 12597 24179 12600
rect 24121 12591 24179 12597
rect 24302 12588 24308 12600
rect 24360 12588 24366 12640
rect 24578 12588 24584 12640
rect 24636 12628 24642 12640
rect 24780 12628 24808 12668
rect 25406 12656 25412 12668
rect 25464 12656 25470 12708
rect 25958 12696 25964 12708
rect 25516 12668 25964 12696
rect 24636 12600 24808 12628
rect 24636 12588 24642 12600
rect 24854 12588 24860 12640
rect 24912 12628 24918 12640
rect 25222 12628 25228 12640
rect 24912 12600 25228 12628
rect 24912 12588 24918 12600
rect 25222 12588 25228 12600
rect 25280 12588 25286 12640
rect 25314 12588 25320 12640
rect 25372 12628 25378 12640
rect 25516 12628 25544 12668
rect 25958 12656 25964 12668
rect 26016 12656 26022 12708
rect 25372 12600 25544 12628
rect 25372 12588 25378 12600
rect 25590 12588 25596 12640
rect 25648 12628 25654 12640
rect 26053 12631 26111 12637
rect 26053 12628 26065 12631
rect 25648 12600 26065 12628
rect 25648 12588 25654 12600
rect 26053 12597 26065 12600
rect 26099 12597 26111 12631
rect 26160 12628 26188 12736
rect 27338 12724 27344 12736
rect 27396 12724 27402 12776
rect 27617 12767 27675 12773
rect 27617 12733 27629 12767
rect 27663 12764 27675 12767
rect 28902 12764 28908 12776
rect 27663 12736 28908 12764
rect 27663 12733 27675 12736
rect 27617 12727 27675 12733
rect 28902 12724 28908 12736
rect 28960 12724 28966 12776
rect 29546 12764 29552 12776
rect 29507 12736 29552 12764
rect 29546 12724 29552 12736
rect 29604 12724 29610 12776
rect 29825 12767 29883 12773
rect 29825 12764 29837 12767
rect 29656 12736 29837 12764
rect 29086 12656 29092 12708
rect 29144 12696 29150 12708
rect 29656 12696 29684 12736
rect 29825 12733 29837 12736
rect 29871 12733 29883 12767
rect 29825 12727 29883 12733
rect 30282 12724 30288 12776
rect 30340 12764 30346 12776
rect 32125 12767 32183 12773
rect 32125 12764 32137 12767
rect 30340 12736 32137 12764
rect 30340 12724 30346 12736
rect 32125 12733 32137 12736
rect 32171 12764 32183 12767
rect 33594 12764 33600 12776
rect 32171 12736 33600 12764
rect 32171 12733 32183 12736
rect 32125 12727 32183 12733
rect 33594 12724 33600 12736
rect 33652 12724 33658 12776
rect 33888 12773 33916 12804
rect 34146 12792 34152 12804
rect 34204 12792 34210 12844
rect 34609 12835 34667 12841
rect 34609 12801 34621 12835
rect 34655 12832 34667 12835
rect 35158 12832 35164 12844
rect 34655 12804 35164 12832
rect 34655 12801 34667 12804
rect 34609 12795 34667 12801
rect 35158 12792 35164 12804
rect 35216 12792 35222 12844
rect 35250 12792 35256 12844
rect 35308 12832 35314 12844
rect 35710 12832 35716 12844
rect 35308 12804 35716 12832
rect 35308 12792 35314 12804
rect 35710 12792 35716 12804
rect 35768 12792 35774 12844
rect 36262 12832 36268 12844
rect 36223 12804 36268 12832
rect 36262 12792 36268 12804
rect 36320 12792 36326 12844
rect 36556 12841 36584 12940
rect 36906 12928 36912 12940
rect 36964 12928 36970 12980
rect 37274 12968 37280 12980
rect 37235 12940 37280 12968
rect 37274 12928 37280 12940
rect 37332 12928 37338 12980
rect 38470 12968 38476 12980
rect 38383 12940 38476 12968
rect 38470 12928 38476 12940
rect 38528 12968 38534 12980
rect 39298 12968 39304 12980
rect 38528 12940 39304 12968
rect 38528 12928 38534 12940
rect 39298 12928 39304 12940
rect 39356 12928 39362 12980
rect 39761 12971 39819 12977
rect 39761 12937 39773 12971
rect 39807 12968 39819 12971
rect 39850 12968 39856 12980
rect 39807 12940 39856 12968
rect 39807 12937 39819 12940
rect 39761 12931 39819 12937
rect 39850 12928 39856 12940
rect 39908 12928 39914 12980
rect 41049 12971 41107 12977
rect 41049 12937 41061 12971
rect 41095 12968 41107 12971
rect 41414 12968 41420 12980
rect 41095 12940 41420 12968
rect 41095 12937 41107 12940
rect 41049 12931 41107 12937
rect 41414 12928 41420 12940
rect 41472 12928 41478 12980
rect 41601 12971 41659 12977
rect 41601 12937 41613 12971
rect 41647 12968 41659 12971
rect 42334 12968 42340 12980
rect 41647 12940 42340 12968
rect 41647 12937 41659 12940
rect 41601 12931 41659 12937
rect 42334 12928 42340 12940
rect 42392 12928 42398 12980
rect 42426 12928 42432 12980
rect 42484 12968 42490 12980
rect 42521 12971 42579 12977
rect 42521 12968 42533 12971
rect 42484 12940 42533 12968
rect 42484 12928 42490 12940
rect 42521 12937 42533 12940
rect 42567 12968 42579 12971
rect 44726 12968 44732 12980
rect 42567 12940 44732 12968
rect 42567 12937 42579 12940
rect 42521 12931 42579 12937
rect 44726 12928 44732 12940
rect 44784 12928 44790 12980
rect 58158 12968 58164 12980
rect 58119 12940 58164 12968
rect 58158 12928 58164 12940
rect 58216 12928 58222 12980
rect 36722 12860 36728 12912
rect 36780 12900 36786 12912
rect 39117 12903 39175 12909
rect 39117 12900 39129 12903
rect 36780 12872 39129 12900
rect 36780 12860 36786 12872
rect 39117 12869 39129 12872
rect 39163 12869 39175 12903
rect 39117 12863 39175 12869
rect 40034 12860 40040 12912
rect 40092 12900 40098 12912
rect 41322 12900 41328 12912
rect 40092 12872 41328 12900
rect 40092 12860 40098 12872
rect 41322 12860 41328 12872
rect 41380 12900 41386 12912
rect 43533 12903 43591 12909
rect 43533 12900 43545 12903
rect 41380 12872 43545 12900
rect 41380 12860 41386 12872
rect 43533 12869 43545 12872
rect 43579 12869 43591 12903
rect 43533 12863 43591 12869
rect 36541 12835 36599 12841
rect 36541 12832 36553 12835
rect 36372 12804 36553 12832
rect 33873 12767 33931 12773
rect 33873 12733 33885 12767
rect 33919 12733 33931 12767
rect 33873 12727 33931 12733
rect 34054 12724 34060 12776
rect 34112 12764 34118 12776
rect 34333 12767 34391 12773
rect 34333 12764 34345 12767
rect 34112 12736 34345 12764
rect 34112 12724 34118 12736
rect 34333 12733 34345 12736
rect 34379 12733 34391 12767
rect 35176 12764 35204 12792
rect 35802 12764 35808 12776
rect 35176 12736 35808 12764
rect 34333 12727 34391 12733
rect 35802 12724 35808 12736
rect 35860 12724 35866 12776
rect 36372 12764 36400 12804
rect 36541 12801 36553 12804
rect 36587 12801 36599 12835
rect 36541 12795 36599 12801
rect 36998 12792 37004 12844
rect 37056 12832 37062 12844
rect 37645 12835 37703 12841
rect 37645 12832 37657 12835
rect 37056 12804 37657 12832
rect 37056 12792 37062 12804
rect 37645 12801 37657 12804
rect 37691 12801 37703 12835
rect 37645 12795 37703 12801
rect 38010 12792 38016 12844
rect 38068 12832 38074 12844
rect 38289 12835 38347 12841
rect 38289 12832 38301 12835
rect 38068 12804 38301 12832
rect 38068 12792 38074 12804
rect 38289 12801 38301 12804
rect 38335 12801 38347 12835
rect 38562 12832 38568 12844
rect 38523 12804 38568 12832
rect 38289 12795 38347 12801
rect 38562 12792 38568 12804
rect 38620 12792 38626 12844
rect 38930 12792 38936 12844
rect 38988 12832 38994 12844
rect 39025 12835 39083 12841
rect 39025 12832 39037 12835
rect 38988 12804 39037 12832
rect 38988 12792 38994 12804
rect 39025 12801 39037 12804
rect 39071 12832 39083 12835
rect 39206 12832 39212 12844
rect 39071 12804 39212 12832
rect 39071 12801 39083 12804
rect 39025 12795 39083 12801
rect 39206 12792 39212 12804
rect 39264 12792 39270 12844
rect 39853 12835 39911 12841
rect 39853 12801 39865 12835
rect 39899 12801 39911 12835
rect 39853 12795 39911 12801
rect 35912 12736 36400 12764
rect 36449 12767 36507 12773
rect 29144 12668 29684 12696
rect 29144 12656 29150 12668
rect 33686 12656 33692 12708
rect 33744 12696 33750 12708
rect 33744 12668 34468 12696
rect 33744 12656 33750 12668
rect 32214 12628 32220 12640
rect 26160 12600 32220 12628
rect 26053 12591 26111 12597
rect 32214 12588 32220 12600
rect 32272 12588 32278 12640
rect 33410 12588 33416 12640
rect 33468 12628 33474 12640
rect 34054 12628 34060 12640
rect 33468 12600 34060 12628
rect 33468 12588 33474 12600
rect 34054 12588 34060 12600
rect 34112 12588 34118 12640
rect 34440 12628 34468 12668
rect 35250 12656 35256 12708
rect 35308 12696 35314 12708
rect 35912 12696 35940 12736
rect 36449 12733 36461 12767
rect 36495 12764 36507 12767
rect 36722 12764 36728 12776
rect 36495 12736 36728 12764
rect 36495 12733 36507 12736
rect 36449 12727 36507 12733
rect 36722 12724 36728 12736
rect 36780 12724 36786 12776
rect 37458 12724 37464 12776
rect 37516 12764 37522 12776
rect 37553 12767 37611 12773
rect 37553 12764 37565 12767
rect 37516 12736 37565 12764
rect 37516 12724 37522 12736
rect 37553 12733 37565 12736
rect 37599 12733 37611 12767
rect 37553 12727 37611 12733
rect 38838 12724 38844 12776
rect 38896 12764 38902 12776
rect 39868 12764 39896 12795
rect 40402 12792 40408 12844
rect 40460 12832 40466 12844
rect 40497 12835 40555 12841
rect 40497 12832 40509 12835
rect 40460 12804 40509 12832
rect 40460 12792 40466 12804
rect 40497 12801 40509 12804
rect 40543 12832 40555 12835
rect 42518 12832 42524 12844
rect 40543 12804 42524 12832
rect 40543 12801 40555 12804
rect 40497 12795 40555 12801
rect 42518 12792 42524 12804
rect 42576 12792 42582 12844
rect 42981 12767 43039 12773
rect 42981 12764 42993 12767
rect 38896 12736 42993 12764
rect 38896 12724 38902 12736
rect 42981 12733 42993 12736
rect 43027 12764 43039 12767
rect 43714 12764 43720 12776
rect 43027 12736 43720 12764
rect 43027 12733 43039 12736
rect 42981 12727 43039 12733
rect 43714 12724 43720 12736
rect 43772 12724 43778 12776
rect 35308 12668 35940 12696
rect 35308 12656 35314 12668
rect 35986 12656 35992 12708
rect 36044 12696 36050 12708
rect 36081 12699 36139 12705
rect 36081 12696 36093 12699
rect 36044 12668 36093 12696
rect 36044 12656 36050 12668
rect 36081 12665 36093 12668
rect 36127 12696 36139 12699
rect 36127 12668 37228 12696
rect 36127 12665 36139 12668
rect 36081 12659 36139 12665
rect 35434 12628 35440 12640
rect 34440 12600 35440 12628
rect 35434 12588 35440 12600
rect 35492 12588 35498 12640
rect 35894 12588 35900 12640
rect 35952 12628 35958 12640
rect 36265 12631 36323 12637
rect 36265 12628 36277 12631
rect 35952 12600 36277 12628
rect 35952 12588 35958 12600
rect 36265 12597 36277 12600
rect 36311 12628 36323 12631
rect 37090 12628 37096 12640
rect 36311 12600 37096 12628
rect 36311 12597 36323 12600
rect 36265 12591 36323 12597
rect 37090 12588 37096 12600
rect 37148 12588 37154 12640
rect 37200 12628 37228 12668
rect 37274 12656 37280 12708
rect 37332 12696 37338 12708
rect 38289 12699 38347 12705
rect 38289 12696 38301 12699
rect 37332 12668 38301 12696
rect 37332 12656 37338 12668
rect 38289 12665 38301 12668
rect 38335 12665 38347 12699
rect 38289 12659 38347 12665
rect 38930 12656 38936 12708
rect 38988 12696 38994 12708
rect 39482 12696 39488 12708
rect 38988 12668 39488 12696
rect 38988 12656 38994 12668
rect 39482 12656 39488 12668
rect 39540 12656 39546 12708
rect 40862 12656 40868 12708
rect 40920 12656 40926 12708
rect 41230 12656 41236 12708
rect 41288 12696 41294 12708
rect 42426 12696 42432 12708
rect 41288 12668 42432 12696
rect 41288 12656 41294 12668
rect 42426 12656 42432 12668
rect 42484 12656 42490 12708
rect 44177 12699 44235 12705
rect 44177 12665 44189 12699
rect 44223 12696 44235 12699
rect 44358 12696 44364 12708
rect 44223 12668 44364 12696
rect 44223 12665 44235 12668
rect 44177 12659 44235 12665
rect 44358 12656 44364 12668
rect 44416 12696 44422 12708
rect 57882 12696 57888 12708
rect 44416 12668 57888 12696
rect 44416 12656 44422 12668
rect 57882 12656 57888 12668
rect 57940 12656 57946 12708
rect 40880 12628 40908 12656
rect 44634 12628 44640 12640
rect 37200 12600 40908 12628
rect 44595 12600 44640 12628
rect 44634 12588 44640 12600
rect 44692 12588 44698 12640
rect 45186 12628 45192 12640
rect 45147 12600 45192 12628
rect 45186 12588 45192 12600
rect 45244 12588 45250 12640
rect 1104 12538 58880 12560
rect 1104 12486 10582 12538
rect 10634 12486 10646 12538
rect 10698 12486 10710 12538
rect 10762 12486 10774 12538
rect 10826 12486 10838 12538
rect 10890 12486 29846 12538
rect 29898 12486 29910 12538
rect 29962 12486 29974 12538
rect 30026 12486 30038 12538
rect 30090 12486 30102 12538
rect 30154 12486 49110 12538
rect 49162 12486 49174 12538
rect 49226 12486 49238 12538
rect 49290 12486 49302 12538
rect 49354 12486 49366 12538
rect 49418 12486 58880 12538
rect 1104 12464 58880 12486
rect 12894 12424 12900 12436
rect 12855 12396 12900 12424
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 18690 12424 18696 12436
rect 18651 12396 18696 12424
rect 18690 12384 18696 12396
rect 18748 12384 18754 12436
rect 19702 12424 19708 12436
rect 19663 12396 19708 12424
rect 19702 12384 19708 12396
rect 19760 12384 19766 12436
rect 20898 12424 20904 12436
rect 20859 12396 20904 12424
rect 20898 12384 20904 12396
rect 20956 12384 20962 12436
rect 21542 12384 21548 12436
rect 21600 12424 21606 12436
rect 21910 12424 21916 12436
rect 21600 12396 21916 12424
rect 21600 12384 21606 12396
rect 21910 12384 21916 12396
rect 21968 12384 21974 12436
rect 24578 12384 24584 12436
rect 24636 12424 24642 12436
rect 25130 12424 25136 12436
rect 24636 12396 25136 12424
rect 24636 12384 24642 12396
rect 25130 12384 25136 12396
rect 25188 12384 25194 12436
rect 25590 12384 25596 12436
rect 25648 12424 25654 12436
rect 25777 12427 25835 12433
rect 25648 12396 25728 12424
rect 25648 12384 25654 12396
rect 20349 12359 20407 12365
rect 20349 12325 20361 12359
rect 20395 12356 20407 12359
rect 22094 12356 22100 12368
rect 20395 12328 22100 12356
rect 20395 12325 20407 12328
rect 20349 12319 20407 12325
rect 22094 12316 22100 12328
rect 22152 12316 22158 12368
rect 22370 12356 22376 12368
rect 22331 12328 22376 12356
rect 22370 12316 22376 12328
rect 22428 12356 22434 12368
rect 24762 12356 24768 12368
rect 22428 12328 24532 12356
rect 24723 12328 24768 12356
rect 22428 12316 22434 12328
rect 19426 12248 19432 12300
rect 19484 12288 19490 12300
rect 23017 12291 23075 12297
rect 23017 12288 23029 12291
rect 19484 12260 23029 12288
rect 19484 12248 19490 12260
rect 23017 12257 23029 12260
rect 23063 12257 23075 12291
rect 23017 12251 23075 12257
rect 24210 12248 24216 12300
rect 24268 12288 24274 12300
rect 24268 12260 24439 12288
rect 24268 12248 24274 12260
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12220 1731 12223
rect 11330 12220 11336 12232
rect 1719 12192 11336 12220
rect 1719 12189 1731 12192
rect 1673 12183 1731 12189
rect 11330 12180 11336 12192
rect 11388 12180 11394 12232
rect 12345 12223 12403 12229
rect 12345 12189 12357 12223
rect 12391 12220 12403 12223
rect 12894 12220 12900 12232
rect 12391 12192 12900 12220
rect 12391 12189 12403 12192
rect 12345 12183 12403 12189
rect 12894 12180 12900 12192
rect 12952 12180 12958 12232
rect 21818 12180 21824 12232
rect 21876 12220 21882 12232
rect 22925 12223 22983 12229
rect 22925 12220 22937 12223
rect 21876 12192 22937 12220
rect 21876 12180 21882 12192
rect 22925 12189 22937 12192
rect 22971 12189 22983 12223
rect 22925 12183 22983 12189
rect 23109 12223 23167 12229
rect 23109 12189 23121 12223
rect 23155 12189 23167 12223
rect 23566 12220 23572 12232
rect 23527 12192 23572 12220
rect 23109 12183 23167 12189
rect 16298 12112 16304 12164
rect 16356 12152 16362 12164
rect 23124 12152 23152 12183
rect 23566 12180 23572 12192
rect 23624 12180 23630 12232
rect 24411 12229 24439 12260
rect 24504 12229 24532 12328
rect 24762 12316 24768 12328
rect 24820 12316 24826 12368
rect 24946 12316 24952 12368
rect 25004 12356 25010 12368
rect 25700 12356 25728 12396
rect 25777 12393 25789 12427
rect 25823 12424 25835 12427
rect 25866 12424 25872 12436
rect 25823 12396 25872 12424
rect 25823 12393 25835 12396
rect 25777 12387 25835 12393
rect 25866 12384 25872 12396
rect 25924 12384 25930 12436
rect 26786 12424 26792 12436
rect 26747 12396 26792 12424
rect 26786 12384 26792 12396
rect 26844 12384 26850 12436
rect 28997 12427 29055 12433
rect 26896 12396 28948 12424
rect 26050 12356 26056 12368
rect 25004 12328 25636 12356
rect 25700 12328 26056 12356
rect 25004 12316 25010 12328
rect 24581 12291 24639 12297
rect 24581 12257 24593 12291
rect 24627 12288 24639 12291
rect 24670 12288 24676 12300
rect 24627 12260 24676 12288
rect 24627 12257 24639 12260
rect 24581 12251 24639 12257
rect 24670 12248 24676 12260
rect 24728 12288 24734 12300
rect 25222 12288 25228 12300
rect 24728 12260 25228 12288
rect 24728 12248 24734 12260
rect 25222 12248 25228 12260
rect 25280 12248 25286 12300
rect 25424 12229 25452 12328
rect 25501 12291 25559 12297
rect 25501 12257 25513 12291
rect 25547 12257 25559 12291
rect 25608 12288 25636 12328
rect 26050 12316 26056 12328
rect 26108 12316 26114 12368
rect 26418 12316 26424 12368
rect 26476 12356 26482 12368
rect 26896 12356 26924 12396
rect 26476 12328 26924 12356
rect 28920 12356 28948 12396
rect 28997 12393 29009 12427
rect 29043 12424 29055 12427
rect 29362 12424 29368 12436
rect 29043 12396 29368 12424
rect 29043 12393 29055 12396
rect 28997 12387 29055 12393
rect 29362 12384 29368 12396
rect 29420 12424 29426 12436
rect 32398 12424 32404 12436
rect 29420 12396 32404 12424
rect 29420 12384 29426 12396
rect 32398 12384 32404 12396
rect 32456 12424 32462 12436
rect 36262 12424 36268 12436
rect 32456 12396 36124 12424
rect 36223 12396 36268 12424
rect 32456 12384 32462 12396
rect 28920 12328 29408 12356
rect 26476 12316 26482 12328
rect 29380 12300 29408 12328
rect 31110 12316 31116 12368
rect 31168 12356 31174 12368
rect 31294 12356 31300 12368
rect 31168 12328 31300 12356
rect 31168 12316 31174 12328
rect 31294 12316 31300 12328
rect 31352 12316 31358 12368
rect 31478 12356 31484 12368
rect 31439 12328 31484 12356
rect 31478 12316 31484 12328
rect 31536 12316 31542 12368
rect 33594 12316 33600 12368
rect 33652 12356 33658 12368
rect 33870 12356 33876 12368
rect 33652 12328 33876 12356
rect 33652 12316 33658 12328
rect 33870 12316 33876 12328
rect 33928 12356 33934 12368
rect 35618 12356 35624 12368
rect 33928 12328 35624 12356
rect 33928 12316 33934 12328
rect 35618 12316 35624 12328
rect 35676 12316 35682 12368
rect 36096 12356 36124 12396
rect 36262 12384 36268 12396
rect 36320 12384 36326 12436
rect 36449 12427 36507 12433
rect 36449 12393 36461 12427
rect 36495 12424 36507 12427
rect 36814 12424 36820 12436
rect 36495 12396 36820 12424
rect 36495 12393 36507 12396
rect 36449 12387 36507 12393
rect 36814 12384 36820 12396
rect 36872 12384 36878 12436
rect 37090 12384 37096 12436
rect 37148 12424 37154 12436
rect 37921 12427 37979 12433
rect 37148 12396 37872 12424
rect 37148 12384 37154 12396
rect 36998 12356 37004 12368
rect 36096 12328 37004 12356
rect 25958 12288 25964 12300
rect 25608 12260 25964 12288
rect 25501 12251 25559 12257
rect 24397 12223 24455 12229
rect 24397 12189 24409 12223
rect 24443 12189 24455 12223
rect 24397 12183 24455 12189
rect 24489 12223 24547 12229
rect 24489 12189 24501 12223
rect 24535 12189 24547 12223
rect 24489 12183 24547 12189
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 25409 12223 25467 12229
rect 25409 12189 25421 12223
rect 25455 12189 25467 12223
rect 25516 12220 25544 12251
rect 25958 12248 25964 12260
rect 26016 12248 26022 12300
rect 26326 12288 26332 12300
rect 26287 12260 26332 12288
rect 26326 12248 26332 12260
rect 26384 12248 26390 12300
rect 26786 12248 26792 12300
rect 26844 12288 26850 12300
rect 27890 12288 27896 12300
rect 26844 12260 27896 12288
rect 26844 12248 26850 12260
rect 27890 12248 27896 12260
rect 27948 12248 27954 12300
rect 29362 12248 29368 12300
rect 29420 12248 29426 12300
rect 29748 12260 31616 12288
rect 25866 12220 25872 12232
rect 25516 12192 25872 12220
rect 25409 12183 25467 12189
rect 23474 12152 23480 12164
rect 16356 12124 23060 12152
rect 23124 12124 23480 12152
rect 16356 12112 16362 12124
rect 1486 12084 1492 12096
rect 1447 12056 1492 12084
rect 1486 12044 1492 12056
rect 1544 12044 1550 12096
rect 11054 12044 11060 12096
rect 11112 12084 11118 12096
rect 12161 12087 12219 12093
rect 12161 12084 12173 12087
rect 11112 12056 12173 12084
rect 11112 12044 11118 12056
rect 12161 12053 12173 12056
rect 12207 12053 12219 12087
rect 18138 12084 18144 12096
rect 18099 12056 18144 12084
rect 12161 12047 12219 12053
rect 18138 12044 18144 12056
rect 18196 12044 18202 12096
rect 23032 12084 23060 12124
rect 23474 12112 23480 12124
rect 23532 12112 23538 12164
rect 24412 12152 24440 12183
rect 24578 12152 24584 12164
rect 24412 12124 24584 12152
rect 24578 12112 24584 12124
rect 24636 12112 24642 12164
rect 24780 12152 24808 12183
rect 25866 12180 25872 12192
rect 25924 12180 25930 12232
rect 26421 12223 26479 12229
rect 26421 12189 26433 12223
rect 26467 12220 26479 12223
rect 26467 12192 27108 12220
rect 26467 12189 26479 12192
rect 26421 12183 26479 12189
rect 26786 12152 26792 12164
rect 24780 12124 26792 12152
rect 26786 12112 26792 12124
rect 26844 12112 26850 12164
rect 23753 12087 23811 12093
rect 23753 12084 23765 12087
rect 23032 12056 23765 12084
rect 23753 12053 23765 12056
rect 23799 12084 23811 12087
rect 25958 12084 25964 12096
rect 23799 12056 25964 12084
rect 23799 12053 23811 12056
rect 23753 12047 23811 12053
rect 25958 12044 25964 12056
rect 26016 12044 26022 12096
rect 27080 12084 27108 12192
rect 27154 12180 27160 12232
rect 27212 12220 27218 12232
rect 27249 12223 27307 12229
rect 27249 12220 27261 12223
rect 27212 12192 27261 12220
rect 27212 12180 27218 12192
rect 27249 12189 27261 12192
rect 27295 12189 27307 12223
rect 27249 12183 27307 12189
rect 29546 12180 29552 12232
rect 29604 12220 29610 12232
rect 29748 12229 29776 12260
rect 29733 12223 29791 12229
rect 29733 12220 29745 12223
rect 29604 12192 29745 12220
rect 29604 12180 29610 12192
rect 29733 12189 29745 12192
rect 29779 12189 29791 12223
rect 31588 12220 31616 12260
rect 31662 12248 31668 12300
rect 31720 12288 31726 12300
rect 36096 12297 36124 12328
rect 36998 12316 37004 12328
rect 37056 12316 37062 12368
rect 37550 12356 37556 12368
rect 37108 12328 37556 12356
rect 36081 12291 36139 12297
rect 31720 12260 36032 12288
rect 31720 12248 31726 12260
rect 31938 12220 31944 12232
rect 31588 12192 31944 12220
rect 29733 12183 29791 12189
rect 31938 12180 31944 12192
rect 31996 12180 32002 12232
rect 33962 12180 33968 12232
rect 34020 12220 34026 12232
rect 34238 12220 34244 12232
rect 34020 12192 34244 12220
rect 34020 12180 34026 12192
rect 34238 12180 34244 12192
rect 34296 12220 34302 12232
rect 34701 12223 34759 12229
rect 34701 12220 34713 12223
rect 34296 12192 34713 12220
rect 34296 12180 34302 12192
rect 34701 12189 34713 12192
rect 34747 12189 34759 12223
rect 34701 12183 34759 12189
rect 34977 12223 35035 12229
rect 34977 12189 34989 12223
rect 35023 12220 35035 12223
rect 35250 12220 35256 12232
rect 35023 12192 35256 12220
rect 35023 12189 35035 12192
rect 34977 12183 35035 12189
rect 35250 12180 35256 12192
rect 35308 12220 35314 12232
rect 35526 12220 35532 12232
rect 35308 12192 35532 12220
rect 35308 12180 35314 12192
rect 35526 12180 35532 12192
rect 35584 12180 35590 12232
rect 36004 12220 36032 12260
rect 36081 12257 36093 12291
rect 36127 12257 36139 12291
rect 36081 12251 36139 12257
rect 36265 12223 36323 12229
rect 36004 12192 36216 12220
rect 27522 12152 27528 12164
rect 27483 12124 27528 12152
rect 27522 12112 27528 12124
rect 27580 12112 27586 12164
rect 28258 12112 28264 12164
rect 28316 12112 28322 12164
rect 29086 12112 29092 12164
rect 29144 12152 29150 12164
rect 30009 12155 30067 12161
rect 30009 12152 30021 12155
rect 29144 12124 30021 12152
rect 29144 12112 29150 12124
rect 30009 12121 30021 12124
rect 30055 12121 30067 12155
rect 31662 12152 31668 12164
rect 31234 12124 31668 12152
rect 30009 12115 30067 12121
rect 31662 12112 31668 12124
rect 31720 12112 31726 12164
rect 32217 12155 32275 12161
rect 32217 12121 32229 12155
rect 32263 12152 32275 12155
rect 32306 12152 32312 12164
rect 32263 12124 32312 12152
rect 32263 12121 32275 12124
rect 32217 12115 32275 12121
rect 32306 12112 32312 12124
rect 32364 12112 32370 12164
rect 32674 12152 32680 12164
rect 32600 12124 32680 12152
rect 30190 12084 30196 12096
rect 27080 12056 30196 12084
rect 30190 12044 30196 12056
rect 30248 12044 30254 12096
rect 31680 12084 31708 12112
rect 32600 12084 32628 12124
rect 32674 12112 32680 12124
rect 32732 12112 32738 12164
rect 35989 12155 36047 12161
rect 35989 12121 36001 12155
rect 36035 12152 36047 12155
rect 36078 12152 36084 12164
rect 36035 12124 36084 12152
rect 36035 12121 36047 12124
rect 35989 12115 36047 12121
rect 36078 12112 36084 12124
rect 36136 12112 36142 12164
rect 36188 12152 36216 12192
rect 36265 12189 36277 12223
rect 36311 12220 36323 12223
rect 37108 12220 37136 12328
rect 37550 12316 37556 12328
rect 37608 12316 37614 12368
rect 37844 12356 37872 12396
rect 37921 12393 37933 12427
rect 37967 12424 37979 12427
rect 38746 12424 38752 12436
rect 37967 12396 38752 12424
rect 37967 12393 37979 12396
rect 37921 12387 37979 12393
rect 38746 12384 38752 12396
rect 38804 12384 38810 12436
rect 40586 12384 40592 12436
rect 40644 12424 40650 12436
rect 41509 12427 41567 12433
rect 41509 12424 41521 12427
rect 40644 12396 41521 12424
rect 40644 12384 40650 12396
rect 41509 12393 41521 12396
rect 41555 12393 41567 12427
rect 41509 12387 41567 12393
rect 43257 12427 43315 12433
rect 43257 12393 43269 12427
rect 43303 12424 43315 12427
rect 45922 12424 45928 12436
rect 43303 12396 45928 12424
rect 43303 12393 43315 12396
rect 43257 12387 43315 12393
rect 45922 12384 45928 12396
rect 45980 12384 45986 12436
rect 39853 12359 39911 12365
rect 39853 12356 39865 12359
rect 37844 12328 39865 12356
rect 39853 12325 39865 12328
rect 39899 12356 39911 12359
rect 39942 12356 39948 12368
rect 39899 12328 39948 12356
rect 39899 12325 39911 12328
rect 39853 12319 39911 12325
rect 39942 12316 39948 12328
rect 40000 12316 40006 12368
rect 40402 12356 40408 12368
rect 40363 12328 40408 12356
rect 40402 12316 40408 12328
rect 40460 12316 40466 12368
rect 42705 12359 42763 12365
rect 42705 12325 42717 12359
rect 42751 12356 42763 12359
rect 43530 12356 43536 12368
rect 42751 12328 43536 12356
rect 42751 12325 42763 12328
rect 42705 12319 42763 12325
rect 43530 12316 43536 12328
rect 43588 12316 43594 12368
rect 38010 12288 38016 12300
rect 37200 12260 38016 12288
rect 37200 12229 37228 12260
rect 38010 12248 38016 12260
rect 38068 12248 38074 12300
rect 36311 12192 37136 12220
rect 37185 12223 37243 12229
rect 36311 12189 36323 12192
rect 36265 12183 36323 12189
rect 37185 12189 37197 12223
rect 37231 12189 37243 12223
rect 37185 12183 37243 12189
rect 37921 12223 37979 12229
rect 37921 12189 37933 12223
rect 37967 12220 37979 12223
rect 38102 12220 38108 12232
rect 37967 12192 38108 12220
rect 37967 12189 37979 12192
rect 37921 12183 37979 12189
rect 38102 12180 38108 12192
rect 38160 12180 38166 12232
rect 38654 12220 38660 12232
rect 38567 12192 38660 12220
rect 38654 12180 38660 12192
rect 38712 12220 38718 12232
rect 39850 12220 39856 12232
rect 38712 12192 39856 12220
rect 38712 12180 38718 12192
rect 39850 12180 39856 12192
rect 39908 12180 39914 12232
rect 38010 12152 38016 12164
rect 36188 12124 38016 12152
rect 38010 12112 38016 12124
rect 38068 12112 38074 12164
rect 31680 12056 32628 12084
rect 33042 12044 33048 12096
rect 33100 12084 33106 12096
rect 33689 12087 33747 12093
rect 33689 12084 33701 12087
rect 33100 12056 33701 12084
rect 33100 12044 33106 12056
rect 33689 12053 33701 12056
rect 33735 12084 33747 12087
rect 35618 12084 35624 12096
rect 33735 12056 35624 12084
rect 33735 12053 33747 12056
rect 33689 12047 33747 12053
rect 35618 12044 35624 12056
rect 35676 12044 35682 12096
rect 36630 12044 36636 12096
rect 36688 12084 36694 12096
rect 37093 12087 37151 12093
rect 37093 12084 37105 12087
rect 36688 12056 37105 12084
rect 36688 12044 36694 12056
rect 37093 12053 37105 12056
rect 37139 12053 37151 12087
rect 37093 12047 37151 12053
rect 37550 12044 37556 12096
rect 37608 12084 37614 12096
rect 38565 12087 38623 12093
rect 38565 12084 38577 12087
rect 37608 12056 38577 12084
rect 37608 12044 37614 12056
rect 38565 12053 38577 12056
rect 38611 12053 38623 12087
rect 38565 12047 38623 12053
rect 38746 12044 38752 12096
rect 38804 12084 38810 12096
rect 38930 12084 38936 12096
rect 38804 12056 38936 12084
rect 38804 12044 38810 12056
rect 38930 12044 38936 12056
rect 38988 12084 38994 12096
rect 39117 12087 39175 12093
rect 39117 12084 39129 12087
rect 38988 12056 39129 12084
rect 38988 12044 38994 12056
rect 39117 12053 39129 12056
rect 39163 12053 39175 12087
rect 39117 12047 39175 12053
rect 40862 12044 40868 12096
rect 40920 12084 40926 12096
rect 40957 12087 41015 12093
rect 40957 12084 40969 12087
rect 40920 12056 40969 12084
rect 40920 12044 40926 12056
rect 40957 12053 40969 12056
rect 41003 12053 41015 12087
rect 42058 12084 42064 12096
rect 42019 12056 42064 12084
rect 40957 12047 41015 12053
rect 42058 12044 42064 12056
rect 42116 12044 42122 12096
rect 43714 12084 43720 12096
rect 43675 12056 43720 12084
rect 43714 12044 43720 12056
rect 43772 12044 43778 12096
rect 44358 12084 44364 12096
rect 44271 12056 44364 12084
rect 44358 12044 44364 12056
rect 44416 12084 44422 12096
rect 45554 12084 45560 12096
rect 44416 12056 45560 12084
rect 44416 12044 44422 12056
rect 45554 12044 45560 12056
rect 45612 12084 45618 12096
rect 46106 12084 46112 12096
rect 45612 12056 46112 12084
rect 45612 12044 45618 12056
rect 46106 12044 46112 12056
rect 46164 12044 46170 12096
rect 1104 11994 58880 12016
rect 1104 11942 20214 11994
rect 20266 11942 20278 11994
rect 20330 11942 20342 11994
rect 20394 11942 20406 11994
rect 20458 11942 20470 11994
rect 20522 11942 39478 11994
rect 39530 11942 39542 11994
rect 39594 11942 39606 11994
rect 39658 11942 39670 11994
rect 39722 11942 39734 11994
rect 39786 11942 58880 11994
rect 1104 11920 58880 11942
rect 15746 11840 15752 11892
rect 15804 11880 15810 11892
rect 16298 11880 16304 11892
rect 15804 11852 16304 11880
rect 15804 11840 15810 11852
rect 16298 11840 16304 11852
rect 16356 11840 16362 11892
rect 21913 11883 21971 11889
rect 21913 11849 21925 11883
rect 21959 11880 21971 11883
rect 22186 11880 22192 11892
rect 21959 11852 22192 11880
rect 21959 11849 21971 11852
rect 21913 11843 21971 11849
rect 22186 11840 22192 11852
rect 22244 11840 22250 11892
rect 22462 11840 22468 11892
rect 22520 11880 22526 11892
rect 23017 11883 23075 11889
rect 23017 11880 23029 11883
rect 22520 11852 23029 11880
rect 22520 11840 22526 11852
rect 23017 11849 23029 11852
rect 23063 11849 23075 11883
rect 23017 11843 23075 11849
rect 23474 11840 23480 11892
rect 23532 11880 23538 11892
rect 23532 11852 23796 11880
rect 23532 11840 23538 11852
rect 20533 11815 20591 11821
rect 20533 11781 20545 11815
rect 20579 11812 20591 11815
rect 22002 11812 22008 11824
rect 20579 11784 22008 11812
rect 20579 11781 20591 11784
rect 20533 11775 20591 11781
rect 22002 11772 22008 11784
rect 22060 11772 22066 11824
rect 23658 11812 23664 11824
rect 23619 11784 23664 11812
rect 23658 11772 23664 11784
rect 23716 11772 23722 11824
rect 20441 11747 20499 11753
rect 20441 11713 20453 11747
rect 20487 11744 20499 11747
rect 20990 11744 20996 11756
rect 20487 11716 20996 11744
rect 20487 11713 20499 11716
rect 20441 11707 20499 11713
rect 20990 11704 20996 11716
rect 21048 11704 21054 11756
rect 22370 11704 22376 11756
rect 22428 11744 22434 11756
rect 22465 11747 22523 11753
rect 22465 11744 22477 11747
rect 22428 11716 22477 11744
rect 22428 11704 22434 11716
rect 22465 11713 22477 11716
rect 22511 11744 22523 11747
rect 22738 11744 22744 11756
rect 22511 11716 22744 11744
rect 22511 11713 22523 11716
rect 22465 11707 22523 11713
rect 22738 11704 22744 11716
rect 22796 11704 22802 11756
rect 22922 11704 22928 11756
rect 22980 11744 22986 11756
rect 23768 11753 23796 11852
rect 24578 11840 24584 11892
rect 24636 11880 24642 11892
rect 26418 11880 26424 11892
rect 24636 11852 26424 11880
rect 24636 11840 24642 11852
rect 26418 11840 26424 11852
rect 26476 11840 26482 11892
rect 28718 11840 28724 11892
rect 28776 11880 28782 11892
rect 36081 11883 36139 11889
rect 28776 11852 36032 11880
rect 28776 11840 28782 11852
rect 25130 11772 25136 11824
rect 25188 11812 25194 11824
rect 26326 11812 26332 11824
rect 25188 11784 26332 11812
rect 25188 11772 25194 11784
rect 26326 11772 26332 11784
rect 26384 11772 26390 11824
rect 26602 11772 26608 11824
rect 26660 11812 26666 11824
rect 26660 11784 28028 11812
rect 26660 11772 26666 11784
rect 23569 11747 23627 11753
rect 23569 11744 23581 11747
rect 22980 11716 23581 11744
rect 22980 11704 22986 11716
rect 23569 11713 23581 11716
rect 23615 11713 23627 11747
rect 23569 11707 23627 11713
rect 23753 11747 23811 11753
rect 23753 11713 23765 11747
rect 23799 11744 23811 11747
rect 24210 11744 24216 11756
rect 23799 11716 24216 11744
rect 23799 11713 23811 11716
rect 23753 11707 23811 11713
rect 24210 11704 24216 11716
rect 24268 11704 24274 11756
rect 24397 11747 24455 11753
rect 24397 11713 24409 11747
rect 24443 11744 24455 11747
rect 24578 11744 24584 11756
rect 24443 11716 24584 11744
rect 24443 11713 24455 11716
rect 24397 11707 24455 11713
rect 17218 11636 17224 11688
rect 17276 11676 17282 11688
rect 19797 11679 19855 11685
rect 19797 11676 19809 11679
rect 17276 11648 19809 11676
rect 17276 11636 17282 11648
rect 19797 11645 19809 11648
rect 19843 11676 19855 11679
rect 24118 11676 24124 11688
rect 19843 11648 24124 11676
rect 19843 11645 19855 11648
rect 19797 11639 19855 11645
rect 24118 11636 24124 11648
rect 24176 11636 24182 11688
rect 19334 11568 19340 11620
rect 19392 11608 19398 11620
rect 24412 11608 24440 11707
rect 24578 11704 24584 11716
rect 24636 11704 24642 11756
rect 25038 11744 25044 11756
rect 24999 11716 25044 11744
rect 25038 11704 25044 11716
rect 25096 11704 25102 11756
rect 25774 11704 25780 11756
rect 25832 11744 25838 11756
rect 26053 11747 26111 11753
rect 26053 11744 26065 11747
rect 25832 11716 26065 11744
rect 25832 11704 25838 11716
rect 26053 11713 26065 11716
rect 26099 11713 26111 11747
rect 26053 11707 26111 11713
rect 26142 11704 26148 11756
rect 26200 11744 26206 11756
rect 27890 11744 27896 11756
rect 26200 11716 27896 11744
rect 26200 11704 26206 11716
rect 27890 11704 27896 11716
rect 27948 11704 27954 11756
rect 28000 11753 28028 11784
rect 31386 11772 31392 11824
rect 31444 11812 31450 11824
rect 32401 11815 32459 11821
rect 32401 11812 32413 11815
rect 31444 11784 32413 11812
rect 31444 11772 31450 11784
rect 32401 11781 32413 11784
rect 32447 11781 32459 11815
rect 32401 11775 32459 11781
rect 32674 11772 32680 11824
rect 32732 11812 32738 11824
rect 32858 11812 32864 11824
rect 32732 11784 32864 11812
rect 32732 11772 32738 11784
rect 32858 11772 32864 11784
rect 32916 11772 32922 11824
rect 27985 11747 28043 11753
rect 27985 11713 27997 11747
rect 28031 11713 28043 11747
rect 27985 11707 28043 11713
rect 28258 11704 28264 11756
rect 28316 11744 28322 11756
rect 28721 11747 28779 11753
rect 28721 11744 28733 11747
rect 28316 11716 28733 11744
rect 28316 11704 28322 11716
rect 28721 11713 28733 11716
rect 28767 11744 28779 11747
rect 28902 11744 28908 11756
rect 28767 11716 28908 11744
rect 28767 11713 28779 11716
rect 28721 11707 28779 11713
rect 28902 11704 28908 11716
rect 28960 11704 28966 11756
rect 29178 11704 29184 11756
rect 29236 11744 29242 11756
rect 29825 11747 29883 11753
rect 29825 11744 29837 11747
rect 29236 11716 29837 11744
rect 29236 11704 29242 11716
rect 29825 11713 29837 11716
rect 29871 11713 29883 11747
rect 29825 11707 29883 11713
rect 24670 11636 24676 11688
rect 24728 11676 24734 11688
rect 25130 11676 25136 11688
rect 24728 11648 25136 11676
rect 24728 11636 24734 11648
rect 25130 11636 25136 11648
rect 25188 11636 25194 11688
rect 25961 11679 26019 11685
rect 25961 11645 25973 11679
rect 26007 11645 26019 11679
rect 25961 11639 26019 11645
rect 30101 11679 30159 11685
rect 30101 11645 30113 11679
rect 30147 11676 30159 11679
rect 30190 11676 30196 11688
rect 30147 11648 30196 11676
rect 30147 11645 30159 11648
rect 30101 11639 30159 11645
rect 19392 11580 24440 11608
rect 19392 11568 19398 11580
rect 24854 11568 24860 11620
rect 24912 11608 24918 11620
rect 25976 11608 26004 11639
rect 30190 11636 30196 11648
rect 30248 11636 30254 11688
rect 31220 11676 31248 11730
rect 31938 11704 31944 11756
rect 31996 11744 32002 11756
rect 32125 11747 32183 11753
rect 32125 11744 32137 11747
rect 31996 11716 32137 11744
rect 31996 11704 32002 11716
rect 32125 11713 32137 11716
rect 32171 11713 32183 11747
rect 32125 11707 32183 11713
rect 34054 11704 34060 11756
rect 34112 11744 34118 11756
rect 34609 11747 34667 11753
rect 34609 11744 34621 11747
rect 34112 11716 34621 11744
rect 34112 11704 34118 11716
rect 34609 11713 34621 11716
rect 34655 11744 34667 11747
rect 34698 11744 34704 11756
rect 34655 11716 34704 11744
rect 34655 11713 34667 11716
rect 34609 11707 34667 11713
rect 34698 11704 34704 11716
rect 34756 11704 34762 11756
rect 35618 11744 35624 11756
rect 35579 11716 35624 11744
rect 35618 11704 35624 11716
rect 35676 11704 35682 11756
rect 35802 11704 35808 11756
rect 35860 11744 35866 11756
rect 35897 11747 35955 11753
rect 35897 11744 35909 11747
rect 35860 11716 35909 11744
rect 35860 11704 35866 11716
rect 35897 11713 35909 11716
rect 35943 11713 35955 11747
rect 36004 11744 36032 11852
rect 36081 11849 36093 11883
rect 36127 11849 36139 11883
rect 36081 11843 36139 11849
rect 36096 11812 36124 11843
rect 36170 11840 36176 11892
rect 36228 11880 36234 11892
rect 36633 11883 36691 11889
rect 36633 11880 36645 11883
rect 36228 11852 36645 11880
rect 36228 11840 36234 11852
rect 36633 11849 36645 11852
rect 36679 11849 36691 11883
rect 38010 11880 38016 11892
rect 37971 11852 38016 11880
rect 36633 11843 36691 11849
rect 38010 11840 38016 11852
rect 38068 11840 38074 11892
rect 38746 11880 38752 11892
rect 38707 11852 38752 11880
rect 38746 11840 38752 11852
rect 38804 11840 38810 11892
rect 39298 11880 39304 11892
rect 39259 11852 39304 11880
rect 39298 11840 39304 11852
rect 39356 11840 39362 11892
rect 40310 11880 40316 11892
rect 40271 11852 40316 11880
rect 40310 11840 40316 11852
rect 40368 11840 40374 11892
rect 40770 11840 40776 11892
rect 40828 11880 40834 11892
rect 40865 11883 40923 11889
rect 40865 11880 40877 11883
rect 40828 11852 40877 11880
rect 40828 11840 40834 11852
rect 40865 11849 40877 11852
rect 40911 11849 40923 11883
rect 41414 11880 41420 11892
rect 41375 11852 41420 11880
rect 40865 11843 40923 11849
rect 41414 11840 41420 11852
rect 41472 11840 41478 11892
rect 42521 11883 42579 11889
rect 42521 11849 42533 11883
rect 42567 11880 42579 11883
rect 42702 11880 42708 11892
rect 42567 11852 42708 11880
rect 42567 11849 42579 11852
rect 42521 11843 42579 11849
rect 42702 11840 42708 11852
rect 42760 11880 42766 11892
rect 44358 11880 44364 11892
rect 42760 11852 44364 11880
rect 42760 11840 42766 11852
rect 44358 11840 44364 11852
rect 44416 11840 44422 11892
rect 36814 11812 36820 11824
rect 36096 11784 36820 11812
rect 36814 11772 36820 11784
rect 36872 11772 36878 11824
rect 37366 11812 37372 11824
rect 36924 11784 37372 11812
rect 36722 11744 36728 11756
rect 36004 11716 36728 11744
rect 35897 11707 35955 11713
rect 31220 11648 34284 11676
rect 26418 11608 26424 11620
rect 24912 11580 26004 11608
rect 26379 11580 26424 11608
rect 24912 11568 24918 11580
rect 26418 11568 26424 11580
rect 26476 11568 26482 11620
rect 27890 11568 27896 11620
rect 27948 11608 27954 11620
rect 28350 11608 28356 11620
rect 27948 11580 28356 11608
rect 27948 11568 27954 11580
rect 28350 11568 28356 11580
rect 28408 11568 28414 11620
rect 28902 11568 28908 11620
rect 28960 11608 28966 11620
rect 34256 11608 34284 11648
rect 34330 11636 34336 11688
rect 34388 11676 34394 11688
rect 35710 11676 35716 11688
rect 34388 11648 34433 11676
rect 35671 11648 35716 11676
rect 34388 11636 34394 11648
rect 35710 11636 35716 11648
rect 35768 11636 35774 11688
rect 35912 11676 35940 11707
rect 36722 11704 36728 11716
rect 36780 11704 36786 11756
rect 36924 11676 36952 11784
rect 37366 11772 37372 11784
rect 37424 11772 37430 11824
rect 43898 11812 43904 11824
rect 37476 11784 43904 11812
rect 37476 11753 37504 11784
rect 43898 11772 43904 11784
rect 43956 11772 43962 11824
rect 37277 11747 37335 11753
rect 37277 11713 37289 11747
rect 37323 11713 37335 11747
rect 37277 11707 37335 11713
rect 37461 11747 37519 11753
rect 37461 11713 37473 11747
rect 37507 11713 37519 11747
rect 37461 11707 37519 11713
rect 38105 11747 38163 11753
rect 38105 11713 38117 11747
rect 38151 11713 38163 11747
rect 38105 11707 38163 11713
rect 35912 11648 36952 11676
rect 37292 11676 37320 11707
rect 38010 11676 38016 11688
rect 37292 11648 38016 11676
rect 38010 11636 38016 11648
rect 38068 11636 38074 11688
rect 36906 11608 36912 11620
rect 28960 11580 29408 11608
rect 28960 11568 28966 11580
rect 14734 11500 14740 11552
rect 14792 11540 14798 11552
rect 18601 11543 18659 11549
rect 18601 11540 18613 11543
rect 14792 11512 18613 11540
rect 14792 11500 14798 11512
rect 18601 11509 18613 11512
rect 18647 11540 18659 11543
rect 19058 11540 19064 11552
rect 18647 11512 19064 11540
rect 18647 11509 18659 11512
rect 18601 11503 18659 11509
rect 19058 11500 19064 11512
rect 19116 11500 19122 11552
rect 19245 11543 19303 11549
rect 19245 11509 19257 11543
rect 19291 11540 19303 11543
rect 19518 11540 19524 11552
rect 19291 11512 19524 11540
rect 19291 11509 19303 11512
rect 19245 11503 19303 11509
rect 19518 11500 19524 11512
rect 19576 11500 19582 11552
rect 20990 11540 20996 11552
rect 20951 11512 20996 11540
rect 20990 11500 20996 11512
rect 21048 11500 21054 11552
rect 24210 11540 24216 11552
rect 24171 11512 24216 11540
rect 24210 11500 24216 11512
rect 24268 11500 24274 11552
rect 25409 11543 25467 11549
rect 25409 11509 25421 11543
rect 25455 11540 25467 11543
rect 26234 11540 26240 11552
rect 25455 11512 26240 11540
rect 25455 11509 25467 11512
rect 25409 11503 25467 11509
rect 26234 11500 26240 11512
rect 26292 11500 26298 11552
rect 26326 11500 26332 11552
rect 26384 11540 26390 11552
rect 28166 11540 28172 11552
rect 26384 11512 28172 11540
rect 26384 11500 26390 11512
rect 28166 11500 28172 11512
rect 28224 11500 28230 11552
rect 29270 11540 29276 11552
rect 29231 11512 29276 11540
rect 29270 11500 29276 11512
rect 29328 11500 29334 11552
rect 29380 11540 29408 11580
rect 31128 11580 31708 11608
rect 31128 11540 31156 11580
rect 31570 11540 31576 11552
rect 29380 11512 31156 11540
rect 31531 11512 31576 11540
rect 31570 11500 31576 11512
rect 31628 11500 31634 11552
rect 31680 11540 31708 11580
rect 33704 11580 34100 11608
rect 34256 11580 36912 11608
rect 33134 11540 33140 11552
rect 31680 11512 33140 11540
rect 33134 11500 33140 11512
rect 33192 11540 33198 11552
rect 33704 11540 33732 11580
rect 33192 11512 33732 11540
rect 33192 11500 33198 11512
rect 33778 11500 33784 11552
rect 33836 11540 33842 11552
rect 33873 11543 33931 11549
rect 33873 11540 33885 11543
rect 33836 11512 33885 11540
rect 33836 11500 33842 11512
rect 33873 11509 33885 11512
rect 33919 11540 33931 11543
rect 33962 11540 33968 11552
rect 33919 11512 33968 11540
rect 33919 11509 33931 11512
rect 33873 11503 33931 11509
rect 33962 11500 33968 11512
rect 34020 11500 34026 11552
rect 34072 11540 34100 11580
rect 36906 11568 36912 11580
rect 36964 11568 36970 11620
rect 38120 11608 38148 11707
rect 38194 11704 38200 11756
rect 38252 11744 38258 11756
rect 38746 11744 38752 11756
rect 38252 11716 38752 11744
rect 38252 11704 38258 11716
rect 38746 11704 38752 11716
rect 38804 11744 38810 11756
rect 41046 11744 41052 11756
rect 38804 11716 41052 11744
rect 38804 11704 38810 11716
rect 41046 11704 41052 11716
rect 41104 11744 41110 11756
rect 42981 11747 43039 11753
rect 42981 11744 42993 11747
rect 41104 11716 42993 11744
rect 41104 11704 41110 11716
rect 42981 11713 42993 11716
rect 43027 11713 43039 11747
rect 43530 11744 43536 11756
rect 43491 11716 43536 11744
rect 42981 11707 43039 11713
rect 38378 11636 38384 11688
rect 38436 11676 38442 11688
rect 42150 11676 42156 11688
rect 38436 11648 42156 11676
rect 38436 11636 38442 11648
rect 42150 11636 42156 11648
rect 42208 11636 42214 11688
rect 42996 11676 43024 11707
rect 43530 11704 43536 11716
rect 43588 11704 43594 11756
rect 44634 11676 44640 11688
rect 42996 11648 44640 11676
rect 44634 11636 44640 11648
rect 44692 11636 44698 11688
rect 38562 11608 38568 11620
rect 37292 11580 37780 11608
rect 38120 11580 38568 11608
rect 35621 11543 35679 11549
rect 35621 11540 35633 11543
rect 34072 11512 35633 11540
rect 35621 11509 35633 11512
rect 35667 11540 35679 11543
rect 37292 11540 37320 11580
rect 35667 11512 37320 11540
rect 37369 11543 37427 11549
rect 35667 11509 35679 11512
rect 35621 11503 35679 11509
rect 37369 11509 37381 11543
rect 37415 11540 37427 11543
rect 37642 11540 37648 11552
rect 37415 11512 37648 11540
rect 37415 11509 37427 11512
rect 37369 11503 37427 11509
rect 37642 11500 37648 11512
rect 37700 11500 37706 11552
rect 37752 11540 37780 11580
rect 38562 11568 38568 11580
rect 38620 11608 38626 11620
rect 38838 11608 38844 11620
rect 38620 11580 38844 11608
rect 38620 11568 38626 11580
rect 38838 11568 38844 11580
rect 38896 11568 38902 11620
rect 39853 11611 39911 11617
rect 39853 11577 39865 11611
rect 39899 11608 39911 11611
rect 42610 11608 42616 11620
rect 39899 11580 42616 11608
rect 39899 11577 39911 11580
rect 39853 11571 39911 11577
rect 39868 11540 39896 11571
rect 42610 11568 42616 11580
rect 42668 11568 42674 11620
rect 37752 11512 39896 11540
rect 1104 11450 58880 11472
rect 1104 11398 10582 11450
rect 10634 11398 10646 11450
rect 10698 11398 10710 11450
rect 10762 11398 10774 11450
rect 10826 11398 10838 11450
rect 10890 11398 29846 11450
rect 29898 11398 29910 11450
rect 29962 11398 29974 11450
rect 30026 11398 30038 11450
rect 30090 11398 30102 11450
rect 30154 11398 49110 11450
rect 49162 11398 49174 11450
rect 49226 11398 49238 11450
rect 49290 11398 49302 11450
rect 49354 11398 49366 11450
rect 49418 11398 58880 11450
rect 1104 11376 58880 11398
rect 19058 11296 19064 11348
rect 19116 11336 19122 11348
rect 19702 11336 19708 11348
rect 19116 11308 19708 11336
rect 19116 11296 19122 11308
rect 19702 11296 19708 11308
rect 19760 11296 19766 11348
rect 19889 11339 19947 11345
rect 19889 11305 19901 11339
rect 19935 11336 19947 11339
rect 21174 11336 21180 11348
rect 19935 11308 21180 11336
rect 19935 11305 19947 11308
rect 19889 11299 19947 11305
rect 21174 11296 21180 11308
rect 21232 11296 21238 11348
rect 21542 11336 21548 11348
rect 21503 11308 21548 11336
rect 21542 11296 21548 11308
rect 21600 11296 21606 11348
rect 22189 11339 22247 11345
rect 22189 11305 22201 11339
rect 22235 11336 22247 11339
rect 22741 11339 22799 11345
rect 22741 11336 22753 11339
rect 22235 11308 22753 11336
rect 22235 11305 22247 11308
rect 22189 11299 22247 11305
rect 22741 11305 22753 11308
rect 22787 11336 22799 11339
rect 22830 11336 22836 11348
rect 22787 11308 22836 11336
rect 22787 11305 22799 11308
rect 22741 11299 22799 11305
rect 22830 11296 22836 11308
rect 22888 11296 22894 11348
rect 23845 11339 23903 11345
rect 23845 11305 23857 11339
rect 23891 11336 23903 11339
rect 23934 11336 23940 11348
rect 23891 11308 23940 11336
rect 23891 11305 23903 11308
rect 23845 11299 23903 11305
rect 23934 11296 23940 11308
rect 23992 11296 23998 11348
rect 24302 11296 24308 11348
rect 24360 11336 24366 11348
rect 25590 11336 25596 11348
rect 24360 11308 24973 11336
rect 25551 11308 25596 11336
rect 24360 11296 24366 11308
rect 20438 11268 20444 11280
rect 20399 11240 20444 11268
rect 20438 11228 20444 11240
rect 20496 11228 20502 11280
rect 20622 11228 20628 11280
rect 20680 11268 20686 11280
rect 24026 11268 24032 11280
rect 20680 11240 24032 11268
rect 20680 11228 20686 11240
rect 24026 11228 24032 11240
rect 24084 11228 24090 11280
rect 24945 11268 24973 11308
rect 25590 11296 25596 11308
rect 25648 11296 25654 11348
rect 25866 11296 25872 11348
rect 25924 11336 25930 11348
rect 27249 11339 27307 11345
rect 27249 11336 27261 11339
rect 25924 11308 27261 11336
rect 25924 11296 25930 11308
rect 27249 11305 27261 11308
rect 27295 11305 27307 11339
rect 27249 11299 27307 11305
rect 27338 11296 27344 11348
rect 27396 11336 27402 11348
rect 27433 11339 27491 11345
rect 27433 11336 27445 11339
rect 27396 11308 27445 11336
rect 27396 11296 27402 11308
rect 27433 11305 27445 11308
rect 27479 11336 27491 11339
rect 27522 11336 27528 11348
rect 27479 11308 27528 11336
rect 27479 11305 27491 11308
rect 27433 11299 27491 11305
rect 27522 11296 27528 11308
rect 27580 11296 27586 11348
rect 28813 11339 28871 11345
rect 28813 11336 28825 11339
rect 28368 11308 28825 11336
rect 26786 11268 26792 11280
rect 24945 11240 26464 11268
rect 26747 11240 26792 11268
rect 23566 11160 23572 11212
rect 23624 11200 23630 11212
rect 26326 11200 26332 11212
rect 23624 11172 25728 11200
rect 26287 11172 26332 11200
rect 23624 11160 23630 11172
rect 19334 11132 19340 11144
rect 19295 11104 19340 11132
rect 19334 11092 19340 11104
rect 19392 11092 19398 11144
rect 20898 11092 20904 11144
rect 20956 11132 20962 11144
rect 23293 11135 23351 11141
rect 23293 11132 23305 11135
rect 20956 11104 23305 11132
rect 20956 11092 20962 11104
rect 23293 11101 23305 11104
rect 23339 11132 23351 11135
rect 24670 11132 24676 11144
rect 23339 11104 24676 11132
rect 23339 11101 23351 11104
rect 23293 11095 23351 11101
rect 24670 11092 24676 11104
rect 24728 11092 24734 11144
rect 25038 11132 25044 11144
rect 24999 11104 25044 11132
rect 25038 11092 25044 11104
rect 25096 11092 25102 11144
rect 25406 11092 25412 11144
rect 25464 11132 25470 11144
rect 25590 11132 25596 11144
rect 25464 11104 25596 11132
rect 25464 11092 25470 11104
rect 25590 11092 25596 11104
rect 25648 11092 25654 11144
rect 21085 11067 21143 11073
rect 21085 11033 21097 11067
rect 21131 11064 21143 11067
rect 22278 11064 22284 11076
rect 21131 11036 22284 11064
rect 21131 11033 21143 11036
rect 21085 11027 21143 11033
rect 22278 11024 22284 11036
rect 22336 11064 22342 11076
rect 23014 11064 23020 11076
rect 22336 11036 23020 11064
rect 22336 11024 22342 11036
rect 23014 11024 23020 11036
rect 23072 11024 23078 11076
rect 24026 11024 24032 11076
rect 24084 11064 24090 11076
rect 25700 11073 25728 11172
rect 26326 11160 26332 11172
rect 26384 11160 26390 11212
rect 26436 11200 26464 11240
rect 26786 11228 26792 11240
rect 26844 11228 26850 11280
rect 27798 11268 27804 11280
rect 27759 11240 27804 11268
rect 27798 11228 27804 11240
rect 27856 11268 27862 11280
rect 28261 11271 28319 11277
rect 28261 11268 28273 11271
rect 27856 11240 28273 11268
rect 27856 11228 27862 11240
rect 28261 11237 28273 11240
rect 28307 11237 28319 11271
rect 28261 11231 28319 11237
rect 27982 11200 27988 11212
rect 26436 11172 27988 11200
rect 27982 11160 27988 11172
rect 28040 11200 28046 11212
rect 28368 11200 28396 11308
rect 28813 11305 28825 11308
rect 28859 11305 28871 11339
rect 34790 11336 34796 11348
rect 28813 11299 28871 11305
rect 28966 11308 32352 11336
rect 34751 11308 34796 11336
rect 28966 11200 28994 11308
rect 32324 11268 32352 11308
rect 34790 11296 34796 11308
rect 34848 11296 34854 11348
rect 35805 11339 35863 11345
rect 35805 11305 35817 11339
rect 35851 11305 35863 11339
rect 35805 11299 35863 11305
rect 32766 11268 32772 11280
rect 32324 11240 32772 11268
rect 32766 11228 32772 11240
rect 32824 11268 32830 11280
rect 35710 11268 35716 11280
rect 32824 11240 35716 11268
rect 32824 11228 32830 11240
rect 35710 11228 35716 11240
rect 35768 11228 35774 11280
rect 35820 11268 35848 11299
rect 36446 11296 36452 11348
rect 36504 11336 36510 11348
rect 36633 11339 36691 11345
rect 36633 11336 36645 11339
rect 36504 11308 36645 11336
rect 36504 11296 36510 11308
rect 36633 11305 36645 11308
rect 36679 11305 36691 11339
rect 36633 11299 36691 11305
rect 36722 11296 36728 11348
rect 36780 11336 36786 11348
rect 36780 11308 37136 11336
rect 36780 11296 36786 11308
rect 36998 11268 37004 11280
rect 35820 11240 37004 11268
rect 36998 11228 37004 11240
rect 37056 11228 37062 11280
rect 37108 11268 37136 11308
rect 37826 11296 37832 11348
rect 37884 11336 37890 11348
rect 38289 11339 38347 11345
rect 38289 11336 38301 11339
rect 37884 11308 38301 11336
rect 37884 11296 37890 11308
rect 38289 11305 38301 11308
rect 38335 11305 38347 11339
rect 38838 11336 38844 11348
rect 38799 11308 38844 11336
rect 38289 11299 38347 11305
rect 38838 11296 38844 11308
rect 38896 11296 38902 11348
rect 39850 11336 39856 11348
rect 39811 11308 39856 11336
rect 39850 11296 39856 11308
rect 39908 11296 39914 11348
rect 41230 11296 41236 11348
rect 41288 11336 41294 11348
rect 42702 11336 42708 11348
rect 41288 11308 42708 11336
rect 41288 11296 41294 11308
rect 42702 11296 42708 11308
rect 42760 11296 42766 11348
rect 37737 11271 37795 11277
rect 37737 11268 37749 11271
rect 37108 11240 37749 11268
rect 37737 11237 37749 11240
rect 37783 11268 37795 11271
rect 37783 11240 38654 11268
rect 37783 11237 37795 11240
rect 37737 11231 37795 11237
rect 30282 11200 30288 11212
rect 28040 11172 28396 11200
rect 28736 11172 28994 11200
rect 30243 11172 30288 11200
rect 28040 11160 28046 11172
rect 28736 11144 28764 11172
rect 30282 11160 30288 11172
rect 30340 11160 30346 11212
rect 30561 11203 30619 11209
rect 30561 11169 30573 11203
rect 30607 11200 30619 11203
rect 31386 11200 31392 11212
rect 30607 11172 31392 11200
rect 30607 11169 30619 11172
rect 30561 11163 30619 11169
rect 31386 11160 31392 11172
rect 31444 11160 31450 11212
rect 31662 11160 31668 11212
rect 31720 11200 31726 11212
rect 34054 11200 34060 11212
rect 31720 11172 34060 11200
rect 31720 11160 31726 11172
rect 34054 11160 34060 11172
rect 34112 11160 34118 11212
rect 34149 11203 34207 11209
rect 34149 11169 34161 11203
rect 34195 11200 34207 11203
rect 34238 11200 34244 11212
rect 34195 11172 34244 11200
rect 34195 11169 34207 11172
rect 34149 11163 34207 11169
rect 34238 11160 34244 11172
rect 34296 11200 34302 11212
rect 34790 11200 34796 11212
rect 34296 11172 34796 11200
rect 34296 11160 34302 11172
rect 34790 11160 34796 11172
rect 34848 11160 34854 11212
rect 35158 11200 35164 11212
rect 35119 11172 35164 11200
rect 35158 11160 35164 11172
rect 35216 11160 35222 11212
rect 35618 11160 35624 11212
rect 35676 11200 35682 11212
rect 36078 11200 36084 11212
rect 35676 11172 36084 11200
rect 35676 11160 35682 11172
rect 36078 11160 36084 11172
rect 36136 11160 36142 11212
rect 38626 11200 38654 11240
rect 39390 11200 39396 11212
rect 38626 11172 39396 11200
rect 39390 11160 39396 11172
rect 39448 11160 39454 11212
rect 41506 11200 41512 11212
rect 41467 11172 41512 11200
rect 41506 11160 41512 11172
rect 41564 11160 41570 11212
rect 26421 11135 26479 11141
rect 26421 11101 26433 11135
rect 26467 11132 26479 11135
rect 26786 11132 26792 11144
rect 26467 11104 26792 11132
rect 26467 11101 26479 11104
rect 26421 11095 26479 11101
rect 26786 11092 26792 11104
rect 26844 11092 26850 11144
rect 27614 11092 27620 11144
rect 27672 11132 27678 11144
rect 28537 11135 28595 11141
rect 28537 11132 28549 11135
rect 27672 11104 28549 11132
rect 27672 11092 27678 11104
rect 28537 11101 28549 11104
rect 28583 11101 28595 11135
rect 28537 11095 28595 11101
rect 28629 11135 28687 11141
rect 28629 11101 28641 11135
rect 28675 11101 28687 11135
rect 28629 11095 28687 11101
rect 24949 11067 25007 11073
rect 24949 11064 24961 11067
rect 24084 11036 24961 11064
rect 24084 11024 24090 11036
rect 24949 11033 24961 11036
rect 24995 11033 25007 11067
rect 24949 11027 25007 11033
rect 25685 11067 25743 11073
rect 25685 11033 25697 11067
rect 25731 11064 25743 11067
rect 26142 11064 26148 11076
rect 25731 11036 26148 11064
rect 25731 11033 25743 11036
rect 25685 11027 25743 11033
rect 26142 11024 26148 11036
rect 26200 11024 26206 11076
rect 26970 11024 26976 11076
rect 27028 11064 27034 11076
rect 27433 11067 27491 11073
rect 27433 11064 27445 11067
rect 27028 11036 27445 11064
rect 27028 11024 27034 11036
rect 27433 11033 27445 11036
rect 27479 11033 27491 11067
rect 27433 11027 27491 11033
rect 27890 11024 27896 11076
rect 27948 11064 27954 11076
rect 28644 11064 28672 11095
rect 28718 11092 28724 11144
rect 28776 11132 28782 11144
rect 28997 11135 29055 11141
rect 28776 11104 28821 11132
rect 28776 11092 28782 11104
rect 28997 11101 29009 11135
rect 29043 11132 29055 11135
rect 29270 11132 29276 11144
rect 29043 11104 29276 11132
rect 29043 11101 29055 11104
rect 28997 11095 29055 11101
rect 29270 11092 29276 11104
rect 29328 11092 29334 11144
rect 31018 11132 31024 11144
rect 30979 11104 31024 11132
rect 31018 11092 31024 11104
rect 31076 11092 31082 11144
rect 33778 11092 33784 11144
rect 33836 11132 33842 11144
rect 33873 11135 33931 11141
rect 33873 11132 33885 11135
rect 33836 11104 33885 11132
rect 33836 11092 33842 11104
rect 33873 11101 33885 11104
rect 33919 11101 33931 11135
rect 33873 11095 33931 11101
rect 33962 11092 33968 11144
rect 34020 11092 34026 11144
rect 34698 11132 34704 11144
rect 34659 11104 34704 11132
rect 34698 11092 34704 11104
rect 34756 11092 34762 11144
rect 34977 11135 35035 11141
rect 34977 11101 34989 11135
rect 35023 11132 35035 11135
rect 35250 11132 35256 11144
rect 35023 11104 35256 11132
rect 35023 11101 35035 11104
rect 34977 11095 35035 11101
rect 35250 11092 35256 11104
rect 35308 11132 35314 11144
rect 35434 11132 35440 11144
rect 35308 11104 35440 11132
rect 35308 11092 35314 11104
rect 35434 11092 35440 11104
rect 35492 11092 35498 11144
rect 35710 11092 35716 11144
rect 35768 11132 35774 11144
rect 35768 11104 36124 11132
rect 35768 11092 35774 11104
rect 27948 11036 28672 11064
rect 28966 11036 31156 11064
rect 27948 11024 27954 11036
rect 17034 10956 17040 11008
rect 17092 10996 17098 11008
rect 23474 10996 23480 11008
rect 17092 10968 23480 10996
rect 17092 10956 17098 10968
rect 23474 10956 23480 10968
rect 23532 10956 23538 11008
rect 25774 10956 25780 11008
rect 25832 10996 25838 11008
rect 28966 10996 28994 11036
rect 25832 10968 28994 10996
rect 25832 10956 25838 10968
rect 30374 10956 30380 11008
rect 30432 10996 30438 11008
rect 30558 10996 30564 11008
rect 30432 10968 30564 10996
rect 30432 10956 30438 10968
rect 30558 10956 30564 10968
rect 30616 10956 30622 11008
rect 31128 10996 31156 11036
rect 31202 11024 31208 11076
rect 31260 11064 31266 11076
rect 31297 11067 31355 11073
rect 31297 11064 31309 11067
rect 31260 11036 31309 11064
rect 31260 11024 31266 11036
rect 31297 11033 31309 11036
rect 31343 11033 31355 11067
rect 31297 11027 31355 11033
rect 31754 11024 31760 11076
rect 31812 11024 31818 11076
rect 33134 11064 33140 11076
rect 32784 11036 33140 11064
rect 31662 10996 31668 11008
rect 31128 10968 31668 10996
rect 31662 10956 31668 10968
rect 31720 10956 31726 11008
rect 32784 11005 32812 11036
rect 33134 11024 33140 11036
rect 33192 11024 33198 11076
rect 33502 11024 33508 11076
rect 33560 11064 33566 11076
rect 33980 11064 34008 11092
rect 35618 11064 35624 11076
rect 33560 11036 35624 11064
rect 33560 11024 33566 11036
rect 35618 11024 35624 11036
rect 35676 11024 35682 11076
rect 32769 10999 32827 11005
rect 32769 10965 32781 10999
rect 32815 10965 32827 10999
rect 32769 10959 32827 10965
rect 33318 10956 33324 11008
rect 33376 10996 33382 11008
rect 33962 10996 33968 11008
rect 33376 10968 33968 10996
rect 33376 10956 33382 10968
rect 33962 10956 33968 10968
rect 34020 10956 34026 11008
rect 34146 10956 34152 11008
rect 34204 10996 34210 11008
rect 34514 10996 34520 11008
rect 34204 10968 34520 10996
rect 34204 10956 34210 10968
rect 34514 10956 34520 10968
rect 34572 10956 34578 11008
rect 34790 10956 34796 11008
rect 34848 10996 34854 11008
rect 35710 10996 35716 11008
rect 34848 10968 35716 10996
rect 34848 10956 34854 10968
rect 35710 10956 35716 10968
rect 35768 10956 35774 11008
rect 35802 10956 35808 11008
rect 35860 11005 35866 11008
rect 35860 10999 35879 11005
rect 35867 10965 35879 10999
rect 35986 10996 35992 11008
rect 35947 10968 35992 10996
rect 35860 10959 35879 10965
rect 35860 10956 35866 10959
rect 35986 10956 35992 10968
rect 36044 10956 36050 11008
rect 36096 10996 36124 11104
rect 36354 11092 36360 11144
rect 36412 11132 36418 11144
rect 36449 11135 36507 11141
rect 36449 11132 36461 11135
rect 36412 11104 36461 11132
rect 36412 11092 36418 11104
rect 36449 11101 36461 11104
rect 36495 11101 36507 11135
rect 36449 11095 36507 11101
rect 37285 11137 37343 11143
rect 37285 11103 37297 11137
rect 37331 11134 37343 11137
rect 37331 11106 37412 11134
rect 37331 11103 37343 11106
rect 37285 11097 37343 11103
rect 36906 11024 36912 11076
rect 36964 11064 36970 11076
rect 37185 11067 37243 11073
rect 37185 11064 37197 11067
rect 36964 11036 37197 11064
rect 36964 11024 36970 11036
rect 37185 11033 37197 11036
rect 37231 11033 37243 11067
rect 37384 11064 37412 11106
rect 37826 11092 37832 11144
rect 37884 11132 37890 11144
rect 40405 11135 40463 11141
rect 40405 11132 40417 11135
rect 37884 11104 40417 11132
rect 37884 11092 37890 11104
rect 40405 11101 40417 11104
rect 40451 11101 40463 11135
rect 40405 11095 40463 11101
rect 41049 11135 41107 11141
rect 41049 11101 41061 11135
rect 41095 11132 41107 11135
rect 46290 11132 46296 11144
rect 41095 11104 46296 11132
rect 41095 11101 41107 11104
rect 41049 11095 41107 11101
rect 46290 11092 46296 11104
rect 46348 11092 46354 11144
rect 58158 11132 58164 11144
rect 58119 11104 58164 11132
rect 58158 11092 58164 11104
rect 58216 11092 58222 11144
rect 37642 11064 37648 11076
rect 37384 11036 37648 11064
rect 37185 11027 37243 11033
rect 37642 11024 37648 11036
rect 37700 11024 37706 11076
rect 42061 11067 42119 11073
rect 42061 11064 42073 11067
rect 38626 11036 42073 11064
rect 38626 10996 38654 11036
rect 42061 11033 42073 11036
rect 42107 11033 42119 11067
rect 42061 11027 42119 11033
rect 42518 11024 42524 11076
rect 42576 11064 42582 11076
rect 57885 11067 57943 11073
rect 57885 11064 57897 11067
rect 42576 11036 57897 11064
rect 42576 11024 42582 11036
rect 57885 11033 57897 11036
rect 57931 11033 57943 11067
rect 57885 11027 57943 11033
rect 36096 10968 38654 10996
rect 1104 10906 58880 10928
rect 1104 10854 20214 10906
rect 20266 10854 20278 10906
rect 20330 10854 20342 10906
rect 20394 10854 20406 10906
rect 20458 10854 20470 10906
rect 20522 10854 39478 10906
rect 39530 10854 39542 10906
rect 39594 10854 39606 10906
rect 39658 10854 39670 10906
rect 39722 10854 39734 10906
rect 39786 10854 58880 10906
rect 1104 10832 58880 10854
rect 19978 10752 19984 10804
rect 20036 10792 20042 10804
rect 20717 10795 20775 10801
rect 20717 10792 20729 10795
rect 20036 10764 20729 10792
rect 20036 10752 20042 10764
rect 20717 10761 20729 10764
rect 20763 10761 20775 10795
rect 20717 10755 20775 10761
rect 21174 10752 21180 10804
rect 21232 10792 21238 10804
rect 21269 10795 21327 10801
rect 21269 10792 21281 10795
rect 21232 10764 21281 10792
rect 21232 10752 21238 10764
rect 21269 10761 21281 10764
rect 21315 10792 21327 10795
rect 21358 10792 21364 10804
rect 21315 10764 21364 10792
rect 21315 10761 21327 10764
rect 21269 10755 21327 10761
rect 21358 10752 21364 10764
rect 21416 10752 21422 10804
rect 22646 10792 22652 10804
rect 22607 10764 22652 10792
rect 22646 10752 22652 10764
rect 22704 10752 22710 10804
rect 23201 10795 23259 10801
rect 23201 10761 23213 10795
rect 23247 10792 23259 10795
rect 23750 10792 23756 10804
rect 23247 10764 23756 10792
rect 23247 10761 23259 10764
rect 23201 10755 23259 10761
rect 23750 10752 23756 10764
rect 23808 10792 23814 10804
rect 24762 10792 24768 10804
rect 23808 10764 24768 10792
rect 23808 10752 23814 10764
rect 24762 10752 24768 10764
rect 24820 10752 24826 10804
rect 28905 10795 28963 10801
rect 28905 10792 28917 10795
rect 25608 10764 28917 10792
rect 24302 10724 24308 10736
rect 24263 10696 24308 10724
rect 24302 10684 24308 10696
rect 24360 10684 24366 10736
rect 25608 10733 25636 10764
rect 28905 10761 28917 10764
rect 28951 10792 28963 10795
rect 34514 10792 34520 10804
rect 28951 10764 34520 10792
rect 28951 10761 28963 10764
rect 28905 10755 28963 10761
rect 34514 10752 34520 10764
rect 34572 10752 34578 10804
rect 36262 10792 36268 10804
rect 34884 10764 36124 10792
rect 36223 10764 36268 10792
rect 25593 10727 25651 10733
rect 25593 10693 25605 10727
rect 25639 10693 25651 10727
rect 25593 10687 25651 10693
rect 26786 10684 26792 10736
rect 26844 10724 26850 10736
rect 31294 10724 31300 10736
rect 26844 10696 31202 10724
rect 31255 10696 31300 10724
rect 26844 10684 26850 10696
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 11054 10656 11060 10668
rect 1719 10628 11060 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 11054 10616 11060 10628
rect 11112 10616 11118 10668
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10656 11759 10659
rect 11747 10628 12296 10656
rect 11747 10625 11759 10628
rect 11701 10619 11759 10625
rect 12268 10597 12296 10628
rect 23474 10616 23480 10668
rect 23532 10656 23538 10668
rect 24210 10656 24216 10668
rect 23532 10628 24216 10656
rect 23532 10616 23538 10628
rect 24210 10616 24216 10628
rect 24268 10656 24274 10668
rect 24765 10659 24823 10665
rect 24765 10656 24777 10659
rect 24268 10628 24777 10656
rect 24268 10616 24274 10628
rect 24765 10625 24777 10628
rect 24811 10625 24823 10659
rect 24946 10656 24952 10668
rect 24907 10628 24952 10656
rect 24765 10619 24823 10625
rect 24946 10616 24952 10628
rect 25004 10616 25010 10668
rect 25774 10656 25780 10668
rect 25240 10628 25780 10656
rect 12253 10591 12311 10597
rect 12253 10557 12265 10591
rect 12299 10588 12311 10591
rect 14918 10588 14924 10600
rect 12299 10560 14924 10588
rect 12299 10557 12311 10560
rect 12253 10551 12311 10557
rect 14918 10548 14924 10560
rect 14976 10588 14982 10600
rect 23382 10588 23388 10600
rect 14976 10560 23388 10588
rect 14976 10548 14982 10560
rect 23382 10548 23388 10560
rect 23440 10548 23446 10600
rect 25240 10588 25268 10628
rect 25774 10616 25780 10628
rect 25832 10616 25838 10668
rect 26142 10616 26148 10668
rect 26200 10656 26206 10668
rect 26329 10659 26387 10665
rect 26329 10656 26341 10659
rect 26200 10628 26341 10656
rect 26200 10616 26206 10628
rect 26329 10625 26341 10628
rect 26375 10625 26387 10659
rect 26329 10619 26387 10625
rect 26694 10616 26700 10668
rect 26752 10656 26758 10668
rect 27617 10659 27675 10665
rect 27617 10656 27629 10659
rect 26752 10628 27629 10656
rect 26752 10616 26758 10628
rect 27617 10625 27629 10628
rect 27663 10656 27675 10659
rect 30193 10659 30251 10665
rect 27663 10628 28672 10656
rect 27663 10625 27675 10628
rect 27617 10619 27675 10625
rect 25406 10588 25412 10600
rect 24412 10560 25268 10588
rect 25319 10560 25412 10588
rect 22097 10523 22155 10529
rect 22097 10489 22109 10523
rect 22143 10520 22155 10523
rect 24412 10520 24440 10560
rect 25406 10548 25412 10560
rect 25464 10588 25470 10600
rect 27246 10588 27252 10600
rect 25464 10560 27252 10588
rect 25464 10548 25470 10560
rect 27246 10548 27252 10560
rect 27304 10548 27310 10600
rect 27706 10588 27712 10600
rect 27667 10560 27712 10588
rect 27706 10548 27712 10560
rect 27764 10548 27770 10600
rect 28644 10588 28672 10628
rect 30193 10625 30205 10659
rect 30239 10656 30251 10659
rect 30282 10656 30288 10668
rect 30239 10628 30288 10656
rect 30239 10625 30251 10628
rect 30193 10619 30251 10625
rect 30282 10616 30288 10628
rect 30340 10616 30346 10668
rect 31174 10656 31202 10696
rect 31294 10684 31300 10696
rect 31352 10684 31358 10736
rect 31386 10684 31392 10736
rect 31444 10724 31450 10736
rect 31444 10696 33272 10724
rect 31444 10684 31450 10696
rect 31478 10656 31484 10668
rect 31174 10628 31484 10656
rect 31478 10616 31484 10628
rect 31536 10616 31542 10668
rect 31573 10659 31631 10665
rect 31573 10625 31585 10659
rect 31619 10656 31631 10659
rect 32401 10659 32459 10665
rect 31619 10628 32168 10656
rect 31619 10625 31631 10628
rect 31573 10619 31631 10625
rect 32030 10588 32036 10600
rect 28644 10560 32036 10588
rect 32030 10548 32036 10560
rect 32088 10548 32094 10600
rect 32140 10597 32168 10628
rect 32401 10625 32413 10659
rect 32447 10656 32459 10659
rect 32490 10656 32496 10668
rect 32447 10628 32496 10656
rect 32447 10625 32459 10628
rect 32401 10619 32459 10625
rect 32490 10616 32496 10628
rect 32548 10616 32554 10668
rect 33045 10659 33103 10665
rect 33045 10625 33057 10659
rect 33091 10625 33103 10659
rect 33244 10656 33272 10696
rect 33318 10684 33324 10736
rect 33376 10724 33382 10736
rect 33686 10724 33692 10736
rect 33376 10696 33692 10724
rect 33376 10684 33382 10696
rect 33686 10684 33692 10696
rect 33744 10684 33750 10736
rect 34884 10699 34912 10764
rect 34839 10693 34912 10699
rect 34839 10668 34851 10693
rect 33965 10659 34023 10665
rect 33965 10656 33977 10659
rect 33244 10628 33977 10656
rect 33045 10619 33103 10625
rect 33965 10625 33977 10628
rect 34011 10656 34023 10659
rect 34146 10656 34152 10668
rect 34011 10628 34152 10656
rect 34011 10625 34023 10628
rect 33965 10619 34023 10625
rect 32125 10591 32183 10597
rect 32125 10557 32137 10591
rect 32171 10557 32183 10591
rect 32125 10551 32183 10557
rect 22143 10492 24440 10520
rect 22143 10489 22155 10492
rect 22097 10483 22155 10489
rect 24762 10480 24768 10532
rect 24820 10520 24826 10532
rect 26145 10523 26203 10529
rect 26145 10520 26157 10523
rect 24820 10492 26157 10520
rect 24820 10480 24826 10492
rect 26145 10489 26157 10492
rect 26191 10489 26203 10523
rect 27982 10520 27988 10532
rect 27943 10492 27988 10520
rect 26145 10483 26203 10489
rect 27982 10480 27988 10492
rect 28040 10480 28046 10532
rect 28350 10480 28356 10532
rect 28408 10520 28414 10532
rect 30374 10520 30380 10532
rect 28408 10492 30380 10520
rect 28408 10480 28414 10492
rect 30374 10480 30380 10492
rect 30432 10480 30438 10532
rect 30837 10523 30895 10529
rect 30837 10489 30849 10523
rect 30883 10520 30895 10523
rect 30883 10492 31754 10520
rect 30883 10489 30895 10492
rect 30837 10483 30895 10489
rect 1486 10452 1492 10464
rect 1447 10424 1492 10452
rect 1486 10412 1492 10424
rect 1544 10412 1550 10464
rect 11514 10452 11520 10464
rect 11475 10424 11520 10452
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 20070 10412 20076 10464
rect 20128 10452 20134 10464
rect 20165 10455 20223 10461
rect 20165 10452 20177 10455
rect 20128 10424 20177 10452
rect 20128 10412 20134 10424
rect 20165 10421 20177 10424
rect 20211 10452 20223 10455
rect 20622 10452 20628 10464
rect 20211 10424 20628 10452
rect 20211 10421 20223 10424
rect 20165 10415 20223 10421
rect 20622 10412 20628 10424
rect 20680 10412 20686 10464
rect 24857 10455 24915 10461
rect 24857 10421 24869 10455
rect 24903 10452 24915 10455
rect 26326 10452 26332 10464
rect 24903 10424 26332 10452
rect 24903 10421 24915 10424
rect 24857 10415 24915 10421
rect 26326 10412 26332 10424
rect 26384 10412 26390 10464
rect 27338 10412 27344 10464
rect 27396 10452 27402 10464
rect 29546 10452 29552 10464
rect 27396 10424 29552 10452
rect 27396 10412 27402 10424
rect 29546 10412 29552 10424
rect 29604 10412 29610 10464
rect 31726 10452 31754 10492
rect 31938 10452 31944 10464
rect 31726 10424 31944 10452
rect 31938 10412 31944 10424
rect 31996 10452 32002 10464
rect 32140 10452 32168 10551
rect 33060 10520 33088 10619
rect 34146 10616 34152 10628
rect 34204 10616 34210 10668
rect 34238 10616 34244 10668
rect 34296 10656 34302 10668
rect 34296 10628 34341 10656
rect 34296 10616 34302 10628
rect 34790 10616 34796 10668
rect 34848 10659 34851 10668
rect 34885 10659 34912 10693
rect 35069 10727 35127 10733
rect 35069 10693 35081 10727
rect 35115 10724 35127 10727
rect 35158 10724 35164 10736
rect 35115 10696 35164 10724
rect 35115 10693 35127 10696
rect 35069 10687 35127 10693
rect 35158 10684 35164 10696
rect 35216 10684 35222 10736
rect 36096 10724 36124 10764
rect 36262 10752 36268 10764
rect 36320 10752 36326 10804
rect 36446 10752 36452 10804
rect 36504 10792 36510 10804
rect 37829 10795 37887 10801
rect 37829 10792 37841 10795
rect 36504 10764 37841 10792
rect 36504 10752 36510 10764
rect 37829 10761 37841 10764
rect 37875 10761 37887 10795
rect 37829 10755 37887 10761
rect 40681 10795 40739 10801
rect 40681 10761 40693 10795
rect 40727 10792 40739 10795
rect 41230 10792 41236 10804
rect 40727 10764 41236 10792
rect 40727 10761 40739 10764
rect 40681 10755 40739 10761
rect 41230 10752 41236 10764
rect 41288 10752 41294 10804
rect 41690 10752 41696 10804
rect 41748 10792 41754 10804
rect 41785 10795 41843 10801
rect 41785 10792 41797 10795
rect 41748 10764 41797 10792
rect 41748 10752 41754 10764
rect 41785 10761 41797 10764
rect 41831 10792 41843 10795
rect 43530 10792 43536 10804
rect 41831 10764 43536 10792
rect 41831 10761 41843 10764
rect 41785 10755 41843 10761
rect 43530 10752 43536 10764
rect 43588 10752 43594 10804
rect 58158 10792 58164 10804
rect 58119 10764 58164 10792
rect 58158 10752 58164 10764
rect 58216 10752 58222 10804
rect 36096 10696 36492 10724
rect 34848 10628 34912 10659
rect 35713 10659 35771 10665
rect 34848 10616 34854 10628
rect 35713 10625 35725 10659
rect 35759 10656 35771 10659
rect 35802 10656 35808 10668
rect 35759 10628 35808 10656
rect 35759 10625 35771 10628
rect 35713 10619 35771 10625
rect 35802 10616 35808 10628
rect 35860 10616 35866 10668
rect 36262 10616 36268 10668
rect 36320 10656 36326 10668
rect 36357 10659 36415 10665
rect 36357 10656 36369 10659
rect 36320 10628 36369 10656
rect 36320 10616 36326 10628
rect 36357 10625 36369 10628
rect 36403 10625 36415 10659
rect 36464 10656 36492 10696
rect 36998 10684 37004 10736
rect 37056 10724 37062 10736
rect 37274 10724 37280 10736
rect 37056 10696 37280 10724
rect 37056 10684 37062 10696
rect 37274 10684 37280 10696
rect 37332 10684 37338 10736
rect 37366 10684 37372 10736
rect 37424 10724 37430 10736
rect 38378 10724 38384 10736
rect 37424 10696 38384 10724
rect 37424 10684 37430 10696
rect 38378 10684 38384 10696
rect 38436 10684 38442 10736
rect 38562 10684 38568 10736
rect 38620 10724 38626 10736
rect 40129 10727 40187 10733
rect 40129 10724 40141 10727
rect 38620 10696 40141 10724
rect 38620 10684 38626 10696
rect 40129 10693 40141 10696
rect 40175 10724 40187 10727
rect 41138 10724 41144 10736
rect 40175 10696 41144 10724
rect 40175 10693 40187 10696
rect 40129 10687 40187 10693
rect 41138 10684 41144 10696
rect 41196 10684 41202 10736
rect 38933 10659 38991 10665
rect 38933 10656 38945 10659
rect 36464 10628 38945 10656
rect 36357 10619 36415 10625
rect 38933 10625 38945 10628
rect 38979 10625 38991 10659
rect 38933 10619 38991 10625
rect 33134 10548 33140 10600
rect 33192 10588 33198 10600
rect 34057 10591 34115 10597
rect 34057 10588 34069 10591
rect 33192 10560 34069 10588
rect 33192 10548 33198 10560
rect 34057 10557 34069 10560
rect 34103 10588 34115 10591
rect 37277 10591 37335 10597
rect 37277 10588 37289 10591
rect 34103 10560 37289 10588
rect 34103 10557 34115 10560
rect 34057 10551 34115 10557
rect 37277 10557 37289 10560
rect 37323 10557 37335 10591
rect 37277 10551 37335 10557
rect 33686 10520 33692 10532
rect 33060 10492 33692 10520
rect 33686 10480 33692 10492
rect 33744 10480 33750 10532
rect 33778 10480 33784 10532
rect 33836 10520 33842 10532
rect 33836 10492 33881 10520
rect 33836 10480 33842 10492
rect 34146 10480 34152 10532
rect 34204 10520 34210 10532
rect 34701 10523 34759 10529
rect 34701 10520 34713 10523
rect 34204 10492 34713 10520
rect 34204 10480 34210 10492
rect 34701 10489 34713 10492
rect 34747 10489 34759 10523
rect 35526 10520 35532 10532
rect 35487 10492 35532 10520
rect 34701 10483 34759 10489
rect 35526 10480 35532 10492
rect 35584 10480 35590 10532
rect 33410 10452 33416 10464
rect 31996 10424 33416 10452
rect 31996 10412 32002 10424
rect 33410 10412 33416 10424
rect 33468 10412 33474 10464
rect 33962 10452 33968 10464
rect 33923 10424 33968 10452
rect 33962 10412 33968 10424
rect 34020 10412 34026 10464
rect 34606 10412 34612 10464
rect 34664 10452 34670 10464
rect 34885 10455 34943 10461
rect 34885 10452 34897 10455
rect 34664 10424 34897 10452
rect 34664 10412 34670 10424
rect 34885 10421 34897 10424
rect 34931 10421 34943 10455
rect 34885 10415 34943 10421
rect 35158 10412 35164 10464
rect 35216 10452 35222 10464
rect 35710 10452 35716 10464
rect 35216 10424 35716 10452
rect 35216 10412 35222 10424
rect 35710 10412 35716 10424
rect 35768 10412 35774 10464
rect 37274 10412 37280 10464
rect 37332 10452 37338 10464
rect 37918 10452 37924 10464
rect 37332 10424 37924 10452
rect 37332 10412 37338 10424
rect 37918 10412 37924 10424
rect 37976 10452 37982 10464
rect 39485 10455 39543 10461
rect 39485 10452 39497 10455
rect 37976 10424 39497 10452
rect 37976 10412 37982 10424
rect 39485 10421 39497 10424
rect 39531 10421 39543 10455
rect 39485 10415 39543 10421
rect 1104 10362 58880 10384
rect 1104 10310 10582 10362
rect 10634 10310 10646 10362
rect 10698 10310 10710 10362
rect 10762 10310 10774 10362
rect 10826 10310 10838 10362
rect 10890 10310 29846 10362
rect 29898 10310 29910 10362
rect 29962 10310 29974 10362
rect 30026 10310 30038 10362
rect 30090 10310 30102 10362
rect 30154 10310 49110 10362
rect 49162 10310 49174 10362
rect 49226 10310 49238 10362
rect 49290 10310 49302 10362
rect 49354 10310 49366 10362
rect 49418 10310 58880 10362
rect 1104 10288 58880 10310
rect 19702 10208 19708 10260
rect 19760 10248 19766 10260
rect 20993 10251 21051 10257
rect 20993 10248 21005 10251
rect 19760 10220 21005 10248
rect 19760 10208 19766 10220
rect 20993 10217 21005 10220
rect 21039 10248 21051 10251
rect 21545 10251 21603 10257
rect 21545 10248 21557 10251
rect 21039 10220 21557 10248
rect 21039 10217 21051 10220
rect 20993 10211 21051 10217
rect 21545 10217 21557 10220
rect 21591 10217 21603 10251
rect 21545 10211 21603 10217
rect 22189 10251 22247 10257
rect 22189 10217 22201 10251
rect 22235 10248 22247 10251
rect 23474 10248 23480 10260
rect 22235 10220 23480 10248
rect 22235 10217 22247 10220
rect 22189 10211 22247 10217
rect 21560 10180 21588 10211
rect 23474 10208 23480 10220
rect 23532 10208 23538 10260
rect 23750 10248 23756 10260
rect 23711 10220 23756 10248
rect 23750 10208 23756 10220
rect 23808 10208 23814 10260
rect 24578 10248 24584 10260
rect 24539 10220 24584 10248
rect 24578 10208 24584 10220
rect 24636 10208 24642 10260
rect 25222 10208 25228 10260
rect 25280 10248 25286 10260
rect 25866 10248 25872 10260
rect 25280 10220 25872 10248
rect 25280 10208 25286 10220
rect 25866 10208 25872 10220
rect 25924 10208 25930 10260
rect 26234 10248 26240 10260
rect 26195 10220 26240 10248
rect 26234 10208 26240 10220
rect 26292 10208 26298 10260
rect 27065 10251 27123 10257
rect 27065 10217 27077 10251
rect 27111 10248 27123 10251
rect 27430 10248 27436 10260
rect 27111 10220 27436 10248
rect 27111 10217 27123 10220
rect 27065 10211 27123 10217
rect 27430 10208 27436 10220
rect 27488 10208 27494 10260
rect 28442 10248 28448 10260
rect 28403 10220 28448 10248
rect 28442 10208 28448 10220
rect 28500 10208 28506 10260
rect 34698 10248 34704 10260
rect 29840 10220 34704 10248
rect 23290 10180 23296 10192
rect 21560 10152 23296 10180
rect 23290 10140 23296 10152
rect 23348 10140 23354 10192
rect 24486 10140 24492 10192
rect 24544 10180 24550 10192
rect 25317 10183 25375 10189
rect 25317 10180 25329 10183
rect 24544 10152 25329 10180
rect 24544 10140 24550 10152
rect 25317 10149 25329 10152
rect 25363 10180 25375 10183
rect 27706 10180 27712 10192
rect 25363 10152 27712 10180
rect 25363 10149 25375 10152
rect 25317 10143 25375 10149
rect 27706 10140 27712 10152
rect 27764 10140 27770 10192
rect 27798 10140 27804 10192
rect 27856 10180 27862 10192
rect 27985 10183 28043 10189
rect 27856 10152 27901 10180
rect 27856 10140 27862 10152
rect 27985 10149 27997 10183
rect 28031 10180 28043 10183
rect 29840 10180 29868 10220
rect 34698 10208 34704 10220
rect 34756 10208 34762 10260
rect 35710 10208 35716 10260
rect 35768 10248 35774 10260
rect 35768 10220 37274 10248
rect 35768 10208 35774 10220
rect 28031 10152 29868 10180
rect 28031 10149 28043 10152
rect 27985 10143 28043 10149
rect 34146 10140 34152 10192
rect 34204 10180 34210 10192
rect 34790 10180 34796 10192
rect 34204 10152 34796 10180
rect 34204 10140 34210 10152
rect 34790 10140 34796 10152
rect 34848 10140 34854 10192
rect 34977 10183 35035 10189
rect 34977 10149 34989 10183
rect 35023 10180 35035 10183
rect 36538 10180 36544 10192
rect 35023 10152 36544 10180
rect 35023 10149 35035 10152
rect 34977 10143 35035 10149
rect 36538 10140 36544 10152
rect 36596 10140 36602 10192
rect 37246 10180 37274 10220
rect 38286 10208 38292 10260
rect 38344 10248 38350 10260
rect 38381 10251 38439 10257
rect 38381 10248 38393 10251
rect 38344 10220 38393 10248
rect 38344 10208 38350 10220
rect 38381 10217 38393 10220
rect 38427 10217 38439 10251
rect 38381 10211 38439 10217
rect 39945 10251 40003 10257
rect 39945 10217 39957 10251
rect 39991 10248 40003 10251
rect 40034 10248 40040 10260
rect 39991 10220 40040 10248
rect 39991 10217 40003 10220
rect 39945 10211 40003 10217
rect 40034 10208 40040 10220
rect 40092 10208 40098 10260
rect 41046 10248 41052 10260
rect 41007 10220 41052 10248
rect 41046 10208 41052 10220
rect 41104 10208 41110 10260
rect 41966 10180 41972 10192
rect 37246 10152 41972 10180
rect 41966 10140 41972 10152
rect 42024 10140 42030 10192
rect 19794 10072 19800 10124
rect 19852 10112 19858 10124
rect 23201 10115 23259 10121
rect 23201 10112 23213 10115
rect 19852 10084 23213 10112
rect 19852 10072 19858 10084
rect 23201 10081 23213 10084
rect 23247 10081 23259 10115
rect 23201 10075 23259 10081
rect 23216 10044 23244 10075
rect 24394 10072 24400 10124
rect 24452 10112 24458 10124
rect 27617 10115 27675 10121
rect 24452 10084 27016 10112
rect 24452 10072 24458 10084
rect 25314 10044 25320 10056
rect 23216 10016 25320 10044
rect 25314 10004 25320 10016
rect 25372 10004 25378 10056
rect 25866 10004 25872 10056
rect 25924 10044 25930 10056
rect 26237 10047 26295 10053
rect 26237 10044 26249 10047
rect 25924 10016 26249 10044
rect 25924 10004 25930 10016
rect 26237 10013 26249 10016
rect 26283 10044 26295 10047
rect 26694 10044 26700 10056
rect 26283 10016 26700 10044
rect 26283 10013 26295 10016
rect 26237 10007 26295 10013
rect 26694 10004 26700 10016
rect 26752 10044 26758 10056
rect 26881 10047 26939 10053
rect 26881 10044 26893 10047
rect 26752 10016 26893 10044
rect 26752 10004 26758 10016
rect 26881 10013 26893 10016
rect 26927 10013 26939 10047
rect 26988 10044 27016 10084
rect 27617 10081 27629 10115
rect 27663 10112 27675 10115
rect 28074 10112 28080 10124
rect 27663 10084 28080 10112
rect 27663 10081 27675 10084
rect 27617 10075 27675 10081
rect 28074 10072 28080 10084
rect 28132 10072 28138 10124
rect 28534 10072 28540 10124
rect 28592 10112 28598 10124
rect 28721 10115 28779 10121
rect 28721 10112 28733 10115
rect 28592 10084 28733 10112
rect 28592 10072 28598 10084
rect 28721 10081 28733 10084
rect 28767 10112 28779 10115
rect 28902 10112 28908 10124
rect 28767 10084 28908 10112
rect 28767 10081 28779 10084
rect 28721 10075 28779 10081
rect 28902 10072 28908 10084
rect 28960 10072 28966 10124
rect 29546 10072 29552 10124
rect 29604 10112 29610 10124
rect 29733 10115 29791 10121
rect 29733 10112 29745 10115
rect 29604 10084 29745 10112
rect 29604 10072 29610 10084
rect 29733 10081 29745 10084
rect 29779 10081 29791 10115
rect 30006 10112 30012 10124
rect 29967 10084 30012 10112
rect 29733 10075 29791 10081
rect 30006 10072 30012 10084
rect 30064 10072 30070 10124
rect 30098 10072 30104 10124
rect 30156 10112 30162 10124
rect 30558 10112 30564 10124
rect 30156 10084 30564 10112
rect 30156 10072 30162 10084
rect 30558 10072 30564 10084
rect 30616 10072 30622 10124
rect 31938 10112 31944 10124
rect 31899 10084 31944 10112
rect 31938 10072 31944 10084
rect 31996 10072 32002 10124
rect 33318 10072 33324 10124
rect 33376 10112 33382 10124
rect 34238 10112 34244 10124
rect 33376 10084 34244 10112
rect 33376 10072 33382 10084
rect 34238 10072 34244 10084
rect 34296 10072 34302 10124
rect 34422 10072 34428 10124
rect 34480 10112 34486 10124
rect 36173 10115 36231 10121
rect 36173 10112 36185 10115
rect 34480 10084 36185 10112
rect 34480 10072 34486 10084
rect 36173 10081 36185 10084
rect 36219 10081 36231 10115
rect 37642 10112 37648 10124
rect 36173 10075 36231 10081
rect 36280 10084 37648 10112
rect 27246 10044 27252 10056
rect 26988 10016 27252 10044
rect 26881 10007 26939 10013
rect 27246 10004 27252 10016
rect 27304 10044 27310 10056
rect 27709 10047 27767 10053
rect 27709 10044 27721 10047
rect 27304 10016 27721 10044
rect 27304 10004 27310 10016
rect 27709 10013 27721 10016
rect 27755 10013 27767 10047
rect 27709 10007 27767 10013
rect 22741 9979 22799 9985
rect 22741 9945 22753 9979
rect 22787 9976 22799 9979
rect 26786 9976 26792 9988
rect 22787 9948 26792 9976
rect 22787 9945 22799 9948
rect 22741 9939 22799 9945
rect 26786 9936 26792 9948
rect 26844 9936 26850 9988
rect 27724 9908 27752 10007
rect 28166 10004 28172 10056
rect 28224 10044 28230 10056
rect 28813 10047 28871 10053
rect 28813 10044 28825 10047
rect 28224 10016 28825 10044
rect 28224 10004 28230 10016
rect 28813 10013 28825 10016
rect 28859 10013 28871 10047
rect 28813 10007 28871 10013
rect 31662 10004 31668 10056
rect 31720 10044 31726 10056
rect 32217 10047 32275 10053
rect 31720 10016 31892 10044
rect 31720 10004 31726 10016
rect 27798 9936 27804 9988
rect 27856 9976 27862 9988
rect 27985 9979 28043 9985
rect 27985 9976 27997 9979
rect 27856 9948 27997 9976
rect 27856 9936 27862 9948
rect 27985 9945 27997 9948
rect 28031 9945 28043 9979
rect 27985 9939 28043 9945
rect 28442 9936 28448 9988
rect 28500 9976 28506 9988
rect 30098 9976 30104 9988
rect 28500 9948 30104 9976
rect 28500 9936 28506 9948
rect 30098 9936 30104 9948
rect 30156 9936 30162 9988
rect 31754 9976 31760 9988
rect 31234 9948 31760 9976
rect 31754 9936 31760 9948
rect 31812 9936 31818 9988
rect 31864 9976 31892 10016
rect 32217 10013 32229 10047
rect 32263 10044 32275 10047
rect 32398 10044 32404 10056
rect 32263 10016 32404 10044
rect 32263 10013 32275 10016
rect 32217 10007 32275 10013
rect 32398 10004 32404 10016
rect 32456 10004 32462 10056
rect 32674 10004 32680 10056
rect 32732 10044 32738 10056
rect 32861 10047 32919 10053
rect 32861 10044 32873 10047
rect 32732 10016 32873 10044
rect 32732 10004 32738 10016
rect 32861 10013 32873 10016
rect 32907 10013 32919 10047
rect 33873 10047 33931 10053
rect 33873 10044 33885 10047
rect 32861 10007 32919 10013
rect 32968 10016 33885 10044
rect 32968 9976 32996 10016
rect 33873 10013 33885 10016
rect 33919 10013 33931 10047
rect 33873 10007 33931 10013
rect 34514 10004 34520 10056
rect 34572 10044 34578 10056
rect 34793 10047 34851 10053
rect 34793 10044 34805 10047
rect 34572 10016 34805 10044
rect 34572 10004 34578 10016
rect 34793 10013 34805 10016
rect 34839 10013 34851 10047
rect 35434 10044 35440 10056
rect 35395 10016 35440 10044
rect 34793 10007 34851 10013
rect 35434 10004 35440 10016
rect 35492 10004 35498 10056
rect 35618 10044 35624 10056
rect 35579 10016 35624 10044
rect 35618 10004 35624 10016
rect 35676 10004 35682 10056
rect 36280 10053 36308 10084
rect 37642 10072 37648 10084
rect 37700 10112 37706 10124
rect 38562 10112 38568 10124
rect 37700 10084 38568 10112
rect 37700 10072 37706 10084
rect 38562 10072 38568 10084
rect 38620 10072 38626 10124
rect 38930 10112 38936 10124
rect 38891 10084 38936 10112
rect 38930 10072 38936 10084
rect 38988 10072 38994 10124
rect 40954 10112 40960 10124
rect 39960 10084 40960 10112
rect 36265 10047 36323 10053
rect 36265 10013 36277 10047
rect 36311 10013 36323 10047
rect 37826 10044 37832 10056
rect 37787 10016 37832 10044
rect 36265 10007 36323 10013
rect 37826 10004 37832 10016
rect 37884 10044 37890 10056
rect 39960 10044 39988 10084
rect 40954 10072 40960 10084
rect 41012 10072 41018 10124
rect 37884 10016 39988 10044
rect 37884 10004 37890 10016
rect 40034 10004 40040 10056
rect 40092 10044 40098 10056
rect 58069 10047 58127 10053
rect 40092 10016 45554 10044
rect 40092 10004 40098 10016
rect 31864 9948 32996 9976
rect 33137 9979 33195 9985
rect 33137 9945 33149 9979
rect 33183 9976 33195 9979
rect 33226 9976 33232 9988
rect 33183 9948 33232 9976
rect 33183 9945 33195 9948
rect 33137 9939 33195 9945
rect 33226 9936 33232 9948
rect 33284 9936 33290 9988
rect 33597 9979 33655 9985
rect 33597 9945 33609 9979
rect 33643 9976 33655 9979
rect 34054 9976 34060 9988
rect 33643 9948 34060 9976
rect 33643 9945 33655 9948
rect 33597 9939 33655 9945
rect 34054 9936 34060 9948
rect 34112 9976 34118 9988
rect 34606 9976 34612 9988
rect 34112 9948 34612 9976
rect 34112 9936 34118 9948
rect 34606 9936 34612 9948
rect 34664 9936 34670 9988
rect 45526 9976 45554 10016
rect 58069 10013 58081 10047
rect 58115 10044 58127 10047
rect 58158 10044 58164 10056
rect 58115 10016 58164 10044
rect 58115 10013 58127 10016
rect 58069 10007 58127 10013
rect 58158 10004 58164 10016
rect 58216 10004 58222 10056
rect 57517 9979 57575 9985
rect 57517 9976 57529 9979
rect 45526 9948 57529 9976
rect 57517 9945 57529 9948
rect 57563 9945 57575 9979
rect 57517 9939 57575 9945
rect 31018 9908 31024 9920
rect 27724 9880 31024 9908
rect 31018 9868 31024 9880
rect 31076 9868 31082 9920
rect 31481 9911 31539 9917
rect 31481 9877 31493 9911
rect 31527 9908 31539 9911
rect 31570 9908 31576 9920
rect 31527 9880 31576 9908
rect 31527 9877 31539 9880
rect 31481 9871 31539 9877
rect 31570 9868 31576 9880
rect 31628 9908 31634 9920
rect 33778 9908 33784 9920
rect 31628 9880 33784 9908
rect 31628 9868 31634 9880
rect 33778 9868 33784 9880
rect 33836 9868 33842 9920
rect 33870 9868 33876 9920
rect 33928 9908 33934 9920
rect 33965 9911 34023 9917
rect 33965 9908 33977 9911
rect 33928 9880 33977 9908
rect 33928 9868 33934 9880
rect 33965 9877 33977 9880
rect 34011 9877 34023 9911
rect 34146 9908 34152 9920
rect 34107 9880 34152 9908
rect 33965 9871 34023 9877
rect 34146 9868 34152 9880
rect 34204 9868 34210 9920
rect 34514 9868 34520 9920
rect 34572 9908 34578 9920
rect 35437 9911 35495 9917
rect 35437 9908 35449 9911
rect 34572 9880 35449 9908
rect 34572 9868 34578 9880
rect 35437 9877 35449 9880
rect 35483 9877 35495 9911
rect 35437 9871 35495 9877
rect 35802 9868 35808 9920
rect 35860 9908 35866 9920
rect 36817 9911 36875 9917
rect 36817 9908 36829 9911
rect 35860 9880 36829 9908
rect 35860 9868 35866 9880
rect 36817 9877 36829 9880
rect 36863 9908 36875 9911
rect 37182 9908 37188 9920
rect 36863 9880 37188 9908
rect 36863 9877 36875 9880
rect 36817 9871 36875 9877
rect 37182 9868 37188 9880
rect 37240 9908 37246 9920
rect 37277 9911 37335 9917
rect 37277 9908 37289 9911
rect 37240 9880 37289 9908
rect 37240 9868 37246 9880
rect 37277 9877 37289 9880
rect 37323 9877 37335 9911
rect 37277 9871 37335 9877
rect 38930 9868 38936 9920
rect 38988 9908 38994 9920
rect 40405 9911 40463 9917
rect 40405 9908 40417 9911
rect 38988 9880 40417 9908
rect 38988 9868 38994 9880
rect 40405 9877 40417 9880
rect 40451 9877 40463 9911
rect 40405 9871 40463 9877
rect 1104 9818 58880 9840
rect 1104 9766 20214 9818
rect 20266 9766 20278 9818
rect 20330 9766 20342 9818
rect 20394 9766 20406 9818
rect 20458 9766 20470 9818
rect 20522 9766 39478 9818
rect 39530 9766 39542 9818
rect 39594 9766 39606 9818
rect 39658 9766 39670 9818
rect 39722 9766 39734 9818
rect 39786 9766 58880 9818
rect 1104 9744 58880 9766
rect 24670 9704 24676 9716
rect 24631 9676 24676 9704
rect 24670 9664 24676 9676
rect 24728 9664 24734 9716
rect 26142 9664 26148 9716
rect 26200 9704 26206 9716
rect 26200 9676 27476 9704
rect 26200 9664 26206 9676
rect 11609 9639 11667 9645
rect 11609 9605 11621 9639
rect 11655 9636 11667 9639
rect 18414 9636 18420 9648
rect 11655 9608 18420 9636
rect 11655 9605 11667 9608
rect 11609 9599 11667 9605
rect 10597 9571 10655 9577
rect 10597 9537 10609 9571
rect 10643 9568 10655 9571
rect 11624 9568 11652 9599
rect 18414 9596 18420 9608
rect 18472 9596 18478 9648
rect 22741 9639 22799 9645
rect 22741 9605 22753 9639
rect 22787 9636 22799 9639
rect 25406 9636 25412 9648
rect 22787 9608 25412 9636
rect 22787 9605 22799 9608
rect 22741 9599 22799 9605
rect 10643 9540 11652 9568
rect 10643 9537 10655 9540
rect 10597 9531 10655 9537
rect 22002 9392 22008 9444
rect 22060 9432 22066 9444
rect 22756 9432 22784 9599
rect 25406 9596 25412 9608
rect 25464 9596 25470 9648
rect 25958 9596 25964 9648
rect 26016 9636 26022 9648
rect 27448 9645 27476 9676
rect 27706 9664 27712 9716
rect 27764 9704 27770 9716
rect 27890 9704 27896 9716
rect 27764 9676 27896 9704
rect 27764 9664 27770 9676
rect 27890 9664 27896 9676
rect 27948 9664 27954 9716
rect 27982 9664 27988 9716
rect 28040 9704 28046 9716
rect 28261 9707 28319 9713
rect 28261 9704 28273 9707
rect 28040 9676 28273 9704
rect 28040 9664 28046 9676
rect 28261 9673 28273 9676
rect 28307 9673 28319 9707
rect 28261 9667 28319 9673
rect 28442 9664 28448 9716
rect 28500 9704 28506 9716
rect 28500 9676 28545 9704
rect 28500 9664 28506 9676
rect 28626 9664 28632 9716
rect 28684 9704 28690 9716
rect 30558 9704 30564 9716
rect 28684 9676 30564 9704
rect 28684 9664 28690 9676
rect 30558 9664 30564 9676
rect 30616 9664 30622 9716
rect 31018 9664 31024 9716
rect 31076 9704 31082 9716
rect 31846 9704 31852 9716
rect 31076 9676 31852 9704
rect 31076 9664 31082 9676
rect 31846 9664 31852 9676
rect 31904 9664 31910 9716
rect 33134 9664 33140 9716
rect 33192 9704 33198 9716
rect 35066 9704 35072 9716
rect 33192 9676 35072 9704
rect 33192 9664 33198 9676
rect 35066 9664 35072 9676
rect 35124 9664 35130 9716
rect 35158 9664 35164 9716
rect 35216 9704 35222 9716
rect 40862 9704 40868 9716
rect 35216 9676 40868 9704
rect 35216 9664 35222 9676
rect 40862 9664 40868 9676
rect 40920 9664 40926 9716
rect 58158 9704 58164 9716
rect 58119 9676 58164 9704
rect 58158 9664 58164 9676
rect 58216 9664 58222 9716
rect 27433 9639 27491 9645
rect 26016 9608 26280 9636
rect 26016 9596 26022 9608
rect 26252 9580 26280 9608
rect 27433 9605 27445 9639
rect 27479 9605 27491 9639
rect 27433 9599 27491 9605
rect 27617 9639 27675 9645
rect 27617 9605 27629 9639
rect 27663 9636 27675 9639
rect 27663 9608 31892 9636
rect 27663 9605 27675 9608
rect 27617 9599 27675 9605
rect 23842 9528 23848 9580
rect 23900 9568 23906 9580
rect 26145 9571 26203 9577
rect 26145 9568 26157 9571
rect 23900 9540 26157 9568
rect 23900 9528 23906 9540
rect 26145 9537 26157 9540
rect 26191 9537 26203 9571
rect 26145 9531 26203 9537
rect 26234 9528 26240 9580
rect 26292 9568 26298 9580
rect 26292 9540 26337 9568
rect 26292 9528 26298 9540
rect 26878 9528 26884 9580
rect 26936 9568 26942 9580
rect 27338 9568 27344 9580
rect 26936 9540 27344 9568
rect 26936 9528 26942 9540
rect 27338 9528 27344 9540
rect 27396 9568 27402 9580
rect 27816 9568 28028 9574
rect 28077 9571 28135 9577
rect 28077 9568 28089 9571
rect 27396 9546 28089 9568
rect 27396 9540 27844 9546
rect 28000 9540 28089 9546
rect 27396 9528 27402 9540
rect 28077 9537 28089 9540
rect 28123 9537 28135 9571
rect 28350 9568 28356 9580
rect 28311 9540 28356 9568
rect 28077 9531 28135 9537
rect 28350 9528 28356 9540
rect 28408 9528 28414 9580
rect 29270 9528 29276 9580
rect 29328 9568 29334 9580
rect 29454 9568 29460 9580
rect 29328 9540 29460 9568
rect 29328 9528 29334 9540
rect 29454 9528 29460 9540
rect 29512 9568 29518 9580
rect 29822 9568 29828 9580
rect 29512 9540 29828 9568
rect 29512 9528 29518 9540
rect 29822 9528 29828 9540
rect 29880 9528 29886 9580
rect 30098 9568 30104 9580
rect 30059 9540 30104 9568
rect 30098 9528 30104 9540
rect 30156 9528 30162 9580
rect 31110 9568 31116 9580
rect 31071 9540 31116 9568
rect 31110 9528 31116 9540
rect 31168 9528 31174 9580
rect 25038 9460 25044 9512
rect 25096 9500 25102 9512
rect 25133 9503 25191 9509
rect 25133 9500 25145 9503
rect 25096 9472 25145 9500
rect 25096 9460 25102 9472
rect 25133 9469 25145 9472
rect 25179 9500 25191 9503
rect 26326 9500 26332 9512
rect 25179 9472 26332 9500
rect 25179 9469 25191 9472
rect 25133 9463 25191 9469
rect 26326 9460 26332 9472
rect 26384 9500 26390 9512
rect 27798 9500 27804 9512
rect 26384 9472 27804 9500
rect 26384 9460 26390 9472
rect 27798 9460 27804 9472
rect 27856 9460 27862 9512
rect 29089 9503 29147 9509
rect 29089 9500 29101 9503
rect 28092 9472 29101 9500
rect 28092 9444 28120 9472
rect 29089 9469 29101 9472
rect 29135 9469 29147 9503
rect 30009 9503 30067 9509
rect 30009 9500 30021 9503
rect 29089 9463 29147 9469
rect 29196 9472 30021 9500
rect 23566 9432 23572 9444
rect 22060 9404 22784 9432
rect 23216 9404 23572 9432
rect 22060 9392 22066 9404
rect 8662 9324 8668 9376
rect 8720 9364 8726 9376
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 8720 9336 10425 9364
rect 8720 9324 8726 9336
rect 10413 9333 10425 9336
rect 10459 9333 10471 9367
rect 10413 9327 10471 9333
rect 22189 9367 22247 9373
rect 22189 9333 22201 9367
rect 22235 9364 22247 9367
rect 23216 9364 23244 9404
rect 23566 9392 23572 9404
rect 23624 9392 23630 9444
rect 24762 9432 24768 9444
rect 24412 9404 24768 9432
rect 24412 9376 24440 9404
rect 24762 9392 24768 9404
rect 24820 9392 24826 9444
rect 26418 9392 26424 9444
rect 26476 9432 26482 9444
rect 27706 9432 27712 9444
rect 26476 9404 27712 9432
rect 26476 9392 26482 9404
rect 27706 9392 27712 9404
rect 27764 9392 27770 9444
rect 28074 9392 28080 9444
rect 28132 9392 28138 9444
rect 22235 9336 23244 9364
rect 23293 9367 23351 9373
rect 22235 9333 22247 9336
rect 22189 9327 22247 9333
rect 23293 9333 23305 9367
rect 23339 9364 23351 9367
rect 23474 9364 23480 9376
rect 23339 9336 23480 9364
rect 23339 9333 23351 9336
rect 23293 9327 23351 9333
rect 23474 9324 23480 9336
rect 23532 9324 23538 9376
rect 24121 9367 24179 9373
rect 24121 9333 24133 9367
rect 24167 9364 24179 9367
rect 24394 9364 24400 9376
rect 24167 9336 24400 9364
rect 24167 9333 24179 9336
rect 24121 9327 24179 9333
rect 24394 9324 24400 9336
rect 24452 9324 24458 9376
rect 28442 9324 28448 9376
rect 28500 9364 28506 9376
rect 29196 9364 29224 9472
rect 30009 9469 30021 9472
rect 30055 9469 30067 9503
rect 31018 9500 31024 9512
rect 30009 9463 30067 9469
rect 30392 9472 30880 9500
rect 30979 9472 31024 9500
rect 29822 9392 29828 9444
rect 29880 9432 29886 9444
rect 30392 9432 30420 9472
rect 29880 9404 30420 9432
rect 30469 9435 30527 9441
rect 29880 9392 29886 9404
rect 30469 9401 30481 9435
rect 30515 9432 30527 9435
rect 30650 9432 30656 9444
rect 30515 9404 30656 9432
rect 30515 9401 30527 9404
rect 30469 9395 30527 9401
rect 30650 9392 30656 9404
rect 30708 9392 30714 9444
rect 30852 9432 30880 9472
rect 31018 9460 31024 9472
rect 31076 9460 31082 9512
rect 31864 9500 31892 9608
rect 31938 9596 31944 9648
rect 31996 9636 32002 9648
rect 32309 9639 32367 9645
rect 32309 9636 32321 9639
rect 31996 9608 32321 9636
rect 31996 9596 32002 9608
rect 32309 9605 32321 9608
rect 32355 9605 32367 9639
rect 32309 9599 32367 9605
rect 32490 9596 32496 9648
rect 32548 9636 32554 9648
rect 32548 9608 32593 9636
rect 32548 9596 32554 9608
rect 33042 9596 33048 9648
rect 33100 9636 33106 9648
rect 33597 9639 33655 9645
rect 33597 9636 33609 9639
rect 33100 9608 33609 9636
rect 33100 9596 33106 9608
rect 33597 9605 33609 9608
rect 33643 9605 33655 9639
rect 33597 9599 33655 9605
rect 33781 9639 33839 9645
rect 33781 9605 33793 9639
rect 33827 9636 33839 9639
rect 34146 9636 34152 9648
rect 33827 9608 34152 9636
rect 33827 9605 33839 9608
rect 33781 9599 33839 9605
rect 34146 9596 34152 9608
rect 34204 9596 34210 9648
rect 35342 9636 35348 9648
rect 34624 9608 35348 9636
rect 32398 9528 32404 9580
rect 32456 9568 32462 9580
rect 33965 9571 34023 9577
rect 32456 9540 32501 9568
rect 32456 9528 32462 9540
rect 33965 9537 33977 9571
rect 34011 9568 34023 9571
rect 34238 9568 34244 9580
rect 34011 9540 34244 9568
rect 34011 9537 34023 9540
rect 33965 9531 34023 9537
rect 34238 9528 34244 9540
rect 34296 9528 34302 9580
rect 34422 9568 34428 9580
rect 34383 9540 34428 9568
rect 34422 9528 34428 9540
rect 34480 9528 34486 9580
rect 34624 9577 34652 9608
rect 35342 9596 35348 9608
rect 35400 9636 35406 9648
rect 35713 9639 35771 9645
rect 35713 9636 35725 9639
rect 35400 9608 35725 9636
rect 35400 9596 35406 9608
rect 35713 9605 35725 9608
rect 35759 9605 35771 9639
rect 35713 9599 35771 9605
rect 36357 9639 36415 9645
rect 36357 9605 36369 9639
rect 36403 9636 36415 9639
rect 37182 9636 37188 9648
rect 36403 9608 37188 9636
rect 36403 9605 36415 9608
rect 36357 9599 36415 9605
rect 37182 9596 37188 9608
rect 37240 9596 37246 9648
rect 34609 9571 34667 9577
rect 34609 9537 34621 9571
rect 34655 9537 34667 9571
rect 34609 9531 34667 9537
rect 34974 9528 34980 9580
rect 35032 9568 35038 9580
rect 35253 9571 35311 9577
rect 35253 9568 35265 9571
rect 35032 9540 35265 9568
rect 35032 9528 35038 9540
rect 35253 9537 35265 9540
rect 35299 9537 35311 9571
rect 35253 9531 35311 9537
rect 36998 9528 37004 9580
rect 37056 9568 37062 9580
rect 43254 9568 43260 9580
rect 37056 9540 43260 9568
rect 37056 9528 37062 9540
rect 43254 9528 43260 9540
rect 43312 9528 43318 9580
rect 36262 9500 36268 9512
rect 31864 9472 36268 9500
rect 36262 9460 36268 9472
rect 36320 9460 36326 9512
rect 38470 9500 38476 9512
rect 36372 9472 38476 9500
rect 31294 9432 31300 9444
rect 30852 9404 31300 9432
rect 31294 9392 31300 9404
rect 31352 9392 31358 9444
rect 31478 9432 31484 9444
rect 31439 9404 31484 9432
rect 31478 9392 31484 9404
rect 31536 9392 31542 9444
rect 32674 9432 32680 9444
rect 32635 9404 32680 9432
rect 32674 9392 32680 9404
rect 32732 9392 32738 9444
rect 34238 9392 34244 9444
rect 34296 9432 34302 9444
rect 36372 9432 36400 9472
rect 38470 9460 38476 9472
rect 38528 9460 38534 9512
rect 41690 9500 41696 9512
rect 41386 9472 41696 9500
rect 34296 9404 36400 9432
rect 34296 9392 34302 9404
rect 36906 9392 36912 9444
rect 36964 9432 36970 9444
rect 39485 9435 39543 9441
rect 39485 9432 39497 9435
rect 36964 9404 39497 9432
rect 36964 9392 36970 9404
rect 39485 9401 39497 9404
rect 39531 9432 39543 9435
rect 40037 9435 40095 9441
rect 40037 9432 40049 9435
rect 39531 9404 40049 9432
rect 39531 9401 39543 9404
rect 39485 9395 39543 9401
rect 40037 9401 40049 9404
rect 40083 9432 40095 9435
rect 41386 9432 41414 9472
rect 41690 9460 41696 9472
rect 41748 9460 41754 9512
rect 40083 9404 41414 9432
rect 40083 9401 40095 9404
rect 40037 9395 40095 9401
rect 29454 9364 29460 9376
rect 28500 9336 29224 9364
rect 29415 9336 29460 9364
rect 28500 9324 28506 9336
rect 29454 9324 29460 9336
rect 29512 9324 29518 9376
rect 32125 9367 32183 9373
rect 32125 9333 32137 9367
rect 32171 9364 32183 9367
rect 32306 9364 32312 9376
rect 32171 9336 32312 9364
rect 32171 9333 32183 9336
rect 32125 9327 32183 9333
rect 32306 9324 32312 9336
rect 32364 9324 32370 9376
rect 34514 9364 34520 9376
rect 34475 9336 34520 9364
rect 34514 9324 34520 9336
rect 34572 9324 34578 9376
rect 35158 9364 35164 9376
rect 35119 9336 35164 9364
rect 35158 9324 35164 9336
rect 35216 9324 35222 9376
rect 36998 9324 37004 9376
rect 37056 9364 37062 9376
rect 37277 9367 37335 9373
rect 37277 9364 37289 9367
rect 37056 9336 37289 9364
rect 37056 9324 37062 9336
rect 37277 9333 37289 9336
rect 37323 9333 37335 9367
rect 37277 9327 37335 9333
rect 37921 9367 37979 9373
rect 37921 9333 37933 9367
rect 37967 9364 37979 9367
rect 38010 9364 38016 9376
rect 37967 9336 38016 9364
rect 37967 9333 37979 9336
rect 37921 9327 37979 9333
rect 38010 9324 38016 9336
rect 38068 9324 38074 9376
rect 38473 9367 38531 9373
rect 38473 9333 38485 9367
rect 38519 9364 38531 9367
rect 38654 9364 38660 9376
rect 38519 9336 38660 9364
rect 38519 9333 38531 9336
rect 38473 9327 38531 9333
rect 38654 9324 38660 9336
rect 38712 9324 38718 9376
rect 38930 9364 38936 9376
rect 38891 9336 38936 9364
rect 38930 9324 38936 9336
rect 38988 9324 38994 9376
rect 1104 9274 58880 9296
rect 1104 9222 10582 9274
rect 10634 9222 10646 9274
rect 10698 9222 10710 9274
rect 10762 9222 10774 9274
rect 10826 9222 10838 9274
rect 10890 9222 29846 9274
rect 29898 9222 29910 9274
rect 29962 9222 29974 9274
rect 30026 9222 30038 9274
rect 30090 9222 30102 9274
rect 30154 9222 49110 9274
rect 49162 9222 49174 9274
rect 49226 9222 49238 9274
rect 49290 9222 49302 9274
rect 49354 9222 49366 9274
rect 49418 9222 58880 9274
rect 1104 9200 58880 9222
rect 24949 9163 25007 9169
rect 24949 9129 24961 9163
rect 24995 9160 25007 9163
rect 25774 9160 25780 9172
rect 24995 9132 25780 9160
rect 24995 9129 25007 9132
rect 24949 9123 25007 9129
rect 25774 9120 25780 9132
rect 25832 9120 25838 9172
rect 26510 9160 26516 9172
rect 26471 9132 26516 9160
rect 26510 9120 26516 9132
rect 26568 9120 26574 9172
rect 27706 9160 27712 9172
rect 27619 9132 27712 9160
rect 27706 9120 27712 9132
rect 27764 9160 27770 9172
rect 27764 9132 28120 9160
rect 27764 9120 27770 9132
rect 23842 9052 23848 9104
rect 23900 9092 23906 9104
rect 25130 9092 25136 9104
rect 23900 9064 25136 9092
rect 23900 9052 23906 9064
rect 25130 9052 25136 9064
rect 25188 9052 25194 9104
rect 26053 9095 26111 9101
rect 26053 9061 26065 9095
rect 26099 9092 26111 9095
rect 28092 9092 28120 9132
rect 28626 9120 28632 9172
rect 28684 9160 28690 9172
rect 28813 9163 28871 9169
rect 28813 9160 28825 9163
rect 28684 9132 28825 9160
rect 28684 9120 28690 9132
rect 28813 9129 28825 9132
rect 28859 9129 28871 9163
rect 28813 9123 28871 9129
rect 29362 9120 29368 9172
rect 29420 9120 29426 9172
rect 29733 9163 29791 9169
rect 29733 9129 29745 9163
rect 29779 9160 29791 9163
rect 30466 9160 30472 9172
rect 29779 9132 30472 9160
rect 29779 9129 29791 9132
rect 29733 9123 29791 9129
rect 30466 9120 30472 9132
rect 30524 9120 30530 9172
rect 31570 9160 31576 9172
rect 31531 9132 31576 9160
rect 31570 9120 31576 9132
rect 31628 9120 31634 9172
rect 32493 9163 32551 9169
rect 32493 9129 32505 9163
rect 32539 9160 32551 9163
rect 32950 9160 32956 9172
rect 32539 9132 32956 9160
rect 32539 9129 32551 9132
rect 32493 9123 32551 9129
rect 32950 9120 32956 9132
rect 33008 9120 33014 9172
rect 33318 9160 33324 9172
rect 33279 9132 33324 9160
rect 33318 9120 33324 9132
rect 33376 9120 33382 9172
rect 33965 9163 34023 9169
rect 33965 9129 33977 9163
rect 34011 9160 34023 9163
rect 34422 9160 34428 9172
rect 34011 9132 34428 9160
rect 34011 9129 34023 9132
rect 33965 9123 34023 9129
rect 34422 9120 34428 9132
rect 34480 9120 34486 9172
rect 35250 9160 35256 9172
rect 35211 9132 35256 9160
rect 35250 9120 35256 9132
rect 35308 9120 35314 9172
rect 36262 9120 36268 9172
rect 36320 9160 36326 9172
rect 37461 9163 37519 9169
rect 37461 9160 37473 9163
rect 36320 9132 37473 9160
rect 36320 9120 36326 9132
rect 37461 9129 37473 9132
rect 37507 9160 37519 9163
rect 38654 9160 38660 9172
rect 37507 9132 38660 9160
rect 37507 9129 37519 9132
rect 37461 9123 37519 9129
rect 38654 9120 38660 9132
rect 38712 9120 38718 9172
rect 28442 9092 28448 9104
rect 26099 9064 28028 9092
rect 28092 9064 28448 9092
rect 26099 9061 26111 9064
rect 26053 9055 26111 9061
rect 21726 8984 21732 9036
rect 21784 9024 21790 9036
rect 27706 9024 27712 9036
rect 21784 8996 27712 9024
rect 21784 8984 21790 8996
rect 27706 8984 27712 8996
rect 27764 8984 27770 9036
rect 28000 9024 28028 9064
rect 28442 9052 28448 9064
rect 28500 9052 28506 9104
rect 29380 9092 29408 9120
rect 30926 9092 30932 9104
rect 28552 9064 29868 9092
rect 30887 9064 30932 9092
rect 28074 9024 28080 9036
rect 28000 8996 28080 9024
rect 28074 8984 28080 8996
rect 28132 8984 28138 9036
rect 28258 9024 28264 9036
rect 28219 8996 28264 9024
rect 28258 8984 28264 8996
rect 28316 8984 28322 9036
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 11514 8956 11520 8968
rect 1719 8928 11520 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 21266 8916 21272 8968
rect 21324 8956 21330 8968
rect 25409 8959 25467 8965
rect 25409 8956 25421 8959
rect 21324 8928 25421 8956
rect 21324 8916 21330 8928
rect 25409 8925 25421 8928
rect 25455 8956 25467 8959
rect 26970 8956 26976 8968
rect 25455 8928 26976 8956
rect 25455 8925 25467 8928
rect 25409 8919 25467 8925
rect 26970 8916 26976 8928
rect 27028 8916 27034 8968
rect 27062 8916 27068 8968
rect 27120 8956 27126 8968
rect 27157 8959 27215 8965
rect 27157 8956 27169 8959
rect 27120 8928 27169 8956
rect 27120 8916 27126 8928
rect 27157 8925 27169 8928
rect 27203 8956 27215 8959
rect 28552 8956 28580 9064
rect 28626 8984 28632 9036
rect 28684 9024 28690 9036
rect 29840 9032 29868 9064
rect 30926 9052 30932 9064
rect 30984 9052 30990 9104
rect 31662 9052 31668 9104
rect 31720 9092 31726 9104
rect 36814 9092 36820 9104
rect 31720 9064 31800 9092
rect 31720 9052 31726 9064
rect 29840 9024 30033 9032
rect 30098 9024 30104 9036
rect 28684 8996 29792 9024
rect 29840 9004 30104 9024
rect 30005 8996 30104 9004
rect 28684 8984 28690 8996
rect 27203 8928 28580 8956
rect 27203 8925 27215 8928
rect 27157 8919 27215 8925
rect 28718 8916 28724 8968
rect 28776 8956 28782 8968
rect 28813 8959 28871 8965
rect 28813 8956 28825 8959
rect 28776 8928 28825 8956
rect 28776 8916 28782 8928
rect 28813 8925 28825 8928
rect 28859 8925 28871 8959
rect 28813 8919 28871 8925
rect 29764 8931 29792 8996
rect 30098 8984 30104 8996
rect 30156 8984 30162 9036
rect 30650 9024 30656 9036
rect 30611 8996 30656 9024
rect 30650 8984 30656 8996
rect 30708 8984 30714 9036
rect 31772 9033 31800 9064
rect 31864 9064 36820 9092
rect 31757 9027 31815 9033
rect 31757 8993 31769 9027
rect 31803 8993 31815 9027
rect 31757 8987 31815 8993
rect 30558 8956 30564 8968
rect 29764 8925 29837 8931
rect 30519 8928 30564 8956
rect 16850 8848 16856 8900
rect 16908 8888 16914 8900
rect 26418 8888 26424 8900
rect 16908 8860 26424 8888
rect 16908 8848 16914 8860
rect 26418 8848 26424 8860
rect 26476 8848 26482 8900
rect 26510 8848 26516 8900
rect 26568 8888 26574 8900
rect 29549 8891 29607 8897
rect 29764 8894 29791 8925
rect 29549 8888 29561 8891
rect 26568 8860 29561 8888
rect 26568 8848 26574 8860
rect 29549 8857 29561 8860
rect 29595 8857 29607 8891
rect 29779 8891 29791 8894
rect 29825 8891 29837 8925
rect 30558 8916 30564 8928
rect 30616 8916 30622 8968
rect 31864 8965 31892 9064
rect 36814 9052 36820 9064
rect 36872 9052 36878 9104
rect 37642 9052 37648 9104
rect 37700 9092 37706 9104
rect 38013 9095 38071 9101
rect 38013 9092 38025 9095
rect 37700 9064 38025 9092
rect 37700 9052 37706 9064
rect 38013 9061 38025 9064
rect 38059 9092 38071 9095
rect 38562 9092 38568 9104
rect 38059 9064 38568 9092
rect 38059 9061 38071 9064
rect 38013 9055 38071 9061
rect 38562 9052 38568 9064
rect 38620 9052 38626 9104
rect 32398 8984 32404 9036
rect 32456 9024 32462 9036
rect 32858 9024 32864 9036
rect 32456 8996 32864 9024
rect 32456 8984 32462 8996
rect 32858 8984 32864 8996
rect 32916 8984 32922 9036
rect 33042 8984 33048 9036
rect 33100 9024 33106 9036
rect 33137 9027 33195 9033
rect 33137 9024 33149 9027
rect 33100 8996 33149 9024
rect 33100 8984 33106 8996
rect 33137 8993 33149 8996
rect 33183 8993 33195 9027
rect 34330 9024 34336 9036
rect 33137 8987 33195 8993
rect 33336 8996 34336 9024
rect 31580 8959 31638 8965
rect 31580 8925 31592 8959
rect 31626 8958 31638 8959
rect 31849 8959 31907 8965
rect 31626 8930 31708 8958
rect 31626 8925 31638 8930
rect 31580 8919 31638 8925
rect 29779 8885 29837 8891
rect 29549 8851 29607 8857
rect 30006 8848 30012 8900
rect 30064 8888 30070 8900
rect 31680 8888 31708 8930
rect 31849 8925 31861 8959
rect 31895 8925 31907 8959
rect 31849 8919 31907 8925
rect 32030 8916 32036 8968
rect 32088 8956 32094 8968
rect 32309 8959 32367 8965
rect 32309 8956 32321 8959
rect 32088 8928 32321 8956
rect 32088 8916 32094 8928
rect 32309 8925 32321 8928
rect 32355 8925 32367 8959
rect 32309 8919 32367 8925
rect 33336 8888 33364 8996
rect 34330 8984 34336 8996
rect 34388 8984 34394 9036
rect 34701 9027 34759 9033
rect 34701 9024 34713 9027
rect 34440 8996 34713 9024
rect 33413 8959 33471 8965
rect 33413 8925 33425 8959
rect 33459 8925 33471 8959
rect 33413 8919 33471 8925
rect 30064 8860 31616 8888
rect 31680 8860 33364 8888
rect 33428 8888 33456 8919
rect 33686 8916 33692 8968
rect 33744 8956 33750 8968
rect 34057 8959 34115 8965
rect 34057 8956 34069 8959
rect 33744 8928 34069 8956
rect 33744 8916 33750 8928
rect 34057 8925 34069 8928
rect 34103 8956 34115 8959
rect 34238 8956 34244 8968
rect 34103 8928 34244 8956
rect 34103 8925 34115 8928
rect 34057 8919 34115 8925
rect 34238 8916 34244 8928
rect 34296 8956 34302 8968
rect 34440 8956 34468 8996
rect 34701 8993 34713 8996
rect 34747 8993 34759 9027
rect 34701 8987 34759 8993
rect 35250 8984 35256 9036
rect 35308 9024 35314 9036
rect 35526 9024 35532 9036
rect 35308 8996 35532 9024
rect 35308 8984 35314 8996
rect 35526 8984 35532 8996
rect 35584 9024 35590 9036
rect 35897 9027 35955 9033
rect 35897 9024 35909 9027
rect 35584 8996 35909 9024
rect 35584 8984 35590 8996
rect 35897 8993 35909 8996
rect 35943 9024 35955 9027
rect 43806 9024 43812 9036
rect 35943 8996 43812 9024
rect 35943 8993 35955 8996
rect 35897 8987 35955 8993
rect 43806 8984 43812 8996
rect 43864 8984 43870 9036
rect 37458 8956 37464 8968
rect 34296 8928 34468 8956
rect 34532 8928 37464 8956
rect 34296 8916 34302 8928
rect 34422 8888 34428 8900
rect 33428 8860 34428 8888
rect 30064 8848 30070 8860
rect 1486 8820 1492 8832
rect 1447 8792 1492 8820
rect 1486 8780 1492 8792
rect 1544 8780 1550 8832
rect 20622 8780 20628 8832
rect 20680 8820 20686 8832
rect 22741 8823 22799 8829
rect 22741 8820 22753 8823
rect 20680 8792 22753 8820
rect 20680 8780 20686 8792
rect 22741 8789 22753 8792
rect 22787 8820 22799 8823
rect 23290 8820 23296 8832
rect 22787 8792 23296 8820
rect 22787 8789 22799 8792
rect 22741 8783 22799 8789
rect 23290 8780 23296 8792
rect 23348 8780 23354 8832
rect 23842 8820 23848 8832
rect 23803 8792 23848 8820
rect 23842 8780 23848 8792
rect 23900 8780 23906 8832
rect 24118 8780 24124 8832
rect 24176 8820 24182 8832
rect 29362 8820 29368 8832
rect 24176 8792 29368 8820
rect 24176 8780 24182 8792
rect 29362 8780 29368 8792
rect 29420 8780 29426 8832
rect 29914 8820 29920 8832
rect 29875 8792 29920 8820
rect 29914 8780 29920 8792
rect 29972 8780 29978 8832
rect 31386 8780 31392 8832
rect 31444 8820 31450 8832
rect 31588 8820 31616 8860
rect 34422 8848 34428 8860
rect 34480 8848 34486 8900
rect 32674 8820 32680 8832
rect 31444 8792 31489 8820
rect 31588 8792 32680 8820
rect 31444 8780 31450 8792
rect 32674 8780 32680 8792
rect 32732 8780 32738 8832
rect 33137 8823 33195 8829
rect 33137 8789 33149 8823
rect 33183 8820 33195 8823
rect 34532 8820 34560 8928
rect 37458 8916 37464 8928
rect 37516 8916 37522 8968
rect 34698 8848 34704 8900
rect 34756 8888 34762 8900
rect 36354 8888 36360 8900
rect 34756 8860 36360 8888
rect 34756 8848 34762 8860
rect 36354 8848 36360 8860
rect 36412 8888 36418 8900
rect 36909 8891 36967 8897
rect 36909 8888 36921 8891
rect 36412 8860 36921 8888
rect 36412 8848 36418 8860
rect 36909 8857 36921 8860
rect 36955 8857 36967 8891
rect 36909 8851 36967 8857
rect 37826 8848 37832 8900
rect 37884 8888 37890 8900
rect 38565 8891 38623 8897
rect 38565 8888 38577 8891
rect 37884 8860 38577 8888
rect 37884 8848 37890 8860
rect 38565 8857 38577 8860
rect 38611 8888 38623 8891
rect 38930 8888 38936 8900
rect 38611 8860 38936 8888
rect 38611 8857 38623 8860
rect 38565 8851 38623 8857
rect 38930 8848 38936 8860
rect 38988 8888 38994 8900
rect 39117 8891 39175 8897
rect 39117 8888 39129 8891
rect 38988 8860 39129 8888
rect 38988 8848 38994 8860
rect 39117 8857 39129 8860
rect 39163 8857 39175 8891
rect 39117 8851 39175 8857
rect 33183 8792 34560 8820
rect 39132 8820 39160 8851
rect 45554 8820 45560 8832
rect 39132 8792 45560 8820
rect 33183 8789 33195 8792
rect 33137 8783 33195 8789
rect 45554 8780 45560 8792
rect 45612 8820 45618 8832
rect 46198 8820 46204 8832
rect 45612 8792 46204 8820
rect 45612 8780 45618 8792
rect 46198 8780 46204 8792
rect 46256 8780 46262 8832
rect 1104 8730 58880 8752
rect 1104 8678 20214 8730
rect 20266 8678 20278 8730
rect 20330 8678 20342 8730
rect 20394 8678 20406 8730
rect 20458 8678 20470 8730
rect 20522 8678 39478 8730
rect 39530 8678 39542 8730
rect 39594 8678 39606 8730
rect 39658 8678 39670 8730
rect 39722 8678 39734 8730
rect 39786 8678 58880 8730
rect 1104 8656 58880 8678
rect 23474 8576 23480 8628
rect 23532 8616 23538 8628
rect 24581 8619 24639 8625
rect 24581 8616 24593 8619
rect 23532 8588 24593 8616
rect 23532 8576 23538 8588
rect 24581 8585 24593 8588
rect 24627 8585 24639 8619
rect 24581 8579 24639 8585
rect 24946 8576 24952 8628
rect 25004 8616 25010 8628
rect 25133 8619 25191 8625
rect 25133 8616 25145 8619
rect 25004 8588 25145 8616
rect 25004 8576 25010 8588
rect 25133 8585 25145 8588
rect 25179 8585 25191 8619
rect 26326 8616 26332 8628
rect 26287 8588 26332 8616
rect 25133 8579 25191 8585
rect 26326 8576 26332 8588
rect 26384 8576 26390 8628
rect 27062 8616 27068 8628
rect 27023 8588 27068 8616
rect 27062 8576 27068 8588
rect 27120 8576 27126 8628
rect 27614 8616 27620 8628
rect 27575 8588 27620 8616
rect 27614 8576 27620 8588
rect 27672 8576 27678 8628
rect 27706 8576 27712 8628
rect 27764 8616 27770 8628
rect 27982 8616 27988 8628
rect 27764 8588 27988 8616
rect 27764 8576 27770 8588
rect 27982 8576 27988 8588
rect 28040 8576 28046 8628
rect 28166 8616 28172 8628
rect 28127 8588 28172 8616
rect 28166 8576 28172 8588
rect 28224 8576 28230 8628
rect 28718 8616 28724 8628
rect 28679 8588 28724 8616
rect 28718 8576 28724 8588
rect 28776 8576 28782 8628
rect 32214 8616 32220 8628
rect 29288 8588 32220 8616
rect 25498 8508 25504 8560
rect 25556 8548 25562 8560
rect 28626 8548 28632 8560
rect 25556 8520 28632 8548
rect 25556 8508 25562 8520
rect 28626 8508 28632 8520
rect 28684 8508 28690 8560
rect 25774 8480 25780 8492
rect 25735 8452 25780 8480
rect 25774 8440 25780 8452
rect 25832 8440 25838 8492
rect 28810 8480 28816 8492
rect 28771 8452 28816 8480
rect 28810 8440 28816 8452
rect 28868 8440 28874 8492
rect 29288 8480 29316 8588
rect 32214 8576 32220 8588
rect 32272 8576 32278 8628
rect 32309 8619 32367 8625
rect 32309 8585 32321 8619
rect 32355 8616 32367 8619
rect 32582 8616 32588 8628
rect 32355 8588 32588 8616
rect 32355 8585 32367 8588
rect 32309 8579 32367 8585
rect 32582 8576 32588 8588
rect 32640 8576 32646 8628
rect 32674 8576 32680 8628
rect 32732 8616 32738 8628
rect 33410 8616 33416 8628
rect 32732 8588 33416 8616
rect 32732 8576 32738 8588
rect 33410 8576 33416 8588
rect 33468 8576 33474 8628
rect 33597 8619 33655 8625
rect 33597 8585 33609 8619
rect 33643 8616 33655 8619
rect 33962 8616 33968 8628
rect 33643 8588 33968 8616
rect 33643 8585 33655 8588
rect 33597 8579 33655 8585
rect 33962 8576 33968 8588
rect 34020 8576 34026 8628
rect 34146 8616 34152 8628
rect 34107 8588 34152 8616
rect 34146 8576 34152 8588
rect 34204 8576 34210 8628
rect 34606 8576 34612 8628
rect 34664 8616 34670 8628
rect 35161 8619 35219 8625
rect 35161 8616 35173 8619
rect 34664 8588 35173 8616
rect 34664 8576 34670 8588
rect 35161 8585 35173 8588
rect 35207 8585 35219 8619
rect 35161 8579 35219 8585
rect 36357 8619 36415 8625
rect 36357 8585 36369 8619
rect 36403 8616 36415 8619
rect 37274 8616 37280 8628
rect 36403 8588 37280 8616
rect 36403 8585 36415 8588
rect 36357 8579 36415 8585
rect 37274 8576 37280 8588
rect 37332 8576 37338 8628
rect 37366 8576 37372 8628
rect 37424 8616 37430 8628
rect 40218 8616 40224 8628
rect 37424 8588 40224 8616
rect 37424 8576 37430 8588
rect 40218 8576 40224 8588
rect 40276 8576 40282 8628
rect 29362 8508 29368 8560
rect 29420 8548 29426 8560
rect 30006 8548 30012 8560
rect 29420 8520 30012 8548
rect 29420 8508 29426 8520
rect 30006 8508 30012 8520
rect 30064 8508 30070 8560
rect 30098 8508 30104 8560
rect 30156 8548 30162 8560
rect 31113 8551 31171 8557
rect 31113 8548 31125 8551
rect 30156 8520 31125 8548
rect 30156 8508 30162 8520
rect 29457 8483 29515 8489
rect 29457 8480 29469 8483
rect 29288 8452 29469 8480
rect 29457 8449 29469 8452
rect 29503 8449 29515 8483
rect 29457 8443 29515 8449
rect 30190 8440 30196 8492
rect 30248 8480 30254 8492
rect 30285 8483 30343 8489
rect 30285 8480 30297 8483
rect 30248 8452 30297 8480
rect 30248 8440 30254 8452
rect 30285 8449 30297 8452
rect 30331 8449 30343 8483
rect 30926 8480 30932 8492
rect 30285 8443 30343 8449
rect 30576 8452 30932 8480
rect 19426 8372 19432 8424
rect 19484 8412 19490 8424
rect 19484 8384 22094 8412
rect 19484 8372 19490 8384
rect 22066 8344 22094 8384
rect 23290 8372 23296 8424
rect 23348 8412 23354 8424
rect 24029 8415 24087 8421
rect 24029 8412 24041 8415
rect 23348 8384 24041 8412
rect 23348 8372 23354 8384
rect 24029 8381 24041 8384
rect 24075 8412 24087 8415
rect 26786 8412 26792 8424
rect 24075 8384 26792 8412
rect 24075 8381 24087 8384
rect 24029 8375 24087 8381
rect 26786 8372 26792 8384
rect 26844 8372 26850 8424
rect 29362 8412 29368 8424
rect 29323 8384 29368 8412
rect 29362 8372 29368 8384
rect 29420 8372 29426 8424
rect 29730 8372 29736 8424
rect 29788 8412 29794 8424
rect 29825 8415 29883 8421
rect 29825 8412 29837 8415
rect 29788 8384 29837 8412
rect 29788 8372 29794 8384
rect 29825 8381 29837 8384
rect 29871 8381 29883 8415
rect 29825 8375 29883 8381
rect 29914 8372 29920 8424
rect 29972 8412 29978 8424
rect 30377 8415 30435 8421
rect 30377 8412 30389 8415
rect 29972 8384 30389 8412
rect 29972 8372 29978 8384
rect 30377 8381 30389 8384
rect 30423 8381 30435 8415
rect 30377 8375 30435 8381
rect 30576 8344 30604 8452
rect 30926 8440 30932 8452
rect 30984 8440 30990 8492
rect 31036 8480 31064 8520
rect 31113 8517 31125 8520
rect 31159 8517 31171 8551
rect 31113 8511 31171 8517
rect 31294 8508 31300 8560
rect 31352 8557 31358 8560
rect 31352 8551 31387 8557
rect 31375 8548 31387 8551
rect 32950 8548 32956 8560
rect 31375 8520 32956 8548
rect 31375 8517 31387 8520
rect 31352 8511 31387 8517
rect 31352 8508 31358 8511
rect 32950 8508 32956 8520
rect 33008 8508 33014 8560
rect 33428 8548 33456 8576
rect 35710 8548 35716 8560
rect 33428 8520 35716 8548
rect 35710 8508 35716 8520
rect 35768 8508 35774 8560
rect 36078 8508 36084 8560
rect 36136 8548 36142 8560
rect 38473 8551 38531 8557
rect 38473 8548 38485 8551
rect 36136 8520 38485 8548
rect 36136 8508 36142 8520
rect 38473 8517 38485 8520
rect 38519 8548 38531 8551
rect 38746 8548 38752 8560
rect 38519 8520 38752 8548
rect 38519 8517 38531 8520
rect 38473 8511 38531 8517
rect 38746 8508 38752 8520
rect 38804 8508 38810 8560
rect 31754 8480 31760 8492
rect 31036 8452 31760 8480
rect 31754 8440 31760 8452
rect 31812 8440 31818 8492
rect 32122 8480 32128 8492
rect 32083 8452 32128 8480
rect 32122 8440 32128 8452
rect 32180 8440 32186 8492
rect 32858 8480 32864 8492
rect 32819 8452 32864 8480
rect 32858 8440 32864 8452
rect 32916 8440 32922 8492
rect 33042 8440 33048 8492
rect 33100 8480 33106 8492
rect 35250 8480 35256 8492
rect 33100 8452 35256 8480
rect 33100 8440 33106 8452
rect 35250 8440 35256 8452
rect 35308 8440 35314 8492
rect 35618 8412 35624 8424
rect 30668 8384 35624 8412
rect 30668 8353 30696 8384
rect 35618 8372 35624 8384
rect 35676 8372 35682 8424
rect 22066 8316 30604 8344
rect 30653 8347 30711 8353
rect 30653 8313 30665 8347
rect 30699 8313 30711 8347
rect 30653 8307 30711 8313
rect 31481 8347 31539 8353
rect 31481 8313 31493 8347
rect 31527 8344 31539 8347
rect 31570 8344 31576 8356
rect 31527 8316 31576 8344
rect 31527 8313 31539 8316
rect 31481 8307 31539 8313
rect 31570 8304 31576 8316
rect 31628 8304 31634 8356
rect 32030 8344 32036 8356
rect 31726 8316 32036 8344
rect 30469 8279 30527 8285
rect 30469 8245 30481 8279
rect 30515 8276 30527 8279
rect 30834 8276 30840 8288
rect 30515 8248 30840 8276
rect 30515 8245 30527 8248
rect 30469 8239 30527 8245
rect 30834 8236 30840 8248
rect 30892 8236 30898 8288
rect 31294 8276 31300 8288
rect 31255 8248 31300 8276
rect 31294 8236 31300 8248
rect 31352 8276 31358 8288
rect 31726 8276 31754 8316
rect 32030 8304 32036 8316
rect 32088 8304 32094 8356
rect 32953 8347 33011 8353
rect 32953 8313 32965 8347
rect 32999 8344 33011 8347
rect 33042 8344 33048 8356
rect 32999 8316 33048 8344
rect 32999 8313 33011 8316
rect 32953 8307 33011 8313
rect 33042 8304 33048 8316
rect 33100 8304 33106 8356
rect 38102 8344 38108 8356
rect 33152 8316 38108 8344
rect 31352 8248 31754 8276
rect 31352 8236 31358 8248
rect 31938 8236 31944 8288
rect 31996 8276 32002 8288
rect 32674 8276 32680 8288
rect 31996 8248 32680 8276
rect 31996 8236 32002 8248
rect 32674 8236 32680 8248
rect 32732 8276 32738 8288
rect 33152 8276 33180 8316
rect 38102 8304 38108 8316
rect 38160 8304 38166 8356
rect 32732 8248 33180 8276
rect 34701 8279 34759 8285
rect 32732 8236 32738 8248
rect 34701 8245 34713 8279
rect 34747 8276 34759 8279
rect 37182 8276 37188 8288
rect 34747 8248 37188 8276
rect 34747 8245 34759 8248
rect 34701 8239 34759 8245
rect 37182 8236 37188 8248
rect 37240 8236 37246 8288
rect 37826 8276 37832 8288
rect 37787 8248 37832 8276
rect 37826 8236 37832 8248
rect 37884 8236 37890 8288
rect 1104 8186 58880 8208
rect 1104 8134 10582 8186
rect 10634 8134 10646 8186
rect 10698 8134 10710 8186
rect 10762 8134 10774 8186
rect 10826 8134 10838 8186
rect 10890 8134 29846 8186
rect 29898 8134 29910 8186
rect 29962 8134 29974 8186
rect 30026 8134 30038 8186
rect 30090 8134 30102 8186
rect 30154 8134 49110 8186
rect 49162 8134 49174 8186
rect 49226 8134 49238 8186
rect 49290 8134 49302 8186
rect 49354 8134 49366 8186
rect 49418 8134 58880 8186
rect 1104 8112 58880 8134
rect 24762 8032 24768 8084
rect 24820 8072 24826 8084
rect 24857 8075 24915 8081
rect 24857 8072 24869 8075
rect 24820 8044 24869 8072
rect 24820 8032 24826 8044
rect 24857 8041 24869 8044
rect 24903 8041 24915 8075
rect 25958 8072 25964 8084
rect 25919 8044 25964 8072
rect 24857 8035 24915 8041
rect 25958 8032 25964 8044
rect 26016 8032 26022 8084
rect 26050 8032 26056 8084
rect 26108 8072 26114 8084
rect 26513 8075 26571 8081
rect 26513 8072 26525 8075
rect 26108 8044 26525 8072
rect 26108 8032 26114 8044
rect 26513 8041 26525 8044
rect 26559 8041 26571 8075
rect 27246 8072 27252 8084
rect 27207 8044 27252 8072
rect 26513 8035 26571 8041
rect 27246 8032 27252 8044
rect 27304 8032 27310 8084
rect 27893 8075 27951 8081
rect 27893 8041 27905 8075
rect 27939 8072 27951 8075
rect 28074 8072 28080 8084
rect 27939 8044 28080 8072
rect 27939 8041 27951 8044
rect 27893 8035 27951 8041
rect 28074 8032 28080 8044
rect 28132 8032 28138 8084
rect 29638 8072 29644 8084
rect 29599 8044 29644 8072
rect 29638 8032 29644 8044
rect 29696 8032 29702 8084
rect 31110 8072 31116 8084
rect 30208 8044 31116 8072
rect 27798 7964 27804 8016
rect 27856 8004 27862 8016
rect 28353 8007 28411 8013
rect 28353 8004 28365 8007
rect 27856 7976 28365 8004
rect 27856 7964 27862 7976
rect 28353 7973 28365 7976
rect 28399 7973 28411 8007
rect 28353 7967 28411 7973
rect 29825 7871 29883 7877
rect 29825 7837 29837 7871
rect 29871 7868 29883 7871
rect 30208 7868 30236 8044
rect 31110 8032 31116 8044
rect 31168 8032 31174 8084
rect 31205 8075 31263 8081
rect 31205 8041 31217 8075
rect 31251 8072 31263 8075
rect 32214 8072 32220 8084
rect 31251 8044 32220 8072
rect 31251 8041 31263 8044
rect 31205 8035 31263 8041
rect 32214 8032 32220 8044
rect 32272 8032 32278 8084
rect 32950 8072 32956 8084
rect 32911 8044 32956 8072
rect 32950 8032 32956 8044
rect 33008 8032 33014 8084
rect 33594 8072 33600 8084
rect 33507 8044 33600 8072
rect 33594 8032 33600 8044
rect 33652 8072 33658 8084
rect 38838 8072 38844 8084
rect 33652 8044 34652 8072
rect 33652 8032 33658 8044
rect 30377 8007 30435 8013
rect 30377 7973 30389 8007
rect 30423 8004 30435 8007
rect 30466 8004 30472 8016
rect 30423 7976 30472 8004
rect 30423 7973 30435 7976
rect 30377 7967 30435 7973
rect 30466 7964 30472 7976
rect 30524 7964 30530 8016
rect 34624 8004 34652 8044
rect 34808 8044 38844 8072
rect 34808 8004 34836 8044
rect 38838 8032 38844 8044
rect 38896 8032 38902 8084
rect 34624 7976 34836 8004
rect 34974 7964 34980 8016
rect 35032 8004 35038 8016
rect 35897 8007 35955 8013
rect 35897 8004 35909 8007
rect 35032 7976 35909 8004
rect 35032 7964 35038 7976
rect 35897 7973 35909 7976
rect 35943 8004 35955 8007
rect 43070 8004 43076 8016
rect 35943 7976 43076 8004
rect 35943 7973 35955 7976
rect 35897 7967 35955 7973
rect 43070 7964 43076 7976
rect 43128 7964 43134 8016
rect 30285 7939 30343 7945
rect 30285 7905 30297 7939
rect 30331 7936 30343 7939
rect 31849 7939 31907 7945
rect 30331 7908 30420 7936
rect 30331 7905 30343 7908
rect 30285 7899 30343 7905
rect 29871 7840 30236 7868
rect 29871 7837 29883 7840
rect 29825 7831 29883 7837
rect 14458 7800 14464 7812
rect 14419 7772 14464 7800
rect 14458 7760 14464 7772
rect 14516 7760 14522 7812
rect 14645 7803 14703 7809
rect 14645 7769 14657 7803
rect 14691 7769 14703 7803
rect 14645 7763 14703 7769
rect 14660 7732 14688 7763
rect 15286 7732 15292 7744
rect 14660 7704 15292 7732
rect 15286 7692 15292 7704
rect 15344 7692 15350 7744
rect 25498 7732 25504 7744
rect 25459 7704 25504 7732
rect 25498 7692 25504 7704
rect 25556 7732 25562 7744
rect 26142 7732 26148 7744
rect 25556 7704 26148 7732
rect 25556 7692 25562 7704
rect 26142 7692 26148 7704
rect 26200 7692 26206 7744
rect 28997 7735 29055 7741
rect 28997 7701 29009 7735
rect 29043 7732 29055 7735
rect 30282 7732 30288 7744
rect 29043 7704 30288 7732
rect 29043 7701 29055 7704
rect 28997 7695 29055 7701
rect 30282 7692 30288 7704
rect 30340 7692 30346 7744
rect 30392 7732 30420 7908
rect 31849 7905 31861 7939
rect 31895 7936 31907 7939
rect 33134 7936 33140 7948
rect 31895 7908 33140 7936
rect 31895 7905 31907 7908
rect 31849 7899 31907 7905
rect 33134 7896 33140 7908
rect 33192 7896 33198 7948
rect 33778 7896 33784 7948
rect 33836 7936 33842 7948
rect 34149 7939 34207 7945
rect 34149 7936 34161 7939
rect 33836 7908 34161 7936
rect 33836 7896 33842 7908
rect 34149 7905 34161 7908
rect 34195 7936 34207 7939
rect 44266 7936 44272 7948
rect 34195 7908 44272 7936
rect 34195 7905 34207 7908
rect 34149 7899 34207 7905
rect 44266 7896 44272 7908
rect 44324 7896 44330 7948
rect 51718 7896 51724 7948
rect 51776 7936 51782 7948
rect 57885 7939 57943 7945
rect 57885 7936 57897 7939
rect 51776 7908 57897 7936
rect 51776 7896 51782 7908
rect 57885 7905 57897 7908
rect 57931 7905 57943 7939
rect 57885 7899 57943 7905
rect 30560 7881 30618 7887
rect 30469 7871 30527 7877
rect 30469 7837 30481 7871
rect 30515 7837 30527 7871
rect 30560 7847 30572 7881
rect 30606 7878 30618 7881
rect 30606 7868 30696 7878
rect 30926 7868 30932 7880
rect 30606 7850 30932 7868
rect 30606 7847 30618 7850
rect 30560 7841 30618 7847
rect 30668 7840 30932 7850
rect 30469 7831 30527 7837
rect 30484 7800 30512 7831
rect 30926 7828 30932 7840
rect 30984 7828 30990 7880
rect 31110 7868 31116 7880
rect 31071 7840 31116 7868
rect 31110 7828 31116 7840
rect 31168 7828 31174 7880
rect 31757 7871 31815 7877
rect 31757 7837 31769 7871
rect 31803 7868 31815 7871
rect 32858 7868 32864 7880
rect 31803 7840 32864 7868
rect 31803 7837 31815 7840
rect 31757 7831 31815 7837
rect 32858 7828 32864 7840
rect 32916 7828 32922 7880
rect 33962 7828 33968 7880
rect 34020 7868 34026 7880
rect 37550 7868 37556 7880
rect 34020 7840 37556 7868
rect 34020 7828 34026 7840
rect 37550 7828 37556 7840
rect 37608 7828 37614 7880
rect 58158 7868 58164 7880
rect 58119 7840 58164 7868
rect 58158 7828 58164 7840
rect 58216 7828 58222 7880
rect 30650 7800 30656 7812
rect 30484 7772 30656 7800
rect 30650 7760 30656 7772
rect 30708 7760 30714 7812
rect 31018 7760 31024 7812
rect 31076 7800 31082 7812
rect 32401 7803 32459 7809
rect 32401 7800 32413 7803
rect 31076 7772 32413 7800
rect 31076 7760 31082 7772
rect 32401 7769 32413 7772
rect 32447 7769 32459 7803
rect 34698 7800 34704 7812
rect 34659 7772 34704 7800
rect 32401 7763 32459 7769
rect 34698 7760 34704 7772
rect 34756 7760 34762 7812
rect 35250 7800 35256 7812
rect 35211 7772 35256 7800
rect 35250 7760 35256 7772
rect 35308 7760 35314 7812
rect 35342 7760 35348 7812
rect 35400 7800 35406 7812
rect 37461 7803 37519 7809
rect 37461 7800 37473 7803
rect 35400 7772 37473 7800
rect 35400 7760 35406 7772
rect 37461 7769 37473 7772
rect 37507 7800 37519 7803
rect 37826 7800 37832 7812
rect 37507 7772 37832 7800
rect 37507 7769 37519 7772
rect 37461 7763 37519 7769
rect 37826 7760 37832 7772
rect 37884 7760 37890 7812
rect 30466 7732 30472 7744
rect 30392 7704 30472 7732
rect 30466 7692 30472 7704
rect 30524 7692 30530 7744
rect 30668 7732 30696 7760
rect 32306 7732 32312 7744
rect 30668 7704 32312 7732
rect 32306 7692 32312 7704
rect 32364 7692 32370 7744
rect 36354 7732 36360 7744
rect 36315 7704 36360 7732
rect 36354 7692 36360 7704
rect 36412 7692 36418 7744
rect 36906 7732 36912 7744
rect 36867 7704 36912 7732
rect 36906 7692 36912 7704
rect 36964 7692 36970 7744
rect 1104 7642 58880 7664
rect 1104 7590 20214 7642
rect 20266 7590 20278 7642
rect 20330 7590 20342 7642
rect 20394 7590 20406 7642
rect 20458 7590 20470 7642
rect 20522 7590 39478 7642
rect 39530 7590 39542 7642
rect 39594 7590 39606 7642
rect 39658 7590 39670 7642
rect 39722 7590 39734 7642
rect 39786 7590 58880 7642
rect 1104 7568 58880 7590
rect 25866 7528 25872 7540
rect 25779 7500 25872 7528
rect 25866 7488 25872 7500
rect 25924 7528 25930 7540
rect 26234 7528 26240 7540
rect 25924 7500 26240 7528
rect 25924 7488 25930 7500
rect 26234 7488 26240 7500
rect 26292 7488 26298 7540
rect 26418 7488 26424 7540
rect 26476 7528 26482 7540
rect 27341 7531 27399 7537
rect 27341 7528 27353 7531
rect 26476 7500 27353 7528
rect 26476 7488 26482 7500
rect 27341 7497 27353 7500
rect 27387 7497 27399 7531
rect 27341 7491 27399 7497
rect 27522 7488 27528 7540
rect 27580 7528 27586 7540
rect 27893 7531 27951 7537
rect 27893 7528 27905 7531
rect 27580 7500 27905 7528
rect 27580 7488 27586 7500
rect 27893 7497 27905 7500
rect 27939 7497 27951 7531
rect 28534 7528 28540 7540
rect 28495 7500 28540 7528
rect 27893 7491 27951 7497
rect 28534 7488 28540 7500
rect 28592 7488 28598 7540
rect 28902 7488 28908 7540
rect 28960 7528 28966 7540
rect 29089 7531 29147 7537
rect 29089 7528 29101 7531
rect 28960 7500 29101 7528
rect 28960 7488 28966 7500
rect 29089 7497 29101 7500
rect 29135 7497 29147 7531
rect 29089 7491 29147 7497
rect 29178 7488 29184 7540
rect 29236 7528 29242 7540
rect 30377 7531 30435 7537
rect 29236 7500 30328 7528
rect 29236 7488 29242 7500
rect 15286 7420 15292 7472
rect 15344 7460 15350 7472
rect 15344 7432 22094 7460
rect 15344 7420 15350 7432
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 8662 7392 8668 7404
rect 1719 7364 8668 7392
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 22066 7324 22094 7432
rect 28994 7420 29000 7472
rect 29052 7460 29058 7472
rect 29733 7463 29791 7469
rect 29733 7460 29745 7463
rect 29052 7432 29745 7460
rect 29052 7420 29058 7432
rect 29733 7429 29745 7432
rect 29779 7429 29791 7463
rect 29733 7423 29791 7429
rect 30300 7404 30328 7500
rect 30377 7497 30389 7531
rect 30423 7528 30435 7531
rect 30742 7528 30748 7540
rect 30423 7500 30748 7528
rect 30423 7497 30435 7500
rect 30377 7491 30435 7497
rect 30742 7488 30748 7500
rect 30800 7488 30806 7540
rect 31018 7528 31024 7540
rect 30979 7500 31024 7528
rect 31018 7488 31024 7500
rect 31076 7488 31082 7540
rect 31754 7488 31760 7540
rect 31812 7528 31818 7540
rect 32125 7531 32183 7537
rect 32125 7528 32137 7531
rect 31812 7500 32137 7528
rect 31812 7488 31818 7500
rect 32125 7497 32137 7500
rect 32171 7497 32183 7531
rect 32674 7528 32680 7540
rect 32635 7500 32680 7528
rect 32125 7491 32183 7497
rect 32674 7488 32680 7500
rect 32732 7488 32738 7540
rect 33870 7528 33876 7540
rect 33831 7500 33876 7528
rect 33870 7488 33876 7500
rect 33928 7488 33934 7540
rect 34974 7528 34980 7540
rect 34935 7500 34980 7528
rect 34974 7488 34980 7500
rect 35032 7488 35038 7540
rect 36078 7528 36084 7540
rect 36039 7500 36084 7528
rect 36078 7488 36084 7500
rect 36136 7488 36142 7540
rect 58158 7528 58164 7540
rect 58119 7500 58164 7528
rect 58158 7488 58164 7500
rect 58216 7488 58222 7540
rect 32582 7420 32588 7472
rect 32640 7460 32646 7472
rect 33229 7463 33287 7469
rect 33229 7460 33241 7463
rect 32640 7432 33241 7460
rect 32640 7420 32646 7432
rect 33229 7429 33241 7432
rect 33275 7429 33287 7463
rect 33229 7423 33287 7429
rect 23382 7352 23388 7404
rect 23440 7392 23446 7404
rect 29638 7392 29644 7404
rect 23440 7364 29644 7392
rect 23440 7352 23446 7364
rect 29638 7352 29644 7364
rect 29696 7392 29702 7404
rect 29825 7395 29883 7401
rect 29825 7392 29837 7395
rect 29696 7364 29837 7392
rect 29696 7352 29702 7364
rect 29825 7361 29837 7364
rect 29871 7361 29883 7395
rect 30282 7392 30288 7404
rect 30195 7364 30288 7392
rect 29825 7355 29883 7361
rect 30282 7352 30288 7364
rect 30340 7352 30346 7404
rect 31113 7395 31171 7401
rect 31113 7361 31125 7395
rect 31159 7392 31171 7395
rect 32766 7392 32772 7404
rect 31159 7364 32772 7392
rect 31159 7361 31171 7364
rect 31113 7355 31171 7361
rect 32766 7352 32772 7364
rect 32824 7392 32830 7404
rect 37642 7392 37648 7404
rect 32824 7364 37648 7392
rect 32824 7352 32830 7364
rect 37642 7352 37648 7364
rect 37700 7352 37706 7404
rect 37182 7324 37188 7336
rect 22066 7296 37188 7324
rect 37182 7284 37188 7296
rect 37240 7284 37246 7336
rect 30466 7216 30472 7268
rect 30524 7256 30530 7268
rect 35250 7256 35256 7268
rect 30524 7228 35256 7256
rect 30524 7216 30530 7228
rect 35250 7216 35256 7228
rect 35308 7216 35314 7268
rect 35894 7216 35900 7268
rect 35952 7256 35958 7268
rect 36541 7259 36599 7265
rect 36541 7256 36553 7259
rect 35952 7228 36553 7256
rect 35952 7216 35958 7228
rect 36541 7225 36553 7228
rect 36587 7256 36599 7259
rect 36906 7256 36912 7268
rect 36587 7228 36912 7256
rect 36587 7225 36599 7228
rect 36541 7219 36599 7225
rect 36906 7216 36912 7228
rect 36964 7216 36970 7268
rect 1486 7188 1492 7200
rect 1447 7160 1492 7188
rect 1486 7148 1492 7160
rect 1544 7148 1550 7200
rect 26421 7191 26479 7197
rect 26421 7157 26433 7191
rect 26467 7188 26479 7191
rect 26694 7188 26700 7200
rect 26467 7160 26700 7188
rect 26467 7157 26479 7160
rect 26421 7151 26479 7157
rect 26694 7148 26700 7160
rect 26752 7188 26758 7200
rect 27246 7188 27252 7200
rect 26752 7160 27252 7188
rect 26752 7148 26758 7160
rect 27246 7148 27252 7160
rect 27304 7148 27310 7200
rect 34422 7188 34428 7200
rect 34383 7160 34428 7188
rect 34422 7148 34428 7160
rect 34480 7148 34486 7200
rect 35342 7148 35348 7200
rect 35400 7188 35406 7200
rect 35437 7191 35495 7197
rect 35437 7188 35449 7191
rect 35400 7160 35449 7188
rect 35400 7148 35406 7160
rect 35437 7157 35449 7160
rect 35483 7157 35495 7191
rect 35437 7151 35495 7157
rect 1104 7098 58880 7120
rect 1104 7046 10582 7098
rect 10634 7046 10646 7098
rect 10698 7046 10710 7098
rect 10762 7046 10774 7098
rect 10826 7046 10838 7098
rect 10890 7046 29846 7098
rect 29898 7046 29910 7098
rect 29962 7046 29974 7098
rect 30026 7046 30038 7098
rect 30090 7046 30102 7098
rect 30154 7046 49110 7098
rect 49162 7046 49174 7098
rect 49226 7046 49238 7098
rect 49290 7046 49302 7098
rect 49354 7046 49366 7098
rect 49418 7046 58880 7098
rect 1104 7024 58880 7046
rect 30834 6944 30840 6996
rect 30892 6984 30898 6996
rect 31021 6987 31079 6993
rect 31021 6984 31033 6987
rect 30892 6956 31033 6984
rect 30892 6944 30898 6956
rect 31021 6953 31033 6956
rect 31067 6953 31079 6987
rect 31021 6947 31079 6953
rect 31294 6944 31300 6996
rect 31352 6984 31358 6996
rect 31573 6987 31631 6993
rect 31573 6984 31585 6987
rect 31352 6956 31585 6984
rect 31352 6944 31358 6956
rect 31573 6953 31585 6956
rect 31619 6953 31631 6987
rect 31573 6947 31631 6953
rect 32582 6944 32588 6996
rect 32640 6984 32646 6996
rect 32677 6987 32735 6993
rect 32677 6984 32689 6987
rect 32640 6956 32689 6984
rect 32640 6944 32646 6956
rect 32677 6953 32689 6956
rect 32723 6953 32735 6987
rect 32677 6947 32735 6953
rect 24578 6808 24584 6860
rect 24636 6848 24642 6860
rect 29362 6848 29368 6860
rect 24636 6820 29368 6848
rect 24636 6808 24642 6820
rect 29362 6808 29368 6820
rect 29420 6808 29426 6860
rect 29730 6808 29736 6860
rect 29788 6848 29794 6860
rect 30469 6851 30527 6857
rect 30469 6848 30481 6851
rect 29788 6820 30481 6848
rect 29788 6808 29794 6820
rect 30469 6817 30481 6820
rect 30515 6817 30527 6851
rect 30469 6811 30527 6817
rect 33873 6851 33931 6857
rect 33873 6817 33885 6851
rect 33919 6848 33931 6851
rect 34054 6848 34060 6860
rect 33919 6820 34060 6848
rect 33919 6817 33931 6820
rect 33873 6811 33931 6817
rect 34054 6808 34060 6820
rect 34112 6808 34118 6860
rect 34238 6808 34244 6860
rect 34296 6848 34302 6860
rect 34701 6851 34759 6857
rect 34701 6848 34713 6851
rect 34296 6820 34713 6848
rect 34296 6808 34302 6820
rect 34701 6817 34713 6820
rect 34747 6817 34759 6851
rect 34701 6811 34759 6817
rect 16298 6740 16304 6792
rect 16356 6780 16362 6792
rect 28350 6780 28356 6792
rect 16356 6752 28356 6780
rect 16356 6740 16362 6752
rect 28350 6740 28356 6752
rect 28408 6780 28414 6792
rect 28902 6780 28908 6792
rect 28408 6752 28908 6780
rect 28408 6740 28414 6752
rect 28902 6740 28908 6752
rect 28960 6740 28966 6792
rect 28997 6783 29055 6789
rect 28997 6749 29009 6783
rect 29043 6780 29055 6783
rect 29270 6780 29276 6792
rect 29043 6752 29276 6780
rect 29043 6749 29055 6752
rect 28997 6743 29055 6749
rect 29270 6740 29276 6752
rect 29328 6740 29334 6792
rect 32217 6783 32275 6789
rect 32217 6749 32229 6783
rect 32263 6780 32275 6783
rect 33778 6780 33784 6792
rect 32263 6752 33784 6780
rect 32263 6749 32275 6752
rect 32217 6743 32275 6749
rect 33778 6740 33784 6752
rect 33836 6740 33842 6792
rect 34422 6740 34428 6792
rect 34480 6780 34486 6792
rect 45646 6780 45652 6792
rect 34480 6752 45652 6780
rect 34480 6740 34486 6752
rect 45646 6740 45652 6752
rect 45704 6740 45710 6792
rect 22738 6672 22744 6724
rect 22796 6712 22802 6724
rect 27246 6712 27252 6724
rect 22796 6684 26924 6712
rect 27207 6684 27252 6712
rect 22796 6672 22802 6684
rect 26234 6644 26240 6656
rect 26195 6616 26240 6644
rect 26234 6604 26240 6616
rect 26292 6604 26298 6656
rect 26786 6644 26792 6656
rect 26747 6616 26792 6644
rect 26786 6604 26792 6616
rect 26844 6604 26850 6656
rect 26896 6644 26924 6684
rect 27246 6672 27252 6684
rect 27304 6672 27310 6724
rect 27338 6672 27344 6724
rect 27396 6712 27402 6724
rect 27893 6715 27951 6721
rect 27893 6712 27905 6715
rect 27396 6684 27905 6712
rect 27396 6672 27402 6684
rect 27893 6681 27905 6684
rect 27939 6681 27951 6715
rect 27893 6675 27951 6681
rect 28626 6672 28632 6724
rect 28684 6712 28690 6724
rect 29917 6715 29975 6721
rect 29917 6712 29929 6715
rect 28684 6684 29929 6712
rect 28684 6672 28690 6684
rect 29917 6681 29929 6684
rect 29963 6681 29975 6715
rect 31938 6712 31944 6724
rect 29917 6675 29975 6681
rect 30024 6684 31944 6712
rect 30024 6644 30052 6684
rect 31938 6672 31944 6684
rect 31996 6672 32002 6724
rect 32030 6672 32036 6724
rect 32088 6712 32094 6724
rect 41874 6712 41880 6724
rect 32088 6684 41880 6712
rect 32088 6672 32094 6684
rect 41874 6672 41880 6684
rect 41932 6672 41938 6724
rect 26896 6616 30052 6644
rect 33321 6647 33379 6653
rect 33321 6613 33333 6647
rect 33367 6644 33379 6647
rect 33410 6644 33416 6656
rect 33367 6616 33416 6644
rect 33367 6613 33379 6616
rect 33321 6607 33379 6613
rect 33410 6604 33416 6616
rect 33468 6604 33474 6656
rect 35342 6644 35348 6656
rect 35303 6616 35348 6644
rect 35342 6604 35348 6616
rect 35400 6604 35406 6656
rect 35894 6644 35900 6656
rect 35855 6616 35900 6644
rect 35894 6604 35900 6616
rect 35952 6604 35958 6656
rect 1104 6554 58880 6576
rect 1104 6502 20214 6554
rect 20266 6502 20278 6554
rect 20330 6502 20342 6554
rect 20394 6502 20406 6554
rect 20458 6502 20470 6554
rect 20522 6502 39478 6554
rect 39530 6502 39542 6554
rect 39594 6502 39606 6554
rect 39658 6502 39670 6554
rect 39722 6502 39734 6554
rect 39786 6502 58880 6554
rect 1104 6480 58880 6502
rect 28261 6443 28319 6449
rect 28261 6409 28273 6443
rect 28307 6440 28319 6443
rect 29362 6440 29368 6452
rect 28307 6412 29368 6440
rect 28307 6409 28319 6412
rect 28261 6403 28319 6409
rect 29362 6400 29368 6412
rect 29420 6400 29426 6452
rect 30190 6440 30196 6452
rect 30151 6412 30196 6440
rect 30190 6400 30196 6412
rect 30248 6400 30254 6452
rect 30558 6400 30564 6452
rect 30616 6440 30622 6452
rect 30653 6443 30711 6449
rect 30653 6440 30665 6443
rect 30616 6412 30665 6440
rect 30616 6400 30622 6412
rect 30653 6409 30665 6412
rect 30699 6409 30711 6443
rect 32122 6440 32128 6452
rect 32083 6412 32128 6440
rect 30653 6403 30711 6409
rect 32122 6400 32128 6412
rect 32180 6400 32186 6452
rect 32766 6440 32772 6452
rect 32727 6412 32772 6440
rect 32766 6400 32772 6412
rect 32824 6400 32830 6452
rect 34425 6443 34483 6449
rect 34425 6409 34437 6443
rect 34471 6440 34483 6443
rect 34977 6443 35035 6449
rect 34977 6440 34989 6443
rect 34471 6412 34989 6440
rect 34471 6409 34483 6412
rect 34425 6403 34483 6409
rect 34977 6409 34989 6412
rect 35023 6440 35035 6443
rect 36078 6440 36084 6452
rect 35023 6412 36084 6440
rect 35023 6409 35035 6412
rect 34977 6403 35035 6409
rect 36078 6400 36084 6412
rect 36136 6400 36142 6452
rect 27982 6332 27988 6384
rect 28040 6372 28046 6384
rect 28721 6375 28779 6381
rect 28721 6372 28733 6375
rect 28040 6344 28733 6372
rect 28040 6332 28046 6344
rect 28721 6341 28733 6344
rect 28767 6341 28779 6375
rect 28721 6335 28779 6341
rect 28902 6332 28908 6384
rect 28960 6372 28966 6384
rect 29273 6375 29331 6381
rect 29273 6372 29285 6375
rect 28960 6344 29285 6372
rect 28960 6332 28966 6344
rect 29273 6341 29285 6344
rect 29319 6341 29331 6375
rect 29273 6335 29331 6341
rect 29638 6332 29644 6384
rect 29696 6372 29702 6384
rect 34238 6372 34244 6384
rect 29696 6344 34244 6372
rect 29696 6332 29702 6344
rect 34238 6332 34244 6344
rect 34296 6332 34302 6384
rect 26786 6264 26792 6316
rect 26844 6304 26850 6316
rect 33229 6307 33287 6313
rect 33229 6304 33241 6307
rect 26844 6276 33241 6304
rect 26844 6264 26850 6276
rect 33229 6273 33241 6276
rect 33275 6304 33287 6307
rect 33781 6307 33839 6313
rect 33781 6304 33793 6307
rect 33275 6276 33793 6304
rect 33275 6273 33287 6276
rect 33229 6267 33287 6273
rect 33781 6273 33793 6276
rect 33827 6304 33839 6307
rect 35342 6304 35348 6316
rect 33827 6276 35348 6304
rect 33827 6273 33839 6276
rect 33781 6267 33839 6273
rect 35342 6264 35348 6276
rect 35400 6304 35406 6316
rect 35437 6307 35495 6313
rect 35437 6304 35449 6307
rect 35400 6276 35449 6304
rect 35400 6264 35406 6276
rect 35437 6273 35449 6276
rect 35483 6273 35495 6307
rect 35437 6267 35495 6273
rect 27246 6196 27252 6248
rect 27304 6236 27310 6248
rect 36630 6236 36636 6248
rect 27304 6208 36636 6236
rect 27304 6196 27310 6208
rect 36630 6196 36636 6208
rect 36688 6196 36694 6248
rect 15746 6128 15752 6180
rect 15804 6168 15810 6180
rect 30650 6168 30656 6180
rect 15804 6140 30656 6168
rect 15804 6128 15810 6140
rect 30650 6128 30656 6140
rect 30708 6168 30714 6180
rect 31205 6171 31263 6177
rect 31205 6168 31217 6171
rect 30708 6140 31217 6168
rect 30708 6128 30714 6140
rect 31205 6137 31217 6140
rect 31251 6137 31263 6171
rect 31205 6131 31263 6137
rect 31938 6128 31944 6180
rect 31996 6168 32002 6180
rect 39114 6168 39120 6180
rect 31996 6140 39120 6168
rect 31996 6128 32002 6140
rect 39114 6128 39120 6140
rect 39172 6128 39178 6180
rect 26234 6060 26240 6112
rect 26292 6100 26298 6112
rect 27338 6100 27344 6112
rect 26292 6072 27344 6100
rect 26292 6060 26298 6072
rect 27338 6060 27344 6072
rect 27396 6060 27402 6112
rect 1104 6010 58880 6032
rect 1104 5958 10582 6010
rect 10634 5958 10646 6010
rect 10698 5958 10710 6010
rect 10762 5958 10774 6010
rect 10826 5958 10838 6010
rect 10890 5958 29846 6010
rect 29898 5958 29910 6010
rect 29962 5958 29974 6010
rect 30026 5958 30038 6010
rect 30090 5958 30102 6010
rect 30154 5958 49110 6010
rect 49162 5958 49174 6010
rect 49226 5958 49238 6010
rect 49290 5958 49302 6010
rect 49354 5958 49366 6010
rect 49418 5958 58880 6010
rect 1104 5936 58880 5958
rect 28442 5896 28448 5908
rect 28403 5868 28448 5896
rect 28442 5856 28448 5868
rect 28500 5856 28506 5908
rect 28810 5856 28816 5908
rect 28868 5896 28874 5908
rect 28997 5899 29055 5905
rect 28997 5896 29009 5899
rect 28868 5868 29009 5896
rect 28868 5856 28874 5868
rect 28997 5865 29009 5868
rect 29043 5865 29055 5899
rect 29638 5896 29644 5908
rect 29599 5868 29644 5896
rect 28997 5859 29055 5865
rect 29638 5856 29644 5868
rect 29696 5856 29702 5908
rect 30193 5899 30251 5905
rect 30193 5865 30205 5899
rect 30239 5896 30251 5899
rect 30282 5896 30288 5908
rect 30239 5868 30288 5896
rect 30239 5865 30251 5868
rect 30193 5859 30251 5865
rect 30282 5856 30288 5868
rect 30340 5856 30346 5908
rect 30466 5856 30472 5908
rect 30524 5896 30530 5908
rect 30653 5899 30711 5905
rect 30653 5896 30665 5899
rect 30524 5868 30665 5896
rect 30524 5856 30530 5868
rect 30653 5865 30665 5868
rect 30699 5865 30711 5899
rect 30653 5859 30711 5865
rect 31110 5856 31116 5908
rect 31168 5896 31174 5908
rect 31205 5899 31263 5905
rect 31205 5896 31217 5899
rect 31168 5868 31217 5896
rect 31168 5856 31174 5868
rect 31205 5865 31217 5868
rect 31251 5865 31263 5899
rect 31205 5859 31263 5865
rect 32214 5856 32220 5908
rect 32272 5896 32278 5908
rect 32401 5899 32459 5905
rect 32401 5896 32413 5899
rect 32272 5868 32413 5896
rect 32272 5856 32278 5868
rect 32401 5865 32413 5868
rect 32447 5896 32459 5899
rect 36354 5896 36360 5908
rect 32447 5868 36360 5896
rect 32447 5865 32459 5868
rect 32401 5859 32459 5865
rect 36354 5856 36360 5868
rect 36412 5856 36418 5908
rect 32858 5828 32864 5840
rect 32819 5800 32864 5828
rect 32858 5788 32864 5800
rect 32916 5788 32922 5840
rect 33502 5828 33508 5840
rect 33463 5800 33508 5828
rect 33502 5788 33508 5800
rect 33560 5788 33566 5840
rect 34057 5831 34115 5837
rect 34057 5797 34069 5831
rect 34103 5828 34115 5831
rect 35894 5828 35900 5840
rect 34103 5800 35900 5828
rect 34103 5797 34115 5800
rect 34057 5791 34115 5797
rect 35894 5788 35900 5800
rect 35952 5788 35958 5840
rect 14458 5760 14464 5772
rect 6886 5732 14464 5760
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5692 1731 5695
rect 6886 5692 6914 5732
rect 14458 5720 14464 5732
rect 14516 5720 14522 5772
rect 31849 5763 31907 5769
rect 31849 5729 31861 5763
rect 31895 5760 31907 5763
rect 32766 5760 32772 5772
rect 31895 5732 32772 5760
rect 31895 5729 31907 5732
rect 31849 5723 31907 5729
rect 32766 5720 32772 5732
rect 32824 5720 32830 5772
rect 1719 5664 6914 5692
rect 13541 5695 13599 5701
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 13541 5661 13553 5695
rect 13587 5692 13599 5695
rect 58158 5692 58164 5704
rect 13587 5664 14228 5692
rect 58119 5664 58164 5692
rect 13587 5661 13599 5664
rect 13541 5655 13599 5661
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 8846 5516 8852 5568
rect 8904 5556 8910 5568
rect 14200 5565 14228 5664
rect 58158 5652 58164 5664
rect 58216 5652 58222 5704
rect 37182 5584 37188 5636
rect 37240 5624 37246 5636
rect 57885 5627 57943 5633
rect 57885 5624 57897 5627
rect 37240 5596 57897 5624
rect 37240 5584 37246 5596
rect 57885 5593 57897 5596
rect 57931 5593 57943 5627
rect 57885 5587 57943 5593
rect 13357 5559 13415 5565
rect 13357 5556 13369 5559
rect 8904 5528 13369 5556
rect 8904 5516 8910 5528
rect 13357 5525 13369 5528
rect 13403 5525 13415 5559
rect 13357 5519 13415 5525
rect 14185 5559 14243 5565
rect 14185 5525 14197 5559
rect 14231 5556 14243 5559
rect 22002 5556 22008 5568
rect 14231 5528 22008 5556
rect 14231 5525 14243 5528
rect 14185 5519 14243 5525
rect 22002 5516 22008 5528
rect 22060 5516 22066 5568
rect 1104 5466 58880 5488
rect 1104 5414 20214 5466
rect 20266 5414 20278 5466
rect 20330 5414 20342 5466
rect 20394 5414 20406 5466
rect 20458 5414 20470 5466
rect 20522 5414 39478 5466
rect 39530 5414 39542 5466
rect 39594 5414 39606 5466
rect 39658 5414 39670 5466
rect 39722 5414 39734 5466
rect 39786 5414 58880 5466
rect 1104 5392 58880 5414
rect 18414 5312 18420 5364
rect 18472 5352 18478 5364
rect 29454 5352 29460 5364
rect 18472 5324 26924 5352
rect 29415 5324 29460 5352
rect 18472 5312 18478 5324
rect 14918 5244 14924 5296
rect 14976 5284 14982 5296
rect 26896 5284 26924 5324
rect 29454 5312 29460 5324
rect 29512 5312 29518 5364
rect 30374 5312 30380 5364
rect 30432 5352 30438 5364
rect 30469 5355 30527 5361
rect 30469 5352 30481 5355
rect 30432 5324 30481 5352
rect 30432 5312 30438 5324
rect 30469 5321 30481 5324
rect 30515 5352 30527 5355
rect 30558 5352 30564 5364
rect 30515 5324 30564 5352
rect 30515 5321 30527 5324
rect 30469 5315 30527 5321
rect 30558 5312 30564 5324
rect 30616 5312 30622 5364
rect 41782 5352 41788 5364
rect 30668 5324 41788 5352
rect 30668 5284 30696 5324
rect 41782 5312 41788 5324
rect 41840 5312 41846 5364
rect 58158 5352 58164 5364
rect 58119 5324 58164 5352
rect 58158 5312 58164 5324
rect 58216 5312 58222 5364
rect 32214 5284 32220 5296
rect 14976 5256 22094 5284
rect 26896 5256 30696 5284
rect 31726 5256 32220 5284
rect 14976 5244 14982 5256
rect 22066 5080 22094 5256
rect 27338 5176 27344 5228
rect 27396 5216 27402 5228
rect 28905 5219 28963 5225
rect 28905 5216 28917 5219
rect 27396 5188 28917 5216
rect 27396 5176 27402 5188
rect 28905 5185 28917 5188
rect 28951 5216 28963 5219
rect 30009 5219 30067 5225
rect 30009 5216 30021 5219
rect 28951 5188 30021 5216
rect 28951 5185 28963 5188
rect 28905 5179 28963 5185
rect 30009 5185 30021 5188
rect 30055 5216 30067 5219
rect 31726 5216 31754 5256
rect 32214 5244 32220 5256
rect 32272 5244 32278 5296
rect 30055 5188 31754 5216
rect 30055 5185 30067 5188
rect 30009 5179 30067 5185
rect 37274 5080 37280 5092
rect 22066 5052 37280 5080
rect 37274 5040 37280 5052
rect 37332 5040 37338 5092
rect 1104 4922 58880 4944
rect 1104 4870 10582 4922
rect 10634 4870 10646 4922
rect 10698 4870 10710 4922
rect 10762 4870 10774 4922
rect 10826 4870 10838 4922
rect 10890 4870 29846 4922
rect 29898 4870 29910 4922
rect 29962 4870 29974 4922
rect 30026 4870 30038 4922
rect 30090 4870 30102 4922
rect 30154 4870 49110 4922
rect 49162 4870 49174 4922
rect 49226 4870 49238 4922
rect 49290 4870 49302 4922
rect 49354 4870 49366 4922
rect 49418 4870 58880 4922
rect 1104 4848 58880 4870
rect 29546 4808 29552 4820
rect 29507 4780 29552 4808
rect 29546 4768 29552 4780
rect 29604 4768 29610 4820
rect 58069 4607 58127 4613
rect 58069 4573 58081 4607
rect 58115 4604 58127 4607
rect 58158 4604 58164 4616
rect 58115 4576 58164 4604
rect 58115 4573 58127 4576
rect 58069 4567 58127 4573
rect 58158 4564 58164 4576
rect 58216 4564 58222 4616
rect 41690 4496 41696 4548
rect 41748 4536 41754 4548
rect 57517 4539 57575 4545
rect 57517 4536 57529 4539
rect 41748 4508 57529 4536
rect 41748 4496 41754 4508
rect 57517 4505 57529 4508
rect 57563 4505 57575 4539
rect 57517 4499 57575 4505
rect 1104 4378 58880 4400
rect 1104 4326 20214 4378
rect 20266 4326 20278 4378
rect 20330 4326 20342 4378
rect 20394 4326 20406 4378
rect 20458 4326 20470 4378
rect 20522 4326 39478 4378
rect 39530 4326 39542 4378
rect 39594 4326 39606 4378
rect 39658 4326 39670 4378
rect 39722 4326 39734 4378
rect 39786 4326 58880 4378
rect 1104 4304 58880 4326
rect 58158 4264 58164 4276
rect 58119 4236 58164 4264
rect 58158 4224 58164 4236
rect 58216 4224 58222 4276
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 1719 4100 2268 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 2240 4001 2268 4100
rect 16114 4088 16120 4140
rect 16172 4128 16178 4140
rect 47118 4128 47124 4140
rect 16172 4100 47124 4128
rect 16172 4088 16178 4100
rect 47118 4088 47124 4100
rect 47176 4088 47182 4140
rect 19242 4020 19248 4072
rect 19300 4060 19306 4072
rect 45094 4060 45100 4072
rect 19300 4032 45100 4060
rect 19300 4020 19306 4032
rect 45094 4020 45100 4032
rect 45152 4020 45158 4072
rect 2225 3995 2283 4001
rect 2225 3961 2237 3995
rect 2271 3992 2283 3995
rect 20990 3992 20996 4004
rect 2271 3964 20996 3992
rect 2271 3961 2283 3964
rect 2225 3955 2283 3961
rect 20990 3952 20996 3964
rect 21048 3952 21054 4004
rect 23566 3952 23572 4004
rect 23624 3992 23630 4004
rect 48498 3992 48504 4004
rect 23624 3964 48504 3992
rect 23624 3952 23630 3964
rect 48498 3952 48504 3964
rect 48556 3952 48562 4004
rect 1486 3924 1492 3936
rect 1447 3896 1492 3924
rect 1486 3884 1492 3896
rect 1544 3884 1550 3936
rect 1104 3834 58880 3856
rect 1104 3782 10582 3834
rect 10634 3782 10646 3834
rect 10698 3782 10710 3834
rect 10762 3782 10774 3834
rect 10826 3782 10838 3834
rect 10890 3782 29846 3834
rect 29898 3782 29910 3834
rect 29962 3782 29974 3834
rect 30026 3782 30038 3834
rect 30090 3782 30102 3834
rect 30154 3782 49110 3834
rect 49162 3782 49174 3834
rect 49226 3782 49238 3834
rect 49290 3782 49302 3834
rect 49354 3782 49366 3834
rect 49418 3782 58880 3834
rect 1104 3760 58880 3782
rect 40037 3655 40095 3661
rect 40037 3621 40049 3655
rect 40083 3652 40095 3655
rect 42426 3652 42432 3664
rect 40083 3624 42432 3652
rect 40083 3621 40095 3624
rect 40037 3615 40095 3621
rect 42426 3612 42432 3624
rect 42484 3612 42490 3664
rect 37826 3476 37832 3528
rect 37884 3516 37890 3528
rect 39853 3519 39911 3525
rect 39853 3516 39865 3519
rect 37884 3488 39865 3516
rect 37884 3476 37890 3488
rect 39853 3485 39865 3488
rect 39899 3516 39911 3519
rect 40497 3519 40555 3525
rect 40497 3516 40509 3519
rect 39899 3488 40509 3516
rect 39899 3485 39911 3488
rect 39853 3479 39911 3485
rect 40497 3485 40509 3488
rect 40543 3485 40555 3519
rect 40497 3479 40555 3485
rect 1104 3290 58880 3312
rect 1104 3238 20214 3290
rect 20266 3238 20278 3290
rect 20330 3238 20342 3290
rect 20394 3238 20406 3290
rect 20458 3238 20470 3290
rect 20522 3238 39478 3290
rect 39530 3238 39542 3290
rect 39594 3238 39606 3290
rect 39658 3238 39670 3290
rect 39722 3238 39734 3290
rect 39786 3238 58880 3290
rect 1104 3216 58880 3238
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3040 1639 3043
rect 8846 3040 8852 3052
rect 1627 3012 8852 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 8846 3000 8852 3012
rect 8904 3000 8910 3052
rect 37734 3040 37740 3052
rect 37695 3012 37740 3040
rect 37734 3000 37740 3012
rect 37792 3000 37798 3052
rect 37918 2904 37924 2916
rect 37879 2876 37924 2904
rect 37918 2864 37924 2876
rect 37976 2864 37982 2916
rect 1394 2836 1400 2848
rect 1355 2808 1400 2836
rect 1394 2796 1400 2808
rect 1452 2796 1458 2848
rect 1104 2746 58880 2768
rect 1104 2694 10582 2746
rect 10634 2694 10646 2746
rect 10698 2694 10710 2746
rect 10762 2694 10774 2746
rect 10826 2694 10838 2746
rect 10890 2694 29846 2746
rect 29898 2694 29910 2746
rect 29962 2694 29974 2746
rect 30026 2694 30038 2746
rect 30090 2694 30102 2746
rect 30154 2694 49110 2746
rect 49162 2694 49174 2746
rect 49226 2694 49238 2746
rect 49290 2694 49302 2746
rect 49354 2694 49366 2746
rect 49418 2694 58880 2746
rect 1104 2672 58880 2694
rect 30558 2592 30564 2644
rect 30616 2632 30622 2644
rect 56502 2632 56508 2644
rect 30616 2604 56508 2632
rect 30616 2592 30622 2604
rect 56502 2592 56508 2604
rect 56560 2592 56566 2644
rect 12894 2564 12900 2576
rect 6886 2536 12900 2564
rect 4525 2499 4583 2505
rect 4525 2465 4537 2499
rect 4571 2496 4583 2499
rect 6886 2496 6914 2536
rect 12894 2524 12900 2536
rect 12952 2524 12958 2576
rect 17954 2524 17960 2576
rect 18012 2564 18018 2576
rect 46934 2564 46940 2576
rect 18012 2536 46940 2564
rect 18012 2524 18018 2536
rect 46934 2524 46940 2536
rect 46992 2524 46998 2576
rect 4571 2468 6914 2496
rect 7193 2499 7251 2505
rect 4571 2465 4583 2468
rect 4525 2459 4583 2465
rect 7193 2465 7205 2499
rect 7239 2496 7251 2499
rect 24854 2496 24860 2508
rect 7239 2468 24860 2496
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2428 1731 2431
rect 3973 2431 4031 2437
rect 1719 2400 3832 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 1486 2292 1492 2304
rect 1447 2264 1492 2292
rect 1486 2252 1492 2264
rect 1544 2252 1550 2304
rect 3804 2301 3832 2400
rect 3973 2397 3985 2431
rect 4019 2428 4031 2431
rect 4540 2428 4568 2459
rect 4019 2400 4568 2428
rect 6641 2431 6699 2437
rect 4019 2397 4031 2400
rect 3973 2391 4031 2397
rect 6641 2397 6653 2431
rect 6687 2428 6699 2431
rect 7208 2428 7236 2459
rect 24854 2456 24860 2468
rect 24912 2456 24918 2508
rect 25866 2456 25872 2508
rect 25924 2496 25930 2508
rect 48774 2496 48780 2508
rect 25924 2468 48780 2496
rect 25924 2456 25930 2468
rect 48774 2456 48780 2468
rect 48832 2456 48838 2508
rect 6687 2400 7236 2428
rect 18325 2431 18383 2437
rect 6687 2397 6699 2400
rect 6641 2391 6699 2397
rect 18325 2397 18337 2431
rect 18371 2428 18383 2431
rect 18371 2400 19380 2428
rect 18371 2397 18383 2400
rect 18325 2391 18383 2397
rect 19352 2369 19380 2400
rect 29914 2388 29920 2440
rect 29972 2428 29978 2440
rect 30009 2431 30067 2437
rect 30009 2428 30021 2431
rect 29972 2400 30021 2428
rect 29972 2388 29978 2400
rect 30009 2397 30021 2400
rect 30055 2428 30067 2431
rect 30653 2431 30711 2437
rect 30653 2428 30665 2431
rect 30055 2400 30665 2428
rect 30055 2397 30067 2400
rect 30009 2391 30067 2397
rect 30653 2397 30665 2400
rect 30699 2397 30711 2431
rect 30653 2391 30711 2397
rect 37553 2431 37611 2437
rect 37553 2397 37565 2431
rect 37599 2428 37611 2431
rect 37734 2428 37740 2440
rect 37599 2400 37740 2428
rect 37599 2397 37611 2400
rect 37553 2391 37611 2397
rect 37734 2388 37740 2400
rect 37792 2388 37798 2440
rect 42426 2428 42432 2440
rect 42387 2400 42432 2428
rect 42426 2388 42432 2400
rect 42484 2388 42490 2440
rect 54021 2431 54079 2437
rect 54021 2428 54033 2431
rect 45526 2400 54033 2428
rect 19337 2363 19395 2369
rect 19337 2329 19349 2363
rect 19383 2360 19395 2363
rect 37826 2360 37832 2372
rect 19383 2332 37832 2360
rect 19383 2329 19395 2332
rect 19337 2323 19395 2329
rect 37826 2320 37832 2332
rect 37884 2320 37890 2372
rect 37918 2320 37924 2372
rect 37976 2360 37982 2372
rect 45526 2360 45554 2400
rect 54021 2397 54033 2400
rect 54067 2397 54079 2431
rect 54021 2391 54079 2397
rect 57333 2431 57391 2437
rect 57333 2397 57345 2431
rect 57379 2428 57391 2431
rect 57379 2400 57928 2428
rect 57379 2397 57391 2400
rect 57333 2391 57391 2397
rect 37976 2332 45554 2360
rect 37976 2320 37982 2332
rect 46198 2320 46204 2372
rect 46256 2360 46262 2372
rect 56137 2363 56195 2369
rect 56137 2360 56149 2363
rect 46256 2332 56149 2360
rect 46256 2320 46262 2332
rect 56137 2329 56149 2332
rect 56183 2329 56195 2363
rect 56137 2323 56195 2329
rect 57900 2304 57928 2400
rect 3789 2295 3847 2301
rect 3789 2261 3801 2295
rect 3835 2261 3847 2295
rect 3789 2255 3847 2261
rect 5994 2252 6000 2304
rect 6052 2292 6058 2304
rect 6457 2295 6515 2301
rect 6457 2292 6469 2295
rect 6052 2264 6469 2292
rect 6052 2252 6058 2264
rect 6457 2261 6469 2264
rect 6503 2261 6515 2295
rect 6457 2255 6515 2261
rect 17954 2252 17960 2304
rect 18012 2292 18018 2304
rect 18141 2295 18199 2301
rect 18141 2292 18153 2295
rect 18012 2264 18153 2292
rect 18012 2252 18018 2264
rect 18141 2261 18153 2264
rect 18187 2261 18199 2295
rect 18141 2255 18199 2261
rect 30193 2295 30251 2301
rect 30193 2261 30205 2295
rect 30239 2292 30251 2295
rect 31202 2292 31208 2304
rect 30239 2264 31208 2292
rect 30239 2261 30251 2264
rect 30193 2255 30251 2261
rect 31202 2252 31208 2264
rect 31260 2252 31266 2304
rect 41966 2252 41972 2304
rect 42024 2292 42030 2304
rect 42613 2295 42671 2301
rect 42613 2292 42625 2295
rect 42024 2264 42625 2292
rect 42024 2252 42030 2264
rect 42613 2261 42625 2264
rect 42659 2261 42671 2295
rect 42613 2255 42671 2261
rect 53926 2252 53932 2304
rect 53984 2292 53990 2304
rect 54205 2295 54263 2301
rect 54205 2292 54217 2295
rect 53984 2264 54217 2292
rect 53984 2252 53990 2264
rect 54205 2261 54217 2264
rect 54251 2261 54263 2295
rect 57882 2292 57888 2304
rect 57843 2264 57888 2292
rect 54205 2255 54263 2261
rect 57882 2252 57888 2264
rect 57940 2252 57946 2304
rect 1104 2202 58880 2224
rect 1104 2150 20214 2202
rect 20266 2150 20278 2202
rect 20330 2150 20342 2202
rect 20394 2150 20406 2202
rect 20458 2150 20470 2202
rect 20522 2150 39478 2202
rect 39530 2150 39542 2202
rect 39594 2150 39606 2202
rect 39658 2150 39670 2202
rect 39722 2150 39734 2202
rect 39786 2150 58880 2202
rect 1104 2128 58880 2150
rect 24394 2048 24400 2100
rect 24452 2088 24458 2100
rect 45370 2088 45376 2100
rect 24452 2060 45376 2088
rect 24452 2048 24458 2060
rect 45370 2048 45376 2060
rect 45428 2048 45434 2100
rect 25498 1980 25504 2032
rect 25556 2020 25562 2032
rect 45462 2020 45468 2032
rect 25556 1992 45468 2020
rect 25556 1980 25562 1992
rect 45462 1980 45468 1992
rect 45520 1980 45526 2032
rect 26050 1912 26056 1964
rect 26108 1952 26114 1964
rect 48406 1952 48412 1964
rect 26108 1924 48412 1952
rect 26108 1912 26114 1924
rect 48406 1912 48412 1924
rect 48464 1912 48470 1964
<< via1 >>
rect 17224 28160 17276 28212
rect 32312 28160 32364 28212
rect 14648 28092 14700 28144
rect 38200 28092 38252 28144
rect 41420 28092 41472 28144
rect 18788 28024 18840 28076
rect 32864 28024 32916 28076
rect 19064 27956 19116 28008
rect 37464 27956 37516 28008
rect 23940 27888 23992 27940
rect 44272 27888 44324 27940
rect 14096 27820 14148 27872
rect 37372 27820 37424 27872
rect 10582 27718 10634 27770
rect 10646 27718 10698 27770
rect 10710 27718 10762 27770
rect 10774 27718 10826 27770
rect 10838 27718 10890 27770
rect 29846 27718 29898 27770
rect 29910 27718 29962 27770
rect 29974 27718 30026 27770
rect 30038 27718 30090 27770
rect 30102 27718 30154 27770
rect 49110 27718 49162 27770
rect 49174 27718 49226 27770
rect 49238 27718 49290 27770
rect 49302 27718 49354 27770
rect 49366 27718 49418 27770
rect 30288 27616 30340 27668
rect 39856 27616 39908 27668
rect 1492 27591 1544 27600
rect 1492 27557 1501 27591
rect 1501 27557 1535 27591
rect 1535 27557 1544 27591
rect 1492 27548 1544 27557
rect 2780 27548 2832 27600
rect 8300 27548 8352 27600
rect 3884 27412 3936 27464
rect 14372 27480 14424 27532
rect 13820 27412 13872 27464
rect 19524 27455 19576 27464
rect 19524 27421 19533 27455
rect 19533 27421 19567 27455
rect 19567 27421 19576 27455
rect 19524 27412 19576 27421
rect 19984 27455 20036 27464
rect 19984 27421 19993 27455
rect 19993 27421 20027 27455
rect 20027 27421 20036 27455
rect 19984 27412 20036 27421
rect 24492 27548 24544 27600
rect 30196 27548 30248 27600
rect 30748 27548 30800 27600
rect 35348 27548 35400 27600
rect 35624 27591 35676 27600
rect 35624 27557 35633 27591
rect 35633 27557 35667 27591
rect 35667 27557 35676 27591
rect 35624 27548 35676 27557
rect 52000 27591 52052 27600
rect 52000 27557 52009 27591
rect 52009 27557 52043 27591
rect 52043 27557 52052 27591
rect 52000 27548 52052 27557
rect 18420 27344 18472 27396
rect 20628 27387 20680 27396
rect 3884 27319 3936 27328
rect 3884 27285 3893 27319
rect 3893 27285 3927 27319
rect 3927 27285 3936 27319
rect 3884 27276 3936 27285
rect 9772 27319 9824 27328
rect 9772 27285 9781 27319
rect 9781 27285 9815 27319
rect 9815 27285 9824 27319
rect 9772 27276 9824 27285
rect 14280 27319 14332 27328
rect 14280 27285 14289 27319
rect 14289 27285 14323 27319
rect 14323 27285 14332 27319
rect 14280 27276 14332 27285
rect 19340 27319 19392 27328
rect 19340 27285 19349 27319
rect 19349 27285 19383 27319
rect 19383 27285 19392 27319
rect 19340 27276 19392 27285
rect 20628 27353 20637 27387
rect 20637 27353 20671 27387
rect 20671 27353 20680 27387
rect 20628 27344 20680 27353
rect 33508 27480 33560 27532
rect 28632 27412 28684 27464
rect 30380 27412 30432 27464
rect 29644 27344 29696 27396
rect 32128 27344 32180 27396
rect 34152 27387 34204 27396
rect 34152 27353 34161 27387
rect 34161 27353 34195 27387
rect 34195 27353 34204 27387
rect 34152 27344 34204 27353
rect 25780 27319 25832 27328
rect 25780 27285 25789 27319
rect 25789 27285 25823 27319
rect 25823 27285 25832 27319
rect 25780 27276 25832 27285
rect 26424 27319 26476 27328
rect 26424 27285 26433 27319
rect 26433 27285 26467 27319
rect 26467 27285 26476 27319
rect 26424 27276 26476 27285
rect 28540 27319 28592 27328
rect 28540 27285 28549 27319
rect 28549 27285 28583 27319
rect 28583 27285 28592 27319
rect 28540 27276 28592 27285
rect 31576 27276 31628 27328
rect 32864 27276 32916 27328
rect 33140 27276 33192 27328
rect 40868 27455 40920 27464
rect 40868 27421 40877 27455
rect 40877 27421 40911 27455
rect 40911 27421 40920 27455
rect 40868 27412 40920 27421
rect 46388 27455 46440 27464
rect 46388 27421 46397 27455
rect 46397 27421 46431 27455
rect 46431 27421 46440 27455
rect 46388 27412 46440 27421
rect 46480 27412 46532 27464
rect 52460 27412 52512 27464
rect 57244 27455 57296 27464
rect 57244 27421 57253 27455
rect 57253 27421 57287 27455
rect 57287 27421 57296 27455
rect 57244 27412 57296 27421
rect 57888 27387 57940 27396
rect 57888 27353 57897 27387
rect 57897 27353 57931 27387
rect 57931 27353 57940 27387
rect 57888 27344 57940 27353
rect 58072 27387 58124 27396
rect 58072 27353 58081 27387
rect 58081 27353 58115 27387
rect 58115 27353 58124 27387
rect 58072 27344 58124 27353
rect 41052 27319 41104 27328
rect 41052 27285 41061 27319
rect 41061 27285 41095 27319
rect 41095 27285 41104 27319
rect 41052 27276 41104 27285
rect 46296 27276 46348 27328
rect 20214 27174 20266 27226
rect 20278 27174 20330 27226
rect 20342 27174 20394 27226
rect 20406 27174 20458 27226
rect 20470 27174 20522 27226
rect 39478 27174 39530 27226
rect 39542 27174 39594 27226
rect 39606 27174 39658 27226
rect 39670 27174 39722 27226
rect 39734 27174 39786 27226
rect 1400 27072 1452 27124
rect 9772 27072 9824 27124
rect 14464 26936 14516 26988
rect 19524 27072 19576 27124
rect 25780 27115 25832 27124
rect 25780 27081 25789 27115
rect 25789 27081 25823 27115
rect 25823 27081 25832 27115
rect 25780 27072 25832 27081
rect 34060 27115 34112 27124
rect 34060 27081 34069 27115
rect 34069 27081 34103 27115
rect 34103 27081 34112 27115
rect 34060 27072 34112 27081
rect 57152 27072 57204 27124
rect 28632 27004 28684 27056
rect 33048 27004 33100 27056
rect 33140 27004 33192 27056
rect 44180 27004 44232 27056
rect 57244 27047 57296 27056
rect 57244 27013 57253 27047
rect 57253 27013 57287 27047
rect 57287 27013 57296 27047
rect 57244 27004 57296 27013
rect 21916 26936 21968 26988
rect 14280 26868 14332 26920
rect 22836 26868 22888 26920
rect 27528 26868 27580 26920
rect 3884 26800 3936 26852
rect 19984 26800 20036 26852
rect 32036 26936 32088 26988
rect 32312 26936 32364 26988
rect 33232 26868 33284 26920
rect 56600 26936 56652 26988
rect 37096 26868 37148 26920
rect 17408 26732 17460 26784
rect 30196 26800 30248 26852
rect 33048 26800 33100 26852
rect 41604 26800 41656 26852
rect 25136 26732 25188 26784
rect 27344 26775 27396 26784
rect 27344 26741 27353 26775
rect 27353 26741 27387 26775
rect 27387 26741 27396 26775
rect 27344 26732 27396 26741
rect 28356 26775 28408 26784
rect 28356 26741 28365 26775
rect 28365 26741 28399 26775
rect 28399 26741 28408 26775
rect 28356 26732 28408 26741
rect 29460 26775 29512 26784
rect 29460 26741 29469 26775
rect 29469 26741 29503 26775
rect 29503 26741 29512 26775
rect 29460 26732 29512 26741
rect 30564 26732 30616 26784
rect 30840 26775 30892 26784
rect 30840 26741 30849 26775
rect 30849 26741 30883 26775
rect 30883 26741 30892 26775
rect 30840 26732 30892 26741
rect 31484 26775 31536 26784
rect 31484 26741 31493 26775
rect 31493 26741 31527 26775
rect 31527 26741 31536 26775
rect 31484 26732 31536 26741
rect 31668 26732 31720 26784
rect 32588 26732 32640 26784
rect 33324 26732 33376 26784
rect 35716 26775 35768 26784
rect 35716 26741 35725 26775
rect 35725 26741 35759 26775
rect 35759 26741 35768 26775
rect 35716 26732 35768 26741
rect 35900 26732 35952 26784
rect 37556 26732 37608 26784
rect 10582 26630 10634 26682
rect 10646 26630 10698 26682
rect 10710 26630 10762 26682
rect 10774 26630 10826 26682
rect 10838 26630 10890 26682
rect 29846 26630 29898 26682
rect 29910 26630 29962 26682
rect 29974 26630 30026 26682
rect 30038 26630 30090 26682
rect 30102 26630 30154 26682
rect 49110 26630 49162 26682
rect 49174 26630 49226 26682
rect 49238 26630 49290 26682
rect 49302 26630 49354 26682
rect 49366 26630 49418 26682
rect 30472 26571 30524 26580
rect 30472 26537 30481 26571
rect 30481 26537 30515 26571
rect 30515 26537 30524 26571
rect 30472 26528 30524 26537
rect 31208 26571 31260 26580
rect 31208 26537 31217 26571
rect 31217 26537 31251 26571
rect 31251 26537 31260 26571
rect 31208 26528 31260 26537
rect 36912 26528 36964 26580
rect 46572 26528 46624 26580
rect 58072 26571 58124 26580
rect 58072 26537 58081 26571
rect 58081 26537 58115 26571
rect 58115 26537 58124 26571
rect 58072 26528 58124 26537
rect 23204 26460 23256 26512
rect 29552 26503 29604 26512
rect 23388 26392 23440 26444
rect 28816 26392 28868 26444
rect 29552 26469 29561 26503
rect 29561 26469 29595 26503
rect 29595 26469 29604 26503
rect 29552 26460 29604 26469
rect 35440 26460 35492 26512
rect 35808 26460 35860 26512
rect 45008 26460 45060 26512
rect 8576 26324 8628 26376
rect 27712 26324 27764 26376
rect 28356 26324 28408 26376
rect 29736 26367 29788 26376
rect 29736 26333 29745 26367
rect 29745 26333 29779 26367
rect 29779 26333 29788 26367
rect 29736 26324 29788 26333
rect 30748 26392 30800 26444
rect 33968 26392 34020 26444
rect 34244 26392 34296 26444
rect 37556 26392 37608 26444
rect 43536 26392 43588 26444
rect 31208 26367 31260 26376
rect 31208 26333 31217 26367
rect 31217 26333 31251 26367
rect 31251 26333 31260 26367
rect 31208 26324 31260 26333
rect 31944 26367 31996 26376
rect 31944 26333 31953 26367
rect 31953 26333 31987 26367
rect 31987 26333 31996 26367
rect 31944 26324 31996 26333
rect 28264 26299 28316 26308
rect 28264 26265 28273 26299
rect 28273 26265 28307 26299
rect 28307 26265 28316 26299
rect 28264 26256 28316 26265
rect 31852 26256 31904 26308
rect 32496 26367 32548 26376
rect 32496 26333 32505 26367
rect 32505 26333 32539 26367
rect 32539 26333 32548 26367
rect 33232 26367 33284 26376
rect 32496 26324 32548 26333
rect 33232 26333 33241 26367
rect 33241 26333 33275 26367
rect 33275 26333 33284 26367
rect 33232 26324 33284 26333
rect 35716 26324 35768 26376
rect 45560 26324 45612 26376
rect 33140 26299 33192 26308
rect 33140 26265 33149 26299
rect 33149 26265 33183 26299
rect 33183 26265 33192 26299
rect 33140 26256 33192 26265
rect 33784 26299 33836 26308
rect 33784 26265 33793 26299
rect 33793 26265 33827 26299
rect 33827 26265 33836 26299
rect 33784 26256 33836 26265
rect 34060 26256 34112 26308
rect 36176 26256 36228 26308
rect 36912 26299 36964 26308
rect 36912 26265 36921 26299
rect 36921 26265 36955 26299
rect 36955 26265 36964 26299
rect 36912 26256 36964 26265
rect 40960 26256 41012 26308
rect 1492 26231 1544 26240
rect 1492 26197 1501 26231
rect 1501 26197 1535 26231
rect 1535 26197 1544 26231
rect 1492 26188 1544 26197
rect 18972 26188 19024 26240
rect 19340 26188 19392 26240
rect 24676 26231 24728 26240
rect 24676 26197 24685 26231
rect 24685 26197 24719 26231
rect 24719 26197 24728 26231
rect 24676 26188 24728 26197
rect 25136 26231 25188 26240
rect 25136 26197 25145 26231
rect 25145 26197 25179 26231
rect 25179 26197 25188 26231
rect 25136 26188 25188 26197
rect 25412 26188 25464 26240
rect 28080 26188 28132 26240
rect 29092 26188 29144 26240
rect 31484 26188 31536 26240
rect 32680 26188 32732 26240
rect 35624 26188 35676 26240
rect 35808 26231 35860 26240
rect 35808 26197 35817 26231
rect 35817 26197 35851 26231
rect 35851 26197 35860 26231
rect 35808 26188 35860 26197
rect 38384 26188 38436 26240
rect 20214 26086 20266 26138
rect 20278 26086 20330 26138
rect 20342 26086 20394 26138
rect 20406 26086 20458 26138
rect 20470 26086 20522 26138
rect 39478 26086 39530 26138
rect 39542 26086 39594 26138
rect 39606 26086 39658 26138
rect 39670 26086 39722 26138
rect 39734 26086 39786 26138
rect 25412 25984 25464 26036
rect 30472 26027 30524 26036
rect 24676 25916 24728 25968
rect 27804 25916 27856 25968
rect 28356 25916 28408 25968
rect 26792 25848 26844 25900
rect 29368 25848 29420 25900
rect 30472 25993 30481 26027
rect 30481 25993 30515 26027
rect 30515 25993 30524 26027
rect 30472 25984 30524 25993
rect 29920 25916 29972 25968
rect 32496 25984 32548 26036
rect 33508 25984 33560 26036
rect 37280 26027 37332 26036
rect 37280 25993 37289 26027
rect 37289 25993 37323 26027
rect 37323 25993 37332 26027
rect 37280 25984 37332 25993
rect 38384 26027 38436 26036
rect 38384 25993 38393 26027
rect 38393 25993 38427 26027
rect 38427 25993 38436 26027
rect 38384 25984 38436 25993
rect 40592 25984 40644 26036
rect 46480 25984 46532 26036
rect 37740 25916 37792 25968
rect 31576 25891 31628 25900
rect 31576 25857 31585 25891
rect 31585 25857 31619 25891
rect 31619 25857 31628 25891
rect 31576 25848 31628 25857
rect 33692 25891 33744 25900
rect 29644 25780 29696 25832
rect 2228 25712 2280 25764
rect 22008 25712 22060 25764
rect 23020 25712 23072 25764
rect 27252 25755 27304 25764
rect 27252 25721 27261 25755
rect 27261 25721 27295 25755
rect 27295 25721 27304 25755
rect 27252 25712 27304 25721
rect 28540 25712 28592 25764
rect 28724 25712 28776 25764
rect 29920 25712 29972 25764
rect 30380 25712 30432 25764
rect 30932 25780 30984 25832
rect 31392 25780 31444 25832
rect 32956 25780 33008 25832
rect 33692 25857 33701 25891
rect 33701 25857 33735 25891
rect 33735 25857 33744 25891
rect 33692 25848 33744 25857
rect 34428 25848 34480 25900
rect 36636 25848 36688 25900
rect 35256 25780 35308 25832
rect 39212 25780 39264 25832
rect 58164 25848 58216 25900
rect 32588 25712 32640 25764
rect 35532 25712 35584 25764
rect 35716 25712 35768 25764
rect 57888 25755 57940 25764
rect 57888 25721 57897 25755
rect 57897 25721 57931 25755
rect 57931 25721 57940 25755
rect 57888 25712 57940 25721
rect 20720 25644 20772 25696
rect 24400 25687 24452 25696
rect 24400 25653 24409 25687
rect 24409 25653 24443 25687
rect 24443 25653 24452 25687
rect 24400 25644 24452 25653
rect 24860 25687 24912 25696
rect 24860 25653 24869 25687
rect 24869 25653 24903 25687
rect 24903 25653 24912 25687
rect 24860 25644 24912 25653
rect 25044 25644 25096 25696
rect 25412 25687 25464 25696
rect 25412 25653 25421 25687
rect 25421 25653 25455 25687
rect 25455 25653 25464 25687
rect 25412 25644 25464 25653
rect 27160 25644 27212 25696
rect 28080 25644 28132 25696
rect 28908 25687 28960 25696
rect 28908 25653 28917 25687
rect 28917 25653 28951 25687
rect 28951 25653 28960 25687
rect 28908 25644 28960 25653
rect 29460 25687 29512 25696
rect 29460 25653 29469 25687
rect 29469 25653 29503 25687
rect 29503 25653 29512 25687
rect 29460 25644 29512 25653
rect 30840 25644 30892 25696
rect 31760 25644 31812 25696
rect 32312 25644 32364 25696
rect 32404 25644 32456 25696
rect 33600 25687 33652 25696
rect 33600 25653 33609 25687
rect 33609 25653 33643 25687
rect 33643 25653 33652 25687
rect 33600 25644 33652 25653
rect 34336 25644 34388 25696
rect 34704 25687 34756 25696
rect 34704 25653 34713 25687
rect 34713 25653 34747 25687
rect 34747 25653 34756 25687
rect 34704 25644 34756 25653
rect 36452 25644 36504 25696
rect 38292 25644 38344 25696
rect 56600 25644 56652 25696
rect 10582 25542 10634 25594
rect 10646 25542 10698 25594
rect 10710 25542 10762 25594
rect 10774 25542 10826 25594
rect 10838 25542 10890 25594
rect 29846 25542 29898 25594
rect 29910 25542 29962 25594
rect 29974 25542 30026 25594
rect 30038 25542 30090 25594
rect 30102 25542 30154 25594
rect 49110 25542 49162 25594
rect 49174 25542 49226 25594
rect 49238 25542 49290 25594
rect 49302 25542 49354 25594
rect 49366 25542 49418 25594
rect 14464 25415 14516 25424
rect 14464 25381 14473 25415
rect 14473 25381 14507 25415
rect 14507 25381 14516 25415
rect 14464 25372 14516 25381
rect 21640 25372 21692 25424
rect 25780 25440 25832 25492
rect 26424 25440 26476 25492
rect 31576 25440 31628 25492
rect 33048 25440 33100 25492
rect 34612 25440 34664 25492
rect 34796 25440 34848 25492
rect 34980 25440 35032 25492
rect 37372 25440 37424 25492
rect 37556 25483 37608 25492
rect 37556 25449 37565 25483
rect 37565 25449 37599 25483
rect 37599 25449 37608 25483
rect 37556 25440 37608 25449
rect 23940 25372 23992 25424
rect 25228 25372 25280 25424
rect 26240 25372 26292 25424
rect 28724 25372 28776 25424
rect 35532 25372 35584 25424
rect 35624 25372 35676 25424
rect 38292 25372 38344 25424
rect 25780 25304 25832 25356
rect 27712 25304 27764 25356
rect 28816 25347 28868 25356
rect 28816 25313 28825 25347
rect 28825 25313 28859 25347
rect 28859 25313 28868 25347
rect 28816 25304 28868 25313
rect 29000 25304 29052 25356
rect 21456 25236 21508 25288
rect 26884 25236 26936 25288
rect 28172 25236 28224 25288
rect 28632 25279 28684 25288
rect 28632 25245 28641 25279
rect 28641 25245 28675 25279
rect 28675 25245 28684 25279
rect 28632 25236 28684 25245
rect 30288 25236 30340 25288
rect 30564 25279 30616 25288
rect 30564 25245 30573 25279
rect 30573 25245 30607 25279
rect 30607 25245 30616 25279
rect 30564 25236 30616 25245
rect 21088 25168 21140 25220
rect 23848 25168 23900 25220
rect 29184 25168 29236 25220
rect 29736 25211 29788 25220
rect 29736 25177 29745 25211
rect 29745 25177 29779 25211
rect 29779 25177 29788 25211
rect 29736 25168 29788 25177
rect 24952 25143 25004 25152
rect 24952 25109 24961 25143
rect 24961 25109 24995 25143
rect 24995 25109 25004 25143
rect 24952 25100 25004 25109
rect 26148 25100 26200 25152
rect 27160 25100 27212 25152
rect 27896 25143 27948 25152
rect 27896 25109 27905 25143
rect 27905 25109 27939 25143
rect 27939 25109 27948 25143
rect 27896 25100 27948 25109
rect 28448 25143 28500 25152
rect 28448 25109 28457 25143
rect 28457 25109 28491 25143
rect 28491 25109 28500 25143
rect 28448 25100 28500 25109
rect 31116 25100 31168 25152
rect 37188 25304 37240 25356
rect 31576 25279 31628 25288
rect 31576 25245 31585 25279
rect 31585 25245 31619 25279
rect 31619 25245 31628 25279
rect 31576 25236 31628 25245
rect 32036 25236 32088 25288
rect 33048 25279 33100 25288
rect 31484 25168 31536 25220
rect 32220 25211 32272 25220
rect 32220 25177 32229 25211
rect 32229 25177 32263 25211
rect 32263 25177 32272 25211
rect 32220 25168 32272 25177
rect 33048 25245 33057 25279
rect 33057 25245 33091 25279
rect 33091 25245 33100 25279
rect 33048 25236 33100 25245
rect 33508 25236 33560 25288
rect 35624 25236 35676 25288
rect 35716 25236 35768 25288
rect 37280 25236 37332 25288
rect 46940 25440 46992 25492
rect 58164 25483 58216 25492
rect 58164 25449 58173 25483
rect 58173 25449 58207 25483
rect 58207 25449 58216 25483
rect 58164 25440 58216 25449
rect 32036 25100 32088 25152
rect 32588 25143 32640 25152
rect 32588 25109 32597 25143
rect 32597 25109 32631 25143
rect 32631 25109 32640 25143
rect 32588 25100 32640 25109
rect 33232 25143 33284 25152
rect 33232 25109 33241 25143
rect 33241 25109 33275 25143
rect 33275 25109 33284 25143
rect 33232 25100 33284 25109
rect 36360 25168 36412 25220
rect 35624 25100 35676 25152
rect 35900 25143 35952 25152
rect 35900 25109 35909 25143
rect 35909 25109 35943 25143
rect 35943 25109 35952 25143
rect 35900 25100 35952 25109
rect 36544 25143 36596 25152
rect 36544 25109 36553 25143
rect 36553 25109 36587 25143
rect 36587 25109 36596 25143
rect 36544 25100 36596 25109
rect 38108 25143 38160 25152
rect 38108 25109 38117 25143
rect 38117 25109 38151 25143
rect 38151 25109 38160 25143
rect 38108 25100 38160 25109
rect 38752 25143 38804 25152
rect 38752 25109 38761 25143
rect 38761 25109 38795 25143
rect 38795 25109 38804 25143
rect 38752 25100 38804 25109
rect 20214 24998 20266 25050
rect 20278 24998 20330 25050
rect 20342 24998 20394 25050
rect 20406 24998 20458 25050
rect 20470 24998 20522 25050
rect 39478 24998 39530 25050
rect 39542 24998 39594 25050
rect 39606 24998 39658 25050
rect 39670 24998 39722 25050
rect 39734 24998 39786 25050
rect 25504 24896 25556 24948
rect 9128 24760 9180 24812
rect 22192 24760 22244 24812
rect 27712 24828 27764 24880
rect 31760 24896 31812 24948
rect 32220 24896 32272 24948
rect 32312 24896 32364 24948
rect 32588 24896 32640 24948
rect 19800 24692 19852 24744
rect 27528 24760 27580 24812
rect 28448 24828 28500 24880
rect 33232 24828 33284 24880
rect 38660 24828 38712 24880
rect 42892 24828 42944 24880
rect 28540 24760 28592 24812
rect 29920 24760 29972 24812
rect 30656 24803 30708 24812
rect 30656 24769 30665 24803
rect 30665 24769 30699 24803
rect 30699 24769 30708 24803
rect 30656 24760 30708 24769
rect 31576 24803 31628 24812
rect 31576 24769 31585 24803
rect 31585 24769 31619 24803
rect 31619 24769 31628 24803
rect 32128 24803 32180 24812
rect 31576 24760 31628 24769
rect 32128 24769 32137 24803
rect 32137 24769 32171 24803
rect 32171 24769 32180 24803
rect 32128 24760 32180 24769
rect 32220 24760 32272 24812
rect 32680 24760 32732 24812
rect 25504 24692 25556 24744
rect 25688 24692 25740 24744
rect 29184 24692 29236 24744
rect 29644 24692 29696 24744
rect 30564 24692 30616 24744
rect 31852 24692 31904 24744
rect 32036 24692 32088 24744
rect 33968 24803 34020 24812
rect 33968 24769 33977 24803
rect 33977 24769 34011 24803
rect 34011 24769 34020 24803
rect 33968 24760 34020 24769
rect 34612 24760 34664 24812
rect 35164 24760 35216 24812
rect 35624 24760 35676 24812
rect 35808 24760 35860 24812
rect 36176 24803 36228 24812
rect 36176 24769 36185 24803
rect 36185 24769 36219 24803
rect 36219 24769 36228 24803
rect 36176 24760 36228 24769
rect 36728 24803 36780 24812
rect 36728 24769 36737 24803
rect 36737 24769 36771 24803
rect 36771 24769 36780 24803
rect 36728 24760 36780 24769
rect 40592 24803 40644 24812
rect 40592 24769 40601 24803
rect 40601 24769 40635 24803
rect 40635 24769 40644 24803
rect 40592 24760 40644 24769
rect 8576 24624 8628 24676
rect 12348 24624 12400 24676
rect 1492 24599 1544 24608
rect 1492 24565 1501 24599
rect 1501 24565 1535 24599
rect 1535 24565 1544 24599
rect 1492 24556 1544 24565
rect 22284 24624 22336 24676
rect 24124 24624 24176 24676
rect 25320 24624 25372 24676
rect 27712 24624 27764 24676
rect 22744 24599 22796 24608
rect 22744 24565 22753 24599
rect 22753 24565 22787 24599
rect 22787 24565 22796 24599
rect 22744 24556 22796 24565
rect 23112 24556 23164 24608
rect 24400 24556 24452 24608
rect 25412 24556 25464 24608
rect 25596 24556 25648 24608
rect 26148 24556 26200 24608
rect 26332 24599 26384 24608
rect 26332 24565 26341 24599
rect 26341 24565 26375 24599
rect 26375 24565 26384 24599
rect 26332 24556 26384 24565
rect 26516 24556 26568 24608
rect 31760 24624 31812 24676
rect 35992 24692 36044 24744
rect 36452 24692 36504 24744
rect 34428 24624 34480 24676
rect 36176 24624 36228 24676
rect 44548 24624 44600 24676
rect 31300 24556 31352 24608
rect 31484 24599 31536 24608
rect 31484 24565 31493 24599
rect 31493 24565 31527 24599
rect 31527 24565 31536 24599
rect 31484 24556 31536 24565
rect 32036 24556 32088 24608
rect 32404 24556 32456 24608
rect 33140 24599 33192 24608
rect 33140 24565 33149 24599
rect 33149 24565 33183 24599
rect 33183 24565 33192 24599
rect 33140 24556 33192 24565
rect 34520 24556 34572 24608
rect 36084 24599 36136 24608
rect 36084 24565 36093 24599
rect 36093 24565 36127 24599
rect 36127 24565 36136 24599
rect 36084 24556 36136 24565
rect 37280 24599 37332 24608
rect 37280 24565 37289 24599
rect 37289 24565 37323 24599
rect 37323 24565 37332 24599
rect 37280 24556 37332 24565
rect 38568 24556 38620 24608
rect 39488 24599 39540 24608
rect 39488 24565 39497 24599
rect 39497 24565 39531 24599
rect 39531 24565 39540 24599
rect 39488 24556 39540 24565
rect 10582 24454 10634 24506
rect 10646 24454 10698 24506
rect 10710 24454 10762 24506
rect 10774 24454 10826 24506
rect 10838 24454 10890 24506
rect 29846 24454 29898 24506
rect 29910 24454 29962 24506
rect 29974 24454 30026 24506
rect 30038 24454 30090 24506
rect 30102 24454 30154 24506
rect 49110 24454 49162 24506
rect 49174 24454 49226 24506
rect 49238 24454 49290 24506
rect 49302 24454 49354 24506
rect 49366 24454 49418 24506
rect 9128 24352 9180 24404
rect 14372 24284 14424 24336
rect 23388 24352 23440 24404
rect 27160 24352 27212 24404
rect 27252 24352 27304 24404
rect 32772 24352 32824 24404
rect 33508 24352 33560 24404
rect 34704 24352 34756 24404
rect 19248 24284 19300 24336
rect 21640 24327 21692 24336
rect 21640 24293 21649 24327
rect 21649 24293 21683 24327
rect 21683 24293 21692 24327
rect 21640 24284 21692 24293
rect 23572 24284 23624 24336
rect 27436 24284 27488 24336
rect 22008 24216 22060 24268
rect 25228 24216 25280 24268
rect 30564 24284 30616 24336
rect 22284 24148 22336 24200
rect 22928 24148 22980 24200
rect 23664 24080 23716 24132
rect 22008 24012 22060 24064
rect 23572 24012 23624 24064
rect 24584 24012 24636 24064
rect 25412 24080 25464 24132
rect 25964 24148 26016 24200
rect 26700 24123 26752 24132
rect 25872 24012 25924 24064
rect 26148 24055 26200 24064
rect 26148 24021 26157 24055
rect 26157 24021 26191 24055
rect 26191 24021 26200 24055
rect 26148 24012 26200 24021
rect 26700 24089 26709 24123
rect 26709 24089 26743 24123
rect 26743 24089 26752 24123
rect 26700 24080 26752 24089
rect 27252 24148 27304 24200
rect 27344 24148 27396 24200
rect 28080 24216 28132 24268
rect 28724 24216 28776 24268
rect 29644 24259 29696 24268
rect 26976 24080 27028 24132
rect 28264 24080 28316 24132
rect 29644 24225 29653 24259
rect 29653 24225 29687 24259
rect 29687 24225 29696 24259
rect 29644 24216 29696 24225
rect 30380 24148 30432 24200
rect 32312 24191 32364 24200
rect 32312 24157 32321 24191
rect 32321 24157 32355 24191
rect 32355 24157 32364 24191
rect 32588 24216 32640 24268
rect 32956 24259 33008 24268
rect 32956 24225 32965 24259
rect 32965 24225 32999 24259
rect 32999 24225 33008 24259
rect 33876 24284 33928 24336
rect 34152 24327 34204 24336
rect 34152 24293 34161 24327
rect 34161 24293 34195 24327
rect 34195 24293 34204 24327
rect 34152 24284 34204 24293
rect 34244 24284 34296 24336
rect 36268 24352 36320 24404
rect 38384 24352 38436 24404
rect 39304 24352 39356 24404
rect 40592 24352 40644 24404
rect 36820 24284 36872 24336
rect 41696 24284 41748 24336
rect 32956 24216 33008 24225
rect 34428 24216 34480 24268
rect 32312 24148 32364 24157
rect 31484 24080 31536 24132
rect 32036 24123 32088 24132
rect 32036 24089 32045 24123
rect 32045 24089 32079 24123
rect 32079 24089 32088 24123
rect 32036 24080 32088 24089
rect 26884 24012 26936 24064
rect 27988 24012 28040 24064
rect 28540 24012 28592 24064
rect 28816 24012 28868 24064
rect 29092 24012 29144 24064
rect 30104 24055 30156 24064
rect 30104 24021 30113 24055
rect 30113 24021 30147 24055
rect 30147 24021 30156 24055
rect 30104 24012 30156 24021
rect 32128 24012 32180 24064
rect 32864 24080 32916 24132
rect 33324 24148 33376 24200
rect 33692 24148 33744 24200
rect 33876 24148 33928 24200
rect 34888 24148 34940 24200
rect 35532 24191 35584 24200
rect 35532 24157 35541 24191
rect 35541 24157 35575 24191
rect 35575 24157 35584 24191
rect 35532 24148 35584 24157
rect 36176 24191 36228 24200
rect 36176 24157 36185 24191
rect 36185 24157 36219 24191
rect 36219 24157 36228 24191
rect 36176 24148 36228 24157
rect 36268 24148 36320 24200
rect 37372 24148 37424 24200
rect 39120 24216 39172 24268
rect 38292 24148 38344 24200
rect 40776 24148 40828 24200
rect 58164 24191 58216 24200
rect 58164 24157 58173 24191
rect 58173 24157 58207 24191
rect 58207 24157 58216 24191
rect 58164 24148 58216 24157
rect 33416 24080 33468 24132
rect 33784 24123 33836 24132
rect 33784 24089 33793 24123
rect 33793 24089 33827 24123
rect 33827 24089 33836 24123
rect 33784 24080 33836 24089
rect 34060 24080 34112 24132
rect 35624 24080 35676 24132
rect 38108 24080 38160 24132
rect 38752 24080 38804 24132
rect 35532 24012 35584 24064
rect 35992 24012 36044 24064
rect 36268 24055 36320 24064
rect 36268 24021 36277 24055
rect 36277 24021 36311 24055
rect 36311 24021 36320 24055
rect 36268 24012 36320 24021
rect 36912 24012 36964 24064
rect 38384 24012 38436 24064
rect 38844 24012 38896 24064
rect 49700 24080 49752 24132
rect 42708 24012 42760 24064
rect 20214 23910 20266 23962
rect 20278 23910 20330 23962
rect 20342 23910 20394 23962
rect 20406 23910 20458 23962
rect 20470 23910 20522 23962
rect 39478 23910 39530 23962
rect 39542 23910 39594 23962
rect 39606 23910 39658 23962
rect 39670 23910 39722 23962
rect 39734 23910 39786 23962
rect 18604 23808 18656 23860
rect 25688 23851 25740 23860
rect 19984 23740 20036 23792
rect 20720 23783 20772 23792
rect 20720 23749 20729 23783
rect 20729 23749 20763 23783
rect 20763 23749 20772 23783
rect 20720 23740 20772 23749
rect 24124 23740 24176 23792
rect 25136 23740 25188 23792
rect 25688 23817 25697 23851
rect 25697 23817 25731 23851
rect 25731 23817 25740 23851
rect 25688 23808 25740 23817
rect 25872 23808 25924 23860
rect 28816 23808 28868 23860
rect 25596 23672 25648 23724
rect 25780 23672 25832 23724
rect 26332 23740 26384 23792
rect 26608 23672 26660 23724
rect 20536 23604 20588 23656
rect 22008 23604 22060 23656
rect 22836 23604 22888 23656
rect 24860 23647 24912 23656
rect 24860 23613 24869 23647
rect 24869 23613 24903 23647
rect 24903 23613 24912 23647
rect 24860 23604 24912 23613
rect 25872 23604 25924 23656
rect 28908 23740 28960 23792
rect 27252 23672 27304 23724
rect 27620 23672 27672 23724
rect 29092 23808 29144 23860
rect 35440 23808 35492 23860
rect 35900 23808 35952 23860
rect 29552 23672 29604 23724
rect 30288 23740 30340 23792
rect 30748 23740 30800 23792
rect 32772 23740 32824 23792
rect 27344 23647 27396 23656
rect 23296 23536 23348 23588
rect 27344 23613 27353 23647
rect 27353 23613 27387 23647
rect 27387 23613 27396 23647
rect 27344 23604 27396 23613
rect 27804 23604 27856 23656
rect 29184 23604 29236 23656
rect 30012 23647 30064 23656
rect 30012 23613 30021 23647
rect 30021 23613 30055 23647
rect 30055 23613 30064 23647
rect 30012 23604 30064 23613
rect 30656 23604 30708 23656
rect 33048 23672 33100 23724
rect 33876 23715 33928 23724
rect 33876 23681 33885 23715
rect 33885 23681 33919 23715
rect 33919 23681 33928 23715
rect 33876 23672 33928 23681
rect 34796 23672 34848 23724
rect 35072 23715 35124 23724
rect 35072 23681 35081 23715
rect 35081 23681 35115 23715
rect 35115 23681 35124 23715
rect 35072 23672 35124 23681
rect 35716 23715 35768 23724
rect 35716 23681 35725 23715
rect 35725 23681 35759 23715
rect 35759 23681 35768 23715
rect 35716 23672 35768 23681
rect 36452 23740 36504 23792
rect 37004 23808 37056 23860
rect 40224 23808 40276 23860
rect 40592 23808 40644 23860
rect 58164 23851 58216 23860
rect 58164 23817 58173 23851
rect 58173 23817 58207 23851
rect 58207 23817 58216 23851
rect 58164 23808 58216 23817
rect 42064 23740 42116 23792
rect 32864 23647 32916 23656
rect 21272 23511 21324 23520
rect 21272 23477 21281 23511
rect 21281 23477 21315 23511
rect 21315 23477 21324 23511
rect 21272 23468 21324 23477
rect 21732 23468 21784 23520
rect 27160 23536 27212 23588
rect 28724 23579 28776 23588
rect 28724 23545 28733 23579
rect 28733 23545 28767 23579
rect 28767 23545 28776 23579
rect 28724 23536 28776 23545
rect 32864 23613 32873 23647
rect 32873 23613 32907 23647
rect 32907 23613 32916 23647
rect 32864 23604 32916 23613
rect 33968 23647 34020 23656
rect 33968 23613 33977 23647
rect 33977 23613 34011 23647
rect 34011 23613 34020 23647
rect 33968 23604 34020 23613
rect 26516 23468 26568 23520
rect 27344 23468 27396 23520
rect 27620 23468 27672 23520
rect 28264 23468 28316 23520
rect 30196 23468 30248 23520
rect 31944 23536 31996 23588
rect 35900 23604 35952 23656
rect 36176 23604 36228 23656
rect 36912 23604 36964 23656
rect 37188 23672 37240 23724
rect 37372 23672 37424 23724
rect 38108 23715 38160 23724
rect 38108 23681 38117 23715
rect 38117 23681 38151 23715
rect 38151 23681 38160 23715
rect 38108 23672 38160 23681
rect 40500 23672 40552 23724
rect 40776 23672 40828 23724
rect 49700 23672 49752 23724
rect 40684 23604 40736 23656
rect 34244 23579 34296 23588
rect 34244 23545 34253 23579
rect 34253 23545 34287 23579
rect 34287 23545 34296 23579
rect 34244 23536 34296 23545
rect 34428 23536 34480 23588
rect 36728 23536 36780 23588
rect 38936 23536 38988 23588
rect 41236 23536 41288 23588
rect 36452 23511 36504 23520
rect 36452 23477 36461 23511
rect 36461 23477 36495 23511
rect 36495 23477 36504 23511
rect 36452 23468 36504 23477
rect 36544 23511 36596 23520
rect 36544 23477 36553 23511
rect 36553 23477 36587 23511
rect 36587 23477 36596 23511
rect 38016 23511 38068 23520
rect 36544 23468 36596 23477
rect 38016 23477 38025 23511
rect 38025 23477 38059 23511
rect 38059 23477 38068 23511
rect 38016 23468 38068 23477
rect 39028 23468 39080 23520
rect 39396 23468 39448 23520
rect 41604 23468 41656 23520
rect 41788 23468 41840 23520
rect 10582 23366 10634 23418
rect 10646 23366 10698 23418
rect 10710 23366 10762 23418
rect 10774 23366 10826 23418
rect 10838 23366 10890 23418
rect 29846 23366 29898 23418
rect 29910 23366 29962 23418
rect 29974 23366 30026 23418
rect 30038 23366 30090 23418
rect 30102 23366 30154 23418
rect 49110 23366 49162 23418
rect 49174 23366 49226 23418
rect 49238 23366 49290 23418
rect 49302 23366 49354 23418
rect 49366 23366 49418 23418
rect 2228 23307 2280 23316
rect 2228 23273 2237 23307
rect 2237 23273 2271 23307
rect 2271 23273 2280 23307
rect 2228 23264 2280 23273
rect 19340 23264 19392 23316
rect 21640 23264 21692 23316
rect 22008 23264 22060 23316
rect 19248 23196 19300 23248
rect 23296 23196 23348 23248
rect 22560 23128 22612 23180
rect 24860 23196 24912 23248
rect 26056 23196 26108 23248
rect 27988 23264 28040 23316
rect 28908 23264 28960 23316
rect 29552 23264 29604 23316
rect 24768 23128 24820 23180
rect 25780 23128 25832 23180
rect 26332 23171 26384 23180
rect 26332 23137 26341 23171
rect 26341 23137 26375 23171
rect 26375 23137 26384 23171
rect 26332 23128 26384 23137
rect 2228 23060 2280 23112
rect 24124 23060 24176 23112
rect 24492 23103 24544 23112
rect 24492 23069 24501 23103
rect 24501 23069 24535 23103
rect 24535 23069 24544 23103
rect 24492 23060 24544 23069
rect 24676 23103 24728 23112
rect 24676 23069 24685 23103
rect 24685 23069 24719 23103
rect 24719 23069 24728 23103
rect 25228 23103 25280 23112
rect 24676 23060 24728 23069
rect 25228 23069 25237 23103
rect 25237 23069 25271 23103
rect 25271 23069 25280 23103
rect 25228 23060 25280 23069
rect 26700 23060 26752 23112
rect 29644 23196 29696 23248
rect 30196 23264 30248 23316
rect 31944 23264 31996 23316
rect 32128 23264 32180 23316
rect 34336 23264 34388 23316
rect 31852 23196 31904 23248
rect 34152 23196 34204 23248
rect 27620 23128 27672 23180
rect 28908 23171 28960 23180
rect 28908 23137 28917 23171
rect 28917 23137 28951 23171
rect 28951 23137 28960 23171
rect 28908 23128 28960 23137
rect 29184 23128 29236 23180
rect 31392 23128 31444 23180
rect 40592 23264 40644 23316
rect 42984 23264 43036 23316
rect 41052 23196 41104 23248
rect 35072 23128 35124 23180
rect 35256 23128 35308 23180
rect 35992 23171 36044 23180
rect 35992 23137 36001 23171
rect 36001 23137 36035 23171
rect 36035 23137 36044 23171
rect 35992 23128 36044 23137
rect 36636 23171 36688 23180
rect 36636 23137 36645 23171
rect 36645 23137 36679 23171
rect 36679 23137 36688 23171
rect 36636 23128 36688 23137
rect 38752 23128 38804 23180
rect 23480 22992 23532 23044
rect 25412 22992 25464 23044
rect 1492 22967 1544 22976
rect 1492 22933 1501 22967
rect 1501 22933 1535 22967
rect 1535 22933 1544 22967
rect 1492 22924 1544 22933
rect 20812 22924 20864 22976
rect 22376 22924 22428 22976
rect 22744 22967 22796 22976
rect 22744 22933 22753 22967
rect 22753 22933 22787 22967
rect 22787 22933 22796 22967
rect 22744 22924 22796 22933
rect 23296 22967 23348 22976
rect 23296 22933 23305 22967
rect 23305 22933 23339 22967
rect 23339 22933 23348 22967
rect 23296 22924 23348 22933
rect 23940 22924 23992 22976
rect 24032 22924 24084 22976
rect 26884 22992 26936 23044
rect 27988 23103 28040 23112
rect 27988 23069 27997 23103
rect 27997 23069 28031 23103
rect 28031 23069 28040 23103
rect 27988 23060 28040 23069
rect 28172 23103 28224 23112
rect 28172 23069 28181 23103
rect 28181 23069 28215 23103
rect 28215 23069 28224 23103
rect 28172 23060 28224 23069
rect 29276 23060 29328 23112
rect 29552 23060 29604 23112
rect 27620 22992 27672 23044
rect 30104 22992 30156 23044
rect 30748 22992 30800 23044
rect 28080 22924 28132 22976
rect 28264 22924 28316 22976
rect 32128 22924 32180 22976
rect 34060 23060 34112 23112
rect 34888 23103 34940 23112
rect 34888 23069 34897 23103
rect 34897 23069 34931 23103
rect 34931 23069 34940 23103
rect 34888 23060 34940 23069
rect 37372 23103 37424 23112
rect 37372 23069 37381 23103
rect 37381 23069 37415 23103
rect 37415 23069 37424 23103
rect 37372 23060 37424 23069
rect 37464 23060 37516 23112
rect 37832 23060 37884 23112
rect 33600 22992 33652 23044
rect 33692 23035 33744 23044
rect 33692 23001 33701 23035
rect 33701 23001 33735 23035
rect 33735 23001 33744 23035
rect 33692 22992 33744 23001
rect 34244 22992 34296 23044
rect 37096 22992 37148 23044
rect 38384 22992 38436 23044
rect 34520 22924 34572 22976
rect 34704 22924 34756 22976
rect 34888 22924 34940 22976
rect 36820 22924 36872 22976
rect 37188 22924 37240 22976
rect 38844 22924 38896 22976
rect 40408 22967 40460 22976
rect 40408 22933 40417 22967
rect 40417 22933 40451 22967
rect 40451 22933 40460 22967
rect 40408 22924 40460 22933
rect 41328 22924 41380 22976
rect 42340 22924 42392 22976
rect 42616 22967 42668 22976
rect 42616 22933 42625 22967
rect 42625 22933 42659 22967
rect 42659 22933 42668 22967
rect 42616 22924 42668 22933
rect 20214 22822 20266 22874
rect 20278 22822 20330 22874
rect 20342 22822 20394 22874
rect 20406 22822 20458 22874
rect 20470 22822 20522 22874
rect 39478 22822 39530 22874
rect 39542 22822 39594 22874
rect 39606 22822 39658 22874
rect 39670 22822 39722 22874
rect 39734 22822 39786 22874
rect 17960 22720 18012 22772
rect 19248 22720 19300 22772
rect 20076 22763 20128 22772
rect 20076 22729 20085 22763
rect 20085 22729 20119 22763
rect 20119 22729 20128 22763
rect 20076 22720 20128 22729
rect 21088 22720 21140 22772
rect 21456 22720 21508 22772
rect 23296 22720 23348 22772
rect 25688 22720 25740 22772
rect 27252 22720 27304 22772
rect 27620 22720 27672 22772
rect 27988 22720 28040 22772
rect 19892 22652 19944 22704
rect 24216 22652 24268 22704
rect 25596 22695 25648 22704
rect 25596 22661 25605 22695
rect 25605 22661 25639 22695
rect 25639 22661 25648 22695
rect 25596 22652 25648 22661
rect 25780 22652 25832 22704
rect 26884 22652 26936 22704
rect 27528 22652 27580 22704
rect 23848 22584 23900 22636
rect 24124 22627 24176 22636
rect 19248 22516 19300 22568
rect 22836 22516 22888 22568
rect 23572 22516 23624 22568
rect 23756 22516 23808 22568
rect 24124 22593 24133 22627
rect 24133 22593 24167 22627
rect 24167 22593 24176 22627
rect 24124 22584 24176 22593
rect 24952 22627 25004 22636
rect 24952 22593 24961 22627
rect 24961 22593 24995 22627
rect 24995 22593 25004 22627
rect 24952 22584 25004 22593
rect 26424 22584 26476 22636
rect 27160 22627 27212 22636
rect 27160 22593 27169 22627
rect 27169 22593 27203 22627
rect 27203 22593 27212 22627
rect 27160 22584 27212 22593
rect 27252 22627 27304 22636
rect 27252 22593 27261 22627
rect 27261 22593 27295 22627
rect 27295 22593 27304 22627
rect 27252 22584 27304 22593
rect 24400 22516 24452 22568
rect 25044 22559 25096 22568
rect 21456 22448 21508 22500
rect 25044 22525 25053 22559
rect 25053 22525 25087 22559
rect 25087 22525 25096 22559
rect 25044 22516 25096 22525
rect 25136 22516 25188 22568
rect 25596 22516 25648 22568
rect 28264 22584 28316 22636
rect 27804 22516 27856 22568
rect 19984 22380 20036 22432
rect 22008 22380 22060 22432
rect 22836 22380 22888 22432
rect 23388 22423 23440 22432
rect 23388 22389 23397 22423
rect 23397 22389 23431 22423
rect 23431 22389 23440 22423
rect 23388 22380 23440 22389
rect 25412 22448 25464 22500
rect 25688 22448 25740 22500
rect 25780 22448 25832 22500
rect 30840 22720 30892 22772
rect 32772 22720 32824 22772
rect 32864 22720 32916 22772
rect 37096 22720 37148 22772
rect 37280 22763 37332 22772
rect 37280 22729 37289 22763
rect 37289 22729 37323 22763
rect 37323 22729 37332 22763
rect 37280 22720 37332 22729
rect 39396 22720 39448 22772
rect 41420 22763 41472 22772
rect 41420 22729 41429 22763
rect 41429 22729 41463 22763
rect 41463 22729 41472 22763
rect 41420 22720 41472 22729
rect 42984 22763 43036 22772
rect 42984 22729 42993 22763
rect 42993 22729 43027 22763
rect 43027 22729 43036 22763
rect 42984 22720 43036 22729
rect 29184 22652 29236 22704
rect 32956 22652 33008 22704
rect 33692 22652 33744 22704
rect 26424 22380 26476 22432
rect 26516 22380 26568 22432
rect 27528 22380 27580 22432
rect 27988 22380 28040 22432
rect 28632 22380 28684 22432
rect 29184 22380 29236 22432
rect 31852 22516 31904 22568
rect 32864 22516 32916 22568
rect 33140 22516 33192 22568
rect 33876 22559 33928 22568
rect 33876 22525 33885 22559
rect 33885 22525 33919 22559
rect 33919 22525 33928 22559
rect 33876 22516 33928 22525
rect 34704 22559 34756 22568
rect 34704 22525 34713 22559
rect 34713 22525 34747 22559
rect 34747 22525 34756 22559
rect 34704 22516 34756 22525
rect 31392 22448 31444 22500
rect 32404 22448 32456 22500
rect 35900 22584 35952 22636
rect 36176 22584 36228 22636
rect 36728 22627 36780 22636
rect 36728 22593 36737 22627
rect 36737 22593 36771 22627
rect 36771 22593 36780 22627
rect 36728 22584 36780 22593
rect 38200 22584 38252 22636
rect 38568 22627 38620 22636
rect 38568 22593 38577 22627
rect 38577 22593 38611 22627
rect 38611 22593 38620 22627
rect 38568 22584 38620 22593
rect 36820 22516 36872 22568
rect 30472 22380 30524 22432
rect 31208 22380 31260 22432
rect 31576 22380 31628 22432
rect 37004 22448 37056 22500
rect 38108 22516 38160 22568
rect 43904 22652 43956 22704
rect 41236 22584 41288 22636
rect 38200 22448 38252 22500
rect 39580 22448 39632 22500
rect 35992 22380 36044 22432
rect 36728 22423 36780 22432
rect 36728 22389 36737 22423
rect 36737 22389 36771 22423
rect 36771 22389 36780 22423
rect 36728 22380 36780 22389
rect 37556 22380 37608 22432
rect 37648 22380 37700 22432
rect 37924 22380 37976 22432
rect 38752 22380 38804 22432
rect 45468 22516 45520 22568
rect 42800 22448 42852 22500
rect 43536 22491 43588 22500
rect 43536 22457 43545 22491
rect 43545 22457 43579 22491
rect 43579 22457 43588 22491
rect 43536 22448 43588 22457
rect 39856 22380 39908 22432
rect 41328 22380 41380 22432
rect 45376 22380 45428 22432
rect 10582 22278 10634 22330
rect 10646 22278 10698 22330
rect 10710 22278 10762 22330
rect 10774 22278 10826 22330
rect 10838 22278 10890 22330
rect 29846 22278 29898 22330
rect 29910 22278 29962 22330
rect 29974 22278 30026 22330
rect 30038 22278 30090 22330
rect 30102 22278 30154 22330
rect 49110 22278 49162 22330
rect 49174 22278 49226 22330
rect 49238 22278 49290 22330
rect 49302 22278 49354 22330
rect 49366 22278 49418 22330
rect 20720 22176 20772 22228
rect 22744 22176 22796 22228
rect 23572 22176 23624 22228
rect 24124 22176 24176 22228
rect 26240 22176 26292 22228
rect 26516 22176 26568 22228
rect 26976 22176 27028 22228
rect 27896 22176 27948 22228
rect 28264 22176 28316 22228
rect 29736 22176 29788 22228
rect 31576 22176 31628 22228
rect 19524 22108 19576 22160
rect 25504 22108 25556 22160
rect 25780 22108 25832 22160
rect 19340 22040 19392 22092
rect 23204 22040 23256 22092
rect 24216 22040 24268 22092
rect 24492 22040 24544 22092
rect 25320 22083 25372 22092
rect 25320 22049 25329 22083
rect 25329 22049 25363 22083
rect 25363 22049 25372 22083
rect 25320 22040 25372 22049
rect 22100 21972 22152 22024
rect 22744 21972 22796 22024
rect 22928 22015 22980 22024
rect 22928 21981 22937 22015
rect 22937 21981 22971 22015
rect 22971 21981 22980 22015
rect 22928 21972 22980 21981
rect 23112 22015 23164 22024
rect 23112 21981 23121 22015
rect 23121 21981 23155 22015
rect 23155 21981 23164 22015
rect 23112 21972 23164 21981
rect 23940 21972 23992 22024
rect 25228 22015 25280 22024
rect 25228 21981 25237 22015
rect 25237 21981 25271 22015
rect 25271 21981 25280 22015
rect 26608 22108 26660 22160
rect 27160 22108 27212 22160
rect 31208 22108 31260 22160
rect 33876 22176 33928 22228
rect 35072 22176 35124 22228
rect 35900 22176 35952 22228
rect 36176 22176 36228 22228
rect 36636 22176 36688 22228
rect 34520 22108 34572 22160
rect 42616 22176 42668 22228
rect 42984 22176 43036 22228
rect 38568 22151 38620 22160
rect 38568 22117 38577 22151
rect 38577 22117 38611 22151
rect 38611 22117 38620 22151
rect 38568 22108 38620 22117
rect 26240 22083 26292 22092
rect 26240 22049 26249 22083
rect 26249 22049 26283 22083
rect 26283 22049 26292 22083
rect 26240 22040 26292 22049
rect 27528 22040 27580 22092
rect 29184 22040 29236 22092
rect 29552 22040 29604 22092
rect 30380 22040 30432 22092
rect 36084 22040 36136 22092
rect 36452 22040 36504 22092
rect 25228 21972 25280 21981
rect 26332 21972 26384 22024
rect 26608 21972 26660 22024
rect 28908 21972 28960 22024
rect 32312 21972 32364 22024
rect 33692 22015 33744 22024
rect 33692 21981 33701 22015
rect 33701 21981 33735 22015
rect 33735 21981 33744 22015
rect 33692 21972 33744 21981
rect 34336 21972 34388 22024
rect 37372 21972 37424 22024
rect 37556 21972 37608 22024
rect 38108 22040 38160 22092
rect 38476 22083 38528 22092
rect 38476 22049 38485 22083
rect 38485 22049 38519 22083
rect 38519 22049 38528 22083
rect 38476 22040 38528 22049
rect 39304 22108 39356 22160
rect 39856 22108 39908 22160
rect 40040 22108 40092 22160
rect 40224 22108 40276 22160
rect 37924 21972 37976 22024
rect 21180 21904 21232 21956
rect 15016 21836 15068 21888
rect 18052 21879 18104 21888
rect 18052 21845 18061 21879
rect 18061 21845 18095 21879
rect 18095 21845 18104 21879
rect 18052 21836 18104 21845
rect 19432 21879 19484 21888
rect 19432 21845 19441 21879
rect 19441 21845 19475 21879
rect 19475 21845 19484 21879
rect 19432 21836 19484 21845
rect 20076 21836 20128 21888
rect 20904 21836 20956 21888
rect 21272 21836 21324 21888
rect 23296 21904 23348 21956
rect 22192 21836 22244 21888
rect 22376 21836 22428 21888
rect 25412 21836 25464 21888
rect 26056 21836 26108 21888
rect 26332 21879 26384 21888
rect 26332 21845 26341 21879
rect 26341 21845 26375 21879
rect 26375 21845 26384 21879
rect 26332 21836 26384 21845
rect 26516 21836 26568 21888
rect 26884 21836 26936 21888
rect 28172 21904 28224 21956
rect 33508 21904 33560 21956
rect 33968 21904 34020 21956
rect 36084 21904 36136 21956
rect 37832 21904 37884 21956
rect 39120 22015 39172 22024
rect 39120 21981 39129 22015
rect 39129 21981 39163 22015
rect 39163 21981 39172 22015
rect 39120 21972 39172 21981
rect 41696 22040 41748 22092
rect 43904 22108 43956 22160
rect 48688 22108 48740 22160
rect 44088 22040 44140 22092
rect 40132 21972 40184 22024
rect 58164 22015 58216 22024
rect 58164 21981 58173 22015
rect 58173 21981 58207 22015
rect 58207 21981 58216 22015
rect 58164 21972 58216 21981
rect 41144 21904 41196 21956
rect 47860 21904 47912 21956
rect 29552 21836 29604 21888
rect 31944 21879 31996 21888
rect 31944 21845 31953 21879
rect 31953 21845 31987 21879
rect 31987 21845 31996 21879
rect 31944 21836 31996 21845
rect 32680 21836 32732 21888
rect 33140 21836 33192 21888
rect 35164 21836 35216 21888
rect 37004 21836 37056 21888
rect 37188 21836 37240 21888
rect 37280 21836 37332 21888
rect 39304 21836 39356 21888
rect 40408 21836 40460 21888
rect 41328 21836 41380 21888
rect 42064 21836 42116 21888
rect 42432 21836 42484 21888
rect 42708 21836 42760 21888
rect 43260 21836 43312 21888
rect 20214 21734 20266 21786
rect 20278 21734 20330 21786
rect 20342 21734 20394 21786
rect 20406 21734 20458 21786
rect 20470 21734 20522 21786
rect 39478 21734 39530 21786
rect 39542 21734 39594 21786
rect 39606 21734 39658 21786
rect 39670 21734 39722 21786
rect 39734 21734 39786 21786
rect 16120 21632 16172 21684
rect 19340 21632 19392 21684
rect 20720 21675 20772 21684
rect 20720 21641 20729 21675
rect 20729 21641 20763 21675
rect 20763 21641 20772 21675
rect 20720 21632 20772 21641
rect 21180 21632 21232 21684
rect 26332 21632 26384 21684
rect 27620 21632 27672 21684
rect 27804 21632 27856 21684
rect 27896 21632 27948 21684
rect 29552 21632 29604 21684
rect 30196 21632 30248 21684
rect 30472 21632 30524 21684
rect 30840 21632 30892 21684
rect 15752 21564 15804 21616
rect 19616 21564 19668 21616
rect 19984 21564 20036 21616
rect 20628 21564 20680 21616
rect 22836 21607 22888 21616
rect 22836 21573 22845 21607
rect 22845 21573 22879 21607
rect 22879 21573 22888 21607
rect 22836 21564 22888 21573
rect 22928 21564 22980 21616
rect 23204 21564 23256 21616
rect 24124 21564 24176 21616
rect 12256 21496 12308 21548
rect 17868 21496 17920 21548
rect 18328 21428 18380 21480
rect 21180 21428 21232 21480
rect 22284 21496 22336 21548
rect 23388 21496 23440 21548
rect 24584 21564 24636 21616
rect 24952 21564 25004 21616
rect 24768 21496 24820 21548
rect 25412 21496 25464 21548
rect 25688 21496 25740 21548
rect 26332 21496 26384 21548
rect 26516 21564 26568 21616
rect 27988 21564 28040 21616
rect 30380 21564 30432 21616
rect 31576 21564 31628 21616
rect 27620 21539 27672 21548
rect 27620 21505 27629 21539
rect 27629 21505 27663 21539
rect 27663 21505 27672 21539
rect 27620 21496 27672 21505
rect 32956 21564 33008 21616
rect 22744 21428 22796 21480
rect 26056 21428 26108 21480
rect 27528 21428 27580 21480
rect 28448 21428 28500 21480
rect 19984 21360 20036 21412
rect 1492 21335 1544 21344
rect 1492 21301 1501 21335
rect 1501 21301 1535 21335
rect 1535 21301 1544 21335
rect 1492 21292 1544 21301
rect 18696 21335 18748 21344
rect 18696 21301 18705 21335
rect 18705 21301 18739 21335
rect 18739 21301 18748 21335
rect 18696 21292 18748 21301
rect 20168 21335 20220 21344
rect 20168 21301 20177 21335
rect 20177 21301 20211 21335
rect 20211 21301 20220 21335
rect 20168 21292 20220 21301
rect 20720 21292 20772 21344
rect 20904 21292 20956 21344
rect 21548 21292 21600 21344
rect 21824 21292 21876 21344
rect 22284 21335 22336 21344
rect 22284 21301 22293 21335
rect 22293 21301 22327 21335
rect 22327 21301 22336 21335
rect 22284 21292 22336 21301
rect 22928 21292 22980 21344
rect 23940 21292 23992 21344
rect 24124 21292 24176 21344
rect 24216 21292 24268 21344
rect 24492 21292 24544 21344
rect 24768 21292 24820 21344
rect 24952 21292 25004 21344
rect 25872 21360 25924 21412
rect 26240 21292 26292 21344
rect 26792 21292 26844 21344
rect 27068 21335 27120 21344
rect 27068 21301 27077 21335
rect 27077 21301 27111 21335
rect 27111 21301 27120 21335
rect 27068 21292 27120 21301
rect 29552 21428 29604 21480
rect 29184 21360 29236 21412
rect 32496 21428 32548 21480
rect 33048 21428 33100 21480
rect 34244 21632 34296 21684
rect 37556 21632 37608 21684
rect 37648 21632 37700 21684
rect 39856 21632 39908 21684
rect 40040 21632 40092 21684
rect 44088 21675 44140 21684
rect 44088 21641 44097 21675
rect 44097 21641 44131 21675
rect 44131 21641 44140 21675
rect 44088 21632 44140 21641
rect 58164 21675 58216 21684
rect 58164 21641 58173 21675
rect 58173 21641 58207 21675
rect 58207 21641 58216 21675
rect 58164 21632 58216 21641
rect 34612 21607 34664 21616
rect 34612 21573 34621 21607
rect 34621 21573 34655 21607
rect 34655 21573 34664 21607
rect 34612 21564 34664 21573
rect 35624 21564 35676 21616
rect 34060 21496 34112 21548
rect 36636 21496 36688 21548
rect 36912 21496 36964 21548
rect 38844 21496 38896 21548
rect 40224 21564 40276 21616
rect 40316 21496 40368 21548
rect 40592 21539 40644 21548
rect 40592 21505 40601 21539
rect 40601 21505 40635 21539
rect 40635 21505 40644 21539
rect 40592 21496 40644 21505
rect 35072 21428 35124 21480
rect 31852 21360 31904 21412
rect 35624 21360 35676 21412
rect 36084 21403 36136 21412
rect 36084 21369 36093 21403
rect 36093 21369 36127 21403
rect 36127 21369 36136 21403
rect 37464 21428 37516 21480
rect 38844 21403 38896 21412
rect 36084 21360 36136 21369
rect 33600 21292 33652 21344
rect 35808 21292 35860 21344
rect 36636 21335 36688 21344
rect 36636 21301 36645 21335
rect 36645 21301 36679 21335
rect 36679 21301 36688 21335
rect 36636 21292 36688 21301
rect 38844 21369 38853 21403
rect 38853 21369 38887 21403
rect 38887 21369 38896 21403
rect 38844 21360 38896 21369
rect 39120 21428 39172 21480
rect 40040 21428 40092 21480
rect 40500 21428 40552 21480
rect 41052 21428 41104 21480
rect 41512 21428 41564 21480
rect 39856 21360 39908 21412
rect 39948 21360 40000 21412
rect 57888 21360 57940 21412
rect 39488 21292 39540 21344
rect 40500 21335 40552 21344
rect 40500 21301 40509 21335
rect 40509 21301 40543 21335
rect 40543 21301 40552 21335
rect 40500 21292 40552 21301
rect 42524 21335 42576 21344
rect 42524 21301 42533 21335
rect 42533 21301 42567 21335
rect 42567 21301 42576 21335
rect 42524 21292 42576 21301
rect 44548 21292 44600 21344
rect 44824 21292 44876 21344
rect 46204 21292 46256 21344
rect 10582 21190 10634 21242
rect 10646 21190 10698 21242
rect 10710 21190 10762 21242
rect 10774 21190 10826 21242
rect 10838 21190 10890 21242
rect 29846 21190 29898 21242
rect 29910 21190 29962 21242
rect 29974 21190 30026 21242
rect 30038 21190 30090 21242
rect 30102 21190 30154 21242
rect 49110 21190 49162 21242
rect 49174 21190 49226 21242
rect 49238 21190 49290 21242
rect 49302 21190 49354 21242
rect 49366 21190 49418 21242
rect 15752 21131 15804 21140
rect 15752 21097 15761 21131
rect 15761 21097 15795 21131
rect 15795 21097 15804 21131
rect 15752 21088 15804 21097
rect 16764 21088 16816 21140
rect 17960 21088 18012 21140
rect 21824 21131 21876 21140
rect 21824 21097 21833 21131
rect 21833 21097 21867 21131
rect 21867 21097 21876 21131
rect 21824 21088 21876 21097
rect 18052 21020 18104 21072
rect 19340 21020 19392 21072
rect 20076 21020 20128 21072
rect 22100 21020 22152 21072
rect 24492 21088 24544 21140
rect 24952 21088 25004 21140
rect 25136 21088 25188 21140
rect 27252 21131 27304 21140
rect 27252 21097 27261 21131
rect 27261 21097 27295 21131
rect 27295 21097 27304 21131
rect 27252 21088 27304 21097
rect 16856 20952 16908 21004
rect 17868 20952 17920 21004
rect 22560 20995 22612 21004
rect 17684 20884 17736 20936
rect 20168 20884 20220 20936
rect 20996 20884 21048 20936
rect 21456 20884 21508 20936
rect 21640 20927 21692 20936
rect 21640 20893 21649 20927
rect 21649 20893 21683 20927
rect 21683 20893 21692 20927
rect 21640 20884 21692 20893
rect 22560 20961 22569 20995
rect 22569 20961 22603 20995
rect 22603 20961 22612 20995
rect 22560 20952 22612 20961
rect 23020 20952 23072 21004
rect 23756 20952 23808 21004
rect 15108 20816 15160 20868
rect 23572 20884 23624 20936
rect 25320 21020 25372 21072
rect 26976 21020 27028 21072
rect 30564 21088 30616 21140
rect 31576 21088 31628 21140
rect 29552 21020 29604 21072
rect 24676 20952 24728 21004
rect 25412 20952 25464 21004
rect 24492 20884 24544 20936
rect 22928 20816 22980 20868
rect 24860 20927 24912 20936
rect 24860 20893 24869 20927
rect 24869 20893 24903 20927
rect 24903 20893 24912 20927
rect 24860 20884 24912 20893
rect 25780 20884 25832 20936
rect 26608 20952 26660 21004
rect 28632 20952 28684 21004
rect 29276 20952 29328 21004
rect 26332 20884 26384 20936
rect 26884 20884 26936 20936
rect 29184 20884 29236 20936
rect 30012 20952 30064 21004
rect 30472 20952 30524 21004
rect 29828 20927 29880 20936
rect 29828 20893 29837 20927
rect 29837 20893 29871 20927
rect 29871 20893 29880 20927
rect 32128 20952 32180 21004
rect 29828 20884 29880 20893
rect 13728 20748 13780 20800
rect 16764 20791 16816 20800
rect 16764 20757 16773 20791
rect 16773 20757 16807 20791
rect 16807 20757 16816 20791
rect 16764 20748 16816 20757
rect 17408 20791 17460 20800
rect 17408 20757 17417 20791
rect 17417 20757 17451 20791
rect 17451 20757 17460 20791
rect 17408 20748 17460 20757
rect 17776 20748 17828 20800
rect 19708 20748 19760 20800
rect 21640 20748 21692 20800
rect 22836 20791 22888 20800
rect 22836 20757 22845 20791
rect 22845 20757 22879 20791
rect 22879 20757 22888 20791
rect 22836 20748 22888 20757
rect 26792 20859 26844 20868
rect 26792 20825 26801 20859
rect 26801 20825 26835 20859
rect 26835 20825 26844 20859
rect 26792 20816 26844 20825
rect 28448 20748 28500 20800
rect 29276 20816 29328 20868
rect 29644 20816 29696 20868
rect 32404 21088 32456 21140
rect 39120 21088 39172 21140
rect 39948 21088 40000 21140
rect 40592 21088 40644 21140
rect 40776 21088 40828 21140
rect 42064 21131 42116 21140
rect 42064 21097 42073 21131
rect 42073 21097 42107 21131
rect 42107 21097 42116 21131
rect 42064 21088 42116 21097
rect 42156 21088 42208 21140
rect 34336 21020 34388 21072
rect 34060 20995 34112 21004
rect 34060 20961 34069 20995
rect 34069 20961 34103 20995
rect 34103 20961 34112 20995
rect 34060 20952 34112 20961
rect 34428 20952 34480 21004
rect 29920 20748 29972 20800
rect 30380 20748 30432 20800
rect 32956 20884 33008 20936
rect 32404 20816 32456 20868
rect 34520 20884 34572 20936
rect 38016 21020 38068 21072
rect 40316 21020 40368 21072
rect 37004 20952 37056 21004
rect 35716 20816 35768 20868
rect 38384 20884 38436 20936
rect 38752 20884 38804 20936
rect 39488 20884 39540 20936
rect 36912 20859 36964 20868
rect 36912 20825 36921 20859
rect 36921 20825 36955 20859
rect 36955 20825 36964 20859
rect 36912 20816 36964 20825
rect 39948 20859 40000 20868
rect 39948 20825 39957 20859
rect 39957 20825 39991 20859
rect 39991 20825 40000 20859
rect 39948 20816 40000 20825
rect 43720 20952 43772 21004
rect 41328 20927 41380 20936
rect 41328 20893 41337 20927
rect 41337 20893 41371 20927
rect 41371 20893 41380 20927
rect 41328 20884 41380 20893
rect 41512 20927 41564 20936
rect 41512 20893 41521 20927
rect 41521 20893 41555 20927
rect 41555 20893 41564 20927
rect 41512 20884 41564 20893
rect 44088 21088 44140 21140
rect 46480 21088 46532 21140
rect 47860 20884 47912 20936
rect 42984 20816 43036 20868
rect 43260 20816 43312 20868
rect 34152 20748 34204 20800
rect 36544 20748 36596 20800
rect 38752 20748 38804 20800
rect 39120 20748 39172 20800
rect 41696 20748 41748 20800
rect 43076 20748 43128 20800
rect 44824 20748 44876 20800
rect 46020 20748 46072 20800
rect 46204 20791 46256 20800
rect 46204 20757 46213 20791
rect 46213 20757 46247 20791
rect 46247 20757 46256 20791
rect 46204 20748 46256 20757
rect 20214 20646 20266 20698
rect 20278 20646 20330 20698
rect 20342 20646 20394 20698
rect 20406 20646 20458 20698
rect 20470 20646 20522 20698
rect 39478 20646 39530 20698
rect 39542 20646 39594 20698
rect 39606 20646 39658 20698
rect 39670 20646 39722 20698
rect 39734 20646 39786 20698
rect 12716 20544 12768 20596
rect 16120 20587 16172 20596
rect 16120 20553 16129 20587
rect 16129 20553 16163 20587
rect 16163 20553 16172 20587
rect 16120 20544 16172 20553
rect 17040 20587 17092 20596
rect 17040 20553 17049 20587
rect 17049 20553 17083 20587
rect 17083 20553 17092 20587
rect 17040 20544 17092 20553
rect 18788 20544 18840 20596
rect 20628 20544 20680 20596
rect 21364 20544 21416 20596
rect 21456 20544 21508 20596
rect 25228 20544 25280 20596
rect 25504 20544 25556 20596
rect 19800 20519 19852 20528
rect 19800 20485 19809 20519
rect 19809 20485 19843 20519
rect 19843 20485 19852 20519
rect 19800 20476 19852 20485
rect 17592 20408 17644 20460
rect 20076 20408 20128 20460
rect 20812 20476 20864 20528
rect 22284 20476 22336 20528
rect 20812 20340 20864 20392
rect 21088 20340 21140 20392
rect 21640 20408 21692 20460
rect 23756 20476 23808 20528
rect 24032 20519 24084 20528
rect 24032 20485 24041 20519
rect 24041 20485 24075 20519
rect 24075 20485 24084 20519
rect 24032 20476 24084 20485
rect 24308 20476 24360 20528
rect 26700 20544 26752 20596
rect 29184 20544 29236 20596
rect 32128 20587 32180 20596
rect 26884 20476 26936 20528
rect 29460 20519 29512 20528
rect 29460 20485 29469 20519
rect 29469 20485 29503 20519
rect 29503 20485 29512 20519
rect 29460 20476 29512 20485
rect 30840 20476 30892 20528
rect 31484 20476 31536 20528
rect 23204 20408 23256 20460
rect 26608 20408 26660 20460
rect 26976 20451 27028 20460
rect 26976 20417 26985 20451
rect 26985 20417 27019 20451
rect 27019 20417 27028 20451
rect 26976 20408 27028 20417
rect 31668 20408 31720 20460
rect 15568 20315 15620 20324
rect 15568 20281 15577 20315
rect 15577 20281 15611 20315
rect 15611 20281 15620 20315
rect 15568 20272 15620 20281
rect 18512 20272 18564 20324
rect 20076 20272 20128 20324
rect 22284 20340 22336 20392
rect 23664 20383 23716 20392
rect 23020 20315 23072 20324
rect 23020 20281 23029 20315
rect 23029 20281 23063 20315
rect 23063 20281 23072 20315
rect 23020 20272 23072 20281
rect 23664 20349 23673 20383
rect 23673 20349 23707 20383
rect 23707 20349 23716 20383
rect 23664 20340 23716 20349
rect 23756 20340 23808 20392
rect 24032 20340 24084 20392
rect 24308 20272 24360 20324
rect 13820 20204 13872 20256
rect 15016 20204 15068 20256
rect 17408 20204 17460 20256
rect 18052 20204 18104 20256
rect 18880 20204 18932 20256
rect 21180 20247 21232 20256
rect 21180 20213 21189 20247
rect 21189 20213 21223 20247
rect 21223 20213 21232 20247
rect 21180 20204 21232 20213
rect 21364 20204 21416 20256
rect 21824 20204 21876 20256
rect 22008 20204 22060 20256
rect 25780 20340 25832 20392
rect 26056 20340 26108 20392
rect 26700 20340 26752 20392
rect 24952 20272 25004 20324
rect 25136 20272 25188 20324
rect 25044 20204 25096 20256
rect 27344 20340 27396 20392
rect 32128 20553 32137 20587
rect 32137 20553 32171 20587
rect 32171 20553 32180 20587
rect 32128 20544 32180 20553
rect 32956 20544 33008 20596
rect 33600 20519 33652 20528
rect 33600 20485 33609 20519
rect 33609 20485 33643 20519
rect 33643 20485 33652 20519
rect 33600 20476 33652 20485
rect 34152 20408 34204 20460
rect 35348 20476 35400 20528
rect 35716 20544 35768 20596
rect 36452 20476 36504 20528
rect 37004 20476 37056 20528
rect 34336 20340 34388 20392
rect 30748 20204 30800 20256
rect 30932 20247 30984 20256
rect 30932 20213 30941 20247
rect 30941 20213 30975 20247
rect 30975 20213 30984 20247
rect 31484 20247 31536 20256
rect 30932 20204 30984 20213
rect 31484 20213 31493 20247
rect 31493 20213 31527 20247
rect 31527 20213 31536 20247
rect 31484 20204 31536 20213
rect 34520 20340 34572 20392
rect 36084 20451 36136 20460
rect 36084 20417 36093 20451
rect 36093 20417 36127 20451
rect 36127 20417 36136 20451
rect 36084 20408 36136 20417
rect 39120 20544 39172 20596
rect 43168 20587 43220 20596
rect 43168 20553 43177 20587
rect 43177 20553 43211 20587
rect 43211 20553 43220 20587
rect 43168 20544 43220 20553
rect 45376 20587 45428 20596
rect 45376 20553 45385 20587
rect 45385 20553 45419 20587
rect 45419 20553 45428 20587
rect 45376 20544 45428 20553
rect 46480 20587 46532 20596
rect 46480 20553 46489 20587
rect 46489 20553 46523 20587
rect 46523 20553 46532 20587
rect 46480 20544 46532 20553
rect 38200 20476 38252 20528
rect 39948 20476 40000 20528
rect 42524 20476 42576 20528
rect 37648 20451 37700 20460
rect 37648 20417 37657 20451
rect 37657 20417 37691 20451
rect 37691 20417 37700 20451
rect 37648 20408 37700 20417
rect 37924 20451 37976 20460
rect 37924 20417 37933 20451
rect 37933 20417 37967 20451
rect 37967 20417 37976 20451
rect 37924 20408 37976 20417
rect 40316 20451 40368 20460
rect 35164 20340 35216 20392
rect 36636 20340 36688 20392
rect 38936 20383 38988 20392
rect 38936 20349 38945 20383
rect 38945 20349 38979 20383
rect 38979 20349 38988 20383
rect 38936 20340 38988 20349
rect 39212 20383 39264 20392
rect 39212 20349 39221 20383
rect 39221 20349 39255 20383
rect 39255 20349 39264 20383
rect 39212 20340 39264 20349
rect 37280 20272 37332 20324
rect 35164 20204 35216 20256
rect 38844 20272 38896 20324
rect 39948 20272 40000 20324
rect 40316 20417 40325 20451
rect 40325 20417 40359 20451
rect 40359 20417 40368 20451
rect 40316 20408 40368 20417
rect 42064 20408 42116 20460
rect 42616 20451 42668 20460
rect 42616 20417 42625 20451
rect 42625 20417 42659 20451
rect 42659 20417 42668 20451
rect 42616 20408 42668 20417
rect 43260 20451 43312 20460
rect 43260 20417 43269 20451
rect 43269 20417 43303 20451
rect 43303 20417 43312 20451
rect 43260 20408 43312 20417
rect 40224 20340 40276 20392
rect 40960 20340 41012 20392
rect 40500 20272 40552 20324
rect 41144 20272 41196 20324
rect 39304 20204 39356 20256
rect 40132 20204 40184 20256
rect 40684 20204 40736 20256
rect 41604 20247 41656 20256
rect 41604 20213 41613 20247
rect 41613 20213 41647 20247
rect 41647 20213 41656 20247
rect 41604 20204 41656 20213
rect 42524 20247 42576 20256
rect 42524 20213 42533 20247
rect 42533 20213 42567 20247
rect 42567 20213 42576 20247
rect 42524 20204 42576 20213
rect 44824 20247 44876 20256
rect 44824 20213 44833 20247
rect 44833 20213 44867 20247
rect 44867 20213 44876 20247
rect 44824 20204 44876 20213
rect 46020 20247 46072 20256
rect 46020 20213 46029 20247
rect 46029 20213 46063 20247
rect 46063 20213 46072 20247
rect 46020 20204 46072 20213
rect 10582 20102 10634 20154
rect 10646 20102 10698 20154
rect 10710 20102 10762 20154
rect 10774 20102 10826 20154
rect 10838 20102 10890 20154
rect 29846 20102 29898 20154
rect 29910 20102 29962 20154
rect 29974 20102 30026 20154
rect 30038 20102 30090 20154
rect 30102 20102 30154 20154
rect 49110 20102 49162 20154
rect 49174 20102 49226 20154
rect 49238 20102 49290 20154
rect 49302 20102 49354 20154
rect 49366 20102 49418 20154
rect 16580 20000 16632 20052
rect 18972 20000 19024 20052
rect 19984 20000 20036 20052
rect 27988 20000 28040 20052
rect 29000 20043 29052 20052
rect 29000 20009 29009 20043
rect 29009 20009 29043 20043
rect 29043 20009 29052 20043
rect 29000 20000 29052 20009
rect 12256 19975 12308 19984
rect 12256 19941 12265 19975
rect 12265 19941 12299 19975
rect 12299 19941 12308 19975
rect 12256 19932 12308 19941
rect 19156 19932 19208 19984
rect 21180 19975 21232 19984
rect 19432 19864 19484 19916
rect 12072 19796 12124 19848
rect 15108 19796 15160 19848
rect 16396 19796 16448 19848
rect 20628 19864 20680 19916
rect 21180 19941 21189 19975
rect 21189 19941 21223 19975
rect 21223 19941 21232 19975
rect 21180 19932 21232 19941
rect 22008 19864 22060 19916
rect 22468 19864 22520 19916
rect 22652 19907 22704 19916
rect 22652 19873 22661 19907
rect 22661 19873 22695 19907
rect 22695 19873 22704 19907
rect 22652 19864 22704 19873
rect 18512 19728 18564 19780
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 12992 19660 13044 19712
rect 13728 19660 13780 19712
rect 14832 19703 14884 19712
rect 14832 19669 14841 19703
rect 14841 19669 14875 19703
rect 14875 19669 14884 19703
rect 14832 19660 14884 19669
rect 16212 19660 16264 19712
rect 17868 19660 17920 19712
rect 19432 19771 19484 19780
rect 19432 19737 19441 19771
rect 19441 19737 19475 19771
rect 19475 19737 19484 19771
rect 19432 19728 19484 19737
rect 21180 19796 21232 19848
rect 22928 19839 22980 19848
rect 22928 19805 22937 19839
rect 22937 19805 22971 19839
rect 22971 19805 22980 19839
rect 22928 19796 22980 19805
rect 23664 19932 23716 19984
rect 24584 19932 24636 19984
rect 27160 19932 27212 19984
rect 28724 19932 28776 19984
rect 20996 19728 21048 19780
rect 25412 19864 25464 19916
rect 26608 19864 26660 19916
rect 26700 19864 26752 19916
rect 28264 19864 28316 19916
rect 30564 19864 30616 19916
rect 32680 19864 32732 19916
rect 33324 19864 33376 19916
rect 33876 19864 33928 19916
rect 36084 20000 36136 20052
rect 37556 20000 37608 20052
rect 37924 20000 37976 20052
rect 38660 20043 38712 20052
rect 38660 20009 38669 20043
rect 38669 20009 38703 20043
rect 38703 20009 38712 20043
rect 38660 20000 38712 20009
rect 39396 20000 39448 20052
rect 40776 20043 40828 20052
rect 40776 20009 40785 20043
rect 40785 20009 40819 20043
rect 40819 20009 40828 20043
rect 40776 20000 40828 20009
rect 41788 20043 41840 20052
rect 41788 20009 41797 20043
rect 41797 20009 41831 20043
rect 41831 20009 41840 20043
rect 41788 20000 41840 20009
rect 34980 19907 35032 19916
rect 34980 19873 34989 19907
rect 34989 19873 35023 19907
rect 35023 19873 35032 19907
rect 34980 19864 35032 19873
rect 39212 19932 39264 19984
rect 40040 19975 40092 19984
rect 40040 19941 40049 19975
rect 40049 19941 40083 19975
rect 40083 19941 40092 19975
rect 40040 19932 40092 19941
rect 40868 19975 40920 19984
rect 40868 19941 40877 19975
rect 40877 19941 40911 19975
rect 40911 19941 40920 19975
rect 40868 19932 40920 19941
rect 24124 19796 24176 19848
rect 24768 19796 24820 19848
rect 28632 19796 28684 19848
rect 29736 19796 29788 19848
rect 22100 19660 22152 19712
rect 23572 19660 23624 19712
rect 25412 19728 25464 19780
rect 26884 19728 26936 19780
rect 33692 19839 33744 19848
rect 33692 19805 33701 19839
rect 33701 19805 33735 19839
rect 33735 19805 33744 19839
rect 33692 19796 33744 19805
rect 24216 19660 24268 19712
rect 26700 19660 26752 19712
rect 29368 19660 29420 19712
rect 30196 19660 30248 19712
rect 32312 19728 32364 19780
rect 38752 19796 38804 19848
rect 38936 19796 38988 19848
rect 34888 19728 34940 19780
rect 35440 19728 35492 19780
rect 37096 19728 37148 19780
rect 37464 19728 37516 19780
rect 38844 19728 38896 19780
rect 39764 19796 39816 19848
rect 40040 19796 40092 19848
rect 30840 19660 30892 19712
rect 31852 19660 31904 19712
rect 36452 19703 36504 19712
rect 36452 19669 36461 19703
rect 36461 19669 36495 19703
rect 36495 19669 36504 19703
rect 36452 19660 36504 19669
rect 37556 19660 37608 19712
rect 39948 19660 40000 19712
rect 41052 19796 41104 19848
rect 41144 19728 41196 19780
rect 42156 19796 42208 19848
rect 42984 19796 43036 19848
rect 43812 19796 43864 19848
rect 44824 20000 44876 20052
rect 46480 20000 46532 20052
rect 46664 20043 46716 20052
rect 46664 20009 46673 20043
rect 46673 20009 46707 20043
rect 46707 20009 46716 20043
rect 46664 20000 46716 20009
rect 46940 19864 46992 19916
rect 46204 19796 46256 19848
rect 44088 19660 44140 19712
rect 44548 19660 44600 19712
rect 45560 19660 45612 19712
rect 46112 19660 46164 19712
rect 46296 19660 46348 19712
rect 47768 19703 47820 19712
rect 47768 19669 47777 19703
rect 47777 19669 47811 19703
rect 47811 19669 47820 19703
rect 47768 19660 47820 19669
rect 58164 19839 58216 19848
rect 58164 19805 58173 19839
rect 58173 19805 58207 19839
rect 58207 19805 58216 19839
rect 58164 19796 58216 19805
rect 51724 19660 51776 19712
rect 20214 19558 20266 19610
rect 20278 19558 20330 19610
rect 20342 19558 20394 19610
rect 20406 19558 20458 19610
rect 20470 19558 20522 19610
rect 39478 19558 39530 19610
rect 39542 19558 39594 19610
rect 39606 19558 39658 19610
rect 39670 19558 39722 19610
rect 39734 19558 39786 19610
rect 12072 19499 12124 19508
rect 12072 19465 12081 19499
rect 12081 19465 12115 19499
rect 12115 19465 12124 19499
rect 12072 19456 12124 19465
rect 20720 19499 20772 19508
rect 17776 19363 17828 19372
rect 17776 19329 17785 19363
rect 17785 19329 17819 19363
rect 17819 19329 17828 19363
rect 17776 19320 17828 19329
rect 18236 19388 18288 19440
rect 12348 19252 12400 19304
rect 15200 19252 15252 19304
rect 17224 19252 17276 19304
rect 16764 19227 16816 19236
rect 15016 19159 15068 19168
rect 15016 19125 15025 19159
rect 15025 19125 15059 19159
rect 15059 19125 15068 19159
rect 15016 19116 15068 19125
rect 16764 19193 16773 19227
rect 16773 19193 16807 19227
rect 16807 19193 16816 19227
rect 16764 19184 16816 19193
rect 17960 19252 18012 19304
rect 18328 19320 18380 19372
rect 19432 19388 19484 19440
rect 18880 19320 18932 19372
rect 19524 19320 19576 19372
rect 20720 19465 20729 19499
rect 20729 19465 20763 19499
rect 20763 19465 20772 19499
rect 20720 19456 20772 19465
rect 20904 19499 20956 19508
rect 20904 19465 20913 19499
rect 20913 19465 20947 19499
rect 20947 19465 20956 19499
rect 20904 19456 20956 19465
rect 21456 19456 21508 19508
rect 22192 19456 22244 19508
rect 23204 19456 23256 19508
rect 23664 19456 23716 19508
rect 19984 19388 20036 19440
rect 20444 19388 20496 19440
rect 19156 19295 19208 19304
rect 19156 19261 19165 19295
rect 19165 19261 19199 19295
rect 19199 19261 19208 19295
rect 19156 19252 19208 19261
rect 19340 19252 19392 19304
rect 19800 19252 19852 19304
rect 20352 19252 20404 19304
rect 20904 19320 20956 19372
rect 21732 19320 21784 19372
rect 22192 19363 22244 19372
rect 22192 19329 22201 19363
rect 22201 19329 22235 19363
rect 22235 19329 22244 19363
rect 22192 19320 22244 19329
rect 22376 19363 22428 19372
rect 22376 19329 22410 19363
rect 22410 19329 22428 19363
rect 22376 19320 22428 19329
rect 22652 19320 22704 19372
rect 22928 19320 22980 19372
rect 25596 19456 25648 19508
rect 25964 19456 26016 19508
rect 30196 19456 30248 19508
rect 26240 19388 26292 19440
rect 29736 19431 29788 19440
rect 29736 19397 29745 19431
rect 29745 19397 29779 19431
rect 29779 19397 29788 19431
rect 29736 19388 29788 19397
rect 36636 19456 36688 19508
rect 34612 19388 34664 19440
rect 35440 19388 35492 19440
rect 35900 19388 35952 19440
rect 24216 19363 24268 19372
rect 24216 19329 24225 19363
rect 24225 19329 24259 19363
rect 24259 19329 24268 19363
rect 24216 19320 24268 19329
rect 24492 19320 24544 19372
rect 27436 19320 27488 19372
rect 29276 19320 29328 19372
rect 29460 19320 29512 19372
rect 31576 19363 31628 19372
rect 31576 19329 31585 19363
rect 31585 19329 31619 19363
rect 31619 19329 31628 19363
rect 31576 19320 31628 19329
rect 34520 19320 34572 19372
rect 38292 19456 38344 19508
rect 39304 19456 39356 19508
rect 37556 19431 37608 19440
rect 37556 19397 37565 19431
rect 37565 19397 37599 19431
rect 37599 19397 37608 19431
rect 37556 19388 37608 19397
rect 46480 19456 46532 19508
rect 46664 19499 46716 19508
rect 46664 19465 46673 19499
rect 46673 19465 46707 19499
rect 46707 19465 46716 19499
rect 46664 19456 46716 19465
rect 58164 19499 58216 19508
rect 58164 19465 58173 19499
rect 58173 19465 58207 19499
rect 58207 19465 58216 19499
rect 58164 19456 58216 19465
rect 40408 19388 40460 19440
rect 40868 19388 40920 19440
rect 41236 19388 41288 19440
rect 44088 19388 44140 19440
rect 48872 19388 48924 19440
rect 39304 19320 39356 19372
rect 40132 19363 40184 19372
rect 40132 19329 40141 19363
rect 40141 19329 40175 19363
rect 40175 19329 40184 19363
rect 40132 19320 40184 19329
rect 42708 19363 42760 19372
rect 42708 19329 42717 19363
rect 42717 19329 42751 19363
rect 42751 19329 42760 19363
rect 42708 19320 42760 19329
rect 42800 19320 42852 19372
rect 42984 19320 43036 19372
rect 43168 19363 43220 19372
rect 43168 19329 43177 19363
rect 43177 19329 43211 19363
rect 43211 19329 43220 19363
rect 43168 19320 43220 19329
rect 43260 19363 43312 19372
rect 43260 19329 43269 19363
rect 43269 19329 43303 19363
rect 43303 19329 43312 19363
rect 43812 19363 43864 19372
rect 43260 19320 43312 19329
rect 43812 19329 43821 19363
rect 43821 19329 43855 19363
rect 43855 19329 43864 19363
rect 43812 19320 43864 19329
rect 44640 19320 44692 19372
rect 21272 19227 21324 19236
rect 18420 19116 18472 19168
rect 18696 19116 18748 19168
rect 19156 19116 19208 19168
rect 20260 19116 20312 19168
rect 21272 19193 21281 19227
rect 21281 19193 21315 19227
rect 21315 19193 21324 19227
rect 21272 19184 21324 19193
rect 22192 19184 22244 19236
rect 24492 19184 24544 19236
rect 26056 19116 26108 19168
rect 30932 19252 30984 19304
rect 32312 19252 32364 19304
rect 33416 19295 33468 19304
rect 33416 19261 33425 19295
rect 33425 19261 33459 19295
rect 33459 19261 33468 19295
rect 33416 19252 33468 19261
rect 35808 19252 35860 19304
rect 29000 19184 29052 19236
rect 36544 19252 36596 19304
rect 39488 19295 39540 19304
rect 39488 19261 39497 19295
rect 39497 19261 39531 19295
rect 39531 19261 39540 19295
rect 39488 19252 39540 19261
rect 39580 19252 39632 19304
rect 48688 19295 48740 19304
rect 48688 19261 48697 19295
rect 48697 19261 48731 19295
rect 48731 19261 48740 19295
rect 48688 19252 48740 19261
rect 41144 19227 41196 19236
rect 29276 19159 29328 19168
rect 29276 19125 29285 19159
rect 29285 19125 29319 19159
rect 29319 19125 29328 19159
rect 29276 19116 29328 19125
rect 29460 19116 29512 19168
rect 30288 19116 30340 19168
rect 30380 19116 30432 19168
rect 34152 19116 34204 19168
rect 34612 19116 34664 19168
rect 41144 19193 41153 19227
rect 41153 19193 41187 19227
rect 41187 19193 41196 19227
rect 41144 19184 41196 19193
rect 41880 19184 41932 19236
rect 42800 19184 42852 19236
rect 49700 19184 49752 19236
rect 36544 19116 36596 19168
rect 36728 19116 36780 19168
rect 39396 19116 39448 19168
rect 40960 19116 41012 19168
rect 41788 19116 41840 19168
rect 42984 19116 43036 19168
rect 43628 19116 43680 19168
rect 46204 19159 46256 19168
rect 46204 19125 46213 19159
rect 46213 19125 46247 19159
rect 46247 19125 46256 19159
rect 46204 19116 46256 19125
rect 10582 19014 10634 19066
rect 10646 19014 10698 19066
rect 10710 19014 10762 19066
rect 10774 19014 10826 19066
rect 10838 19014 10890 19066
rect 29846 19014 29898 19066
rect 29910 19014 29962 19066
rect 29974 19014 30026 19066
rect 30038 19014 30090 19066
rect 30102 19014 30154 19066
rect 49110 19014 49162 19066
rect 49174 19014 49226 19066
rect 49238 19014 49290 19066
rect 49302 19014 49354 19066
rect 49366 19014 49418 19066
rect 12256 18912 12308 18964
rect 15752 18912 15804 18964
rect 16120 18912 16172 18964
rect 17132 18912 17184 18964
rect 17592 18955 17644 18964
rect 17592 18921 17601 18955
rect 17601 18921 17635 18955
rect 17635 18921 17644 18955
rect 17592 18912 17644 18921
rect 16488 18844 16540 18896
rect 17040 18844 17092 18896
rect 18052 18844 18104 18896
rect 14188 18819 14240 18828
rect 14188 18785 14197 18819
rect 14197 18785 14231 18819
rect 14231 18785 14240 18819
rect 14188 18776 14240 18785
rect 14556 18776 14608 18828
rect 15660 18776 15712 18828
rect 17316 18776 17368 18828
rect 17408 18776 17460 18828
rect 17592 18776 17644 18828
rect 16580 18708 16632 18760
rect 15476 18572 15528 18624
rect 16304 18615 16356 18624
rect 16304 18581 16313 18615
rect 16313 18581 16347 18615
rect 16347 18581 16356 18615
rect 16304 18572 16356 18581
rect 16948 18615 17000 18624
rect 16948 18581 16957 18615
rect 16957 18581 16991 18615
rect 16991 18581 17000 18615
rect 17408 18640 17460 18692
rect 20260 18912 20312 18964
rect 20444 18955 20496 18964
rect 20444 18921 20453 18955
rect 20453 18921 20487 18955
rect 20487 18921 20496 18955
rect 20444 18912 20496 18921
rect 20536 18912 20588 18964
rect 26056 18912 26108 18964
rect 29000 18955 29052 18964
rect 19248 18844 19300 18896
rect 19892 18844 19944 18896
rect 21272 18844 21324 18896
rect 22008 18844 22060 18896
rect 29000 18921 29009 18955
rect 29009 18921 29043 18955
rect 29043 18921 29052 18955
rect 29000 18912 29052 18921
rect 33692 18912 33744 18964
rect 31208 18844 31260 18896
rect 34428 18844 34480 18896
rect 19984 18776 20036 18828
rect 20904 18776 20956 18828
rect 21088 18776 21140 18828
rect 21364 18776 21416 18828
rect 21732 18776 21784 18828
rect 21916 18776 21968 18828
rect 23848 18819 23900 18828
rect 23848 18785 23857 18819
rect 23857 18785 23891 18819
rect 23891 18785 23900 18819
rect 23848 18776 23900 18785
rect 23940 18776 23992 18828
rect 24216 18776 24268 18828
rect 31760 18776 31812 18828
rect 36544 18844 36596 18896
rect 18328 18751 18380 18760
rect 18328 18717 18337 18751
rect 18337 18717 18371 18751
rect 18371 18717 18380 18751
rect 18328 18708 18380 18717
rect 18696 18708 18748 18760
rect 19432 18708 19484 18760
rect 20352 18708 20404 18760
rect 20444 18708 20496 18760
rect 21272 18751 21324 18760
rect 21272 18717 21281 18751
rect 21281 18717 21315 18751
rect 21315 18717 21324 18751
rect 21272 18708 21324 18717
rect 21456 18708 21508 18760
rect 24584 18751 24636 18760
rect 24584 18717 24593 18751
rect 24593 18717 24627 18751
rect 24627 18717 24636 18751
rect 24584 18708 24636 18717
rect 24676 18708 24728 18760
rect 27252 18751 27304 18760
rect 27252 18717 27261 18751
rect 27261 18717 27295 18751
rect 27295 18717 27304 18751
rect 27252 18708 27304 18717
rect 29460 18708 29512 18760
rect 19248 18640 19300 18692
rect 20720 18640 20772 18692
rect 22376 18683 22428 18692
rect 22376 18649 22385 18683
rect 22385 18649 22419 18683
rect 22419 18649 22428 18683
rect 22376 18640 22428 18649
rect 24952 18640 25004 18692
rect 16948 18572 17000 18581
rect 18236 18572 18288 18624
rect 21088 18572 21140 18624
rect 21364 18615 21416 18624
rect 21364 18581 21373 18615
rect 21373 18581 21407 18615
rect 21407 18581 21416 18615
rect 21364 18572 21416 18581
rect 21640 18572 21692 18624
rect 21824 18572 21876 18624
rect 26976 18640 27028 18692
rect 25596 18572 25648 18624
rect 29736 18640 29788 18692
rect 31208 18708 31260 18760
rect 31024 18640 31076 18692
rect 34612 18776 34664 18828
rect 36360 18776 36412 18828
rect 38752 18844 38804 18896
rect 38568 18776 38620 18828
rect 34704 18751 34756 18760
rect 34704 18717 34713 18751
rect 34713 18717 34747 18751
rect 34747 18717 34756 18751
rect 34704 18708 34756 18717
rect 38476 18708 38528 18760
rect 39580 18844 39632 18896
rect 41972 18912 42024 18964
rect 42524 18844 42576 18896
rect 39212 18776 39264 18828
rect 40592 18776 40644 18828
rect 43628 18844 43680 18896
rect 46664 18844 46716 18896
rect 47860 18887 47912 18896
rect 47860 18853 47869 18887
rect 47869 18853 47903 18887
rect 47903 18853 47912 18887
rect 47860 18844 47912 18853
rect 39120 18751 39172 18760
rect 39120 18717 39129 18751
rect 39129 18717 39163 18751
rect 39163 18717 39172 18751
rect 39120 18708 39172 18717
rect 41236 18708 41288 18760
rect 32404 18683 32456 18692
rect 32404 18649 32413 18683
rect 32413 18649 32447 18683
rect 32447 18649 32456 18683
rect 32404 18640 32456 18649
rect 33968 18640 34020 18692
rect 35256 18640 35308 18692
rect 35440 18640 35492 18692
rect 36268 18640 36320 18692
rect 38200 18640 38252 18692
rect 27896 18572 27948 18624
rect 29828 18572 29880 18624
rect 30380 18572 30432 18624
rect 32128 18572 32180 18624
rect 34704 18572 34756 18624
rect 35072 18572 35124 18624
rect 35808 18572 35860 18624
rect 40408 18640 40460 18692
rect 39212 18615 39264 18624
rect 39212 18581 39221 18615
rect 39221 18581 39255 18615
rect 39255 18581 39264 18615
rect 39212 18572 39264 18581
rect 40316 18572 40368 18624
rect 43076 18776 43128 18828
rect 44456 18776 44508 18828
rect 48688 18776 48740 18828
rect 43260 18751 43312 18760
rect 43260 18717 43269 18751
rect 43269 18717 43303 18751
rect 43303 18717 43312 18751
rect 43260 18708 43312 18717
rect 43720 18751 43772 18760
rect 43720 18717 43729 18751
rect 43729 18717 43763 18751
rect 43763 18717 43772 18751
rect 43720 18708 43772 18717
rect 42892 18640 42944 18692
rect 58164 18751 58216 18760
rect 58164 18717 58173 18751
rect 58173 18717 58207 18751
rect 58207 18717 58216 18751
rect 58164 18708 58216 18717
rect 46296 18640 46348 18692
rect 57888 18683 57940 18692
rect 57888 18649 57897 18683
rect 57897 18649 57931 18683
rect 57931 18649 57940 18683
rect 57888 18640 57940 18649
rect 42984 18615 43036 18624
rect 42984 18581 42993 18615
rect 42993 18581 43027 18615
rect 43027 18581 43036 18615
rect 42984 18572 43036 18581
rect 43076 18572 43128 18624
rect 43628 18572 43680 18624
rect 43812 18615 43864 18624
rect 43812 18581 43821 18615
rect 43821 18581 43855 18615
rect 43855 18581 43864 18615
rect 43812 18572 43864 18581
rect 44548 18572 44600 18624
rect 45192 18572 45244 18624
rect 45652 18615 45704 18624
rect 45652 18581 45661 18615
rect 45661 18581 45695 18615
rect 45695 18581 45704 18615
rect 45652 18572 45704 18581
rect 20214 18470 20266 18522
rect 20278 18470 20330 18522
rect 20342 18470 20394 18522
rect 20406 18470 20458 18522
rect 20470 18470 20522 18522
rect 39478 18470 39530 18522
rect 39542 18470 39594 18522
rect 39606 18470 39658 18522
rect 39670 18470 39722 18522
rect 39734 18470 39786 18522
rect 12716 18343 12768 18352
rect 12716 18309 12725 18343
rect 12725 18309 12759 18343
rect 12759 18309 12768 18343
rect 12716 18300 12768 18309
rect 15200 18232 15252 18284
rect 16672 18275 16724 18284
rect 16672 18241 16681 18275
rect 16681 18241 16715 18275
rect 16715 18241 16724 18275
rect 16672 18232 16724 18241
rect 20996 18368 21048 18420
rect 21272 18368 21324 18420
rect 23020 18368 23072 18420
rect 23664 18368 23716 18420
rect 25596 18368 25648 18420
rect 25872 18368 25924 18420
rect 17316 18343 17368 18352
rect 17316 18309 17325 18343
rect 17325 18309 17359 18343
rect 17359 18309 17368 18343
rect 17316 18300 17368 18309
rect 18420 18300 18472 18352
rect 17408 18232 17460 18284
rect 18052 18232 18104 18284
rect 18512 18232 18564 18284
rect 18972 18232 19024 18284
rect 19616 18232 19668 18284
rect 20352 18275 20404 18284
rect 20352 18241 20361 18275
rect 20361 18241 20395 18275
rect 20395 18241 20404 18275
rect 20352 18232 20404 18241
rect 17316 18164 17368 18216
rect 17776 18164 17828 18216
rect 18880 18164 18932 18216
rect 20904 18232 20956 18284
rect 21732 18300 21784 18352
rect 21456 18232 21508 18284
rect 24952 18343 25004 18352
rect 24952 18309 24961 18343
rect 24961 18309 24995 18343
rect 24995 18309 25004 18343
rect 24952 18300 25004 18309
rect 25412 18300 25464 18352
rect 29092 18343 29144 18352
rect 29092 18309 29101 18343
rect 29101 18309 29135 18343
rect 29135 18309 29144 18343
rect 29092 18300 29144 18309
rect 30380 18368 30432 18420
rect 33784 18368 33836 18420
rect 38844 18368 38896 18420
rect 39028 18411 39080 18420
rect 39028 18377 39037 18411
rect 39037 18377 39071 18411
rect 39071 18377 39080 18411
rect 39028 18368 39080 18377
rect 39304 18368 39356 18420
rect 40132 18368 40184 18420
rect 22468 18275 22520 18284
rect 22468 18241 22477 18275
rect 22477 18241 22511 18275
rect 22511 18241 22520 18275
rect 22468 18232 22520 18241
rect 23848 18232 23900 18284
rect 31024 18232 31076 18284
rect 31392 18232 31444 18284
rect 16764 18139 16816 18148
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 12164 18071 12216 18080
rect 12164 18037 12173 18071
rect 12173 18037 12207 18071
rect 12207 18037 12216 18071
rect 12164 18028 12216 18037
rect 13820 18028 13872 18080
rect 14372 18071 14424 18080
rect 14372 18037 14381 18071
rect 14381 18037 14415 18071
rect 14415 18037 14424 18071
rect 14372 18028 14424 18037
rect 15016 18071 15068 18080
rect 15016 18037 15025 18071
rect 15025 18037 15059 18071
rect 15059 18037 15068 18071
rect 15016 18028 15068 18037
rect 16488 18028 16540 18080
rect 16764 18105 16773 18139
rect 16773 18105 16807 18139
rect 16807 18105 16816 18139
rect 16764 18096 16816 18105
rect 17592 18096 17644 18148
rect 18144 18028 18196 18080
rect 18328 18028 18380 18080
rect 18512 18071 18564 18080
rect 18512 18037 18521 18071
rect 18521 18037 18555 18071
rect 18555 18037 18564 18071
rect 18512 18028 18564 18037
rect 19616 18096 19668 18148
rect 19800 18096 19852 18148
rect 24216 18164 24268 18216
rect 27160 18164 27212 18216
rect 20720 18096 20772 18148
rect 29368 18164 29420 18216
rect 29460 18164 29512 18216
rect 30380 18164 30432 18216
rect 31208 18164 31260 18216
rect 32312 18164 32364 18216
rect 32772 18164 32824 18216
rect 33416 18207 33468 18216
rect 33416 18173 33425 18207
rect 33425 18173 33459 18207
rect 33459 18173 33468 18207
rect 33416 18164 33468 18173
rect 33784 18207 33836 18216
rect 33784 18173 33793 18207
rect 33793 18173 33827 18207
rect 33827 18173 33836 18207
rect 33784 18164 33836 18173
rect 21640 18028 21692 18080
rect 21916 18071 21968 18080
rect 21916 18037 21925 18071
rect 21925 18037 21959 18071
rect 21959 18037 21968 18071
rect 21916 18028 21968 18037
rect 23480 18028 23532 18080
rect 27896 18028 27948 18080
rect 32036 18096 32088 18148
rect 32496 18096 32548 18148
rect 32680 18096 32732 18148
rect 34704 18207 34756 18216
rect 34704 18173 34713 18207
rect 34713 18173 34747 18207
rect 34747 18173 34756 18207
rect 34704 18164 34756 18173
rect 35072 18164 35124 18216
rect 36268 18207 36320 18216
rect 33048 18028 33100 18080
rect 33416 18028 33468 18080
rect 33968 18028 34020 18080
rect 36268 18173 36277 18207
rect 36277 18173 36311 18207
rect 36311 18173 36320 18207
rect 36268 18164 36320 18173
rect 37464 18300 37516 18352
rect 37648 18300 37700 18352
rect 39212 18300 39264 18352
rect 41604 18368 41656 18420
rect 42432 18368 42484 18420
rect 44180 18368 44232 18420
rect 44456 18368 44508 18420
rect 45008 18411 45060 18420
rect 45008 18377 45017 18411
rect 45017 18377 45051 18411
rect 45051 18377 45060 18411
rect 45008 18368 45060 18377
rect 45100 18368 45152 18420
rect 45560 18411 45612 18420
rect 45560 18377 45569 18411
rect 45569 18377 45603 18411
rect 45603 18377 45612 18411
rect 45560 18368 45612 18377
rect 46112 18411 46164 18420
rect 46112 18377 46121 18411
rect 46121 18377 46155 18411
rect 46155 18377 46164 18411
rect 46112 18368 46164 18377
rect 46940 18368 46992 18420
rect 48688 18411 48740 18420
rect 48688 18377 48697 18411
rect 48697 18377 48731 18411
rect 48731 18377 48740 18411
rect 48688 18368 48740 18377
rect 58164 18411 58216 18420
rect 58164 18377 58173 18411
rect 58173 18377 58207 18411
rect 58207 18377 58216 18411
rect 58164 18368 58216 18377
rect 43812 18300 43864 18352
rect 38660 18232 38712 18284
rect 41328 18232 41380 18284
rect 41880 18275 41932 18284
rect 41880 18241 41889 18275
rect 41889 18241 41923 18275
rect 41923 18241 41932 18275
rect 41880 18232 41932 18241
rect 42800 18275 42852 18284
rect 42800 18241 42809 18275
rect 42809 18241 42843 18275
rect 42843 18241 42852 18275
rect 42800 18232 42852 18241
rect 43168 18232 43220 18284
rect 44916 18300 44968 18352
rect 38568 18096 38620 18148
rect 42064 18164 42116 18216
rect 42708 18164 42760 18216
rect 42892 18207 42944 18216
rect 42892 18173 42901 18207
rect 42901 18173 42935 18207
rect 42935 18173 42944 18207
rect 42892 18164 42944 18173
rect 43904 18164 43956 18216
rect 45008 18232 45060 18284
rect 46204 18232 46256 18284
rect 46572 18232 46624 18284
rect 48320 18232 48372 18284
rect 39396 18028 39448 18080
rect 39488 18071 39540 18080
rect 39488 18037 39497 18071
rect 39497 18037 39531 18071
rect 39531 18037 39540 18071
rect 45560 18096 45612 18148
rect 57888 18164 57940 18216
rect 39488 18028 39540 18037
rect 41328 18028 41380 18080
rect 41420 18028 41472 18080
rect 42708 18028 42760 18080
rect 49608 18028 49660 18080
rect 10582 17926 10634 17978
rect 10646 17926 10698 17978
rect 10710 17926 10762 17978
rect 10774 17926 10826 17978
rect 10838 17926 10890 17978
rect 29846 17926 29898 17978
rect 29910 17926 29962 17978
rect 29974 17926 30026 17978
rect 30038 17926 30090 17978
rect 30102 17926 30154 17978
rect 49110 17926 49162 17978
rect 49174 17926 49226 17978
rect 49238 17926 49290 17978
rect 49302 17926 49354 17978
rect 49366 17926 49418 17978
rect 13912 17824 13964 17876
rect 14556 17824 14608 17876
rect 15936 17867 15988 17876
rect 15936 17833 15945 17867
rect 15945 17833 15979 17867
rect 15979 17833 15988 17867
rect 15936 17824 15988 17833
rect 16120 17824 16172 17876
rect 18052 17824 18104 17876
rect 18144 17756 18196 17808
rect 18604 17824 18656 17876
rect 20720 17824 20772 17876
rect 21548 17867 21600 17876
rect 21548 17833 21557 17867
rect 21557 17833 21591 17867
rect 21591 17833 21600 17867
rect 21548 17824 21600 17833
rect 21732 17824 21784 17876
rect 22100 17824 22152 17876
rect 17408 17731 17460 17740
rect 17408 17697 17417 17731
rect 17417 17697 17451 17731
rect 17451 17697 17460 17731
rect 17408 17688 17460 17697
rect 19432 17756 19484 17808
rect 24584 17824 24636 17876
rect 16396 17620 16448 17672
rect 16488 17663 16540 17672
rect 16488 17629 16497 17663
rect 16497 17629 16531 17663
rect 16531 17629 16540 17663
rect 16488 17620 16540 17629
rect 16672 17620 16724 17672
rect 19064 17688 19116 17740
rect 16856 17552 16908 17604
rect 16948 17552 17000 17604
rect 17592 17620 17644 17672
rect 18788 17620 18840 17672
rect 19432 17663 19484 17672
rect 19432 17629 19441 17663
rect 19441 17629 19475 17663
rect 19475 17629 19484 17663
rect 19432 17620 19484 17629
rect 19616 17688 19668 17740
rect 21180 17688 21232 17740
rect 22468 17688 22520 17740
rect 22928 17688 22980 17740
rect 25688 17824 25740 17876
rect 26056 17688 26108 17740
rect 28540 17824 28592 17876
rect 28908 17824 28960 17876
rect 30656 17824 30708 17876
rect 31576 17824 31628 17876
rect 31760 17824 31812 17876
rect 39764 17824 39816 17876
rect 33692 17756 33744 17808
rect 35900 17756 35952 17808
rect 36728 17756 36780 17808
rect 38936 17756 38988 17808
rect 39304 17756 39356 17808
rect 44180 17824 44232 17876
rect 44272 17824 44324 17876
rect 45100 17867 45152 17876
rect 45100 17833 45109 17867
rect 45109 17833 45143 17867
rect 45143 17833 45152 17867
rect 45100 17824 45152 17833
rect 46480 17867 46532 17876
rect 46480 17833 46489 17867
rect 46489 17833 46523 17867
rect 46523 17833 46532 17867
rect 46480 17824 46532 17833
rect 48688 17824 48740 17876
rect 42248 17756 42300 17808
rect 43260 17799 43312 17808
rect 12992 17484 13044 17536
rect 18604 17484 18656 17536
rect 19248 17552 19300 17604
rect 20352 17620 20404 17672
rect 20720 17663 20772 17672
rect 20720 17629 20729 17663
rect 20729 17629 20763 17663
rect 20763 17629 20772 17663
rect 20720 17620 20772 17629
rect 20904 17620 20956 17672
rect 20996 17552 21048 17604
rect 23664 17620 23716 17672
rect 24400 17620 24452 17672
rect 27988 17688 28040 17740
rect 21272 17484 21324 17536
rect 22376 17552 22428 17604
rect 22836 17552 22888 17604
rect 24308 17552 24360 17604
rect 23020 17484 23072 17536
rect 24768 17484 24820 17536
rect 25136 17552 25188 17604
rect 27068 17552 27120 17604
rect 27528 17484 27580 17536
rect 29460 17620 29512 17672
rect 29552 17552 29604 17604
rect 30840 17484 30892 17536
rect 30932 17484 30984 17536
rect 35992 17688 36044 17740
rect 36820 17688 36872 17740
rect 37004 17731 37056 17740
rect 37004 17697 37013 17731
rect 37013 17697 37047 17731
rect 37047 17697 37056 17731
rect 37004 17688 37056 17697
rect 37280 17731 37332 17740
rect 37280 17697 37289 17731
rect 37289 17697 37323 17731
rect 37323 17697 37332 17731
rect 37280 17688 37332 17697
rect 37372 17688 37424 17740
rect 40960 17688 41012 17740
rect 43260 17765 43269 17799
rect 43269 17765 43303 17799
rect 43303 17765 43312 17799
rect 43260 17756 43312 17765
rect 42616 17688 42668 17740
rect 44640 17688 44692 17740
rect 44824 17688 44876 17740
rect 31668 17620 31720 17672
rect 41788 17620 41840 17672
rect 44088 17620 44140 17672
rect 31852 17552 31904 17604
rect 33048 17552 33100 17604
rect 34704 17595 34756 17604
rect 34704 17561 34713 17595
rect 34713 17561 34747 17595
rect 34747 17561 34756 17595
rect 34704 17552 34756 17561
rect 35072 17552 35124 17604
rect 37372 17552 37424 17604
rect 31392 17484 31444 17536
rect 32496 17484 32548 17536
rect 34888 17484 34940 17536
rect 39028 17484 39080 17536
rect 40592 17552 40644 17604
rect 41328 17595 41380 17604
rect 41328 17561 41337 17595
rect 41337 17561 41371 17595
rect 41371 17561 41380 17595
rect 41328 17552 41380 17561
rect 41880 17552 41932 17604
rect 44548 17620 44600 17672
rect 48228 17688 48280 17740
rect 46480 17620 46532 17672
rect 46664 17620 46716 17672
rect 41696 17484 41748 17536
rect 42064 17527 42116 17536
rect 42064 17493 42073 17527
rect 42073 17493 42107 17527
rect 42107 17493 42116 17527
rect 42064 17484 42116 17493
rect 42432 17527 42484 17536
rect 42432 17493 42441 17527
rect 42441 17493 42475 17527
rect 42475 17493 42484 17527
rect 42432 17484 42484 17493
rect 42800 17484 42852 17536
rect 47032 17527 47084 17536
rect 47032 17493 47041 17527
rect 47041 17493 47075 17527
rect 47075 17493 47084 17527
rect 47032 17484 47084 17493
rect 48228 17527 48280 17536
rect 48228 17493 48237 17527
rect 48237 17493 48271 17527
rect 48271 17493 48280 17527
rect 48228 17484 48280 17493
rect 50160 17527 50212 17536
rect 50160 17493 50169 17527
rect 50169 17493 50203 17527
rect 50203 17493 50212 17527
rect 50160 17484 50212 17493
rect 20214 17382 20266 17434
rect 20278 17382 20330 17434
rect 20342 17382 20394 17434
rect 20406 17382 20458 17434
rect 20470 17382 20522 17434
rect 39478 17382 39530 17434
rect 39542 17382 39594 17434
rect 39606 17382 39658 17434
rect 39670 17382 39722 17434
rect 39734 17382 39786 17434
rect 12716 17280 12768 17332
rect 16028 17280 16080 17332
rect 21180 17280 21232 17332
rect 21916 17280 21968 17332
rect 22836 17280 22888 17332
rect 14280 17144 14332 17196
rect 18972 17212 19024 17264
rect 19340 17255 19392 17264
rect 19340 17221 19349 17255
rect 19349 17221 19383 17255
rect 19383 17221 19392 17255
rect 19340 17212 19392 17221
rect 19432 17212 19484 17264
rect 12624 17076 12676 17128
rect 16856 17144 16908 17196
rect 19064 17144 19116 17196
rect 19984 17212 20036 17264
rect 22100 17212 22152 17264
rect 27712 17280 27764 17332
rect 28632 17280 28684 17332
rect 28908 17280 28960 17332
rect 29552 17280 29604 17332
rect 31668 17280 31720 17332
rect 23020 17212 23072 17264
rect 25044 17212 25096 17264
rect 27344 17255 27396 17264
rect 27344 17221 27353 17255
rect 27353 17221 27387 17255
rect 27387 17221 27396 17255
rect 27344 17212 27396 17221
rect 27804 17212 27856 17264
rect 30656 17212 30708 17264
rect 31484 17212 31536 17264
rect 20260 17144 20312 17196
rect 20444 17144 20496 17196
rect 20628 17144 20680 17196
rect 21088 17144 21140 17196
rect 21824 17187 21876 17196
rect 21824 17153 21833 17187
rect 21833 17153 21867 17187
rect 21867 17153 21876 17187
rect 21824 17144 21876 17153
rect 24676 17187 24728 17196
rect 24676 17153 24685 17187
rect 24685 17153 24719 17187
rect 24719 17153 24728 17187
rect 24676 17144 24728 17153
rect 26056 17144 26108 17196
rect 26608 17144 26660 17196
rect 26792 17144 26844 17196
rect 31852 17280 31904 17332
rect 33232 17280 33284 17332
rect 36728 17280 36780 17332
rect 37832 17280 37884 17332
rect 33048 17212 33100 17264
rect 37556 17212 37608 17264
rect 37648 17212 37700 17264
rect 39948 17212 40000 17264
rect 40592 17212 40644 17264
rect 41236 17280 41288 17332
rect 42708 17280 42760 17332
rect 41788 17212 41840 17264
rect 42156 17144 42208 17196
rect 44180 17212 44232 17264
rect 14832 17076 14884 17128
rect 11888 17008 11940 17060
rect 14004 17008 14056 17060
rect 14372 17008 14424 17060
rect 12624 16983 12676 16992
rect 12624 16949 12633 16983
rect 12633 16949 12667 16983
rect 12667 16949 12676 16983
rect 12624 16940 12676 16949
rect 13084 16983 13136 16992
rect 13084 16949 13093 16983
rect 13093 16949 13127 16983
rect 13127 16949 13136 16983
rect 13084 16940 13136 16949
rect 14096 16983 14148 16992
rect 14096 16949 14105 16983
rect 14105 16949 14139 16983
rect 14139 16949 14148 16983
rect 14096 16940 14148 16949
rect 14648 16983 14700 16992
rect 14648 16949 14657 16983
rect 14657 16949 14691 16983
rect 14691 16949 14700 16983
rect 14648 16940 14700 16949
rect 15292 16983 15344 16992
rect 15292 16949 15301 16983
rect 15301 16949 15335 16983
rect 15335 16949 15344 16983
rect 15292 16940 15344 16949
rect 15936 16983 15988 16992
rect 15936 16949 15945 16983
rect 15945 16949 15979 16983
rect 15979 16949 15988 16983
rect 15936 16940 15988 16949
rect 16396 16940 16448 16992
rect 18788 17076 18840 17128
rect 18880 17076 18932 17128
rect 19156 17076 19208 17128
rect 17500 17051 17552 17060
rect 17500 17017 17509 17051
rect 17509 17017 17543 17051
rect 17543 17017 17552 17051
rect 17500 17008 17552 17017
rect 19432 17119 19484 17128
rect 19432 17085 19466 17119
rect 19466 17085 19484 17119
rect 19432 17076 19484 17085
rect 19616 17076 19668 17128
rect 19800 17008 19852 17060
rect 18696 16940 18748 16992
rect 19616 16983 19668 16992
rect 19616 16949 19625 16983
rect 19625 16949 19659 16983
rect 19659 16949 19668 16983
rect 19616 16940 19668 16949
rect 20352 16940 20404 16992
rect 22376 17076 22428 17128
rect 23296 17076 23348 17128
rect 28540 17076 28592 17128
rect 31668 17076 31720 17128
rect 31760 17076 31812 17128
rect 21916 17051 21968 17060
rect 21916 17017 21925 17051
rect 21925 17017 21959 17051
rect 21959 17017 21968 17051
rect 21916 17008 21968 17017
rect 28908 17008 28960 17060
rect 21640 16940 21692 16992
rect 26240 16940 26292 16992
rect 29276 16940 29328 16992
rect 29460 16983 29512 16992
rect 29460 16949 29469 16983
rect 29469 16949 29503 16983
rect 29503 16949 29512 16983
rect 29460 16940 29512 16949
rect 31392 17008 31444 17060
rect 31852 16940 31904 16992
rect 34336 17076 34388 17128
rect 34888 17076 34940 17128
rect 33968 17008 34020 17060
rect 37556 17076 37608 17128
rect 39028 17076 39080 17128
rect 39304 17076 39356 17128
rect 35808 17008 35860 17060
rect 38108 17008 38160 17060
rect 43996 17119 44048 17128
rect 43996 17085 44005 17119
rect 44005 17085 44039 17119
rect 44039 17085 44048 17119
rect 43996 17076 44048 17085
rect 44180 17076 44232 17128
rect 45284 17144 45336 17196
rect 47032 17280 47084 17332
rect 48136 17280 48188 17332
rect 46020 17212 46072 17264
rect 48596 17212 48648 17264
rect 49608 17212 49660 17264
rect 45100 17076 45152 17128
rect 32772 16940 32824 16992
rect 32956 16940 33008 16992
rect 34152 16940 34204 16992
rect 38292 16940 38344 16992
rect 38660 16940 38712 16992
rect 42616 17008 42668 17060
rect 43260 17008 43312 17060
rect 46204 17144 46256 17196
rect 41512 16940 41564 16992
rect 41880 16940 41932 16992
rect 44916 16940 44968 16992
rect 45192 16983 45244 16992
rect 45192 16949 45201 16983
rect 45201 16949 45235 16983
rect 45235 16949 45244 16983
rect 45192 16940 45244 16949
rect 45652 16983 45704 16992
rect 45652 16949 45661 16983
rect 45661 16949 45695 16983
rect 45695 16949 45704 16983
rect 45652 16940 45704 16949
rect 46480 16983 46532 16992
rect 46480 16949 46489 16983
rect 46489 16949 46523 16983
rect 46523 16949 46532 16983
rect 46480 16940 46532 16949
rect 48964 16940 49016 16992
rect 10582 16838 10634 16890
rect 10646 16838 10698 16890
rect 10710 16838 10762 16890
rect 10774 16838 10826 16890
rect 10838 16838 10890 16890
rect 29846 16838 29898 16890
rect 29910 16838 29962 16890
rect 29974 16838 30026 16890
rect 30038 16838 30090 16890
rect 30102 16838 30154 16890
rect 49110 16838 49162 16890
rect 49174 16838 49226 16890
rect 49238 16838 49290 16890
rect 49302 16838 49354 16890
rect 49366 16838 49418 16890
rect 11888 16779 11940 16788
rect 11888 16745 11897 16779
rect 11897 16745 11931 16779
rect 11931 16745 11940 16779
rect 11888 16736 11940 16745
rect 14096 16736 14148 16788
rect 14648 16736 14700 16788
rect 14924 16736 14976 16788
rect 15384 16779 15436 16788
rect 15384 16745 15393 16779
rect 15393 16745 15427 16779
rect 15427 16745 15436 16779
rect 15384 16736 15436 16745
rect 16672 16736 16724 16788
rect 19432 16736 19484 16788
rect 20444 16736 20496 16788
rect 20904 16736 20956 16788
rect 22192 16736 22244 16788
rect 16764 16668 16816 16720
rect 16948 16668 17000 16720
rect 18696 16711 18748 16720
rect 18696 16677 18705 16711
rect 18705 16677 18739 16711
rect 18739 16677 18748 16711
rect 18696 16668 18748 16677
rect 18880 16668 18932 16720
rect 14832 16600 14884 16652
rect 16672 16600 16724 16652
rect 13084 16532 13136 16584
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 16028 16532 16080 16584
rect 16304 16532 16356 16584
rect 16488 16575 16540 16584
rect 16488 16541 16497 16575
rect 16497 16541 16531 16575
rect 16531 16541 16540 16575
rect 16488 16532 16540 16541
rect 17316 16575 17368 16584
rect 17316 16541 17325 16575
rect 17325 16541 17359 16575
rect 17359 16541 17368 16575
rect 17316 16532 17368 16541
rect 15200 16464 15252 16516
rect 15752 16464 15804 16516
rect 20536 16668 20588 16720
rect 20720 16668 20772 16720
rect 24952 16736 25004 16788
rect 29092 16736 29144 16788
rect 29276 16736 29328 16788
rect 31392 16736 31444 16788
rect 33140 16736 33192 16788
rect 33784 16736 33836 16788
rect 19340 16600 19392 16652
rect 21640 16643 21692 16652
rect 19800 16532 19852 16584
rect 19340 16464 19392 16516
rect 21640 16609 21649 16643
rect 21649 16609 21683 16643
rect 21683 16609 21692 16643
rect 21640 16600 21692 16609
rect 21732 16600 21784 16652
rect 23940 16600 23992 16652
rect 24952 16643 25004 16652
rect 24952 16609 24961 16643
rect 24961 16609 24995 16643
rect 24995 16609 25004 16643
rect 24952 16600 25004 16609
rect 27528 16668 27580 16720
rect 29000 16668 29052 16720
rect 29184 16668 29236 16720
rect 29920 16668 29972 16720
rect 31760 16668 31812 16720
rect 25596 16600 25648 16652
rect 25964 16600 26016 16652
rect 27804 16600 27856 16652
rect 21180 16575 21232 16584
rect 21180 16541 21189 16575
rect 21189 16541 21223 16575
rect 21223 16541 21232 16575
rect 21180 16532 21232 16541
rect 21272 16532 21324 16584
rect 22008 16532 22060 16584
rect 20260 16464 20312 16516
rect 20352 16464 20404 16516
rect 21548 16464 21600 16516
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 14648 16396 14700 16448
rect 18880 16396 18932 16448
rect 19708 16396 19760 16448
rect 19800 16439 19852 16448
rect 19800 16405 19809 16439
rect 19809 16405 19843 16439
rect 19843 16405 19852 16439
rect 20076 16439 20128 16448
rect 19800 16396 19852 16405
rect 20076 16405 20085 16439
rect 20085 16405 20119 16439
rect 20119 16405 20128 16439
rect 20076 16396 20128 16405
rect 21272 16396 21324 16448
rect 23756 16532 23808 16584
rect 24676 16532 24728 16584
rect 27160 16575 27212 16584
rect 27160 16541 27169 16575
rect 27169 16541 27203 16575
rect 27203 16541 27212 16575
rect 27160 16532 27212 16541
rect 29092 16600 29144 16652
rect 31852 16600 31904 16652
rect 33876 16668 33928 16720
rect 35440 16668 35492 16720
rect 34704 16643 34756 16652
rect 34704 16609 34713 16643
rect 34713 16609 34747 16643
rect 34747 16609 34756 16643
rect 34704 16600 34756 16609
rect 35072 16600 35124 16652
rect 29552 16532 29604 16584
rect 22284 16464 22336 16516
rect 25136 16464 25188 16516
rect 22560 16396 22612 16448
rect 23848 16439 23900 16448
rect 23848 16405 23857 16439
rect 23857 16405 23891 16439
rect 23891 16405 23900 16439
rect 23848 16396 23900 16405
rect 23940 16396 23992 16448
rect 26700 16439 26752 16448
rect 26700 16405 26709 16439
rect 26709 16405 26743 16439
rect 26743 16405 26752 16439
rect 26700 16396 26752 16405
rect 28724 16464 28776 16516
rect 29276 16464 29328 16516
rect 31208 16532 31260 16584
rect 36452 16532 36504 16584
rect 37648 16736 37700 16788
rect 38844 16736 38896 16788
rect 44272 16779 44324 16788
rect 44272 16745 44281 16779
rect 44281 16745 44315 16779
rect 44315 16745 44324 16779
rect 44272 16736 44324 16745
rect 45284 16736 45336 16788
rect 45744 16736 45796 16788
rect 48688 16779 48740 16788
rect 48688 16745 48697 16779
rect 48697 16745 48731 16779
rect 48731 16745 48740 16779
rect 48688 16736 48740 16745
rect 49608 16736 49660 16788
rect 38936 16668 38988 16720
rect 37280 16643 37332 16652
rect 37280 16609 37289 16643
rect 37289 16609 37323 16643
rect 37323 16609 37332 16643
rect 37280 16600 37332 16609
rect 37648 16600 37700 16652
rect 41604 16668 41656 16720
rect 43076 16711 43128 16720
rect 39212 16532 39264 16584
rect 31484 16464 31536 16516
rect 32496 16507 32548 16516
rect 32496 16473 32505 16507
rect 32505 16473 32539 16507
rect 32539 16473 32548 16507
rect 32496 16464 32548 16473
rect 32956 16464 33008 16516
rect 34520 16464 34572 16516
rect 35256 16464 35308 16516
rect 41972 16600 42024 16652
rect 42248 16600 42300 16652
rect 43076 16677 43085 16711
rect 43085 16677 43119 16711
rect 43119 16677 43128 16711
rect 43076 16668 43128 16677
rect 44640 16668 44692 16720
rect 45008 16643 45060 16652
rect 45008 16609 45017 16643
rect 45017 16609 45051 16643
rect 45051 16609 45060 16643
rect 45008 16600 45060 16609
rect 41788 16532 41840 16584
rect 33876 16396 33928 16448
rect 34336 16396 34388 16448
rect 40592 16464 40644 16516
rect 41420 16464 41472 16516
rect 42708 16532 42760 16584
rect 44548 16532 44600 16584
rect 47584 16532 47636 16584
rect 58164 16575 58216 16584
rect 58164 16541 58173 16575
rect 58173 16541 58207 16575
rect 58207 16541 58216 16575
rect 58164 16532 58216 16541
rect 39856 16396 39908 16448
rect 43904 16396 43956 16448
rect 45008 16396 45060 16448
rect 48964 16464 49016 16516
rect 45836 16439 45888 16448
rect 45836 16405 45845 16439
rect 45845 16405 45879 16439
rect 45879 16405 45888 16439
rect 45836 16396 45888 16405
rect 48596 16396 48648 16448
rect 20214 16294 20266 16346
rect 20278 16294 20330 16346
rect 20342 16294 20394 16346
rect 20406 16294 20458 16346
rect 20470 16294 20522 16346
rect 39478 16294 39530 16346
rect 39542 16294 39594 16346
rect 39606 16294 39658 16346
rect 39670 16294 39722 16346
rect 39734 16294 39786 16346
rect 12256 16235 12308 16244
rect 12256 16201 12265 16235
rect 12265 16201 12299 16235
rect 12299 16201 12308 16235
rect 12256 16192 12308 16201
rect 15200 16192 15252 16244
rect 15568 16167 15620 16176
rect 15568 16133 15577 16167
rect 15577 16133 15611 16167
rect 15611 16133 15620 16167
rect 15568 16124 15620 16133
rect 17316 16192 17368 16244
rect 17776 16124 17828 16176
rect 17040 16056 17092 16108
rect 12900 15988 12952 16040
rect 16120 15988 16172 16040
rect 17684 15988 17736 16040
rect 15200 15920 15252 15972
rect 17868 16099 17920 16108
rect 17868 16065 17877 16099
rect 17877 16065 17911 16099
rect 17911 16065 17920 16099
rect 17868 16056 17920 16065
rect 18420 16056 18472 16108
rect 18880 16124 18932 16176
rect 19064 16124 19116 16176
rect 20536 16124 20588 16176
rect 18696 16031 18748 16040
rect 18696 15997 18705 16031
rect 18705 15997 18739 16031
rect 18739 15997 18748 16031
rect 18696 15988 18748 15997
rect 19156 16031 19208 16040
rect 19156 15997 19165 16031
rect 19165 15997 19199 16031
rect 19199 15997 19208 16031
rect 19156 15988 19208 15997
rect 19892 16056 19944 16108
rect 20076 16056 20128 16108
rect 20720 16056 20772 16108
rect 19708 16031 19760 16040
rect 19708 15997 19717 16031
rect 19717 15997 19751 16031
rect 19751 15997 19760 16031
rect 19708 15988 19760 15997
rect 20168 15988 20220 16040
rect 24492 16124 24544 16176
rect 21640 16056 21692 16108
rect 21732 16056 21784 16108
rect 15108 15852 15160 15904
rect 16120 15895 16172 15904
rect 16120 15861 16129 15895
rect 16129 15861 16163 15895
rect 16163 15861 16172 15895
rect 16120 15852 16172 15861
rect 16304 15852 16356 15904
rect 20720 15920 20772 15972
rect 17868 15852 17920 15904
rect 18144 15895 18196 15904
rect 18144 15861 18153 15895
rect 18153 15861 18187 15895
rect 18187 15861 18196 15895
rect 18144 15852 18196 15861
rect 19156 15852 19208 15904
rect 19892 15852 19944 15904
rect 21088 16031 21140 16040
rect 21088 15997 21122 16031
rect 21122 15997 21140 16031
rect 22468 16031 22520 16040
rect 21088 15988 21140 15997
rect 22468 15997 22477 16031
rect 22477 15997 22511 16031
rect 22511 15997 22520 16031
rect 22468 15988 22520 15997
rect 22744 16031 22796 16040
rect 22744 15997 22753 16031
rect 22753 15997 22787 16031
rect 22787 15997 22796 16031
rect 22744 15988 22796 15997
rect 23112 15988 23164 16040
rect 25228 16192 25280 16244
rect 25504 16192 25556 16244
rect 27528 16192 27580 16244
rect 31576 16192 31628 16244
rect 32956 16192 33008 16244
rect 34612 16192 34664 16244
rect 35256 16192 35308 16244
rect 35348 16192 35400 16244
rect 38660 16192 38712 16244
rect 39396 16192 39448 16244
rect 41052 16192 41104 16244
rect 44548 16192 44600 16244
rect 44732 16192 44784 16244
rect 47584 16235 47636 16244
rect 47584 16201 47593 16235
rect 47593 16201 47627 16235
rect 47627 16201 47636 16235
rect 47584 16192 47636 16201
rect 48688 16192 48740 16244
rect 58164 16235 58216 16244
rect 58164 16201 58173 16235
rect 58173 16201 58207 16235
rect 58207 16201 58216 16235
rect 58164 16192 58216 16201
rect 26148 16167 26200 16176
rect 26148 16133 26157 16167
rect 26157 16133 26191 16167
rect 26191 16133 26200 16167
rect 26148 16124 26200 16133
rect 26424 16099 26476 16108
rect 26424 16065 26433 16099
rect 26433 16065 26467 16099
rect 26467 16065 26476 16099
rect 26424 16056 26476 16065
rect 29460 16124 29512 16176
rect 27160 16056 27212 16108
rect 29920 16124 29972 16176
rect 30748 16124 30800 16176
rect 34152 16124 34204 16176
rect 37464 16124 37516 16176
rect 45836 16124 45888 16176
rect 48136 16124 48188 16176
rect 30196 16099 30248 16108
rect 30196 16065 30205 16099
rect 30205 16065 30239 16099
rect 30239 16065 30248 16099
rect 30196 16056 30248 16065
rect 31208 16056 31260 16108
rect 33508 16056 33560 16108
rect 33784 16056 33836 16108
rect 39028 16099 39080 16108
rect 39028 16065 39037 16099
rect 39037 16065 39071 16099
rect 39071 16065 39080 16099
rect 39856 16099 39908 16108
rect 39028 16056 39080 16065
rect 39856 16065 39865 16099
rect 39865 16065 39899 16099
rect 39899 16065 39908 16099
rect 39856 16056 39908 16065
rect 40132 16099 40184 16108
rect 40132 16065 40141 16099
rect 40141 16065 40175 16099
rect 40175 16065 40184 16099
rect 40132 16056 40184 16065
rect 22376 15920 22428 15972
rect 24216 15963 24268 15972
rect 24216 15929 24225 15963
rect 24225 15929 24259 15963
rect 24259 15929 24268 15963
rect 24216 15920 24268 15929
rect 21640 15852 21692 15904
rect 24860 15920 24912 15972
rect 24768 15852 24820 15904
rect 28724 15852 28776 15904
rect 30840 15988 30892 16040
rect 31576 15988 31628 16040
rect 33876 15988 33928 16040
rect 33968 16031 34020 16040
rect 33968 15997 33977 16031
rect 33977 15997 34011 16031
rect 34011 15997 34020 16031
rect 33968 15988 34020 15997
rect 34796 15988 34848 16040
rect 33692 15920 33744 15972
rect 34152 15920 34204 15972
rect 35072 15988 35124 16040
rect 38752 16031 38804 16040
rect 38752 15997 38761 16031
rect 38761 15997 38795 16031
rect 38795 15997 38804 16031
rect 38752 15988 38804 15997
rect 42248 16056 42300 16108
rect 40960 15988 41012 16040
rect 40224 15920 40276 15972
rect 42800 16099 42852 16108
rect 42800 16065 42809 16099
rect 42809 16065 42843 16099
rect 42843 16065 42852 16099
rect 42800 16056 42852 16065
rect 42892 16099 42944 16108
rect 42892 16065 42901 16099
rect 42901 16065 42935 16099
rect 42935 16065 42944 16099
rect 42892 16056 42944 16065
rect 42524 15988 42576 16040
rect 43444 16099 43496 16108
rect 43444 16065 43453 16099
rect 43453 16065 43487 16099
rect 43487 16065 43496 16099
rect 44364 16099 44416 16108
rect 43444 16056 43496 16065
rect 44364 16065 44373 16099
rect 44373 16065 44407 16099
rect 44407 16065 44416 16099
rect 44364 16056 44416 16065
rect 43628 16031 43680 16040
rect 43628 15997 43637 16031
rect 43637 15997 43671 16031
rect 43671 15997 43680 16031
rect 43628 15988 43680 15997
rect 43812 15988 43864 16040
rect 48320 16056 48372 16108
rect 49792 16099 49844 16108
rect 49792 16065 49801 16099
rect 49801 16065 49835 16099
rect 49835 16065 49844 16099
rect 49792 16056 49844 16065
rect 43168 15920 43220 15972
rect 43444 15920 43496 15972
rect 43720 15920 43772 15972
rect 46388 15988 46440 16040
rect 30288 15852 30340 15904
rect 30840 15852 30892 15904
rect 35348 15852 35400 15904
rect 39028 15852 39080 15904
rect 40960 15852 41012 15904
rect 41880 15852 41932 15904
rect 42432 15895 42484 15904
rect 42432 15861 42441 15895
rect 42441 15861 42475 15895
rect 42475 15861 42484 15895
rect 42432 15852 42484 15861
rect 43996 15852 44048 15904
rect 44180 15895 44232 15904
rect 44180 15861 44189 15895
rect 44189 15861 44223 15895
rect 44223 15861 44232 15895
rect 44180 15852 44232 15861
rect 44548 15852 44600 15904
rect 44916 15895 44968 15904
rect 44916 15861 44925 15895
rect 44925 15861 44959 15895
rect 44959 15861 44968 15895
rect 44916 15852 44968 15861
rect 45744 15852 45796 15904
rect 46020 15895 46072 15904
rect 46020 15861 46029 15895
rect 46029 15861 46063 15895
rect 46063 15861 46072 15895
rect 46020 15852 46072 15861
rect 10582 15750 10634 15802
rect 10646 15750 10698 15802
rect 10710 15750 10762 15802
rect 10774 15750 10826 15802
rect 10838 15750 10890 15802
rect 29846 15750 29898 15802
rect 29910 15750 29962 15802
rect 29974 15750 30026 15802
rect 30038 15750 30090 15802
rect 30102 15750 30154 15802
rect 49110 15750 49162 15802
rect 49174 15750 49226 15802
rect 49238 15750 49290 15802
rect 49302 15750 49354 15802
rect 49366 15750 49418 15802
rect 14280 15648 14332 15700
rect 15200 15648 15252 15700
rect 15660 15691 15712 15700
rect 15660 15657 15669 15691
rect 15669 15657 15703 15691
rect 15703 15657 15712 15691
rect 15660 15648 15712 15657
rect 20076 15648 20128 15700
rect 21088 15648 21140 15700
rect 21272 15648 21324 15700
rect 15844 15580 15896 15632
rect 21180 15580 21232 15632
rect 15660 15512 15712 15564
rect 16212 15512 16264 15564
rect 18328 15512 18380 15564
rect 17684 15444 17736 15496
rect 20904 15555 20956 15564
rect 19708 15444 19760 15496
rect 20904 15521 20913 15555
rect 20913 15521 20947 15555
rect 20947 15521 20956 15555
rect 20904 15512 20956 15521
rect 20168 15444 20220 15496
rect 20536 15444 20588 15496
rect 20720 15487 20772 15496
rect 20720 15453 20729 15487
rect 20729 15453 20763 15487
rect 20763 15453 20772 15487
rect 21548 15512 21600 15564
rect 21364 15487 21416 15496
rect 20720 15444 20772 15453
rect 21364 15453 21373 15487
rect 21373 15453 21407 15487
rect 21407 15453 21416 15487
rect 21364 15444 21416 15453
rect 22652 15648 22704 15700
rect 23480 15648 23532 15700
rect 24032 15648 24084 15700
rect 25412 15648 25464 15700
rect 21732 15580 21784 15632
rect 24124 15580 24176 15632
rect 24584 15580 24636 15632
rect 25136 15580 25188 15632
rect 29552 15580 29604 15632
rect 32312 15580 32364 15632
rect 32772 15580 32824 15632
rect 39856 15580 39908 15632
rect 22192 15444 22244 15496
rect 15108 15376 15160 15428
rect 18512 15419 18564 15428
rect 18512 15385 18521 15419
rect 18521 15385 18555 15419
rect 18555 15385 18564 15419
rect 18512 15376 18564 15385
rect 11244 15351 11296 15360
rect 11244 15317 11253 15351
rect 11253 15317 11287 15351
rect 11287 15317 11296 15351
rect 11244 15308 11296 15317
rect 12992 15351 13044 15360
rect 12992 15317 13001 15351
rect 13001 15317 13035 15351
rect 13035 15317 13044 15351
rect 12992 15308 13044 15317
rect 17316 15351 17368 15360
rect 17316 15317 17325 15351
rect 17325 15317 17359 15351
rect 17359 15317 17368 15351
rect 17316 15308 17368 15317
rect 17868 15351 17920 15360
rect 17868 15317 17877 15351
rect 17877 15317 17911 15351
rect 17911 15317 17920 15351
rect 17868 15308 17920 15317
rect 18420 15308 18472 15360
rect 20076 15308 20128 15360
rect 20904 15308 20956 15360
rect 22100 15376 22152 15428
rect 26424 15512 26476 15564
rect 26792 15555 26844 15564
rect 26792 15521 26801 15555
rect 26801 15521 26835 15555
rect 26835 15521 26844 15555
rect 26792 15512 26844 15521
rect 28540 15512 28592 15564
rect 36544 15512 36596 15564
rect 36820 15512 36872 15564
rect 38384 15512 38436 15564
rect 41052 15648 41104 15700
rect 41512 15648 41564 15700
rect 42524 15691 42576 15700
rect 42524 15657 42533 15691
rect 42533 15657 42567 15691
rect 42567 15657 42576 15691
rect 42524 15648 42576 15657
rect 43352 15691 43404 15700
rect 43352 15657 43361 15691
rect 43361 15657 43395 15691
rect 43395 15657 43404 15691
rect 43352 15648 43404 15657
rect 43444 15648 43496 15700
rect 45192 15648 45244 15700
rect 45560 15691 45612 15700
rect 45560 15657 45569 15691
rect 45569 15657 45603 15691
rect 45603 15657 45612 15691
rect 45560 15648 45612 15657
rect 47584 15648 47636 15700
rect 48688 15648 48740 15700
rect 42340 15580 42392 15632
rect 42616 15623 42668 15632
rect 42616 15589 42625 15623
rect 42625 15589 42659 15623
rect 42659 15589 42668 15623
rect 42616 15580 42668 15589
rect 44456 15580 44508 15632
rect 41696 15512 41748 15564
rect 23572 15376 23624 15428
rect 23296 15308 23348 15360
rect 24676 15444 24728 15496
rect 27252 15487 27304 15496
rect 27252 15453 27261 15487
rect 27261 15453 27295 15487
rect 27295 15453 27304 15487
rect 27252 15444 27304 15453
rect 32312 15487 32364 15496
rect 32312 15453 32321 15487
rect 32321 15453 32355 15487
rect 32355 15453 32364 15487
rect 32312 15444 32364 15453
rect 34612 15444 34664 15496
rect 36452 15487 36504 15496
rect 36452 15453 36461 15487
rect 36461 15453 36495 15487
rect 36495 15453 36504 15487
rect 36452 15444 36504 15453
rect 38936 15444 38988 15496
rect 39396 15444 39448 15496
rect 25964 15376 26016 15428
rect 26148 15308 26200 15360
rect 27988 15376 28040 15428
rect 29552 15376 29604 15428
rect 30288 15376 30340 15428
rect 31576 15419 31628 15428
rect 28448 15308 28500 15360
rect 29644 15308 29696 15360
rect 30196 15308 30248 15360
rect 30656 15308 30708 15360
rect 30840 15308 30892 15360
rect 31576 15385 31585 15419
rect 31585 15385 31619 15419
rect 31619 15385 31628 15419
rect 31576 15376 31628 15385
rect 31944 15376 31996 15428
rect 32588 15376 32640 15428
rect 33048 15376 33100 15428
rect 33140 15376 33192 15428
rect 33968 15376 34020 15428
rect 36176 15419 36228 15428
rect 31484 15308 31536 15360
rect 32312 15308 32364 15360
rect 34612 15308 34664 15360
rect 36176 15385 36185 15419
rect 36185 15385 36219 15419
rect 36219 15385 36228 15419
rect 36176 15376 36228 15385
rect 37280 15376 37332 15428
rect 38844 15376 38896 15428
rect 39948 15376 40000 15428
rect 40592 15444 40644 15496
rect 41972 15487 42024 15496
rect 41972 15453 41981 15487
rect 41981 15453 42015 15487
rect 42015 15453 42024 15487
rect 41972 15444 42024 15453
rect 41144 15376 41196 15428
rect 43168 15487 43220 15496
rect 43168 15453 43177 15487
rect 43177 15453 43211 15487
rect 43211 15453 43220 15487
rect 43168 15444 43220 15453
rect 43720 15444 43772 15496
rect 58164 15487 58216 15496
rect 58164 15453 58173 15487
rect 58173 15453 58207 15487
rect 58207 15453 58216 15487
rect 58164 15444 58216 15453
rect 42524 15376 42576 15428
rect 43352 15376 43404 15428
rect 57888 15419 57940 15428
rect 57888 15385 57897 15419
rect 57897 15385 57931 15419
rect 57931 15385 57940 15419
rect 57888 15376 57940 15385
rect 39304 15308 39356 15360
rect 41880 15308 41932 15360
rect 42340 15308 42392 15360
rect 42984 15308 43036 15360
rect 43628 15308 43680 15360
rect 43996 15351 44048 15360
rect 43996 15317 44005 15351
rect 44005 15317 44039 15351
rect 44039 15317 44048 15351
rect 43996 15308 44048 15317
rect 46388 15308 46440 15360
rect 48320 15351 48372 15360
rect 48320 15317 48329 15351
rect 48329 15317 48363 15351
rect 48363 15317 48372 15351
rect 48320 15308 48372 15317
rect 48596 15308 48648 15360
rect 20214 15206 20266 15258
rect 20278 15206 20330 15258
rect 20342 15206 20394 15258
rect 20406 15206 20458 15258
rect 20470 15206 20522 15258
rect 39478 15206 39530 15258
rect 39542 15206 39594 15258
rect 39606 15206 39658 15258
rect 39670 15206 39722 15258
rect 39734 15206 39786 15258
rect 12716 15104 12768 15156
rect 13636 15104 13688 15156
rect 15200 15104 15252 15156
rect 18512 15104 18564 15156
rect 19248 15104 19300 15156
rect 17684 15036 17736 15088
rect 18052 15036 18104 15088
rect 20904 15104 20956 15156
rect 21732 15104 21784 15156
rect 21824 15104 21876 15156
rect 22284 15104 22336 15156
rect 23112 15104 23164 15156
rect 23848 15104 23900 15156
rect 25688 15104 25740 15156
rect 30564 15104 30616 15156
rect 31024 15104 31076 15156
rect 31576 15104 31628 15156
rect 31852 15104 31904 15156
rect 34428 15104 34480 15156
rect 35716 15104 35768 15156
rect 37372 15104 37424 15156
rect 38200 15104 38252 15156
rect 40592 15104 40644 15156
rect 43536 15147 43588 15156
rect 43536 15113 43545 15147
rect 43545 15113 43579 15147
rect 43579 15113 43588 15147
rect 43536 15104 43588 15113
rect 43628 15104 43680 15156
rect 44180 15147 44232 15156
rect 11244 14968 11296 15020
rect 17316 15011 17368 15020
rect 17316 14977 17325 15011
rect 17325 14977 17359 15011
rect 17359 14977 17368 15011
rect 17316 14968 17368 14977
rect 18144 14968 18196 15020
rect 19064 15011 19116 15020
rect 19064 14977 19073 15011
rect 19073 14977 19107 15011
rect 19107 14977 19116 15011
rect 19064 14968 19116 14977
rect 19248 15011 19300 15020
rect 19248 14977 19257 15011
rect 19257 14977 19291 15011
rect 19291 14977 19300 15011
rect 19248 14968 19300 14977
rect 20076 14968 20128 15020
rect 16120 14900 16172 14952
rect 1492 14875 1544 14884
rect 1492 14841 1501 14875
rect 1501 14841 1535 14875
rect 1535 14841 1544 14875
rect 1492 14832 1544 14841
rect 17224 14832 17276 14884
rect 18880 14832 18932 14884
rect 18972 14832 19024 14884
rect 19340 14832 19392 14884
rect 20260 14900 20312 14952
rect 21548 15036 21600 15088
rect 23940 15036 23992 15088
rect 24860 15036 24912 15088
rect 28540 15036 28592 15088
rect 29000 15079 29052 15088
rect 29000 15045 29009 15079
rect 29009 15045 29043 15079
rect 29043 15045 29052 15079
rect 29000 15036 29052 15045
rect 21732 14968 21784 15020
rect 22100 14968 22152 15020
rect 22652 14968 22704 15020
rect 22928 14968 22980 15020
rect 23204 14968 23256 15020
rect 23480 14968 23532 15020
rect 23756 14968 23808 15020
rect 24400 14968 24452 15020
rect 23388 14943 23440 14952
rect 23388 14909 23397 14943
rect 23397 14909 23431 14943
rect 23431 14909 23440 14943
rect 24676 14943 24728 14952
rect 23388 14900 23440 14909
rect 24676 14909 24685 14943
rect 24685 14909 24719 14943
rect 24719 14909 24728 14943
rect 24676 14900 24728 14909
rect 24952 14943 25004 14952
rect 24952 14909 24961 14943
rect 24961 14909 24995 14943
rect 24995 14909 25004 14943
rect 24952 14900 25004 14909
rect 25320 14900 25372 14952
rect 26792 14968 26844 15020
rect 29552 15036 29604 15088
rect 30840 15036 30892 15088
rect 31668 15036 31720 15088
rect 32864 15036 32916 15088
rect 32128 15011 32180 15020
rect 26240 14900 26292 14952
rect 32128 14977 32137 15011
rect 32137 14977 32171 15011
rect 32171 14977 32180 15011
rect 32128 14968 32180 14977
rect 35256 15036 35308 15088
rect 36544 15036 36596 15088
rect 37648 14968 37700 15020
rect 38200 15011 38252 15020
rect 30380 14943 30432 14952
rect 21824 14832 21876 14884
rect 21916 14832 21968 14884
rect 20168 14807 20220 14816
rect 20168 14773 20177 14807
rect 20177 14773 20211 14807
rect 20211 14773 20220 14807
rect 20168 14764 20220 14773
rect 20352 14764 20404 14816
rect 20628 14764 20680 14816
rect 21548 14764 21600 14816
rect 22100 14764 22152 14816
rect 22284 14832 22336 14884
rect 22744 14764 22796 14816
rect 22928 14807 22980 14816
rect 22928 14773 22937 14807
rect 22937 14773 22971 14807
rect 22971 14773 22980 14807
rect 22928 14764 22980 14773
rect 26700 14764 26752 14816
rect 27528 14807 27580 14816
rect 27528 14773 27537 14807
rect 27537 14773 27571 14807
rect 27571 14773 27580 14807
rect 27528 14764 27580 14773
rect 29552 14832 29604 14884
rect 30380 14909 30389 14943
rect 30389 14909 30423 14943
rect 30423 14909 30432 14943
rect 30380 14900 30432 14909
rect 32680 14900 32732 14952
rect 34152 14900 34204 14952
rect 34704 14943 34756 14952
rect 34704 14909 34713 14943
rect 34713 14909 34747 14943
rect 34747 14909 34756 14943
rect 34704 14900 34756 14909
rect 36820 14900 36872 14952
rect 38200 14977 38209 15011
rect 38209 14977 38243 15011
rect 38243 14977 38252 15011
rect 38200 14968 38252 14977
rect 39396 14968 39448 15020
rect 39948 14968 40000 15020
rect 40224 14968 40276 15020
rect 41052 14968 41104 15020
rect 41788 15036 41840 15088
rect 44180 15113 44189 15147
rect 44189 15113 44223 15147
rect 44223 15113 44232 15147
rect 44180 15104 44232 15113
rect 46388 15147 46440 15156
rect 46388 15113 46397 15147
rect 46397 15113 46431 15147
rect 46431 15113 46440 15147
rect 46388 15104 46440 15113
rect 46480 15104 46532 15156
rect 47584 15147 47636 15156
rect 47584 15113 47593 15147
rect 47593 15113 47627 15147
rect 47627 15113 47636 15147
rect 47584 15104 47636 15113
rect 44088 15036 44140 15088
rect 46664 15036 46716 15088
rect 46940 15079 46992 15088
rect 46940 15045 46949 15079
rect 46949 15045 46983 15079
rect 46983 15045 46992 15079
rect 46940 15036 46992 15045
rect 58164 15079 58216 15088
rect 58164 15045 58173 15079
rect 58173 15045 58207 15079
rect 58207 15045 58216 15079
rect 58164 15036 58216 15045
rect 32036 14832 32088 14884
rect 33692 14832 33744 14884
rect 40592 14900 40644 14952
rect 40868 14943 40920 14952
rect 40868 14909 40877 14943
rect 40877 14909 40911 14943
rect 40911 14909 40920 14943
rect 40868 14900 40920 14909
rect 41788 14900 41840 14952
rect 33416 14764 33468 14816
rect 36176 14807 36228 14816
rect 36176 14773 36185 14807
rect 36185 14773 36219 14807
rect 36219 14773 36228 14807
rect 36176 14764 36228 14773
rect 36636 14807 36688 14816
rect 36636 14773 36645 14807
rect 36645 14773 36679 14807
rect 36679 14773 36688 14807
rect 36636 14764 36688 14773
rect 37924 14764 37976 14816
rect 38108 14764 38160 14816
rect 38844 14764 38896 14816
rect 40776 14832 40828 14884
rect 40040 14764 40092 14816
rect 40408 14764 40460 14816
rect 40684 14807 40736 14816
rect 40684 14773 40693 14807
rect 40693 14773 40727 14807
rect 40727 14773 40736 14807
rect 40684 14764 40736 14773
rect 41788 14807 41840 14816
rect 41788 14773 41797 14807
rect 41797 14773 41831 14807
rect 41831 14773 41840 14807
rect 42156 14900 42208 14952
rect 42524 14900 42576 14952
rect 44180 14900 44232 14952
rect 44640 14900 44692 14952
rect 45284 14875 45336 14884
rect 45284 14841 45293 14875
rect 45293 14841 45327 14875
rect 45327 14841 45336 14875
rect 45284 14832 45336 14841
rect 41788 14764 41840 14773
rect 42892 14764 42944 14816
rect 43076 14764 43128 14816
rect 44088 14764 44140 14816
rect 48136 14807 48188 14816
rect 48136 14773 48145 14807
rect 48145 14773 48179 14807
rect 48179 14773 48188 14807
rect 48136 14764 48188 14773
rect 10582 14662 10634 14714
rect 10646 14662 10698 14714
rect 10710 14662 10762 14714
rect 10774 14662 10826 14714
rect 10838 14662 10890 14714
rect 29846 14662 29898 14714
rect 29910 14662 29962 14714
rect 29974 14662 30026 14714
rect 30038 14662 30090 14714
rect 30102 14662 30154 14714
rect 49110 14662 49162 14714
rect 49174 14662 49226 14714
rect 49238 14662 49290 14714
rect 49302 14662 49354 14714
rect 49366 14662 49418 14714
rect 14280 14603 14332 14612
rect 14280 14569 14289 14603
rect 14289 14569 14323 14603
rect 14323 14569 14332 14603
rect 14280 14560 14332 14569
rect 15384 14603 15436 14612
rect 15384 14569 15393 14603
rect 15393 14569 15427 14603
rect 15427 14569 15436 14603
rect 15384 14560 15436 14569
rect 15476 14560 15528 14612
rect 19524 14560 19576 14612
rect 24492 14603 24544 14612
rect 19064 14492 19116 14544
rect 19248 14492 19300 14544
rect 19616 14492 19668 14544
rect 20352 14535 20404 14544
rect 20352 14501 20361 14535
rect 20361 14501 20395 14535
rect 20395 14501 20404 14535
rect 20352 14492 20404 14501
rect 20444 14535 20496 14544
rect 20444 14501 20453 14535
rect 20453 14501 20487 14535
rect 20487 14501 20496 14535
rect 20444 14492 20496 14501
rect 20628 14492 20680 14544
rect 20720 14492 20772 14544
rect 20076 14424 20128 14476
rect 20812 14424 20864 14476
rect 21272 14492 21324 14544
rect 22836 14492 22888 14544
rect 24492 14569 24501 14603
rect 24501 14569 24535 14603
rect 24535 14569 24544 14603
rect 24492 14560 24544 14569
rect 25136 14560 25188 14612
rect 29644 14560 29696 14612
rect 32588 14560 32640 14612
rect 33876 14560 33928 14612
rect 25044 14492 25096 14544
rect 26424 14492 26476 14544
rect 26884 14492 26936 14544
rect 27344 14492 27396 14544
rect 29828 14492 29880 14544
rect 10600 14263 10652 14272
rect 10600 14229 10609 14263
rect 10609 14229 10643 14263
rect 10643 14229 10652 14263
rect 10600 14220 10652 14229
rect 19524 14356 19576 14408
rect 19984 14356 20036 14408
rect 20168 14356 20220 14408
rect 18328 14288 18380 14340
rect 20352 14288 20404 14340
rect 20536 14399 20588 14408
rect 20536 14365 20544 14399
rect 20544 14365 20578 14399
rect 20578 14365 20588 14399
rect 20536 14356 20588 14365
rect 20904 14356 20956 14408
rect 21548 14424 21600 14476
rect 21824 14424 21876 14476
rect 22284 14467 22336 14476
rect 22284 14433 22293 14467
rect 22293 14433 22327 14467
rect 22327 14433 22336 14467
rect 22284 14424 22336 14433
rect 21272 14399 21324 14408
rect 21272 14365 21301 14399
rect 21301 14365 21324 14399
rect 21272 14356 21324 14365
rect 21364 14356 21416 14408
rect 21916 14288 21968 14340
rect 22100 14356 22152 14408
rect 23204 14356 23256 14408
rect 23388 14356 23440 14408
rect 24584 14399 24636 14408
rect 24584 14365 24593 14399
rect 24593 14365 24627 14399
rect 24627 14365 24636 14399
rect 24584 14356 24636 14365
rect 22468 14288 22520 14340
rect 23296 14288 23348 14340
rect 25320 14288 25372 14340
rect 25964 14288 26016 14340
rect 12624 14220 12676 14272
rect 13728 14220 13780 14272
rect 14924 14220 14976 14272
rect 16396 14263 16448 14272
rect 16396 14229 16405 14263
rect 16405 14229 16439 14263
rect 16439 14229 16448 14263
rect 16396 14220 16448 14229
rect 19064 14220 19116 14272
rect 19340 14220 19392 14272
rect 20720 14220 20772 14272
rect 21548 14263 21600 14272
rect 21548 14229 21557 14263
rect 21557 14229 21591 14263
rect 21591 14229 21600 14263
rect 21548 14220 21600 14229
rect 22100 14220 22152 14272
rect 24216 14220 24268 14272
rect 24492 14220 24544 14272
rect 28264 14288 28316 14340
rect 28632 14288 28684 14340
rect 30748 14424 30800 14476
rect 31116 14424 31168 14476
rect 31760 14492 31812 14544
rect 34520 14492 34572 14544
rect 36452 14535 36504 14544
rect 36452 14501 36461 14535
rect 36461 14501 36495 14535
rect 36495 14501 36504 14535
rect 36452 14492 36504 14501
rect 37924 14492 37976 14544
rect 40224 14560 40276 14612
rect 40592 14560 40644 14612
rect 40868 14560 40920 14612
rect 41052 14603 41104 14612
rect 41052 14569 41061 14603
rect 41061 14569 41095 14603
rect 41095 14569 41104 14603
rect 41052 14560 41104 14569
rect 41328 14560 41380 14612
rect 41512 14560 41564 14612
rect 36360 14424 36412 14476
rect 38568 14424 38620 14476
rect 39396 14424 39448 14476
rect 40132 14492 40184 14544
rect 40960 14492 41012 14544
rect 42984 14492 43036 14544
rect 44364 14560 44416 14612
rect 45192 14560 45244 14612
rect 46204 14492 46256 14544
rect 29552 14399 29604 14408
rect 29552 14365 29561 14399
rect 29561 14365 29595 14399
rect 29595 14365 29604 14399
rect 29552 14356 29604 14365
rect 29920 14356 29972 14408
rect 30656 14356 30708 14408
rect 33140 14356 33192 14408
rect 33968 14399 34020 14408
rect 33968 14365 33977 14399
rect 33977 14365 34011 14399
rect 34011 14365 34020 14399
rect 33968 14356 34020 14365
rect 34520 14356 34572 14408
rect 36084 14356 36136 14408
rect 36820 14356 36872 14408
rect 37096 14356 37148 14408
rect 37648 14356 37700 14408
rect 34152 14288 34204 14340
rect 34980 14331 35032 14340
rect 34980 14297 34989 14331
rect 34989 14297 35023 14331
rect 35023 14297 35032 14331
rect 34980 14288 35032 14297
rect 27160 14220 27212 14272
rect 30380 14220 30432 14272
rect 30656 14220 30708 14272
rect 32404 14220 32456 14272
rect 33784 14220 33836 14272
rect 37372 14288 37424 14340
rect 38200 14356 38252 14408
rect 37924 14288 37976 14340
rect 38108 14331 38160 14340
rect 38108 14297 38117 14331
rect 38117 14297 38151 14331
rect 38151 14297 38160 14331
rect 38108 14288 38160 14297
rect 38752 14288 38804 14340
rect 39764 14356 39816 14408
rect 40868 14424 40920 14476
rect 40408 14356 40460 14408
rect 40960 14399 41012 14408
rect 40960 14365 40969 14399
rect 40969 14365 41003 14399
rect 41003 14365 41012 14399
rect 40960 14356 41012 14365
rect 41696 14399 41748 14408
rect 41696 14365 41705 14399
rect 41705 14365 41739 14399
rect 41739 14365 41748 14399
rect 41696 14356 41748 14365
rect 42248 14399 42300 14408
rect 42248 14365 42257 14399
rect 42257 14365 42291 14399
rect 42291 14365 42300 14399
rect 42248 14356 42300 14365
rect 40776 14288 40828 14340
rect 46572 14356 46624 14408
rect 41512 14220 41564 14272
rect 44640 14288 44692 14340
rect 48136 14288 48188 14340
rect 42340 14263 42392 14272
rect 42340 14229 42349 14263
rect 42349 14229 42383 14263
rect 42383 14229 42392 14263
rect 42340 14220 42392 14229
rect 45560 14263 45612 14272
rect 45560 14229 45569 14263
rect 45569 14229 45603 14263
rect 45603 14229 45612 14263
rect 45560 14220 45612 14229
rect 45928 14220 45980 14272
rect 48320 14424 48372 14476
rect 20214 14118 20266 14170
rect 20278 14118 20330 14170
rect 20342 14118 20394 14170
rect 20406 14118 20458 14170
rect 20470 14118 20522 14170
rect 39478 14118 39530 14170
rect 39542 14118 39594 14170
rect 39606 14118 39658 14170
rect 39670 14118 39722 14170
rect 39734 14118 39786 14170
rect 14464 14016 14516 14068
rect 15108 14016 15160 14068
rect 16488 14016 16540 14068
rect 16672 14016 16724 14068
rect 17776 14059 17828 14068
rect 17776 14025 17785 14059
rect 17785 14025 17819 14059
rect 17819 14025 17828 14059
rect 17776 14016 17828 14025
rect 18328 14059 18380 14068
rect 18328 14025 18337 14059
rect 18337 14025 18371 14059
rect 18371 14025 18380 14059
rect 18328 14016 18380 14025
rect 19616 14016 19668 14068
rect 20996 14016 21048 14068
rect 16396 13948 16448 14000
rect 17960 13948 18012 14000
rect 21180 13948 21232 14000
rect 10600 13880 10652 13932
rect 13728 13880 13780 13932
rect 13636 13812 13688 13864
rect 14740 13812 14792 13864
rect 19984 13880 20036 13932
rect 20536 13923 20588 13932
rect 20536 13889 20545 13923
rect 20545 13889 20579 13923
rect 20579 13889 20588 13923
rect 20536 13880 20588 13889
rect 20996 13923 21048 13932
rect 20996 13889 21005 13923
rect 21005 13889 21039 13923
rect 21039 13889 21048 13923
rect 20996 13880 21048 13889
rect 20444 13855 20496 13864
rect 20444 13821 20453 13855
rect 20453 13821 20487 13855
rect 20487 13821 20496 13855
rect 20444 13812 20496 13821
rect 20812 13812 20864 13864
rect 24492 14016 24544 14068
rect 24584 14016 24636 14068
rect 22192 13923 22244 13932
rect 22192 13889 22201 13923
rect 22201 13889 22235 13923
rect 22235 13889 22244 13923
rect 22836 13923 22888 13932
rect 22192 13880 22244 13889
rect 22836 13889 22845 13923
rect 22845 13889 22879 13923
rect 22879 13889 22888 13923
rect 22836 13880 22888 13889
rect 23020 13880 23072 13932
rect 23848 13923 23900 13932
rect 21548 13744 21600 13796
rect 22008 13744 22060 13796
rect 22376 13812 22428 13864
rect 23204 13855 23256 13864
rect 23204 13821 23213 13855
rect 23213 13821 23247 13855
rect 23247 13821 23256 13855
rect 23204 13812 23256 13821
rect 23848 13889 23857 13923
rect 23857 13889 23891 13923
rect 23891 13889 23900 13923
rect 23848 13880 23900 13889
rect 23940 13923 23992 13932
rect 23940 13889 23949 13923
rect 23949 13889 23983 13923
rect 23983 13889 23992 13923
rect 24124 13923 24176 13932
rect 23940 13880 23992 13889
rect 24124 13889 24133 13923
rect 24133 13889 24167 13923
rect 24167 13889 24176 13923
rect 24124 13880 24176 13889
rect 24216 13923 24268 13932
rect 24216 13889 24225 13923
rect 24225 13889 24259 13923
rect 24259 13889 24268 13923
rect 24216 13880 24268 13889
rect 25228 13948 25280 14000
rect 25964 14016 26016 14068
rect 27896 14016 27948 14068
rect 28540 14016 28592 14068
rect 29644 14059 29696 14068
rect 27344 13948 27396 14000
rect 26792 13880 26844 13932
rect 27160 13880 27212 13932
rect 29644 14025 29653 14059
rect 29653 14025 29687 14059
rect 29687 14025 29696 14059
rect 29644 14016 29696 14025
rect 36636 14016 36688 14068
rect 36912 14016 36964 14068
rect 39212 14016 39264 14068
rect 40132 14016 40184 14068
rect 42984 14059 43036 14068
rect 42984 14025 42993 14059
rect 42993 14025 43027 14059
rect 43027 14025 43036 14059
rect 42984 14016 43036 14025
rect 44272 14016 44324 14068
rect 44456 14016 44508 14068
rect 45284 14016 45336 14068
rect 29184 13948 29236 14000
rect 31484 13948 31536 14000
rect 32864 13948 32916 14000
rect 26424 13855 26476 13864
rect 22468 13744 22520 13796
rect 24584 13744 24636 13796
rect 26424 13821 26433 13855
rect 26433 13821 26467 13855
rect 26467 13821 26476 13855
rect 26424 13812 26476 13821
rect 29644 13812 29696 13864
rect 29828 13812 29880 13864
rect 29920 13812 29972 13864
rect 30564 13812 30616 13864
rect 31668 13880 31720 13932
rect 31852 13812 31904 13864
rect 33600 13812 33652 13864
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 17592 13676 17644 13728
rect 20904 13676 20956 13728
rect 21272 13676 21324 13728
rect 22376 13676 22428 13728
rect 22744 13676 22796 13728
rect 26056 13676 26108 13728
rect 30748 13676 30800 13728
rect 30932 13676 30984 13728
rect 31944 13676 31996 13728
rect 32036 13676 32088 13728
rect 32956 13676 33008 13728
rect 35072 13948 35124 14000
rect 34152 13880 34204 13932
rect 35348 13812 35400 13864
rect 38660 13948 38712 14000
rect 36544 13923 36596 13932
rect 36544 13889 36553 13923
rect 36553 13889 36587 13923
rect 36587 13889 36596 13923
rect 36544 13880 36596 13889
rect 37096 13880 37148 13932
rect 37924 13880 37976 13932
rect 36268 13812 36320 13864
rect 36820 13812 36872 13864
rect 39120 13880 39172 13932
rect 39488 13880 39540 13932
rect 39212 13855 39264 13864
rect 39212 13821 39221 13855
rect 39221 13821 39255 13855
rect 39255 13821 39264 13855
rect 39212 13812 39264 13821
rect 39396 13812 39448 13864
rect 41420 13948 41472 14000
rect 41512 13948 41564 14000
rect 40132 13880 40184 13932
rect 40776 13923 40828 13932
rect 40776 13889 40785 13923
rect 40785 13889 40819 13923
rect 40819 13889 40828 13923
rect 40776 13880 40828 13889
rect 41144 13880 41196 13932
rect 42800 13948 42852 14000
rect 45744 13948 45796 14000
rect 46480 13948 46532 14000
rect 35992 13744 36044 13796
rect 36452 13744 36504 13796
rect 36728 13744 36780 13796
rect 40224 13744 40276 13796
rect 40776 13744 40828 13796
rect 37648 13676 37700 13728
rect 38108 13676 38160 13728
rect 39212 13676 39264 13728
rect 39580 13676 39632 13728
rect 40132 13719 40184 13728
rect 40132 13685 40141 13719
rect 40141 13685 40175 13719
rect 40175 13685 40184 13719
rect 42708 13880 42760 13932
rect 44180 13880 44232 13932
rect 41512 13855 41564 13864
rect 41512 13821 41521 13855
rect 41521 13821 41555 13855
rect 41555 13821 41564 13855
rect 41512 13812 41564 13821
rect 41696 13812 41748 13864
rect 43536 13812 43588 13864
rect 43812 13812 43864 13864
rect 45008 13744 45060 13796
rect 40132 13676 40184 13685
rect 41696 13676 41748 13728
rect 41972 13676 42024 13728
rect 42524 13719 42576 13728
rect 42524 13685 42533 13719
rect 42533 13685 42567 13719
rect 42567 13685 42576 13719
rect 42524 13676 42576 13685
rect 45560 13676 45612 13728
rect 10582 13574 10634 13626
rect 10646 13574 10698 13626
rect 10710 13574 10762 13626
rect 10774 13574 10826 13626
rect 10838 13574 10890 13626
rect 29846 13574 29898 13626
rect 29910 13574 29962 13626
rect 29974 13574 30026 13626
rect 30038 13574 30090 13626
rect 30102 13574 30154 13626
rect 49110 13574 49162 13626
rect 49174 13574 49226 13626
rect 49238 13574 49290 13626
rect 49302 13574 49354 13626
rect 49366 13574 49418 13626
rect 14188 13472 14240 13524
rect 16764 13472 16816 13524
rect 19340 13472 19392 13524
rect 20076 13472 20128 13524
rect 22008 13472 22060 13524
rect 22192 13472 22244 13524
rect 25596 13472 25648 13524
rect 27344 13472 27396 13524
rect 12164 13404 12216 13456
rect 17132 13447 17184 13456
rect 17132 13413 17141 13447
rect 17141 13413 17175 13447
rect 17175 13413 17184 13447
rect 17132 13404 17184 13413
rect 21732 13404 21784 13456
rect 24676 13404 24728 13456
rect 28080 13472 28132 13524
rect 28356 13472 28408 13524
rect 30196 13472 30248 13524
rect 31208 13472 31260 13524
rect 19156 13336 19208 13388
rect 18052 13268 18104 13320
rect 20812 13268 20864 13320
rect 21364 13311 21416 13320
rect 21364 13277 21373 13311
rect 21373 13277 21407 13311
rect 21407 13277 21416 13311
rect 21364 13268 21416 13277
rect 22008 13336 22060 13388
rect 23572 13379 23624 13388
rect 23572 13345 23581 13379
rect 23581 13345 23615 13379
rect 23615 13345 23624 13379
rect 23572 13336 23624 13345
rect 25780 13336 25832 13388
rect 29276 13404 29328 13456
rect 29552 13404 29604 13456
rect 31116 13404 31168 13456
rect 32036 13472 32088 13524
rect 28264 13336 28316 13388
rect 33508 13472 33560 13524
rect 33784 13515 33836 13524
rect 33784 13481 33793 13515
rect 33793 13481 33827 13515
rect 33827 13481 33836 13515
rect 33784 13472 33836 13481
rect 22192 13268 22244 13320
rect 23848 13311 23900 13320
rect 23848 13277 23857 13311
rect 23857 13277 23891 13311
rect 23891 13277 23900 13311
rect 23848 13268 23900 13277
rect 24768 13268 24820 13320
rect 18328 13200 18380 13252
rect 19616 13200 19668 13252
rect 11336 13175 11388 13184
rect 11336 13141 11345 13175
rect 11345 13141 11379 13175
rect 11379 13141 11388 13175
rect 11336 13132 11388 13141
rect 18420 13132 18472 13184
rect 20996 13200 21048 13252
rect 23020 13200 23072 13252
rect 24952 13200 25004 13252
rect 26148 13268 26200 13320
rect 26976 13268 27028 13320
rect 29000 13311 29052 13320
rect 29000 13277 29009 13311
rect 29009 13277 29043 13311
rect 29043 13277 29052 13311
rect 29828 13311 29880 13320
rect 29000 13268 29052 13277
rect 29828 13277 29837 13311
rect 29837 13277 29871 13311
rect 29871 13277 29880 13311
rect 29828 13268 29880 13277
rect 31208 13268 31260 13320
rect 26240 13200 26292 13252
rect 28172 13200 28224 13252
rect 28724 13243 28776 13252
rect 28724 13209 28733 13243
rect 28733 13209 28767 13243
rect 28767 13209 28776 13243
rect 28724 13200 28776 13209
rect 41236 13515 41288 13524
rect 41236 13481 41245 13515
rect 41245 13481 41279 13515
rect 41279 13481 41288 13515
rect 41236 13472 41288 13481
rect 42616 13472 42668 13524
rect 43536 13472 43588 13524
rect 38016 13447 38068 13456
rect 38016 13413 38025 13447
rect 38025 13413 38059 13447
rect 38059 13413 38068 13447
rect 38016 13404 38068 13413
rect 38476 13404 38528 13456
rect 46112 13472 46164 13524
rect 46480 13472 46532 13524
rect 45560 13447 45612 13456
rect 31852 13268 31904 13320
rect 34060 13268 34112 13320
rect 21272 13132 21324 13184
rect 21916 13132 21968 13184
rect 24124 13132 24176 13184
rect 25136 13175 25188 13184
rect 25136 13141 25145 13175
rect 25145 13141 25179 13175
rect 25179 13141 25188 13175
rect 25136 13132 25188 13141
rect 25964 13132 26016 13184
rect 34244 13200 34296 13252
rect 35164 13268 35216 13320
rect 36268 13336 36320 13388
rect 38108 13336 38160 13388
rect 38292 13379 38344 13388
rect 38292 13345 38301 13379
rect 38301 13345 38335 13379
rect 38335 13345 38344 13379
rect 38292 13336 38344 13345
rect 38660 13336 38712 13388
rect 45560 13413 45569 13447
rect 45569 13413 45603 13447
rect 45603 13413 45612 13447
rect 45560 13404 45612 13413
rect 35716 13268 35768 13320
rect 35808 13268 35860 13320
rect 37096 13268 37148 13320
rect 37372 13268 37424 13320
rect 37924 13268 37976 13320
rect 38384 13311 38436 13320
rect 38384 13277 38393 13311
rect 38393 13277 38427 13311
rect 38427 13277 38436 13311
rect 38384 13268 38436 13277
rect 40040 13311 40092 13320
rect 40040 13277 40049 13311
rect 40049 13277 40083 13311
rect 40083 13277 40092 13311
rect 40040 13268 40092 13277
rect 42800 13336 42852 13388
rect 46204 13336 46256 13388
rect 41604 13268 41656 13320
rect 43352 13311 43404 13320
rect 43352 13277 43361 13311
rect 43361 13277 43395 13311
rect 43395 13277 43404 13311
rect 43352 13268 43404 13277
rect 58164 13311 58216 13320
rect 58164 13277 58173 13311
rect 58173 13277 58207 13311
rect 58207 13277 58216 13311
rect 58164 13268 58216 13277
rect 35440 13200 35492 13252
rect 37648 13200 37700 13252
rect 38844 13200 38896 13252
rect 38936 13132 38988 13184
rect 39120 13175 39172 13184
rect 39120 13141 39129 13175
rect 39129 13141 39163 13175
rect 39163 13141 39172 13175
rect 39120 13132 39172 13141
rect 39488 13200 39540 13252
rect 41236 13200 41288 13252
rect 41328 13200 41380 13252
rect 57888 13243 57940 13252
rect 57888 13209 57897 13243
rect 57897 13209 57931 13243
rect 57931 13209 57940 13243
rect 57888 13200 57940 13209
rect 40224 13132 40276 13184
rect 41420 13132 41472 13184
rect 41604 13132 41656 13184
rect 42892 13132 42944 13184
rect 20214 13030 20266 13082
rect 20278 13030 20330 13082
rect 20342 13030 20394 13082
rect 20406 13030 20458 13082
rect 20470 13030 20522 13082
rect 39478 13030 39530 13082
rect 39542 13030 39594 13082
rect 39606 13030 39658 13082
rect 39670 13030 39722 13082
rect 39734 13030 39786 13082
rect 18512 12971 18564 12980
rect 18512 12937 18521 12971
rect 18521 12937 18555 12971
rect 18555 12937 18564 12971
rect 18512 12928 18564 12937
rect 20076 12971 20128 12980
rect 20076 12937 20085 12971
rect 20085 12937 20119 12971
rect 20119 12937 20128 12971
rect 20076 12928 20128 12937
rect 21916 12928 21968 12980
rect 22652 12928 22704 12980
rect 17960 12903 18012 12912
rect 17960 12869 17969 12903
rect 17969 12869 18003 12903
rect 18003 12869 18012 12903
rect 17960 12860 18012 12869
rect 19248 12860 19300 12912
rect 18420 12792 18472 12844
rect 19708 12860 19760 12912
rect 21824 12860 21876 12912
rect 22192 12860 22244 12912
rect 24584 12928 24636 12980
rect 24768 12928 24820 12980
rect 26424 12971 26476 12980
rect 20720 12835 20772 12844
rect 20720 12801 20729 12835
rect 20729 12801 20763 12835
rect 20763 12801 20772 12835
rect 20720 12792 20772 12801
rect 22284 12792 22336 12844
rect 22836 12792 22888 12844
rect 23480 12792 23532 12844
rect 24124 12792 24176 12844
rect 15476 12724 15528 12776
rect 23388 12724 23440 12776
rect 23756 12767 23808 12776
rect 23756 12733 23765 12767
rect 23765 12733 23799 12767
rect 23799 12733 23808 12767
rect 23756 12724 23808 12733
rect 24952 12767 25004 12776
rect 24952 12733 24961 12767
rect 24961 12733 24995 12767
rect 24995 12733 25004 12767
rect 24952 12724 25004 12733
rect 21640 12656 21692 12708
rect 25412 12860 25464 12912
rect 25228 12792 25280 12844
rect 26424 12937 26433 12971
rect 26433 12937 26467 12971
rect 26467 12937 26476 12971
rect 26424 12928 26476 12937
rect 26976 12928 27028 12980
rect 27344 12928 27396 12980
rect 27804 12928 27856 12980
rect 29092 12971 29144 12980
rect 29092 12937 29101 12971
rect 29101 12937 29135 12971
rect 29135 12937 29144 12971
rect 29092 12928 29144 12937
rect 31116 12928 31168 12980
rect 31300 12971 31352 12980
rect 31300 12937 31309 12971
rect 31309 12937 31343 12971
rect 31343 12937 31352 12971
rect 31300 12928 31352 12937
rect 36176 12928 36228 12980
rect 32404 12903 32456 12912
rect 32404 12869 32413 12903
rect 32413 12869 32447 12903
rect 32447 12869 32456 12903
rect 32404 12860 32456 12869
rect 34428 12860 34480 12912
rect 31208 12792 31260 12844
rect 31668 12792 31720 12844
rect 27344 12767 27396 12776
rect 12992 12588 13044 12640
rect 20076 12588 20128 12640
rect 23020 12588 23072 12640
rect 23204 12631 23256 12640
rect 23204 12597 23213 12631
rect 23213 12597 23247 12631
rect 23247 12597 23256 12631
rect 23204 12588 23256 12597
rect 23664 12588 23716 12640
rect 24032 12588 24084 12640
rect 24308 12588 24360 12640
rect 24584 12588 24636 12640
rect 25412 12656 25464 12708
rect 25964 12699 26016 12708
rect 24860 12588 24912 12640
rect 25228 12588 25280 12640
rect 25320 12588 25372 12640
rect 25964 12665 25973 12699
rect 25973 12665 26007 12699
rect 26007 12665 26016 12699
rect 25964 12656 26016 12665
rect 25596 12588 25648 12640
rect 27344 12733 27353 12767
rect 27353 12733 27387 12767
rect 27387 12733 27396 12767
rect 27344 12724 27396 12733
rect 28908 12724 28960 12776
rect 29552 12767 29604 12776
rect 29552 12733 29561 12767
rect 29561 12733 29595 12767
rect 29595 12733 29604 12767
rect 29552 12724 29604 12733
rect 29092 12656 29144 12708
rect 30288 12724 30340 12776
rect 33600 12724 33652 12776
rect 34152 12792 34204 12844
rect 35164 12792 35216 12844
rect 35256 12835 35308 12844
rect 35256 12801 35265 12835
rect 35265 12801 35299 12835
rect 35299 12801 35308 12835
rect 35256 12792 35308 12801
rect 35716 12792 35768 12844
rect 36268 12835 36320 12844
rect 36268 12801 36277 12835
rect 36277 12801 36311 12835
rect 36311 12801 36320 12835
rect 36268 12792 36320 12801
rect 36912 12928 36964 12980
rect 37280 12971 37332 12980
rect 37280 12937 37289 12971
rect 37289 12937 37323 12971
rect 37323 12937 37332 12971
rect 37280 12928 37332 12937
rect 38476 12971 38528 12980
rect 38476 12937 38485 12971
rect 38485 12937 38519 12971
rect 38519 12937 38528 12971
rect 38476 12928 38528 12937
rect 39304 12928 39356 12980
rect 39856 12928 39908 12980
rect 41420 12928 41472 12980
rect 42340 12928 42392 12980
rect 42432 12928 42484 12980
rect 44732 12928 44784 12980
rect 58164 12971 58216 12980
rect 58164 12937 58173 12971
rect 58173 12937 58207 12971
rect 58207 12937 58216 12971
rect 58164 12928 58216 12937
rect 36728 12860 36780 12912
rect 40040 12860 40092 12912
rect 41328 12860 41380 12912
rect 34060 12724 34112 12776
rect 35808 12724 35860 12776
rect 37004 12792 37056 12844
rect 38016 12792 38068 12844
rect 38568 12835 38620 12844
rect 38568 12801 38577 12835
rect 38577 12801 38611 12835
rect 38611 12801 38620 12835
rect 38568 12792 38620 12801
rect 38936 12792 38988 12844
rect 39212 12792 39264 12844
rect 33692 12656 33744 12708
rect 32220 12588 32272 12640
rect 33416 12588 33468 12640
rect 34060 12588 34112 12640
rect 35256 12656 35308 12708
rect 36728 12724 36780 12776
rect 37464 12724 37516 12776
rect 38844 12724 38896 12776
rect 40408 12792 40460 12844
rect 42524 12792 42576 12844
rect 43720 12724 43772 12776
rect 35992 12656 36044 12708
rect 35440 12631 35492 12640
rect 35440 12597 35449 12631
rect 35449 12597 35483 12631
rect 35483 12597 35492 12631
rect 35440 12588 35492 12597
rect 35900 12588 35952 12640
rect 37096 12588 37148 12640
rect 37280 12656 37332 12708
rect 38936 12656 38988 12708
rect 39488 12656 39540 12708
rect 40868 12656 40920 12708
rect 41236 12656 41288 12708
rect 42432 12656 42484 12708
rect 44364 12656 44416 12708
rect 57888 12656 57940 12708
rect 44640 12631 44692 12640
rect 44640 12597 44649 12631
rect 44649 12597 44683 12631
rect 44683 12597 44692 12631
rect 44640 12588 44692 12597
rect 45192 12631 45244 12640
rect 45192 12597 45201 12631
rect 45201 12597 45235 12631
rect 45235 12597 45244 12631
rect 45192 12588 45244 12597
rect 10582 12486 10634 12538
rect 10646 12486 10698 12538
rect 10710 12486 10762 12538
rect 10774 12486 10826 12538
rect 10838 12486 10890 12538
rect 29846 12486 29898 12538
rect 29910 12486 29962 12538
rect 29974 12486 30026 12538
rect 30038 12486 30090 12538
rect 30102 12486 30154 12538
rect 49110 12486 49162 12538
rect 49174 12486 49226 12538
rect 49238 12486 49290 12538
rect 49302 12486 49354 12538
rect 49366 12486 49418 12538
rect 12900 12427 12952 12436
rect 12900 12393 12909 12427
rect 12909 12393 12943 12427
rect 12943 12393 12952 12427
rect 12900 12384 12952 12393
rect 18696 12427 18748 12436
rect 18696 12393 18705 12427
rect 18705 12393 18739 12427
rect 18739 12393 18748 12427
rect 18696 12384 18748 12393
rect 19708 12427 19760 12436
rect 19708 12393 19717 12427
rect 19717 12393 19751 12427
rect 19751 12393 19760 12427
rect 19708 12384 19760 12393
rect 20904 12427 20956 12436
rect 20904 12393 20913 12427
rect 20913 12393 20947 12427
rect 20947 12393 20956 12427
rect 20904 12384 20956 12393
rect 21548 12384 21600 12436
rect 21916 12427 21968 12436
rect 21916 12393 21925 12427
rect 21925 12393 21959 12427
rect 21959 12393 21968 12427
rect 21916 12384 21968 12393
rect 24584 12384 24636 12436
rect 25136 12384 25188 12436
rect 25596 12384 25648 12436
rect 22100 12316 22152 12368
rect 22376 12359 22428 12368
rect 22376 12325 22385 12359
rect 22385 12325 22419 12359
rect 22419 12325 22428 12359
rect 24768 12359 24820 12368
rect 22376 12316 22428 12325
rect 19432 12248 19484 12300
rect 24216 12248 24268 12300
rect 11336 12180 11388 12232
rect 12900 12180 12952 12232
rect 21824 12180 21876 12232
rect 23572 12223 23624 12232
rect 16304 12112 16356 12164
rect 23572 12189 23581 12223
rect 23581 12189 23615 12223
rect 23615 12189 23624 12223
rect 23572 12180 23624 12189
rect 24768 12325 24777 12359
rect 24777 12325 24811 12359
rect 24811 12325 24820 12359
rect 24768 12316 24820 12325
rect 24952 12316 25004 12368
rect 25872 12384 25924 12436
rect 26792 12427 26844 12436
rect 26792 12393 26801 12427
rect 26801 12393 26835 12427
rect 26835 12393 26844 12427
rect 26792 12384 26844 12393
rect 24676 12248 24728 12300
rect 25228 12248 25280 12300
rect 26056 12316 26108 12368
rect 26424 12316 26476 12368
rect 29368 12384 29420 12436
rect 32404 12384 32456 12436
rect 36268 12427 36320 12436
rect 31116 12316 31168 12368
rect 31300 12316 31352 12368
rect 31484 12359 31536 12368
rect 31484 12325 31493 12359
rect 31493 12325 31527 12359
rect 31527 12325 31536 12359
rect 31484 12316 31536 12325
rect 33600 12316 33652 12368
rect 33876 12316 33928 12368
rect 35624 12316 35676 12368
rect 36268 12393 36277 12427
rect 36277 12393 36311 12427
rect 36311 12393 36320 12427
rect 36268 12384 36320 12393
rect 36820 12384 36872 12436
rect 37096 12384 37148 12436
rect 25964 12248 26016 12300
rect 26332 12291 26384 12300
rect 26332 12257 26341 12291
rect 26341 12257 26375 12291
rect 26375 12257 26384 12291
rect 26332 12248 26384 12257
rect 26792 12248 26844 12300
rect 27896 12248 27948 12300
rect 29368 12248 29420 12300
rect 1492 12087 1544 12096
rect 1492 12053 1501 12087
rect 1501 12053 1535 12087
rect 1535 12053 1544 12087
rect 1492 12044 1544 12053
rect 11060 12044 11112 12096
rect 18144 12087 18196 12096
rect 18144 12053 18153 12087
rect 18153 12053 18187 12087
rect 18187 12053 18196 12087
rect 18144 12044 18196 12053
rect 23480 12112 23532 12164
rect 24584 12112 24636 12164
rect 25872 12180 25924 12232
rect 26792 12112 26844 12164
rect 25964 12044 26016 12096
rect 27160 12180 27212 12232
rect 29552 12180 29604 12232
rect 31668 12248 31720 12300
rect 37004 12316 37056 12368
rect 31944 12223 31996 12232
rect 31944 12189 31953 12223
rect 31953 12189 31987 12223
rect 31987 12189 31996 12223
rect 31944 12180 31996 12189
rect 33968 12180 34020 12232
rect 34244 12180 34296 12232
rect 35256 12180 35308 12232
rect 35532 12180 35584 12232
rect 27528 12155 27580 12164
rect 27528 12121 27537 12155
rect 27537 12121 27571 12155
rect 27571 12121 27580 12155
rect 27528 12112 27580 12121
rect 28264 12112 28316 12164
rect 29092 12112 29144 12164
rect 31668 12112 31720 12164
rect 32312 12112 32364 12164
rect 30196 12044 30248 12096
rect 32680 12112 32732 12164
rect 36084 12112 36136 12164
rect 37556 12316 37608 12368
rect 38752 12384 38804 12436
rect 40592 12384 40644 12436
rect 45928 12384 45980 12436
rect 39948 12316 40000 12368
rect 40408 12359 40460 12368
rect 40408 12325 40417 12359
rect 40417 12325 40451 12359
rect 40451 12325 40460 12359
rect 40408 12316 40460 12325
rect 43536 12316 43588 12368
rect 38016 12248 38068 12300
rect 38108 12180 38160 12232
rect 38660 12223 38712 12232
rect 38660 12189 38669 12223
rect 38669 12189 38703 12223
rect 38703 12189 38712 12223
rect 38660 12180 38712 12189
rect 39856 12180 39908 12232
rect 38016 12112 38068 12164
rect 33048 12044 33100 12096
rect 35624 12044 35676 12096
rect 36636 12044 36688 12096
rect 37556 12044 37608 12096
rect 38752 12044 38804 12096
rect 38936 12044 38988 12096
rect 40868 12044 40920 12096
rect 42064 12087 42116 12096
rect 42064 12053 42073 12087
rect 42073 12053 42107 12087
rect 42107 12053 42116 12087
rect 42064 12044 42116 12053
rect 43720 12087 43772 12096
rect 43720 12053 43729 12087
rect 43729 12053 43763 12087
rect 43763 12053 43772 12087
rect 43720 12044 43772 12053
rect 44364 12087 44416 12096
rect 44364 12053 44373 12087
rect 44373 12053 44407 12087
rect 44407 12053 44416 12087
rect 44364 12044 44416 12053
rect 45560 12044 45612 12096
rect 46112 12044 46164 12096
rect 20214 11942 20266 11994
rect 20278 11942 20330 11994
rect 20342 11942 20394 11994
rect 20406 11942 20458 11994
rect 20470 11942 20522 11994
rect 39478 11942 39530 11994
rect 39542 11942 39594 11994
rect 39606 11942 39658 11994
rect 39670 11942 39722 11994
rect 39734 11942 39786 11994
rect 15752 11840 15804 11892
rect 16304 11840 16356 11892
rect 22192 11840 22244 11892
rect 22468 11840 22520 11892
rect 23480 11840 23532 11892
rect 22008 11772 22060 11824
rect 23664 11815 23716 11824
rect 23664 11781 23673 11815
rect 23673 11781 23707 11815
rect 23707 11781 23716 11815
rect 23664 11772 23716 11781
rect 20996 11704 21048 11756
rect 22376 11704 22428 11756
rect 22744 11704 22796 11756
rect 22928 11704 22980 11756
rect 24584 11840 24636 11892
rect 26424 11840 26476 11892
rect 28724 11840 28776 11892
rect 25136 11772 25188 11824
rect 26332 11772 26384 11824
rect 26608 11772 26660 11824
rect 24216 11704 24268 11756
rect 17224 11636 17276 11688
rect 24124 11636 24176 11688
rect 19340 11568 19392 11620
rect 24584 11704 24636 11756
rect 25044 11747 25096 11756
rect 25044 11713 25053 11747
rect 25053 11713 25087 11747
rect 25087 11713 25096 11747
rect 25044 11704 25096 11713
rect 25780 11704 25832 11756
rect 26148 11704 26200 11756
rect 27896 11704 27948 11756
rect 31392 11772 31444 11824
rect 32680 11772 32732 11824
rect 32864 11772 32916 11824
rect 28264 11704 28316 11756
rect 28908 11704 28960 11756
rect 29184 11704 29236 11756
rect 24676 11636 24728 11688
rect 25136 11679 25188 11688
rect 25136 11645 25145 11679
rect 25145 11645 25179 11679
rect 25179 11645 25188 11679
rect 25136 11636 25188 11645
rect 24860 11568 24912 11620
rect 30196 11636 30248 11688
rect 31944 11704 31996 11756
rect 34060 11704 34112 11756
rect 34704 11704 34756 11756
rect 35624 11747 35676 11756
rect 35624 11713 35633 11747
rect 35633 11713 35667 11747
rect 35667 11713 35676 11747
rect 35624 11704 35676 11713
rect 35808 11704 35860 11756
rect 36176 11840 36228 11892
rect 38016 11883 38068 11892
rect 38016 11849 38025 11883
rect 38025 11849 38059 11883
rect 38059 11849 38068 11883
rect 38016 11840 38068 11849
rect 38752 11883 38804 11892
rect 38752 11849 38761 11883
rect 38761 11849 38795 11883
rect 38795 11849 38804 11883
rect 38752 11840 38804 11849
rect 39304 11883 39356 11892
rect 39304 11849 39313 11883
rect 39313 11849 39347 11883
rect 39347 11849 39356 11883
rect 39304 11840 39356 11849
rect 40316 11883 40368 11892
rect 40316 11849 40325 11883
rect 40325 11849 40359 11883
rect 40359 11849 40368 11883
rect 40316 11840 40368 11849
rect 40776 11840 40828 11892
rect 41420 11883 41472 11892
rect 41420 11849 41429 11883
rect 41429 11849 41463 11883
rect 41463 11849 41472 11883
rect 41420 11840 41472 11849
rect 42708 11840 42760 11892
rect 44364 11840 44416 11892
rect 36820 11772 36872 11824
rect 36728 11747 36780 11756
rect 26424 11611 26476 11620
rect 26424 11577 26433 11611
rect 26433 11577 26467 11611
rect 26467 11577 26476 11611
rect 26424 11568 26476 11577
rect 27896 11568 27948 11620
rect 28356 11568 28408 11620
rect 28908 11568 28960 11620
rect 34336 11679 34388 11688
rect 34336 11645 34345 11679
rect 34345 11645 34379 11679
rect 34379 11645 34388 11679
rect 35716 11679 35768 11688
rect 34336 11636 34388 11645
rect 35716 11645 35725 11679
rect 35725 11645 35759 11679
rect 35759 11645 35768 11679
rect 35716 11636 35768 11645
rect 36728 11713 36737 11747
rect 36737 11713 36771 11747
rect 36771 11713 36780 11747
rect 36728 11704 36780 11713
rect 37372 11772 37424 11824
rect 43904 11772 43956 11824
rect 38016 11636 38068 11688
rect 14740 11500 14792 11552
rect 19064 11500 19116 11552
rect 19524 11500 19576 11552
rect 20996 11543 21048 11552
rect 20996 11509 21005 11543
rect 21005 11509 21039 11543
rect 21039 11509 21048 11543
rect 20996 11500 21048 11509
rect 24216 11543 24268 11552
rect 24216 11509 24225 11543
rect 24225 11509 24259 11543
rect 24259 11509 24268 11543
rect 24216 11500 24268 11509
rect 26240 11500 26292 11552
rect 26332 11500 26384 11552
rect 28172 11500 28224 11552
rect 29276 11543 29328 11552
rect 29276 11509 29285 11543
rect 29285 11509 29319 11543
rect 29319 11509 29328 11543
rect 29276 11500 29328 11509
rect 31576 11543 31628 11552
rect 31576 11509 31585 11543
rect 31585 11509 31619 11543
rect 31619 11509 31628 11543
rect 31576 11500 31628 11509
rect 33140 11500 33192 11552
rect 33784 11500 33836 11552
rect 33968 11500 34020 11552
rect 36912 11568 36964 11620
rect 38200 11704 38252 11756
rect 38752 11704 38804 11756
rect 41052 11704 41104 11756
rect 43536 11747 43588 11756
rect 38384 11636 38436 11688
rect 42156 11636 42208 11688
rect 43536 11713 43545 11747
rect 43545 11713 43579 11747
rect 43579 11713 43588 11747
rect 43536 11704 43588 11713
rect 44640 11636 44692 11688
rect 37648 11500 37700 11552
rect 38568 11568 38620 11620
rect 38844 11568 38896 11620
rect 42616 11568 42668 11620
rect 10582 11398 10634 11450
rect 10646 11398 10698 11450
rect 10710 11398 10762 11450
rect 10774 11398 10826 11450
rect 10838 11398 10890 11450
rect 29846 11398 29898 11450
rect 29910 11398 29962 11450
rect 29974 11398 30026 11450
rect 30038 11398 30090 11450
rect 30102 11398 30154 11450
rect 49110 11398 49162 11450
rect 49174 11398 49226 11450
rect 49238 11398 49290 11450
rect 49302 11398 49354 11450
rect 49366 11398 49418 11450
rect 19064 11296 19116 11348
rect 19708 11296 19760 11348
rect 21180 11296 21232 11348
rect 21548 11339 21600 11348
rect 21548 11305 21557 11339
rect 21557 11305 21591 11339
rect 21591 11305 21600 11339
rect 21548 11296 21600 11305
rect 22836 11296 22888 11348
rect 23940 11296 23992 11348
rect 24308 11296 24360 11348
rect 25596 11339 25648 11348
rect 20444 11271 20496 11280
rect 20444 11237 20453 11271
rect 20453 11237 20487 11271
rect 20487 11237 20496 11271
rect 20444 11228 20496 11237
rect 20628 11228 20680 11280
rect 24032 11228 24084 11280
rect 25596 11305 25605 11339
rect 25605 11305 25639 11339
rect 25639 11305 25648 11339
rect 25596 11296 25648 11305
rect 25872 11296 25924 11348
rect 27344 11296 27396 11348
rect 27528 11296 27580 11348
rect 26792 11271 26844 11280
rect 23572 11160 23624 11212
rect 26332 11203 26384 11212
rect 19340 11135 19392 11144
rect 19340 11101 19349 11135
rect 19349 11101 19383 11135
rect 19383 11101 19392 11135
rect 19340 11092 19392 11101
rect 20904 11092 20956 11144
rect 24676 11092 24728 11144
rect 25044 11135 25096 11144
rect 25044 11101 25053 11135
rect 25053 11101 25087 11135
rect 25087 11101 25096 11135
rect 25044 11092 25096 11101
rect 25412 11092 25464 11144
rect 25596 11092 25648 11144
rect 22284 11024 22336 11076
rect 23020 11024 23072 11076
rect 24032 11024 24084 11076
rect 26332 11169 26341 11203
rect 26341 11169 26375 11203
rect 26375 11169 26384 11203
rect 26332 11160 26384 11169
rect 26792 11237 26801 11271
rect 26801 11237 26835 11271
rect 26835 11237 26844 11271
rect 26792 11228 26844 11237
rect 27804 11271 27856 11280
rect 27804 11237 27813 11271
rect 27813 11237 27847 11271
rect 27847 11237 27856 11271
rect 27804 11228 27856 11237
rect 27988 11160 28040 11212
rect 34796 11339 34848 11348
rect 34796 11305 34805 11339
rect 34805 11305 34839 11339
rect 34839 11305 34848 11339
rect 34796 11296 34848 11305
rect 32772 11228 32824 11280
rect 35716 11228 35768 11280
rect 36452 11296 36504 11348
rect 36728 11296 36780 11348
rect 37004 11228 37056 11280
rect 37832 11296 37884 11348
rect 38844 11339 38896 11348
rect 38844 11305 38853 11339
rect 38853 11305 38887 11339
rect 38887 11305 38896 11339
rect 38844 11296 38896 11305
rect 39856 11339 39908 11348
rect 39856 11305 39865 11339
rect 39865 11305 39899 11339
rect 39899 11305 39908 11339
rect 39856 11296 39908 11305
rect 41236 11296 41288 11348
rect 42708 11339 42760 11348
rect 42708 11305 42717 11339
rect 42717 11305 42751 11339
rect 42751 11305 42760 11339
rect 42708 11296 42760 11305
rect 30288 11203 30340 11212
rect 30288 11169 30297 11203
rect 30297 11169 30331 11203
rect 30331 11169 30340 11203
rect 30288 11160 30340 11169
rect 31392 11160 31444 11212
rect 31668 11160 31720 11212
rect 34060 11160 34112 11212
rect 34244 11160 34296 11212
rect 34796 11160 34848 11212
rect 35164 11203 35216 11212
rect 35164 11169 35173 11203
rect 35173 11169 35207 11203
rect 35207 11169 35216 11203
rect 35164 11160 35216 11169
rect 35624 11160 35676 11212
rect 36084 11160 36136 11212
rect 39396 11160 39448 11212
rect 41512 11203 41564 11212
rect 41512 11169 41521 11203
rect 41521 11169 41555 11203
rect 41555 11169 41564 11203
rect 41512 11160 41564 11169
rect 26792 11092 26844 11144
rect 27620 11092 27672 11144
rect 26148 11024 26200 11076
rect 26976 11024 27028 11076
rect 27896 11024 27948 11076
rect 28724 11135 28776 11144
rect 28724 11101 28733 11135
rect 28733 11101 28767 11135
rect 28767 11101 28776 11135
rect 28724 11092 28776 11101
rect 29276 11092 29328 11144
rect 31024 11135 31076 11144
rect 31024 11101 31033 11135
rect 31033 11101 31067 11135
rect 31067 11101 31076 11135
rect 31024 11092 31076 11101
rect 33784 11092 33836 11144
rect 33968 11092 34020 11144
rect 34704 11135 34756 11144
rect 34704 11101 34713 11135
rect 34713 11101 34747 11135
rect 34747 11101 34756 11135
rect 34704 11092 34756 11101
rect 35256 11092 35308 11144
rect 35440 11092 35492 11144
rect 35716 11092 35768 11144
rect 17040 10956 17092 11008
rect 23480 10956 23532 11008
rect 25780 10956 25832 11008
rect 30380 10956 30432 11008
rect 30564 10956 30616 11008
rect 31208 11024 31260 11076
rect 31760 11024 31812 11076
rect 31668 10956 31720 11008
rect 33140 11024 33192 11076
rect 33508 11024 33560 11076
rect 35624 11067 35676 11076
rect 35624 11033 35633 11067
rect 35633 11033 35667 11067
rect 35667 11033 35676 11067
rect 35624 11024 35676 11033
rect 33324 10956 33376 11008
rect 33968 10956 34020 11008
rect 34152 10956 34204 11008
rect 34520 10956 34572 11008
rect 34796 10956 34848 11008
rect 35716 10956 35768 11008
rect 35808 10999 35860 11008
rect 35808 10965 35833 10999
rect 35833 10965 35860 10999
rect 35992 10999 36044 11008
rect 35808 10956 35860 10965
rect 35992 10965 36001 10999
rect 36001 10965 36035 10999
rect 36035 10965 36044 10999
rect 35992 10956 36044 10965
rect 36360 11092 36412 11144
rect 36912 11024 36964 11076
rect 37832 11092 37884 11144
rect 46296 11092 46348 11144
rect 58164 11135 58216 11144
rect 58164 11101 58173 11135
rect 58173 11101 58207 11135
rect 58207 11101 58216 11135
rect 58164 11092 58216 11101
rect 37648 11024 37700 11076
rect 42524 11024 42576 11076
rect 20214 10854 20266 10906
rect 20278 10854 20330 10906
rect 20342 10854 20394 10906
rect 20406 10854 20458 10906
rect 20470 10854 20522 10906
rect 39478 10854 39530 10906
rect 39542 10854 39594 10906
rect 39606 10854 39658 10906
rect 39670 10854 39722 10906
rect 39734 10854 39786 10906
rect 19984 10752 20036 10804
rect 21180 10752 21232 10804
rect 21364 10752 21416 10804
rect 22652 10795 22704 10804
rect 22652 10761 22661 10795
rect 22661 10761 22695 10795
rect 22695 10761 22704 10795
rect 22652 10752 22704 10761
rect 23756 10795 23808 10804
rect 23756 10761 23765 10795
rect 23765 10761 23799 10795
rect 23799 10761 23808 10795
rect 23756 10752 23808 10761
rect 24768 10752 24820 10804
rect 24308 10727 24360 10736
rect 24308 10693 24317 10727
rect 24317 10693 24351 10727
rect 24351 10693 24360 10727
rect 24308 10684 24360 10693
rect 34520 10752 34572 10804
rect 36268 10795 36320 10804
rect 26792 10684 26844 10736
rect 31300 10727 31352 10736
rect 11060 10616 11112 10668
rect 23480 10616 23532 10668
rect 24216 10616 24268 10668
rect 24952 10659 25004 10668
rect 24952 10625 24961 10659
rect 24961 10625 24995 10659
rect 24995 10625 25004 10659
rect 24952 10616 25004 10625
rect 14924 10548 14976 10600
rect 23388 10548 23440 10600
rect 25780 10616 25832 10668
rect 26148 10616 26200 10668
rect 26700 10616 26752 10668
rect 25412 10591 25464 10600
rect 25412 10557 25421 10591
rect 25421 10557 25455 10591
rect 25455 10557 25464 10591
rect 25412 10548 25464 10557
rect 27252 10548 27304 10600
rect 27712 10591 27764 10600
rect 27712 10557 27721 10591
rect 27721 10557 27755 10591
rect 27755 10557 27764 10591
rect 27712 10548 27764 10557
rect 30288 10616 30340 10668
rect 31300 10693 31309 10727
rect 31309 10693 31343 10727
rect 31343 10693 31352 10727
rect 31300 10684 31352 10693
rect 31392 10684 31444 10736
rect 31484 10616 31536 10668
rect 32036 10548 32088 10600
rect 32496 10616 32548 10668
rect 33324 10727 33376 10736
rect 33324 10693 33333 10727
rect 33333 10693 33367 10727
rect 33367 10693 33376 10727
rect 33324 10684 33376 10693
rect 33692 10684 33744 10736
rect 24768 10480 24820 10532
rect 27988 10523 28040 10532
rect 27988 10489 27997 10523
rect 27997 10489 28031 10523
rect 28031 10489 28040 10523
rect 27988 10480 28040 10489
rect 28356 10480 28408 10532
rect 30380 10480 30432 10532
rect 1492 10455 1544 10464
rect 1492 10421 1501 10455
rect 1501 10421 1535 10455
rect 1535 10421 1544 10455
rect 1492 10412 1544 10421
rect 11520 10455 11572 10464
rect 11520 10421 11529 10455
rect 11529 10421 11563 10455
rect 11563 10421 11572 10455
rect 11520 10412 11572 10421
rect 20076 10412 20128 10464
rect 20628 10412 20680 10464
rect 26332 10412 26384 10464
rect 27344 10412 27396 10464
rect 29552 10412 29604 10464
rect 31944 10412 31996 10464
rect 34152 10616 34204 10668
rect 34244 10659 34296 10668
rect 34244 10625 34253 10659
rect 34253 10625 34287 10659
rect 34287 10625 34296 10659
rect 34244 10616 34296 10625
rect 34796 10616 34848 10668
rect 35164 10684 35216 10736
rect 36268 10761 36277 10795
rect 36277 10761 36311 10795
rect 36311 10761 36320 10795
rect 36268 10752 36320 10761
rect 36452 10752 36504 10804
rect 41236 10795 41288 10804
rect 41236 10761 41245 10795
rect 41245 10761 41279 10795
rect 41279 10761 41288 10795
rect 41236 10752 41288 10761
rect 41696 10752 41748 10804
rect 43536 10752 43588 10804
rect 58164 10795 58216 10804
rect 58164 10761 58173 10795
rect 58173 10761 58207 10795
rect 58207 10761 58216 10795
rect 58164 10752 58216 10761
rect 35808 10616 35860 10668
rect 36268 10616 36320 10668
rect 37004 10684 37056 10736
rect 37280 10684 37332 10736
rect 37372 10684 37424 10736
rect 38384 10727 38436 10736
rect 38384 10693 38393 10727
rect 38393 10693 38427 10727
rect 38427 10693 38436 10727
rect 38384 10684 38436 10693
rect 38568 10684 38620 10736
rect 41144 10684 41196 10736
rect 33140 10548 33192 10600
rect 33692 10480 33744 10532
rect 33784 10523 33836 10532
rect 33784 10489 33793 10523
rect 33793 10489 33827 10523
rect 33827 10489 33836 10523
rect 33784 10480 33836 10489
rect 34152 10480 34204 10532
rect 35532 10523 35584 10532
rect 35532 10489 35541 10523
rect 35541 10489 35575 10523
rect 35575 10489 35584 10523
rect 35532 10480 35584 10489
rect 33416 10412 33468 10464
rect 33968 10455 34020 10464
rect 33968 10421 33977 10455
rect 33977 10421 34011 10455
rect 34011 10421 34020 10455
rect 33968 10412 34020 10421
rect 34612 10412 34664 10464
rect 35164 10412 35216 10464
rect 35716 10412 35768 10464
rect 37280 10412 37332 10464
rect 37924 10412 37976 10464
rect 10582 10310 10634 10362
rect 10646 10310 10698 10362
rect 10710 10310 10762 10362
rect 10774 10310 10826 10362
rect 10838 10310 10890 10362
rect 29846 10310 29898 10362
rect 29910 10310 29962 10362
rect 29974 10310 30026 10362
rect 30038 10310 30090 10362
rect 30102 10310 30154 10362
rect 49110 10310 49162 10362
rect 49174 10310 49226 10362
rect 49238 10310 49290 10362
rect 49302 10310 49354 10362
rect 49366 10310 49418 10362
rect 19708 10208 19760 10260
rect 23480 10208 23532 10260
rect 23756 10251 23808 10260
rect 23756 10217 23765 10251
rect 23765 10217 23799 10251
rect 23799 10217 23808 10251
rect 23756 10208 23808 10217
rect 24584 10251 24636 10260
rect 24584 10217 24593 10251
rect 24593 10217 24627 10251
rect 24627 10217 24636 10251
rect 24584 10208 24636 10217
rect 25228 10208 25280 10260
rect 25872 10208 25924 10260
rect 26240 10251 26292 10260
rect 26240 10217 26249 10251
rect 26249 10217 26283 10251
rect 26283 10217 26292 10251
rect 26240 10208 26292 10217
rect 27436 10208 27488 10260
rect 28448 10251 28500 10260
rect 28448 10217 28457 10251
rect 28457 10217 28491 10251
rect 28491 10217 28500 10251
rect 28448 10208 28500 10217
rect 23296 10140 23348 10192
rect 24492 10140 24544 10192
rect 27712 10140 27764 10192
rect 27804 10183 27856 10192
rect 27804 10149 27813 10183
rect 27813 10149 27847 10183
rect 27847 10149 27856 10183
rect 27804 10140 27856 10149
rect 34704 10208 34756 10260
rect 35716 10208 35768 10260
rect 34152 10140 34204 10192
rect 34796 10140 34848 10192
rect 36544 10140 36596 10192
rect 38292 10208 38344 10260
rect 40040 10208 40092 10260
rect 41052 10251 41104 10260
rect 41052 10217 41061 10251
rect 41061 10217 41095 10251
rect 41095 10217 41104 10251
rect 41052 10208 41104 10217
rect 41972 10140 42024 10192
rect 19800 10072 19852 10124
rect 24400 10072 24452 10124
rect 25320 10004 25372 10056
rect 25872 10004 25924 10056
rect 26700 10004 26752 10056
rect 28080 10072 28132 10124
rect 28540 10072 28592 10124
rect 28908 10072 28960 10124
rect 29552 10072 29604 10124
rect 30012 10115 30064 10124
rect 30012 10081 30021 10115
rect 30021 10081 30055 10115
rect 30055 10081 30064 10115
rect 30012 10072 30064 10081
rect 30104 10072 30156 10124
rect 30564 10072 30616 10124
rect 31944 10115 31996 10124
rect 31944 10081 31953 10115
rect 31953 10081 31987 10115
rect 31987 10081 31996 10115
rect 31944 10072 31996 10081
rect 33324 10072 33376 10124
rect 34244 10072 34296 10124
rect 34428 10072 34480 10124
rect 27252 10004 27304 10056
rect 26792 9936 26844 9988
rect 28172 10004 28224 10056
rect 31668 10004 31720 10056
rect 27804 9936 27856 9988
rect 28448 9936 28500 9988
rect 30104 9936 30156 9988
rect 31760 9936 31812 9988
rect 32404 10004 32456 10056
rect 32680 10004 32732 10056
rect 34520 10004 34572 10056
rect 35440 10047 35492 10056
rect 35440 10013 35449 10047
rect 35449 10013 35483 10047
rect 35483 10013 35492 10047
rect 35440 10004 35492 10013
rect 35624 10047 35676 10056
rect 35624 10013 35633 10047
rect 35633 10013 35667 10047
rect 35667 10013 35676 10047
rect 35624 10004 35676 10013
rect 37648 10072 37700 10124
rect 38568 10072 38620 10124
rect 38936 10115 38988 10124
rect 38936 10081 38945 10115
rect 38945 10081 38979 10115
rect 38979 10081 38988 10115
rect 38936 10072 38988 10081
rect 37832 10047 37884 10056
rect 37832 10013 37841 10047
rect 37841 10013 37875 10047
rect 37875 10013 37884 10047
rect 40960 10072 41012 10124
rect 37832 10004 37884 10013
rect 40040 10004 40092 10056
rect 33232 9936 33284 9988
rect 34060 9936 34112 9988
rect 34612 9936 34664 9988
rect 58164 10004 58216 10056
rect 31024 9868 31076 9920
rect 31576 9868 31628 9920
rect 33784 9911 33836 9920
rect 33784 9877 33793 9911
rect 33793 9877 33827 9911
rect 33827 9877 33836 9911
rect 33784 9868 33836 9877
rect 33876 9868 33928 9920
rect 34152 9911 34204 9920
rect 34152 9877 34161 9911
rect 34161 9877 34195 9911
rect 34195 9877 34204 9911
rect 34152 9868 34204 9877
rect 34520 9868 34572 9920
rect 35808 9868 35860 9920
rect 37188 9868 37240 9920
rect 38936 9868 38988 9920
rect 20214 9766 20266 9818
rect 20278 9766 20330 9818
rect 20342 9766 20394 9818
rect 20406 9766 20458 9818
rect 20470 9766 20522 9818
rect 39478 9766 39530 9818
rect 39542 9766 39594 9818
rect 39606 9766 39658 9818
rect 39670 9766 39722 9818
rect 39734 9766 39786 9818
rect 24676 9707 24728 9716
rect 24676 9673 24685 9707
rect 24685 9673 24719 9707
rect 24719 9673 24728 9707
rect 24676 9664 24728 9673
rect 26148 9664 26200 9716
rect 18420 9596 18472 9648
rect 22008 9392 22060 9444
rect 25412 9596 25464 9648
rect 25964 9596 26016 9648
rect 27712 9664 27764 9716
rect 27896 9664 27948 9716
rect 27988 9664 28040 9716
rect 28448 9707 28500 9716
rect 28448 9673 28457 9707
rect 28457 9673 28491 9707
rect 28491 9673 28500 9707
rect 28448 9664 28500 9673
rect 28632 9707 28684 9716
rect 28632 9673 28641 9707
rect 28641 9673 28675 9707
rect 28675 9673 28684 9707
rect 28632 9664 28684 9673
rect 30564 9664 30616 9716
rect 31024 9664 31076 9716
rect 31852 9664 31904 9716
rect 33140 9664 33192 9716
rect 35072 9664 35124 9716
rect 35164 9664 35216 9716
rect 40868 9664 40920 9716
rect 58164 9707 58216 9716
rect 58164 9673 58173 9707
rect 58173 9673 58207 9707
rect 58207 9673 58216 9707
rect 58164 9664 58216 9673
rect 23848 9528 23900 9580
rect 26240 9571 26292 9580
rect 26240 9537 26249 9571
rect 26249 9537 26283 9571
rect 26283 9537 26292 9571
rect 26240 9528 26292 9537
rect 26884 9528 26936 9580
rect 27344 9528 27396 9580
rect 28356 9571 28408 9580
rect 28356 9537 28365 9571
rect 28365 9537 28399 9571
rect 28399 9537 28408 9571
rect 28356 9528 28408 9537
rect 29276 9571 29328 9580
rect 29276 9537 29285 9571
rect 29285 9537 29319 9571
rect 29319 9537 29328 9571
rect 29276 9528 29328 9537
rect 29460 9528 29512 9580
rect 29828 9528 29880 9580
rect 30104 9571 30156 9580
rect 30104 9537 30113 9571
rect 30113 9537 30147 9571
rect 30147 9537 30156 9571
rect 30104 9528 30156 9537
rect 31116 9571 31168 9580
rect 31116 9537 31125 9571
rect 31125 9537 31159 9571
rect 31159 9537 31168 9571
rect 31116 9528 31168 9537
rect 25044 9460 25096 9512
rect 26332 9460 26384 9512
rect 27804 9460 27856 9512
rect 8668 9324 8720 9376
rect 23572 9392 23624 9444
rect 24768 9392 24820 9444
rect 26424 9392 26476 9444
rect 27712 9392 27764 9444
rect 28080 9392 28132 9444
rect 23480 9324 23532 9376
rect 24400 9324 24452 9376
rect 28448 9324 28500 9376
rect 31024 9503 31076 9512
rect 29828 9392 29880 9444
rect 30656 9392 30708 9444
rect 31024 9469 31033 9503
rect 31033 9469 31067 9503
rect 31067 9469 31076 9503
rect 31024 9460 31076 9469
rect 31944 9596 31996 9648
rect 32496 9639 32548 9648
rect 32496 9605 32505 9639
rect 32505 9605 32539 9639
rect 32539 9605 32548 9639
rect 32496 9596 32548 9605
rect 33048 9596 33100 9648
rect 34152 9596 34204 9648
rect 32404 9571 32456 9580
rect 32404 9537 32413 9571
rect 32413 9537 32447 9571
rect 32447 9537 32456 9571
rect 32404 9528 32456 9537
rect 34244 9528 34296 9580
rect 34428 9571 34480 9580
rect 34428 9537 34437 9571
rect 34437 9537 34471 9571
rect 34471 9537 34480 9571
rect 34428 9528 34480 9537
rect 35348 9596 35400 9648
rect 37188 9596 37240 9648
rect 34980 9528 35032 9580
rect 37004 9528 37056 9580
rect 43260 9528 43312 9580
rect 36268 9460 36320 9512
rect 31300 9392 31352 9444
rect 31484 9435 31536 9444
rect 31484 9401 31493 9435
rect 31493 9401 31527 9435
rect 31527 9401 31536 9435
rect 31484 9392 31536 9401
rect 32680 9435 32732 9444
rect 32680 9401 32689 9435
rect 32689 9401 32723 9435
rect 32723 9401 32732 9435
rect 32680 9392 32732 9401
rect 34244 9392 34296 9444
rect 38476 9460 38528 9512
rect 36912 9392 36964 9444
rect 41696 9460 41748 9512
rect 29460 9367 29512 9376
rect 29460 9333 29469 9367
rect 29469 9333 29503 9367
rect 29503 9333 29512 9367
rect 29460 9324 29512 9333
rect 32312 9324 32364 9376
rect 34520 9367 34572 9376
rect 34520 9333 34529 9367
rect 34529 9333 34563 9367
rect 34563 9333 34572 9367
rect 34520 9324 34572 9333
rect 35164 9367 35216 9376
rect 35164 9333 35173 9367
rect 35173 9333 35207 9367
rect 35207 9333 35216 9367
rect 35164 9324 35216 9333
rect 37004 9324 37056 9376
rect 38016 9324 38068 9376
rect 38660 9324 38712 9376
rect 38936 9367 38988 9376
rect 38936 9333 38945 9367
rect 38945 9333 38979 9367
rect 38979 9333 38988 9367
rect 38936 9324 38988 9333
rect 10582 9222 10634 9274
rect 10646 9222 10698 9274
rect 10710 9222 10762 9274
rect 10774 9222 10826 9274
rect 10838 9222 10890 9274
rect 29846 9222 29898 9274
rect 29910 9222 29962 9274
rect 29974 9222 30026 9274
rect 30038 9222 30090 9274
rect 30102 9222 30154 9274
rect 49110 9222 49162 9274
rect 49174 9222 49226 9274
rect 49238 9222 49290 9274
rect 49302 9222 49354 9274
rect 49366 9222 49418 9274
rect 25780 9120 25832 9172
rect 26516 9163 26568 9172
rect 26516 9129 26525 9163
rect 26525 9129 26559 9163
rect 26559 9129 26568 9163
rect 26516 9120 26568 9129
rect 27712 9163 27764 9172
rect 27712 9129 27721 9163
rect 27721 9129 27755 9163
rect 27755 9129 27764 9163
rect 27712 9120 27764 9129
rect 23848 9052 23900 9104
rect 25136 9052 25188 9104
rect 28632 9120 28684 9172
rect 29368 9120 29420 9172
rect 30472 9120 30524 9172
rect 31576 9163 31628 9172
rect 31576 9129 31585 9163
rect 31585 9129 31619 9163
rect 31619 9129 31628 9163
rect 31576 9120 31628 9129
rect 32956 9120 33008 9172
rect 33324 9163 33376 9172
rect 33324 9129 33333 9163
rect 33333 9129 33367 9163
rect 33367 9129 33376 9163
rect 33324 9120 33376 9129
rect 34428 9120 34480 9172
rect 35256 9163 35308 9172
rect 35256 9129 35265 9163
rect 35265 9129 35299 9163
rect 35299 9129 35308 9163
rect 35256 9120 35308 9129
rect 36268 9120 36320 9172
rect 38660 9120 38712 9172
rect 21732 8984 21784 9036
rect 27712 8984 27764 9036
rect 28448 9052 28500 9104
rect 30932 9095 30984 9104
rect 28080 8984 28132 9036
rect 28264 9027 28316 9036
rect 28264 8993 28273 9027
rect 28273 8993 28307 9027
rect 28307 8993 28316 9027
rect 28264 8984 28316 8993
rect 11520 8916 11572 8968
rect 21272 8916 21324 8968
rect 26976 8916 27028 8968
rect 27068 8916 27120 8968
rect 28632 8984 28684 9036
rect 30932 9061 30941 9095
rect 30941 9061 30975 9095
rect 30975 9061 30984 9095
rect 30932 9052 30984 9061
rect 31668 9052 31720 9104
rect 28724 8916 28776 8968
rect 30104 8984 30156 9036
rect 30656 9027 30708 9036
rect 30656 8993 30665 9027
rect 30665 8993 30699 9027
rect 30699 8993 30708 9027
rect 30656 8984 30708 8993
rect 30564 8959 30616 8968
rect 16856 8848 16908 8900
rect 26424 8848 26476 8900
rect 26516 8848 26568 8900
rect 30564 8925 30573 8959
rect 30573 8925 30607 8959
rect 30607 8925 30616 8959
rect 30564 8916 30616 8925
rect 36820 9052 36872 9104
rect 37648 9052 37700 9104
rect 38568 9052 38620 9104
rect 32404 8984 32456 9036
rect 32864 8984 32916 9036
rect 33048 8984 33100 9036
rect 30012 8848 30064 8900
rect 32036 8916 32088 8968
rect 34336 8984 34388 9036
rect 33692 8916 33744 8968
rect 34244 8916 34296 8968
rect 35256 8984 35308 9036
rect 35532 8984 35584 9036
rect 43812 8984 43864 9036
rect 1492 8823 1544 8832
rect 1492 8789 1501 8823
rect 1501 8789 1535 8823
rect 1535 8789 1544 8823
rect 1492 8780 1544 8789
rect 20628 8780 20680 8832
rect 23296 8823 23348 8832
rect 23296 8789 23305 8823
rect 23305 8789 23339 8823
rect 23339 8789 23348 8823
rect 23296 8780 23348 8789
rect 23848 8823 23900 8832
rect 23848 8789 23857 8823
rect 23857 8789 23891 8823
rect 23891 8789 23900 8823
rect 23848 8780 23900 8789
rect 24124 8780 24176 8832
rect 29368 8780 29420 8832
rect 29920 8823 29972 8832
rect 29920 8789 29929 8823
rect 29929 8789 29963 8823
rect 29963 8789 29972 8823
rect 29920 8780 29972 8789
rect 31392 8823 31444 8832
rect 31392 8789 31401 8823
rect 31401 8789 31435 8823
rect 31435 8789 31444 8823
rect 34428 8848 34480 8900
rect 31392 8780 31444 8789
rect 32680 8780 32732 8832
rect 37464 8916 37516 8968
rect 34704 8848 34756 8900
rect 36360 8891 36412 8900
rect 36360 8857 36369 8891
rect 36369 8857 36403 8891
rect 36403 8857 36412 8891
rect 36360 8848 36412 8857
rect 37832 8848 37884 8900
rect 38936 8848 38988 8900
rect 45560 8780 45612 8832
rect 46204 8780 46256 8832
rect 20214 8678 20266 8730
rect 20278 8678 20330 8730
rect 20342 8678 20394 8730
rect 20406 8678 20458 8730
rect 20470 8678 20522 8730
rect 39478 8678 39530 8730
rect 39542 8678 39594 8730
rect 39606 8678 39658 8730
rect 39670 8678 39722 8730
rect 39734 8678 39786 8730
rect 23480 8576 23532 8628
rect 24952 8576 25004 8628
rect 26332 8619 26384 8628
rect 26332 8585 26341 8619
rect 26341 8585 26375 8619
rect 26375 8585 26384 8619
rect 26332 8576 26384 8585
rect 27068 8619 27120 8628
rect 27068 8585 27077 8619
rect 27077 8585 27111 8619
rect 27111 8585 27120 8619
rect 27068 8576 27120 8585
rect 27620 8619 27672 8628
rect 27620 8585 27629 8619
rect 27629 8585 27663 8619
rect 27663 8585 27672 8619
rect 27620 8576 27672 8585
rect 27712 8576 27764 8628
rect 27988 8576 28040 8628
rect 28172 8619 28224 8628
rect 28172 8585 28181 8619
rect 28181 8585 28215 8619
rect 28215 8585 28224 8619
rect 28172 8576 28224 8585
rect 28724 8619 28776 8628
rect 28724 8585 28733 8619
rect 28733 8585 28767 8619
rect 28767 8585 28776 8619
rect 28724 8576 28776 8585
rect 25504 8508 25556 8560
rect 28632 8508 28684 8560
rect 25780 8483 25832 8492
rect 25780 8449 25789 8483
rect 25789 8449 25823 8483
rect 25823 8449 25832 8483
rect 25780 8440 25832 8449
rect 28816 8483 28868 8492
rect 28816 8449 28825 8483
rect 28825 8449 28859 8483
rect 28859 8449 28868 8483
rect 28816 8440 28868 8449
rect 32220 8576 32272 8628
rect 32588 8576 32640 8628
rect 32680 8576 32732 8628
rect 33416 8576 33468 8628
rect 33968 8576 34020 8628
rect 34152 8619 34204 8628
rect 34152 8585 34161 8619
rect 34161 8585 34195 8619
rect 34195 8585 34204 8619
rect 34152 8576 34204 8585
rect 34612 8576 34664 8628
rect 37280 8576 37332 8628
rect 37372 8619 37424 8628
rect 37372 8585 37381 8619
rect 37381 8585 37415 8619
rect 37415 8585 37424 8619
rect 37372 8576 37424 8585
rect 40224 8576 40276 8628
rect 29368 8508 29420 8560
rect 30012 8508 30064 8560
rect 30104 8508 30156 8560
rect 30196 8440 30248 8492
rect 19432 8372 19484 8424
rect 23296 8372 23348 8424
rect 26792 8372 26844 8424
rect 29368 8415 29420 8424
rect 29368 8381 29377 8415
rect 29377 8381 29411 8415
rect 29411 8381 29420 8415
rect 29368 8372 29420 8381
rect 29736 8372 29788 8424
rect 29920 8372 29972 8424
rect 30932 8440 30984 8492
rect 31300 8551 31352 8560
rect 31300 8517 31341 8551
rect 31341 8517 31352 8551
rect 31300 8508 31352 8517
rect 32956 8508 33008 8560
rect 35716 8551 35768 8560
rect 35716 8517 35725 8551
rect 35725 8517 35759 8551
rect 35759 8517 35768 8551
rect 35716 8508 35768 8517
rect 36084 8508 36136 8560
rect 38752 8508 38804 8560
rect 31760 8440 31812 8492
rect 32128 8483 32180 8492
rect 32128 8449 32137 8483
rect 32137 8449 32171 8483
rect 32171 8449 32180 8483
rect 32128 8440 32180 8449
rect 32864 8483 32916 8492
rect 32864 8449 32873 8483
rect 32873 8449 32907 8483
rect 32907 8449 32916 8483
rect 32864 8440 32916 8449
rect 33048 8440 33100 8492
rect 35256 8440 35308 8492
rect 35624 8372 35676 8424
rect 31576 8304 31628 8356
rect 30840 8236 30892 8288
rect 31300 8279 31352 8288
rect 31300 8245 31309 8279
rect 31309 8245 31343 8279
rect 31343 8245 31352 8279
rect 32036 8304 32088 8356
rect 33048 8304 33100 8356
rect 31300 8236 31352 8245
rect 31944 8236 31996 8288
rect 32680 8236 32732 8288
rect 38108 8304 38160 8356
rect 37188 8236 37240 8288
rect 37832 8279 37884 8288
rect 37832 8245 37841 8279
rect 37841 8245 37875 8279
rect 37875 8245 37884 8279
rect 37832 8236 37884 8245
rect 10582 8134 10634 8186
rect 10646 8134 10698 8186
rect 10710 8134 10762 8186
rect 10774 8134 10826 8186
rect 10838 8134 10890 8186
rect 29846 8134 29898 8186
rect 29910 8134 29962 8186
rect 29974 8134 30026 8186
rect 30038 8134 30090 8186
rect 30102 8134 30154 8186
rect 49110 8134 49162 8186
rect 49174 8134 49226 8186
rect 49238 8134 49290 8186
rect 49302 8134 49354 8186
rect 49366 8134 49418 8186
rect 24768 8032 24820 8084
rect 25964 8075 26016 8084
rect 25964 8041 25973 8075
rect 25973 8041 26007 8075
rect 26007 8041 26016 8075
rect 25964 8032 26016 8041
rect 26056 8032 26108 8084
rect 27252 8075 27304 8084
rect 27252 8041 27261 8075
rect 27261 8041 27295 8075
rect 27295 8041 27304 8075
rect 27252 8032 27304 8041
rect 28080 8032 28132 8084
rect 29644 8075 29696 8084
rect 29644 8041 29653 8075
rect 29653 8041 29687 8075
rect 29687 8041 29696 8075
rect 29644 8032 29696 8041
rect 27804 7964 27856 8016
rect 31116 8032 31168 8084
rect 32220 8032 32272 8084
rect 32956 8075 33008 8084
rect 32956 8041 32965 8075
rect 32965 8041 32999 8075
rect 32999 8041 33008 8075
rect 32956 8032 33008 8041
rect 33600 8075 33652 8084
rect 33600 8041 33609 8075
rect 33609 8041 33643 8075
rect 33643 8041 33652 8075
rect 33600 8032 33652 8041
rect 30472 7964 30524 8016
rect 38844 8032 38896 8084
rect 34980 7964 35032 8016
rect 43076 7964 43128 8016
rect 14464 7803 14516 7812
rect 14464 7769 14473 7803
rect 14473 7769 14507 7803
rect 14507 7769 14516 7803
rect 14464 7760 14516 7769
rect 15292 7735 15344 7744
rect 15292 7701 15301 7735
rect 15301 7701 15335 7735
rect 15335 7701 15344 7735
rect 15292 7692 15344 7701
rect 25504 7735 25556 7744
rect 25504 7701 25513 7735
rect 25513 7701 25547 7735
rect 25547 7701 25556 7735
rect 25504 7692 25556 7701
rect 26148 7692 26200 7744
rect 30288 7692 30340 7744
rect 33140 7896 33192 7948
rect 33784 7896 33836 7948
rect 44272 7896 44324 7948
rect 51724 7896 51776 7948
rect 30932 7828 30984 7880
rect 31116 7871 31168 7880
rect 31116 7837 31125 7871
rect 31125 7837 31159 7871
rect 31159 7837 31168 7871
rect 31116 7828 31168 7837
rect 32864 7828 32916 7880
rect 33968 7828 34020 7880
rect 37556 7828 37608 7880
rect 58164 7871 58216 7880
rect 58164 7837 58173 7871
rect 58173 7837 58207 7871
rect 58207 7837 58216 7871
rect 58164 7828 58216 7837
rect 30656 7760 30708 7812
rect 31024 7760 31076 7812
rect 34704 7803 34756 7812
rect 34704 7769 34713 7803
rect 34713 7769 34747 7803
rect 34747 7769 34756 7803
rect 34704 7760 34756 7769
rect 35256 7803 35308 7812
rect 35256 7769 35265 7803
rect 35265 7769 35299 7803
rect 35299 7769 35308 7803
rect 35256 7760 35308 7769
rect 35348 7760 35400 7812
rect 37832 7760 37884 7812
rect 30472 7692 30524 7744
rect 32312 7692 32364 7744
rect 36360 7735 36412 7744
rect 36360 7701 36369 7735
rect 36369 7701 36403 7735
rect 36403 7701 36412 7735
rect 36360 7692 36412 7701
rect 36912 7735 36964 7744
rect 36912 7701 36921 7735
rect 36921 7701 36955 7735
rect 36955 7701 36964 7735
rect 36912 7692 36964 7701
rect 20214 7590 20266 7642
rect 20278 7590 20330 7642
rect 20342 7590 20394 7642
rect 20406 7590 20458 7642
rect 20470 7590 20522 7642
rect 39478 7590 39530 7642
rect 39542 7590 39594 7642
rect 39606 7590 39658 7642
rect 39670 7590 39722 7642
rect 39734 7590 39786 7642
rect 25872 7531 25924 7540
rect 25872 7497 25881 7531
rect 25881 7497 25915 7531
rect 25915 7497 25924 7531
rect 25872 7488 25924 7497
rect 26240 7488 26292 7540
rect 26424 7488 26476 7540
rect 27528 7488 27580 7540
rect 28540 7531 28592 7540
rect 28540 7497 28549 7531
rect 28549 7497 28583 7531
rect 28583 7497 28592 7531
rect 28540 7488 28592 7497
rect 28908 7488 28960 7540
rect 29184 7488 29236 7540
rect 15292 7420 15344 7472
rect 8668 7352 8720 7404
rect 29000 7420 29052 7472
rect 30748 7488 30800 7540
rect 31024 7531 31076 7540
rect 31024 7497 31033 7531
rect 31033 7497 31067 7531
rect 31067 7497 31076 7531
rect 31024 7488 31076 7497
rect 31760 7488 31812 7540
rect 32680 7531 32732 7540
rect 32680 7497 32689 7531
rect 32689 7497 32723 7531
rect 32723 7497 32732 7531
rect 32680 7488 32732 7497
rect 33876 7531 33928 7540
rect 33876 7497 33885 7531
rect 33885 7497 33919 7531
rect 33919 7497 33928 7531
rect 33876 7488 33928 7497
rect 34980 7531 35032 7540
rect 34980 7497 34989 7531
rect 34989 7497 35023 7531
rect 35023 7497 35032 7531
rect 34980 7488 35032 7497
rect 36084 7531 36136 7540
rect 36084 7497 36093 7531
rect 36093 7497 36127 7531
rect 36127 7497 36136 7531
rect 36084 7488 36136 7497
rect 58164 7531 58216 7540
rect 58164 7497 58173 7531
rect 58173 7497 58207 7531
rect 58207 7497 58216 7531
rect 58164 7488 58216 7497
rect 32588 7420 32640 7472
rect 23388 7352 23440 7404
rect 29644 7352 29696 7404
rect 30288 7395 30340 7404
rect 30288 7361 30297 7395
rect 30297 7361 30331 7395
rect 30331 7361 30340 7395
rect 30288 7352 30340 7361
rect 32772 7352 32824 7404
rect 37648 7352 37700 7404
rect 37188 7284 37240 7336
rect 30472 7216 30524 7268
rect 35256 7216 35308 7268
rect 35900 7216 35952 7268
rect 36912 7216 36964 7268
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 26700 7148 26752 7200
rect 27252 7148 27304 7200
rect 34428 7191 34480 7200
rect 34428 7157 34437 7191
rect 34437 7157 34471 7191
rect 34471 7157 34480 7191
rect 34428 7148 34480 7157
rect 35348 7148 35400 7200
rect 10582 7046 10634 7098
rect 10646 7046 10698 7098
rect 10710 7046 10762 7098
rect 10774 7046 10826 7098
rect 10838 7046 10890 7098
rect 29846 7046 29898 7098
rect 29910 7046 29962 7098
rect 29974 7046 30026 7098
rect 30038 7046 30090 7098
rect 30102 7046 30154 7098
rect 49110 7046 49162 7098
rect 49174 7046 49226 7098
rect 49238 7046 49290 7098
rect 49302 7046 49354 7098
rect 49366 7046 49418 7098
rect 30840 6944 30892 6996
rect 31300 6944 31352 6996
rect 32588 6944 32640 6996
rect 24584 6808 24636 6860
rect 29368 6808 29420 6860
rect 29736 6808 29788 6860
rect 34060 6808 34112 6860
rect 34244 6808 34296 6860
rect 16304 6740 16356 6792
rect 28356 6740 28408 6792
rect 28908 6740 28960 6792
rect 29276 6740 29328 6792
rect 33784 6740 33836 6792
rect 34428 6740 34480 6792
rect 45652 6740 45704 6792
rect 22744 6672 22796 6724
rect 27252 6715 27304 6724
rect 26240 6647 26292 6656
rect 26240 6613 26249 6647
rect 26249 6613 26283 6647
rect 26283 6613 26292 6647
rect 26240 6604 26292 6613
rect 26792 6647 26844 6656
rect 26792 6613 26801 6647
rect 26801 6613 26835 6647
rect 26835 6613 26844 6647
rect 26792 6604 26844 6613
rect 27252 6681 27261 6715
rect 27261 6681 27295 6715
rect 27295 6681 27304 6715
rect 27252 6672 27304 6681
rect 27344 6672 27396 6724
rect 28632 6672 28684 6724
rect 31944 6672 31996 6724
rect 32036 6672 32088 6724
rect 41880 6672 41932 6724
rect 33416 6604 33468 6656
rect 35348 6647 35400 6656
rect 35348 6613 35357 6647
rect 35357 6613 35391 6647
rect 35391 6613 35400 6647
rect 35348 6604 35400 6613
rect 35900 6647 35952 6656
rect 35900 6613 35909 6647
rect 35909 6613 35943 6647
rect 35943 6613 35952 6647
rect 35900 6604 35952 6613
rect 20214 6502 20266 6554
rect 20278 6502 20330 6554
rect 20342 6502 20394 6554
rect 20406 6502 20458 6554
rect 20470 6502 20522 6554
rect 39478 6502 39530 6554
rect 39542 6502 39594 6554
rect 39606 6502 39658 6554
rect 39670 6502 39722 6554
rect 39734 6502 39786 6554
rect 29368 6400 29420 6452
rect 30196 6443 30248 6452
rect 30196 6409 30205 6443
rect 30205 6409 30239 6443
rect 30239 6409 30248 6443
rect 30196 6400 30248 6409
rect 30564 6400 30616 6452
rect 32128 6443 32180 6452
rect 32128 6409 32137 6443
rect 32137 6409 32171 6443
rect 32171 6409 32180 6443
rect 32128 6400 32180 6409
rect 32772 6443 32824 6452
rect 32772 6409 32781 6443
rect 32781 6409 32815 6443
rect 32815 6409 32824 6443
rect 32772 6400 32824 6409
rect 36084 6400 36136 6452
rect 27988 6332 28040 6384
rect 28908 6332 28960 6384
rect 29644 6332 29696 6384
rect 34244 6332 34296 6384
rect 26792 6264 26844 6316
rect 35348 6264 35400 6316
rect 27252 6196 27304 6248
rect 36636 6196 36688 6248
rect 15752 6128 15804 6180
rect 30656 6128 30708 6180
rect 31944 6128 31996 6180
rect 39120 6128 39172 6180
rect 26240 6060 26292 6112
rect 27344 6103 27396 6112
rect 27344 6069 27353 6103
rect 27353 6069 27387 6103
rect 27387 6069 27396 6103
rect 27344 6060 27396 6069
rect 10582 5958 10634 6010
rect 10646 5958 10698 6010
rect 10710 5958 10762 6010
rect 10774 5958 10826 6010
rect 10838 5958 10890 6010
rect 29846 5958 29898 6010
rect 29910 5958 29962 6010
rect 29974 5958 30026 6010
rect 30038 5958 30090 6010
rect 30102 5958 30154 6010
rect 49110 5958 49162 6010
rect 49174 5958 49226 6010
rect 49238 5958 49290 6010
rect 49302 5958 49354 6010
rect 49366 5958 49418 6010
rect 28448 5899 28500 5908
rect 28448 5865 28457 5899
rect 28457 5865 28491 5899
rect 28491 5865 28500 5899
rect 28448 5856 28500 5865
rect 28816 5856 28868 5908
rect 29644 5899 29696 5908
rect 29644 5865 29653 5899
rect 29653 5865 29687 5899
rect 29687 5865 29696 5899
rect 29644 5856 29696 5865
rect 30288 5856 30340 5908
rect 30472 5856 30524 5908
rect 31116 5856 31168 5908
rect 32220 5856 32272 5908
rect 36360 5856 36412 5908
rect 32864 5831 32916 5840
rect 32864 5797 32873 5831
rect 32873 5797 32907 5831
rect 32907 5797 32916 5831
rect 32864 5788 32916 5797
rect 33508 5831 33560 5840
rect 33508 5797 33517 5831
rect 33517 5797 33551 5831
rect 33551 5797 33560 5831
rect 33508 5788 33560 5797
rect 35900 5788 35952 5840
rect 14464 5720 14516 5772
rect 32772 5720 32824 5772
rect 58164 5695 58216 5704
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 8852 5516 8904 5568
rect 58164 5661 58173 5695
rect 58173 5661 58207 5695
rect 58207 5661 58216 5695
rect 58164 5652 58216 5661
rect 37188 5584 37240 5636
rect 22008 5516 22060 5568
rect 20214 5414 20266 5466
rect 20278 5414 20330 5466
rect 20342 5414 20394 5466
rect 20406 5414 20458 5466
rect 20470 5414 20522 5466
rect 39478 5414 39530 5466
rect 39542 5414 39594 5466
rect 39606 5414 39658 5466
rect 39670 5414 39722 5466
rect 39734 5414 39786 5466
rect 18420 5312 18472 5364
rect 29460 5355 29512 5364
rect 14924 5244 14976 5296
rect 29460 5321 29469 5355
rect 29469 5321 29503 5355
rect 29503 5321 29512 5355
rect 29460 5312 29512 5321
rect 30380 5312 30432 5364
rect 30564 5312 30616 5364
rect 41788 5312 41840 5364
rect 58164 5355 58216 5364
rect 58164 5321 58173 5355
rect 58173 5321 58207 5355
rect 58207 5321 58216 5355
rect 58164 5312 58216 5321
rect 32220 5287 32272 5296
rect 27344 5176 27396 5228
rect 32220 5253 32229 5287
rect 32229 5253 32263 5287
rect 32263 5253 32272 5287
rect 32220 5244 32272 5253
rect 37280 5040 37332 5092
rect 10582 4870 10634 4922
rect 10646 4870 10698 4922
rect 10710 4870 10762 4922
rect 10774 4870 10826 4922
rect 10838 4870 10890 4922
rect 29846 4870 29898 4922
rect 29910 4870 29962 4922
rect 29974 4870 30026 4922
rect 30038 4870 30090 4922
rect 30102 4870 30154 4922
rect 49110 4870 49162 4922
rect 49174 4870 49226 4922
rect 49238 4870 49290 4922
rect 49302 4870 49354 4922
rect 49366 4870 49418 4922
rect 29552 4811 29604 4820
rect 29552 4777 29561 4811
rect 29561 4777 29595 4811
rect 29595 4777 29604 4811
rect 29552 4768 29604 4777
rect 58164 4564 58216 4616
rect 41696 4496 41748 4548
rect 20214 4326 20266 4378
rect 20278 4326 20330 4378
rect 20342 4326 20394 4378
rect 20406 4326 20458 4378
rect 20470 4326 20522 4378
rect 39478 4326 39530 4378
rect 39542 4326 39594 4378
rect 39606 4326 39658 4378
rect 39670 4326 39722 4378
rect 39734 4326 39786 4378
rect 58164 4267 58216 4276
rect 58164 4233 58173 4267
rect 58173 4233 58207 4267
rect 58207 4233 58216 4267
rect 58164 4224 58216 4233
rect 16120 4088 16172 4140
rect 47124 4088 47176 4140
rect 19248 4020 19300 4072
rect 45100 4020 45152 4072
rect 20996 3952 21048 4004
rect 23572 3952 23624 4004
rect 48504 3952 48556 4004
rect 1492 3927 1544 3936
rect 1492 3893 1501 3927
rect 1501 3893 1535 3927
rect 1535 3893 1544 3927
rect 1492 3884 1544 3893
rect 10582 3782 10634 3834
rect 10646 3782 10698 3834
rect 10710 3782 10762 3834
rect 10774 3782 10826 3834
rect 10838 3782 10890 3834
rect 29846 3782 29898 3834
rect 29910 3782 29962 3834
rect 29974 3782 30026 3834
rect 30038 3782 30090 3834
rect 30102 3782 30154 3834
rect 49110 3782 49162 3834
rect 49174 3782 49226 3834
rect 49238 3782 49290 3834
rect 49302 3782 49354 3834
rect 49366 3782 49418 3834
rect 42432 3612 42484 3664
rect 37832 3476 37884 3528
rect 20214 3238 20266 3290
rect 20278 3238 20330 3290
rect 20342 3238 20394 3290
rect 20406 3238 20458 3290
rect 20470 3238 20522 3290
rect 39478 3238 39530 3290
rect 39542 3238 39594 3290
rect 39606 3238 39658 3290
rect 39670 3238 39722 3290
rect 39734 3238 39786 3290
rect 8852 3000 8904 3052
rect 37740 3043 37792 3052
rect 37740 3009 37749 3043
rect 37749 3009 37783 3043
rect 37783 3009 37792 3043
rect 37740 3000 37792 3009
rect 37924 2907 37976 2916
rect 37924 2873 37933 2907
rect 37933 2873 37967 2907
rect 37967 2873 37976 2907
rect 37924 2864 37976 2873
rect 1400 2839 1452 2848
rect 1400 2805 1409 2839
rect 1409 2805 1443 2839
rect 1443 2805 1452 2839
rect 1400 2796 1452 2805
rect 10582 2694 10634 2746
rect 10646 2694 10698 2746
rect 10710 2694 10762 2746
rect 10774 2694 10826 2746
rect 10838 2694 10890 2746
rect 29846 2694 29898 2746
rect 29910 2694 29962 2746
rect 29974 2694 30026 2746
rect 30038 2694 30090 2746
rect 30102 2694 30154 2746
rect 49110 2694 49162 2746
rect 49174 2694 49226 2746
rect 49238 2694 49290 2746
rect 49302 2694 49354 2746
rect 49366 2694 49418 2746
rect 30564 2592 30616 2644
rect 56508 2592 56560 2644
rect 12900 2524 12952 2576
rect 17960 2524 18012 2576
rect 46940 2524 46992 2576
rect 1492 2295 1544 2304
rect 1492 2261 1501 2295
rect 1501 2261 1535 2295
rect 1535 2261 1544 2295
rect 1492 2252 1544 2261
rect 24860 2456 24912 2508
rect 25872 2456 25924 2508
rect 48780 2456 48832 2508
rect 29920 2388 29972 2440
rect 37740 2388 37792 2440
rect 42432 2431 42484 2440
rect 42432 2397 42441 2431
rect 42441 2397 42475 2431
rect 42475 2397 42484 2431
rect 42432 2388 42484 2397
rect 37832 2320 37884 2372
rect 37924 2320 37976 2372
rect 46204 2320 46256 2372
rect 6000 2252 6052 2304
rect 17960 2252 18012 2304
rect 31208 2252 31260 2304
rect 41972 2252 42024 2304
rect 53932 2252 53984 2304
rect 57888 2295 57940 2304
rect 57888 2261 57897 2295
rect 57897 2261 57931 2295
rect 57931 2261 57940 2295
rect 57888 2252 57940 2261
rect 20214 2150 20266 2202
rect 20278 2150 20330 2202
rect 20342 2150 20394 2202
rect 20406 2150 20458 2202
rect 20470 2150 20522 2202
rect 39478 2150 39530 2202
rect 39542 2150 39594 2202
rect 39606 2150 39658 2202
rect 39670 2150 39722 2202
rect 39734 2150 39786 2202
rect 24400 2048 24452 2100
rect 45376 2048 45428 2100
rect 25504 1980 25556 2032
rect 45468 1980 45520 2032
rect 26056 1912 26108 1964
rect 48412 1912 48464 1964
<< metal2 >>
rect 1398 29200 1454 29209
rect 2686 29200 2742 30000
rect 8114 29322 8170 30000
rect 13542 29322 13598 30000
rect 18326 29608 18382 29617
rect 18326 29543 18382 29552
rect 8114 29294 8248 29322
rect 8114 29200 8170 29294
rect 1398 29135 1454 29144
rect 1412 27130 1440 29135
rect 1492 27600 1544 27606
rect 1490 27568 1492 27577
rect 1544 27568 1546 27577
rect 2700 27554 2728 29200
rect 2780 27600 2832 27606
rect 2700 27548 2780 27554
rect 2700 27542 2832 27548
rect 8220 27554 8248 29294
rect 13542 29294 13768 29322
rect 13542 29200 13598 29294
rect 10582 27772 10890 27792
rect 10582 27770 10588 27772
rect 10644 27770 10668 27772
rect 10724 27770 10748 27772
rect 10804 27770 10828 27772
rect 10884 27770 10890 27772
rect 10644 27718 10646 27770
rect 10826 27718 10828 27770
rect 10582 27716 10588 27718
rect 10644 27716 10668 27718
rect 10724 27716 10748 27718
rect 10804 27716 10828 27718
rect 10884 27716 10890 27718
rect 10582 27696 10890 27716
rect 8300 27600 8352 27606
rect 8220 27548 8300 27554
rect 8220 27542 8352 27548
rect 13740 27554 13768 29294
rect 14830 28792 14886 28801
rect 14830 28727 14886 28736
rect 14738 28656 14794 28665
rect 14738 28591 14794 28600
rect 14554 28384 14610 28393
rect 14554 28319 14610 28328
rect 14096 27872 14148 27878
rect 14096 27814 14148 27820
rect 2700 27526 2820 27542
rect 8220 27526 8340 27542
rect 13740 27526 13860 27554
rect 1490 27503 1546 27512
rect 13832 27470 13860 27526
rect 3884 27464 3936 27470
rect 3884 27406 3936 27412
rect 13820 27464 13872 27470
rect 13820 27406 13872 27412
rect 3896 27334 3924 27406
rect 3884 27328 3936 27334
rect 3884 27270 3936 27276
rect 9772 27328 9824 27334
rect 9772 27270 9824 27276
rect 1400 27124 1452 27130
rect 1400 27066 1452 27072
rect 3896 26858 3924 27270
rect 9784 27130 9812 27270
rect 9772 27124 9824 27130
rect 9772 27066 9824 27072
rect 3884 26852 3936 26858
rect 3884 26794 3936 26800
rect 10582 26684 10890 26704
rect 10582 26682 10588 26684
rect 10644 26682 10668 26684
rect 10724 26682 10748 26684
rect 10804 26682 10828 26684
rect 10884 26682 10890 26684
rect 10644 26630 10646 26682
rect 10826 26630 10828 26682
rect 10582 26628 10588 26630
rect 10644 26628 10668 26630
rect 10724 26628 10748 26630
rect 10804 26628 10828 26630
rect 10884 26628 10890 26630
rect 10582 26608 10890 26628
rect 8576 26376 8628 26382
rect 8576 26318 8628 26324
rect 1492 26240 1544 26246
rect 1492 26182 1544 26188
rect 1504 26081 1532 26182
rect 1490 26072 1546 26081
rect 1490 26007 1546 26016
rect 2228 25764 2280 25770
rect 2228 25706 2280 25712
rect 1492 24608 1544 24614
rect 1492 24550 1544 24556
rect 1504 24449 1532 24550
rect 1490 24440 1546 24449
rect 1490 24375 1546 24384
rect 2240 23322 2268 25706
rect 8588 24682 8616 26318
rect 10582 25596 10890 25616
rect 10582 25594 10588 25596
rect 10644 25594 10668 25596
rect 10724 25594 10748 25596
rect 10804 25594 10828 25596
rect 10884 25594 10890 25596
rect 10644 25542 10646 25594
rect 10826 25542 10828 25594
rect 10582 25540 10588 25542
rect 10644 25540 10668 25542
rect 10724 25540 10748 25542
rect 10804 25540 10828 25542
rect 10884 25540 10890 25542
rect 10582 25520 10890 25540
rect 9128 24812 9180 24818
rect 9128 24754 9180 24760
rect 8576 24676 8628 24682
rect 8576 24618 8628 24624
rect 9140 24410 9168 24754
rect 12348 24676 12400 24682
rect 12348 24618 12400 24624
rect 10582 24508 10890 24528
rect 10582 24506 10588 24508
rect 10644 24506 10668 24508
rect 10724 24506 10748 24508
rect 10804 24506 10828 24508
rect 10884 24506 10890 24508
rect 10644 24454 10646 24506
rect 10826 24454 10828 24506
rect 10582 24452 10588 24454
rect 10644 24452 10668 24454
rect 10724 24452 10748 24454
rect 10804 24452 10828 24454
rect 10884 24452 10890 24454
rect 10582 24432 10890 24452
rect 9128 24404 9180 24410
rect 9128 24346 9180 24352
rect 10582 23420 10890 23440
rect 10582 23418 10588 23420
rect 10644 23418 10668 23420
rect 10724 23418 10748 23420
rect 10804 23418 10828 23420
rect 10884 23418 10890 23420
rect 10644 23366 10646 23418
rect 10826 23366 10828 23418
rect 10582 23364 10588 23366
rect 10644 23364 10668 23366
rect 10724 23364 10748 23366
rect 10804 23364 10828 23366
rect 10884 23364 10890 23366
rect 10582 23344 10890 23364
rect 2228 23316 2280 23322
rect 2228 23258 2280 23264
rect 2240 23118 2268 23258
rect 2228 23112 2280 23118
rect 2228 23054 2280 23060
rect 1492 22976 1544 22982
rect 1492 22918 1544 22924
rect 1504 22817 1532 22918
rect 1490 22808 1546 22817
rect 1490 22743 1546 22752
rect 10582 22332 10890 22352
rect 10582 22330 10588 22332
rect 10644 22330 10668 22332
rect 10724 22330 10748 22332
rect 10804 22330 10828 22332
rect 10884 22330 10890 22332
rect 10644 22278 10646 22330
rect 10826 22278 10828 22330
rect 10582 22276 10588 22278
rect 10644 22276 10668 22278
rect 10724 22276 10748 22278
rect 10804 22276 10828 22278
rect 10884 22276 10890 22278
rect 10582 22256 10890 22276
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 1492 21344 1544 21350
rect 1490 21312 1492 21321
rect 1544 21312 1546 21321
rect 1490 21247 1546 21256
rect 10582 21244 10890 21264
rect 10582 21242 10588 21244
rect 10644 21242 10668 21244
rect 10724 21242 10748 21244
rect 10804 21242 10828 21244
rect 10884 21242 10890 21244
rect 10644 21190 10646 21242
rect 10826 21190 10828 21242
rect 10582 21188 10588 21190
rect 10644 21188 10668 21190
rect 10724 21188 10748 21190
rect 10804 21188 10828 21190
rect 10884 21188 10890 21190
rect 10582 21168 10890 21188
rect 10582 20156 10890 20176
rect 10582 20154 10588 20156
rect 10644 20154 10668 20156
rect 10724 20154 10748 20156
rect 10804 20154 10828 20156
rect 10884 20154 10890 20156
rect 10644 20102 10646 20154
rect 10826 20102 10828 20154
rect 10582 20100 10588 20102
rect 10644 20100 10668 20102
rect 10724 20100 10748 20102
rect 10804 20100 10828 20102
rect 10884 20100 10890 20102
rect 10582 20080 10890 20100
rect 12268 19990 12296 21490
rect 12256 19984 12308 19990
rect 12256 19926 12308 19932
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 1492 19712 1544 19718
rect 1490 19680 1492 19689
rect 1544 19680 1546 19689
rect 1490 19615 1546 19624
rect 12084 19514 12112 19790
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 12360 19310 12388 24618
rect 13910 21992 13966 22001
rect 13910 21927 13966 21936
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 10582 19068 10890 19088
rect 10582 19066 10588 19068
rect 10644 19066 10668 19068
rect 10724 19066 10748 19068
rect 10804 19066 10828 19068
rect 10884 19066 10890 19068
rect 10644 19014 10646 19066
rect 10826 19014 10828 19066
rect 10582 19012 10588 19014
rect 10644 19012 10668 19014
rect 10724 19012 10748 19014
rect 10804 19012 10828 19014
rect 10884 19012 10890 19014
rect 10582 18992 10890 19012
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 1492 18080 1544 18086
rect 1490 18048 1492 18057
rect 12164 18080 12216 18086
rect 1544 18048 1546 18057
rect 12164 18022 12216 18028
rect 1490 17983 1546 17992
rect 10582 17980 10890 18000
rect 10582 17978 10588 17980
rect 10644 17978 10668 17980
rect 10724 17978 10748 17980
rect 10804 17978 10828 17980
rect 10884 17978 10890 17980
rect 10644 17926 10646 17978
rect 10826 17926 10828 17978
rect 10582 17924 10588 17926
rect 10644 17924 10668 17926
rect 10724 17924 10748 17926
rect 10804 17924 10828 17926
rect 10884 17924 10890 17926
rect 10582 17904 10890 17924
rect 11888 17060 11940 17066
rect 11888 17002 11940 17008
rect 10582 16892 10890 16912
rect 10582 16890 10588 16892
rect 10644 16890 10668 16892
rect 10724 16890 10748 16892
rect 10804 16890 10828 16892
rect 10884 16890 10890 16892
rect 10644 16838 10646 16890
rect 10826 16838 10828 16890
rect 10582 16836 10588 16838
rect 10644 16836 10668 16838
rect 10724 16836 10748 16838
rect 10804 16836 10828 16838
rect 10884 16836 10890 16838
rect 10582 16816 10890 16836
rect 11900 16794 11928 17002
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 1490 16552 1546 16561
rect 1490 16487 1546 16496
rect 1504 16454 1532 16487
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 10582 15804 10890 15824
rect 10582 15802 10588 15804
rect 10644 15802 10668 15804
rect 10724 15802 10748 15804
rect 10804 15802 10828 15804
rect 10884 15802 10890 15804
rect 10644 15750 10646 15802
rect 10826 15750 10828 15802
rect 10582 15748 10588 15750
rect 10644 15748 10668 15750
rect 10724 15748 10748 15750
rect 10804 15748 10828 15750
rect 10884 15748 10890 15750
rect 10582 15728 10890 15748
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 11256 15026 11284 15302
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 1490 14920 1546 14929
rect 1490 14855 1492 14864
rect 1544 14855 1546 14864
rect 1492 14826 1544 14832
rect 10582 14716 10890 14736
rect 10582 14714 10588 14716
rect 10644 14714 10668 14716
rect 10724 14714 10748 14716
rect 10804 14714 10828 14716
rect 10884 14714 10890 14716
rect 10644 14662 10646 14714
rect 10826 14662 10828 14714
rect 10582 14660 10588 14662
rect 10644 14660 10668 14662
rect 10724 14660 10748 14662
rect 10804 14660 10828 14662
rect 10884 14660 10890 14662
rect 10582 14640 10890 14660
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10612 13938 10640 14214
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 1492 13728 1544 13734
rect 1492 13670 1544 13676
rect 1504 13433 1532 13670
rect 10582 13628 10890 13648
rect 10582 13626 10588 13628
rect 10644 13626 10668 13628
rect 10724 13626 10748 13628
rect 10804 13626 10828 13628
rect 10884 13626 10890 13628
rect 10644 13574 10646 13626
rect 10826 13574 10828 13626
rect 10582 13572 10588 13574
rect 10644 13572 10668 13574
rect 10724 13572 10748 13574
rect 10804 13572 10828 13574
rect 10884 13572 10890 13574
rect 10582 13552 10890 13572
rect 12176 13462 12204 18022
rect 12268 16250 12296 18906
rect 12728 18358 12756 20538
rect 13740 19718 13768 20742
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 12716 18352 12768 18358
rect 12716 18294 12768 18300
rect 12728 17338 12756 18294
rect 13004 17542 13032 19654
rect 13832 18086 13860 20198
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13924 17882 13952 21927
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 14108 17785 14136 27814
rect 14372 27532 14424 27538
rect 14372 27474 14424 27480
rect 14280 27328 14332 27334
rect 14280 27270 14332 27276
rect 14292 26926 14320 27270
rect 14280 26920 14332 26926
rect 14280 26862 14332 26868
rect 14384 24342 14412 27474
rect 14464 26988 14516 26994
rect 14464 26930 14516 26936
rect 14476 25430 14504 26930
rect 14464 25424 14516 25430
rect 14464 25366 14516 25372
rect 14372 24336 14424 24342
rect 14372 24278 14424 24284
rect 14462 21584 14518 21593
rect 14462 21519 14518 21528
rect 14278 19680 14334 19689
rect 14278 19615 14334 19624
rect 14186 18864 14242 18873
rect 14186 18799 14188 18808
rect 14240 18799 14242 18808
rect 14188 18770 14240 18776
rect 14094 17776 14150 17785
rect 14094 17711 14150 17720
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12636 16998 12664 17070
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12636 14278 12664 16934
rect 12728 15162 12756 17274
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12164 13456 12216 13462
rect 1490 13424 1546 13433
rect 12164 13398 12216 13404
rect 1490 13359 1546 13368
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 10582 12540 10890 12560
rect 10582 12538 10588 12540
rect 10644 12538 10668 12540
rect 10724 12538 10748 12540
rect 10804 12538 10828 12540
rect 10884 12538 10890 12540
rect 10644 12486 10646 12538
rect 10826 12486 10828 12538
rect 10582 12484 10588 12486
rect 10644 12484 10668 12486
rect 10724 12484 10748 12486
rect 10804 12484 10828 12486
rect 10884 12484 10890 12486
rect 10582 12464 10890 12484
rect 11348 12238 11376 13126
rect 12912 12442 12940 15982
rect 13004 15366 13032 17478
rect 14002 17368 14058 17377
rect 14002 17303 14058 17312
rect 14016 17066 14044 17303
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 14108 16998 14136 17711
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 13096 16590 13124 16934
rect 14108 16794 14136 16934
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 13004 12646 13032 15302
rect 13636 15156 13688 15162
rect 13636 15098 13688 15104
rect 13648 13870 13676 15098
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13740 13938 13768 14214
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 14200 13530 14228 18770
rect 14292 17202 14320 19615
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14384 17066 14412 18022
rect 14372 17060 14424 17066
rect 14372 17002 14424 17008
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14292 14618 14320 15642
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 12912 12238 12940 12378
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 1504 11801 1532 12038
rect 1490 11792 1546 11801
rect 1490 11727 1546 11736
rect 10582 11452 10890 11472
rect 10582 11450 10588 11452
rect 10644 11450 10668 11452
rect 10724 11450 10748 11452
rect 10804 11450 10828 11452
rect 10884 11450 10890 11452
rect 10644 11398 10646 11450
rect 10826 11398 10828 11450
rect 10582 11396 10588 11398
rect 10644 11396 10668 11398
rect 10724 11396 10748 11398
rect 10804 11396 10828 11398
rect 10884 11396 10890 11398
rect 10582 11376 10890 11396
rect 11072 10674 11100 12038
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 1492 10464 1544 10470
rect 1492 10406 1544 10412
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 1504 10169 1532 10406
rect 10582 10364 10890 10384
rect 10582 10362 10588 10364
rect 10644 10362 10668 10364
rect 10724 10362 10748 10364
rect 10804 10362 10828 10364
rect 10884 10362 10890 10364
rect 10644 10310 10646 10362
rect 10826 10310 10828 10362
rect 10582 10308 10588 10310
rect 10644 10308 10668 10310
rect 10724 10308 10748 10310
rect 10804 10308 10828 10310
rect 10884 10308 10890 10310
rect 10582 10288 10890 10308
rect 1490 10160 1546 10169
rect 1490 10095 1546 10104
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1504 8673 1532 8774
rect 1490 8664 1546 8673
rect 1490 8599 1546 8608
rect 8680 7410 8708 9318
rect 10582 9276 10890 9296
rect 10582 9274 10588 9276
rect 10644 9274 10668 9276
rect 10724 9274 10748 9276
rect 10804 9274 10828 9276
rect 10884 9274 10890 9276
rect 10644 9222 10646 9274
rect 10826 9222 10828 9274
rect 10582 9220 10588 9222
rect 10644 9220 10668 9222
rect 10724 9220 10748 9222
rect 10804 9220 10828 9222
rect 10884 9220 10890 9222
rect 10582 9200 10890 9220
rect 11532 8974 11560 10406
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 10582 8188 10890 8208
rect 10582 8186 10588 8188
rect 10644 8186 10668 8188
rect 10724 8186 10748 8188
rect 10804 8186 10828 8188
rect 10884 8186 10890 8188
rect 10644 8134 10646 8186
rect 10826 8134 10828 8186
rect 10582 8132 10588 8134
rect 10644 8132 10668 8134
rect 10724 8132 10748 8134
rect 10804 8132 10828 8134
rect 10884 8132 10890 8134
rect 10582 8112 10890 8132
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 7041 1532 7142
rect 10582 7100 10890 7120
rect 10582 7098 10588 7100
rect 10644 7098 10668 7100
rect 10724 7098 10748 7100
rect 10804 7098 10828 7100
rect 10884 7098 10890 7100
rect 10644 7046 10646 7098
rect 10826 7046 10828 7098
rect 10582 7044 10588 7046
rect 10644 7044 10668 7046
rect 10724 7044 10748 7046
rect 10804 7044 10828 7046
rect 10884 7044 10890 7046
rect 1490 7032 1546 7041
rect 10582 7024 10890 7044
rect 1490 6967 1546 6976
rect 13004 6914 13032 12582
rect 12912 6886 13032 6914
rect 10582 6012 10890 6032
rect 10582 6010 10588 6012
rect 10644 6010 10668 6012
rect 10724 6010 10748 6012
rect 10804 6010 10828 6012
rect 10884 6010 10890 6012
rect 10644 5958 10646 6010
rect 10826 5958 10828 6010
rect 10582 5956 10588 5958
rect 10644 5956 10668 5958
rect 10724 5956 10748 5958
rect 10804 5956 10828 5958
rect 10884 5956 10890 5958
rect 10582 5936 10890 5956
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 8852 5568 8904 5574
rect 8852 5510 8904 5516
rect 1504 5409 1532 5510
rect 1490 5400 1546 5409
rect 1490 5335 1546 5344
rect 1492 3936 1544 3942
rect 1490 3904 1492 3913
rect 1544 3904 1546 3913
rect 1490 3839 1546 3848
rect 8864 3058 8892 5510
rect 10582 4924 10890 4944
rect 10582 4922 10588 4924
rect 10644 4922 10668 4924
rect 10724 4922 10748 4924
rect 10804 4922 10828 4924
rect 10884 4922 10890 4924
rect 10644 4870 10646 4922
rect 10826 4870 10828 4922
rect 10582 4868 10588 4870
rect 10644 4868 10668 4870
rect 10724 4868 10748 4870
rect 10804 4868 10828 4870
rect 10884 4868 10890 4870
rect 10582 4848 10890 4868
rect 10582 3836 10890 3856
rect 10582 3834 10588 3836
rect 10644 3834 10668 3836
rect 10724 3834 10748 3836
rect 10804 3834 10828 3836
rect 10884 3834 10890 3836
rect 10644 3782 10646 3834
rect 10826 3782 10828 3834
rect 10582 3780 10588 3782
rect 10644 3780 10668 3782
rect 10724 3780 10748 3782
rect 10804 3780 10828 3782
rect 10884 3780 10890 3782
rect 10582 3760 10890 3780
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1412 2281 1440 2790
rect 10582 2748 10890 2768
rect 10582 2746 10588 2748
rect 10644 2746 10668 2748
rect 10724 2746 10748 2748
rect 10804 2746 10828 2748
rect 10884 2746 10890 2748
rect 10644 2694 10646 2746
rect 10826 2694 10828 2746
rect 10582 2692 10588 2694
rect 10644 2692 10668 2694
rect 10724 2692 10748 2694
rect 10804 2692 10828 2694
rect 10884 2692 10890 2694
rect 10582 2672 10890 2692
rect 12912 2582 12940 6886
rect 14384 4729 14412 17002
rect 14476 14074 14504 21519
rect 14568 18834 14596 28319
rect 14648 28144 14700 28150
rect 14648 28086 14700 28092
rect 14556 18828 14608 18834
rect 14556 18770 14608 18776
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14464 7812 14516 7818
rect 14464 7754 14516 7760
rect 14476 5778 14504 7754
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14370 4720 14426 4729
rect 14370 4655 14426 4664
rect 12900 2576 12952 2582
rect 12900 2518 12952 2524
rect 1492 2304 1544 2310
rect 1398 2272 1454 2281
rect 1492 2246 1544 2252
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 1398 2207 1454 2216
rect 1504 785 1532 2246
rect 6012 800 6040 2246
rect 14568 2009 14596 17818
rect 14660 16998 14688 28086
rect 14752 17377 14780 28591
rect 14844 22094 14872 28727
rect 17224 28212 17276 28218
rect 17224 28154 17276 28160
rect 15198 25528 15254 25537
rect 15198 25463 15254 25472
rect 14844 22066 14964 22094
rect 14832 19712 14884 19718
rect 14832 19654 14884 19660
rect 14844 19417 14872 19654
rect 14830 19408 14886 19417
rect 14830 19343 14886 19352
rect 14738 17368 14794 17377
rect 14738 17303 14794 17312
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14660 16794 14688 16934
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14660 16454 14688 16730
rect 14844 16658 14872 17070
rect 14936 16794 14964 22066
rect 15016 21888 15068 21894
rect 15016 21830 15068 21836
rect 15028 20262 15056 21830
rect 15108 20868 15160 20874
rect 15108 20810 15160 20816
rect 15016 20256 15068 20262
rect 15016 20198 15068 20204
rect 15120 19854 15148 20810
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 15212 19310 15240 25463
rect 17130 25392 17186 25401
rect 17130 25327 17186 25336
rect 16578 24848 16634 24857
rect 16578 24783 16634 24792
rect 16486 23488 16542 23497
rect 16486 23423 16542 23432
rect 16120 21684 16172 21690
rect 16120 21626 16172 21632
rect 15752 21616 15804 21622
rect 15752 21558 15804 21564
rect 15764 21146 15792 21558
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 15566 20360 15622 20369
rect 15566 20295 15568 20304
rect 15620 20295 15622 20304
rect 15568 20266 15620 20272
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 15028 18737 15056 19110
rect 15014 18728 15070 18737
rect 15014 18663 15070 18672
rect 15014 18456 15070 18465
rect 15014 18391 15070 18400
rect 15028 18086 15056 18391
rect 15212 18290 15240 19246
rect 15764 18970 15792 21082
rect 16132 20602 16160 21626
rect 16120 20596 16172 20602
rect 16120 20538 16172 20544
rect 16396 19848 16448 19854
rect 16396 19790 16448 19796
rect 16212 19712 16264 19718
rect 16212 19654 16264 19660
rect 16224 19145 16252 19654
rect 16210 19136 16266 19145
rect 16210 19071 16266 19080
rect 15752 18964 15804 18970
rect 15752 18906 15804 18912
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 15660 18828 15712 18834
rect 15660 18770 15712 18776
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 15016 18080 15068 18086
rect 15016 18022 15068 18028
rect 14924 16788 14976 16794
rect 14924 16730 14976 16736
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14752 11558 14780 13806
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14844 5137 14872 16594
rect 14936 16425 14964 16730
rect 14922 16416 14978 16425
rect 14922 16351 14978 16360
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14936 10606 14964 14214
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 15028 6914 15056 18022
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15304 16697 15332 16934
rect 15382 16824 15438 16833
rect 15382 16759 15384 16768
rect 15436 16759 15438 16768
rect 15384 16730 15436 16736
rect 15290 16688 15346 16697
rect 15290 16623 15346 16632
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 15212 16250 15240 16458
rect 15200 16244 15252 16250
rect 15200 16186 15252 16192
rect 15200 15972 15252 15978
rect 15200 15914 15252 15920
rect 15108 15904 15160 15910
rect 15106 15872 15108 15881
rect 15160 15872 15162 15881
rect 15106 15807 15162 15816
rect 15212 15706 15240 15914
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15198 15464 15254 15473
rect 15108 15428 15160 15434
rect 15198 15399 15254 15408
rect 15108 15370 15160 15376
rect 15120 14385 15148 15370
rect 15212 15162 15240 15399
rect 15382 15192 15438 15201
rect 15200 15156 15252 15162
rect 15382 15127 15438 15136
rect 15200 15098 15252 15104
rect 15396 14618 15424 15127
rect 15488 14618 15516 18566
rect 15672 17513 15700 18770
rect 15934 18048 15990 18057
rect 15934 17983 15990 17992
rect 15948 17882 15976 17983
rect 16132 17882 16160 18906
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 15658 17504 15714 17513
rect 15658 17439 15714 17448
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 15844 16584 15896 16590
rect 15842 16552 15844 16561
rect 15896 16552 15898 16561
rect 15752 16516 15804 16522
rect 15842 16487 15898 16496
rect 15752 16458 15804 16464
rect 15568 16176 15620 16182
rect 15566 16144 15568 16153
rect 15620 16144 15622 16153
rect 15566 16079 15622 16088
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15106 14376 15162 14385
rect 15106 14311 15162 14320
rect 15108 14068 15160 14074
rect 15108 14010 15160 14016
rect 14936 6886 15056 6914
rect 14936 5302 14964 6886
rect 14924 5296 14976 5302
rect 14924 5238 14976 5244
rect 14830 5128 14886 5137
rect 14830 5063 14886 5072
rect 15120 4593 15148 14010
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15304 7478 15332 7686
rect 15292 7472 15344 7478
rect 15292 7414 15344 7420
rect 15106 4584 15162 4593
rect 15106 4519 15162 4528
rect 15396 3505 15424 14554
rect 15488 12782 15516 14554
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15580 12434 15608 16079
rect 15658 16008 15714 16017
rect 15658 15943 15714 15952
rect 15672 15706 15700 15943
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15488 12406 15608 12434
rect 15488 5273 15516 12406
rect 15672 6914 15700 15506
rect 15764 11898 15792 16458
rect 15856 15638 15884 16487
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 15948 12073 15976 16934
rect 16040 16590 16068 17274
rect 16118 17096 16174 17105
rect 16118 17031 16174 17040
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 16132 16046 16160 17031
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16132 14958 16160 15846
rect 16224 15570 16252 19071
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 16408 18578 16436 19790
rect 16500 19009 16528 23423
rect 16592 20058 16620 24783
rect 16946 23352 17002 23361
rect 16946 23287 17002 23296
rect 16670 21312 16726 21321
rect 16670 21247 16726 21256
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16486 19000 16542 19009
rect 16486 18935 16542 18944
rect 16500 18902 16528 18935
rect 16488 18896 16540 18902
rect 16488 18838 16540 18844
rect 16592 18766 16620 19994
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16316 17649 16344 18566
rect 16408 18550 16528 18578
rect 16500 18086 16528 18550
rect 16578 18320 16634 18329
rect 16684 18290 16712 21247
rect 16764 21140 16816 21146
rect 16764 21082 16816 21088
rect 16776 20806 16804 21082
rect 16856 21004 16908 21010
rect 16856 20946 16908 20952
rect 16764 20800 16816 20806
rect 16764 20742 16816 20748
rect 16762 19272 16818 19281
rect 16762 19207 16764 19216
rect 16816 19207 16818 19216
rect 16764 19178 16816 19184
rect 16578 18255 16634 18264
rect 16672 18284 16724 18290
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16500 17678 16528 18022
rect 16592 17762 16620 18255
rect 16776 18272 16804 19178
rect 16868 18340 16896 20946
rect 16960 18630 16988 23287
rect 17038 21040 17094 21049
rect 17038 20975 17094 20984
rect 17052 20602 17080 20975
rect 17040 20596 17092 20602
rect 17040 20538 17092 20544
rect 17052 18902 17080 20538
rect 17144 18970 17172 25327
rect 17236 19310 17264 28154
rect 17408 26784 17460 26790
rect 17408 26726 17460 26732
rect 17420 20806 17448 26726
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 17880 21010 17908 21490
rect 17972 21146 18000 22714
rect 18052 21888 18104 21894
rect 18052 21830 18104 21836
rect 17960 21140 18012 21146
rect 17960 21082 18012 21088
rect 18064 21078 18092 21830
rect 18340 21486 18368 29543
rect 18970 29200 19026 30000
rect 19890 29336 19946 29345
rect 19890 29271 19946 29280
rect 18788 28076 18840 28082
rect 18788 28018 18840 28024
rect 18420 27396 18472 27402
rect 18420 27338 18472 27344
rect 18432 22094 18460 27338
rect 18604 23860 18656 23866
rect 18604 23802 18656 23808
rect 18432 22066 18552 22094
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 18052 21072 18104 21078
rect 18052 21014 18104 21020
rect 17868 21004 17920 21010
rect 17868 20946 17920 20952
rect 17684 20936 17736 20942
rect 17684 20878 17736 20884
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17408 20256 17460 20262
rect 17408 20198 17460 20204
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 17040 18896 17092 18902
rect 17040 18838 17092 18844
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 17236 18442 17264 19246
rect 17314 19000 17370 19009
rect 17314 18935 17370 18944
rect 17328 18834 17356 18935
rect 17420 18834 17448 20198
rect 17604 19122 17632 20402
rect 17696 19281 17724 20878
rect 17776 20800 17828 20806
rect 17776 20742 17828 20748
rect 17788 19378 17816 20742
rect 17958 20496 18014 20505
rect 17958 20431 18014 20440
rect 17868 19712 17920 19718
rect 17868 19654 17920 19660
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17682 19272 17738 19281
rect 17682 19207 17738 19216
rect 17604 19094 17724 19122
rect 17590 19000 17646 19009
rect 17590 18935 17592 18944
rect 17644 18935 17646 18944
rect 17592 18906 17644 18912
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 17408 18828 17460 18834
rect 17408 18770 17460 18776
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 17314 18728 17370 18737
rect 17408 18692 17460 18698
rect 17370 18672 17408 18680
rect 17314 18663 17408 18672
rect 17328 18652 17408 18663
rect 17408 18634 17460 18640
rect 17236 18414 17448 18442
rect 17316 18352 17368 18358
rect 16868 18312 16988 18340
rect 16960 18306 16988 18312
rect 17144 18312 17316 18340
rect 17144 18306 17172 18312
rect 16960 18278 17172 18306
rect 17316 18294 17368 18300
rect 17420 18290 17448 18414
rect 16776 18244 16896 18272
rect 16672 18226 16724 18232
rect 16762 18184 16818 18193
rect 16762 18119 16764 18128
rect 16816 18119 16818 18128
rect 16764 18090 16816 18096
rect 16868 17762 16896 18244
rect 16592 17734 16804 17762
rect 16868 17734 16988 17762
rect 16396 17672 16448 17678
rect 16302 17640 16358 17649
rect 16396 17614 16448 17620
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 16302 17575 16358 17584
rect 16408 17241 16436 17614
rect 16394 17232 16450 17241
rect 16394 17167 16450 17176
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16304 16584 16356 16590
rect 16304 16526 16356 16532
rect 16316 15910 16344 16526
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16210 15464 16266 15473
rect 16210 15399 16266 15408
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 15934 12064 15990 12073
rect 15934 11999 15990 12008
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 16224 6914 16252 15399
rect 16316 12170 16344 15846
rect 16408 14278 16436 16934
rect 16500 16590 16528 17614
rect 16684 16946 16712 17614
rect 16592 16918 16712 16946
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16408 14006 16436 14214
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 16500 12345 16528 14010
rect 16486 12336 16542 12345
rect 16486 12271 16542 12280
rect 16304 12164 16356 12170
rect 16304 12106 16356 12112
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 15672 6886 15792 6914
rect 15764 6186 15792 6886
rect 16132 6886 16252 6914
rect 15752 6180 15804 6186
rect 15752 6122 15804 6128
rect 15474 5264 15530 5273
rect 15474 5199 15530 5208
rect 16132 4146 16160 6886
rect 16316 6798 16344 11834
rect 16592 11121 16620 16918
rect 16776 16810 16804 17734
rect 16960 17610 16988 17734
rect 16856 17604 16908 17610
rect 16856 17546 16908 17552
rect 16948 17604 17000 17610
rect 16948 17546 17000 17552
rect 16868 17202 16896 17546
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16684 16794 16804 16810
rect 16672 16788 16804 16794
rect 16724 16782 16804 16788
rect 16672 16730 16724 16736
rect 16764 16720 16816 16726
rect 16764 16662 16816 16668
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16684 14074 16712 16594
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16776 13530 16804 16662
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16578 11112 16634 11121
rect 16578 11047 16634 11056
rect 16868 8906 16896 17138
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 16960 9489 16988 16662
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 17052 11014 17080 16050
rect 17144 13462 17172 18278
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 17316 18216 17368 18222
rect 17316 18158 17368 18164
rect 17328 17921 17356 18158
rect 17604 18154 17632 18770
rect 17696 18306 17724 19094
rect 17880 18714 17908 19654
rect 17972 19310 18000 20431
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 18064 19961 18092 20198
rect 18234 20088 18290 20097
rect 18234 20023 18290 20032
rect 18050 19952 18106 19961
rect 18050 19887 18106 19896
rect 18248 19446 18276 20023
rect 18236 19440 18288 19446
rect 18236 19382 18288 19388
rect 18340 19378 18368 21422
rect 18524 20330 18552 22066
rect 18512 20324 18564 20330
rect 18512 20266 18564 20272
rect 18512 19780 18564 19786
rect 18512 19722 18564 19728
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 17960 19304 18012 19310
rect 18524 19258 18552 19722
rect 17960 19246 18012 19252
rect 18340 19230 18552 19258
rect 18234 19136 18290 19145
rect 18234 19071 18290 19080
rect 18142 19000 18198 19009
rect 18142 18935 18198 18944
rect 18052 18896 18104 18902
rect 18052 18838 18104 18844
rect 17880 18686 18000 18714
rect 17696 18278 17908 18306
rect 17776 18216 17828 18222
rect 17696 18176 17776 18204
rect 17592 18148 17644 18154
rect 17592 18090 17644 18096
rect 17314 17912 17370 17921
rect 17314 17847 17370 17856
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 17328 16250 17356 16526
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17314 15736 17370 15745
rect 17314 15671 17370 15680
rect 17328 15366 17356 15671
rect 17316 15360 17368 15366
rect 17314 15328 17316 15337
rect 17368 15328 17370 15337
rect 17314 15263 17370 15272
rect 17314 15056 17370 15065
rect 17314 14991 17316 15000
rect 17368 14991 17370 15000
rect 17316 14962 17368 14968
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17132 13456 17184 13462
rect 17132 13398 17184 13404
rect 17236 11694 17264 14826
rect 17328 14657 17356 14962
rect 17314 14648 17370 14657
rect 17314 14583 17370 14592
rect 17420 11801 17448 17682
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17500 17060 17552 17066
rect 17500 17002 17552 17008
rect 17512 16697 17540 17002
rect 17498 16688 17554 16697
rect 17498 16623 17554 16632
rect 17604 13734 17632 17614
rect 17696 16046 17724 18176
rect 17776 18158 17828 18164
rect 17776 16176 17828 16182
rect 17776 16118 17828 16124
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17696 15094 17724 15438
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 17592 13728 17644 13734
rect 17696 13705 17724 15030
rect 17788 14074 17816 16118
rect 17880 16114 17908 18278
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17880 15910 17908 16050
rect 17868 15904 17920 15910
rect 17972 15881 18000 18686
rect 18064 18290 18092 18838
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 18156 18086 18184 18935
rect 18248 18737 18276 19071
rect 18340 18766 18368 19230
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 18328 18760 18380 18766
rect 18234 18728 18290 18737
rect 18432 18748 18460 19110
rect 18432 18720 18552 18748
rect 18328 18702 18380 18708
rect 18234 18663 18290 18672
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 17868 15846 17920 15852
rect 17958 15872 18014 15881
rect 17958 15807 18014 15816
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17592 13670 17644 13676
rect 17682 13696 17738 13705
rect 17682 13631 17738 13640
rect 17880 12889 17908 15302
rect 18064 15094 18092 17818
rect 18156 17814 18184 18022
rect 18144 17808 18196 17814
rect 18144 17750 18196 17756
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 18156 15337 18184 15846
rect 18142 15328 18198 15337
rect 18142 15263 18198 15272
rect 18052 15088 18104 15094
rect 18052 15030 18104 15036
rect 17958 14784 18014 14793
rect 17958 14719 18014 14728
rect 17972 14006 18000 14719
rect 17960 14000 18012 14006
rect 17960 13942 18012 13948
rect 18064 13326 18092 15030
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 17960 12912 18012 12918
rect 17866 12880 17922 12889
rect 17960 12854 18012 12860
rect 17866 12815 17922 12824
rect 17406 11792 17462 11801
rect 17406 11727 17462 11736
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 16946 9480 17002 9489
rect 16946 9415 17002 9424
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 15382 3496 15438 3505
rect 15382 3431 15438 3440
rect 17972 2582 18000 12854
rect 18156 12102 18184 14962
rect 18248 12617 18276 18566
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 18340 15570 18368 18022
rect 18432 17513 18460 18294
rect 18524 18290 18552 18720
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18418 17504 18474 17513
rect 18418 17439 18474 17448
rect 18524 17218 18552 18022
rect 18616 17882 18644 23802
rect 18800 22094 18828 28018
rect 18984 26246 19012 29200
rect 19064 28008 19116 28014
rect 19064 27950 19116 27956
rect 18972 26240 19024 26246
rect 18972 26182 19024 26188
rect 18708 22066 18828 22094
rect 18708 21350 18736 22066
rect 18696 21344 18748 21350
rect 18696 21286 18748 21292
rect 18708 19174 18736 21286
rect 18788 20596 18840 20602
rect 18788 20538 18840 20544
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18694 19000 18750 19009
rect 18694 18935 18750 18944
rect 18708 18766 18736 18935
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18604 17876 18656 17882
rect 18604 17818 18656 17824
rect 18800 17678 18828 20538
rect 18880 20256 18932 20262
rect 18880 20198 18932 20204
rect 18970 20224 19026 20233
rect 18892 19689 18920 20198
rect 18970 20159 19026 20168
rect 18984 20058 19012 20159
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 18878 19680 18934 19689
rect 18878 19615 18934 19624
rect 18892 19378 18920 19615
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18984 19281 19012 19994
rect 19076 19553 19104 27950
rect 19524 27464 19576 27470
rect 19524 27406 19576 27412
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19352 26246 19380 27270
rect 19536 27130 19564 27406
rect 19524 27124 19576 27130
rect 19524 27066 19576 27072
rect 19340 26240 19392 26246
rect 19340 26182 19392 26188
rect 19800 24744 19852 24750
rect 19800 24686 19852 24692
rect 19248 24336 19300 24342
rect 19248 24278 19300 24284
rect 19260 23254 19288 24278
rect 19340 23316 19392 23322
rect 19340 23258 19392 23264
rect 19248 23248 19300 23254
rect 19248 23190 19300 23196
rect 19260 22778 19288 23190
rect 19248 22772 19300 22778
rect 19248 22714 19300 22720
rect 19154 22672 19210 22681
rect 19154 22607 19210 22616
rect 19168 19990 19196 22607
rect 19248 22568 19300 22574
rect 19248 22510 19300 22516
rect 19156 19984 19208 19990
rect 19156 19926 19208 19932
rect 19062 19544 19118 19553
rect 19062 19479 19118 19488
rect 19260 19334 19288 22510
rect 19352 22098 19380 23258
rect 19524 22160 19576 22166
rect 19524 22102 19576 22108
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19352 21690 19380 22034
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 19340 21072 19392 21078
rect 19340 21014 19392 21020
rect 19168 19310 19288 19334
rect 19352 19310 19380 21014
rect 19444 19922 19472 21830
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19430 19816 19486 19825
rect 19430 19751 19432 19760
rect 19484 19751 19486 19760
rect 19432 19722 19484 19728
rect 19536 19666 19564 22102
rect 19616 21616 19668 21622
rect 19616 21558 19668 21564
rect 19444 19638 19564 19666
rect 19444 19446 19472 19638
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19156 19306 19288 19310
rect 19156 19304 19208 19306
rect 18970 19272 19026 19281
rect 19156 19246 19208 19252
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 18970 19207 19026 19216
rect 18878 19136 18934 19145
rect 18878 19071 18934 19080
rect 18892 18222 18920 19071
rect 18984 18290 19012 19207
rect 19156 19168 19208 19174
rect 19156 19110 19208 19116
rect 19168 18601 19196 19110
rect 19248 18896 19300 18902
rect 19248 18838 19300 18844
rect 19260 18698 19288 18838
rect 19444 18766 19472 19382
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19248 18692 19300 18698
rect 19248 18634 19300 18640
rect 19444 18601 19472 18702
rect 19154 18592 19210 18601
rect 19154 18527 19210 18536
rect 19430 18592 19486 18601
rect 19430 18527 19486 18536
rect 19338 18456 19394 18465
rect 19338 18391 19394 18400
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 18984 17954 19012 18226
rect 18984 17926 19104 17954
rect 19076 17746 19104 17926
rect 19154 17776 19210 17785
rect 19064 17740 19116 17746
rect 19154 17711 19210 17720
rect 19064 17682 19116 17688
rect 18788 17672 18840 17678
rect 18602 17640 18658 17649
rect 18788 17614 18840 17620
rect 18602 17575 18658 17584
rect 18616 17542 18644 17575
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18972 17264 19024 17270
rect 18524 17190 18644 17218
rect 18972 17206 19024 17212
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18328 15564 18380 15570
rect 18328 15506 18380 15512
rect 18432 15366 18460 16050
rect 18512 15428 18564 15434
rect 18512 15370 18564 15376
rect 18420 15360 18472 15366
rect 18420 15302 18472 15308
rect 18328 14340 18380 14346
rect 18328 14282 18380 14288
rect 18340 14074 18368 14282
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18328 13252 18380 13258
rect 18328 13194 18380 13200
rect 18234 12608 18290 12617
rect 18234 12543 18290 12552
rect 18340 12434 18368 13194
rect 18432 13190 18460 15302
rect 18524 15162 18552 15370
rect 18512 15156 18564 15162
rect 18512 15098 18564 15104
rect 18510 13288 18566 13297
rect 18510 13223 18566 13232
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18432 12850 18460 13126
rect 18524 12986 18552 13223
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18340 12406 18460 12434
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18156 7993 18184 12038
rect 18432 9654 18460 12406
rect 18616 10033 18644 17190
rect 18788 17128 18840 17134
rect 18788 17070 18840 17076
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18696 16992 18748 16998
rect 18694 16960 18696 16969
rect 18748 16960 18750 16969
rect 18694 16895 18750 16904
rect 18800 16833 18828 17070
rect 18786 16824 18842 16833
rect 18786 16759 18842 16768
rect 18696 16720 18748 16726
rect 18694 16688 18696 16697
rect 18748 16688 18750 16697
rect 18694 16623 18750 16632
rect 18694 16552 18750 16561
rect 18694 16487 18750 16496
rect 18708 16046 18736 16487
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18708 12442 18736 15982
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18602 10024 18658 10033
rect 18602 9959 18658 9968
rect 18420 9648 18472 9654
rect 18420 9590 18472 9596
rect 18142 7984 18198 7993
rect 18142 7919 18198 7928
rect 18800 6914 18828 16759
rect 18892 16726 18920 17070
rect 18880 16720 18932 16726
rect 18880 16662 18932 16668
rect 18892 16454 18920 16662
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18880 16176 18932 16182
rect 18880 16118 18932 16124
rect 18892 14890 18920 16118
rect 18984 14890 19012 17206
rect 19064 17196 19116 17202
rect 19064 17138 19116 17144
rect 19076 16182 19104 17138
rect 19168 17134 19196 17711
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 19154 16824 19210 16833
rect 19154 16759 19210 16768
rect 19064 16176 19116 16182
rect 19064 16118 19116 16124
rect 19168 16046 19196 16759
rect 19156 16040 19208 16046
rect 19156 15982 19208 15988
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 19064 15020 19116 15026
rect 19064 14962 19116 14968
rect 19076 14929 19104 14962
rect 19062 14920 19118 14929
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18972 14884 19024 14890
rect 19062 14855 19118 14864
rect 18972 14826 19024 14832
rect 19076 14550 19104 14855
rect 19064 14544 19116 14550
rect 19062 14512 19064 14521
rect 19116 14512 19118 14521
rect 19062 14447 19118 14456
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 19076 13841 19104 14214
rect 19062 13832 19118 13841
rect 19062 13767 19118 13776
rect 19062 13696 19118 13705
rect 19062 13631 19118 13640
rect 19076 13433 19104 13631
rect 19062 13424 19118 13433
rect 19168 13394 19196 15846
rect 19260 15162 19288 17546
rect 19352 17270 19380 18391
rect 19432 17808 19484 17814
rect 19432 17750 19484 17756
rect 19444 17678 19472 17750
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19444 17270 19472 17614
rect 19340 17264 19392 17270
rect 19340 17206 19392 17212
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 19444 16794 19472 17070
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19444 16674 19472 16730
rect 19352 16658 19472 16674
rect 19340 16652 19472 16658
rect 19392 16646 19472 16652
rect 19340 16594 19392 16600
rect 19340 16516 19392 16522
rect 19392 16476 19472 16504
rect 19340 16458 19392 16464
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 19248 15020 19300 15026
rect 19248 14962 19300 14968
rect 19260 14550 19288 14962
rect 19340 14884 19392 14890
rect 19340 14826 19392 14832
rect 19248 14544 19300 14550
rect 19248 14486 19300 14492
rect 19352 14278 19380 14826
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19338 13968 19394 13977
rect 19338 13903 19394 13912
rect 19352 13818 19380 13903
rect 19260 13790 19380 13818
rect 19062 13359 19118 13368
rect 19156 13388 19208 13394
rect 19076 12434 19104 13359
rect 19156 13330 19208 13336
rect 19260 12918 19288 13790
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19248 12912 19300 12918
rect 19248 12854 19300 12860
rect 19076 12406 19196 12434
rect 19064 11552 19116 11558
rect 19064 11494 19116 11500
rect 19076 11354 19104 11494
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 18432 6886 18828 6914
rect 19168 6914 19196 12406
rect 19352 11626 19380 13466
rect 19444 12306 19472 16476
rect 19536 15065 19564 19314
rect 19628 18290 19656 21558
rect 19706 20904 19762 20913
rect 19706 20839 19762 20848
rect 19720 20806 19748 20839
rect 19708 20800 19760 20806
rect 19708 20742 19760 20748
rect 19616 18284 19668 18290
rect 19616 18226 19668 18232
rect 19616 18148 19668 18154
rect 19616 18090 19668 18096
rect 19628 17746 19656 18090
rect 19616 17740 19668 17746
rect 19616 17682 19668 17688
rect 19628 17134 19656 17682
rect 19720 17592 19748 20742
rect 19812 20618 19840 24686
rect 19904 22710 19932 29271
rect 24490 29200 24546 30000
rect 29918 29322 29974 30000
rect 34978 29744 35034 29753
rect 34978 29679 35034 29688
rect 34610 29608 34666 29617
rect 34610 29543 34666 29552
rect 29918 29294 30236 29322
rect 29918 29200 29974 29294
rect 24214 28520 24270 28529
rect 24214 28455 24270 28464
rect 23940 27940 23992 27946
rect 23940 27882 23992 27888
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 19996 26858 20024 27406
rect 20628 27396 20680 27402
rect 20628 27338 20680 27344
rect 20214 27228 20522 27248
rect 20214 27226 20220 27228
rect 20276 27226 20300 27228
rect 20356 27226 20380 27228
rect 20436 27226 20460 27228
rect 20516 27226 20522 27228
rect 20276 27174 20278 27226
rect 20458 27174 20460 27226
rect 20214 27172 20220 27174
rect 20276 27172 20300 27174
rect 20356 27172 20380 27174
rect 20436 27172 20460 27174
rect 20516 27172 20522 27174
rect 20214 27152 20522 27172
rect 19984 26852 20036 26858
rect 19984 26794 20036 26800
rect 20074 26480 20130 26489
rect 20074 26415 20130 26424
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 19892 22704 19944 22710
rect 19892 22646 19944 22652
rect 19904 22137 19932 22646
rect 19996 22438 20024 23734
rect 20088 22778 20116 26415
rect 20214 26140 20522 26160
rect 20214 26138 20220 26140
rect 20276 26138 20300 26140
rect 20356 26138 20380 26140
rect 20436 26138 20460 26140
rect 20516 26138 20522 26140
rect 20276 26086 20278 26138
rect 20458 26086 20460 26138
rect 20214 26084 20220 26086
rect 20276 26084 20300 26086
rect 20356 26084 20380 26086
rect 20436 26084 20460 26086
rect 20516 26084 20522 26086
rect 20214 26064 20522 26084
rect 20214 25052 20522 25072
rect 20214 25050 20220 25052
rect 20276 25050 20300 25052
rect 20356 25050 20380 25052
rect 20436 25050 20460 25052
rect 20516 25050 20522 25052
rect 20276 24998 20278 25050
rect 20458 24998 20460 25050
rect 20214 24996 20220 24998
rect 20276 24996 20300 24998
rect 20356 24996 20380 24998
rect 20436 24996 20460 24998
rect 20516 24996 20522 24998
rect 20214 24976 20522 24996
rect 20214 23964 20522 23984
rect 20214 23962 20220 23964
rect 20276 23962 20300 23964
rect 20356 23962 20380 23964
rect 20436 23962 20460 23964
rect 20516 23962 20522 23964
rect 20276 23910 20278 23962
rect 20458 23910 20460 23962
rect 20214 23908 20220 23910
rect 20276 23908 20300 23910
rect 20356 23908 20380 23910
rect 20436 23908 20460 23910
rect 20516 23908 20522 23910
rect 20214 23888 20522 23908
rect 20536 23656 20588 23662
rect 20536 23598 20588 23604
rect 20548 23225 20576 23598
rect 20534 23216 20590 23225
rect 20534 23151 20590 23160
rect 20214 22876 20522 22896
rect 20214 22874 20220 22876
rect 20276 22874 20300 22876
rect 20356 22874 20380 22876
rect 20436 22874 20460 22876
rect 20516 22874 20522 22876
rect 20276 22822 20278 22874
rect 20458 22822 20460 22874
rect 20214 22820 20220 22822
rect 20276 22820 20300 22822
rect 20356 22820 20380 22822
rect 20436 22820 20460 22822
rect 20516 22820 20522 22822
rect 20214 22800 20522 22820
rect 20076 22772 20128 22778
rect 20076 22714 20128 22720
rect 19984 22432 20036 22438
rect 19984 22374 20036 22380
rect 19890 22128 19946 22137
rect 19890 22063 19946 22072
rect 19996 21622 20024 22374
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 19984 21412 20036 21418
rect 19984 21354 20036 21360
rect 19812 20590 19932 20618
rect 19800 20528 19852 20534
rect 19798 20496 19800 20505
rect 19852 20496 19854 20505
rect 19798 20431 19854 20440
rect 19904 19428 19932 20590
rect 19996 20058 20024 21354
rect 20088 21162 20116 21830
rect 20214 21788 20522 21808
rect 20214 21786 20220 21788
rect 20276 21786 20300 21788
rect 20356 21786 20380 21788
rect 20436 21786 20460 21788
rect 20516 21786 20522 21788
rect 20276 21734 20278 21786
rect 20458 21734 20460 21786
rect 20214 21732 20220 21734
rect 20276 21732 20300 21734
rect 20356 21732 20380 21734
rect 20436 21732 20460 21734
rect 20516 21732 20522 21734
rect 20214 21712 20522 21732
rect 20640 21729 20668 27338
rect 21916 26988 21968 26994
rect 21916 26930 21968 26936
rect 21822 25800 21878 25809
rect 21822 25735 21878 25744
rect 20720 25696 20772 25702
rect 20720 25638 20772 25644
rect 20732 23798 20760 25638
rect 21640 25424 21692 25430
rect 21640 25366 21692 25372
rect 21456 25288 21508 25294
rect 21456 25230 21508 25236
rect 21088 25220 21140 25226
rect 21088 25162 21140 25168
rect 20720 23792 20772 23798
rect 20720 23734 20772 23740
rect 21100 23633 21128 25162
rect 21362 23896 21418 23905
rect 21362 23831 21418 23840
rect 21086 23624 21142 23633
rect 21086 23559 21142 23568
rect 21272 23520 21324 23526
rect 21270 23488 21272 23497
rect 21324 23488 21326 23497
rect 21270 23423 21326 23432
rect 20812 22976 20864 22982
rect 20812 22918 20864 22924
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 20626 21720 20682 21729
rect 20732 21690 20760 22170
rect 20626 21655 20682 21664
rect 20720 21684 20772 21690
rect 20720 21626 20772 21632
rect 20628 21616 20680 21622
rect 20628 21558 20680 21564
rect 20166 21448 20222 21457
rect 20166 21383 20222 21392
rect 20180 21350 20208 21383
rect 20168 21344 20220 21350
rect 20168 21286 20220 21292
rect 20088 21134 20208 21162
rect 20076 21072 20128 21078
rect 20076 21014 20128 21020
rect 20088 20466 20116 21014
rect 20180 20942 20208 21134
rect 20168 20936 20220 20942
rect 20168 20878 20220 20884
rect 20214 20700 20522 20720
rect 20214 20698 20220 20700
rect 20276 20698 20300 20700
rect 20356 20698 20380 20700
rect 20436 20698 20460 20700
rect 20516 20698 20522 20700
rect 20276 20646 20278 20698
rect 20458 20646 20460 20698
rect 20214 20644 20220 20646
rect 20276 20644 20300 20646
rect 20356 20644 20380 20646
rect 20436 20644 20460 20646
rect 20516 20644 20522 20646
rect 20214 20624 20522 20644
rect 20640 20602 20668 21558
rect 20732 21350 20760 21626
rect 20720 21344 20772 21350
rect 20720 21286 20772 21292
rect 20824 20777 20852 22918
rect 21088 22772 21140 22778
rect 21088 22714 21140 22720
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20916 21593 20944 21830
rect 20902 21584 20958 21593
rect 20902 21519 20958 21528
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20810 20768 20866 20777
rect 20810 20703 20866 20712
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 20076 20324 20128 20330
rect 20076 20266 20128 20272
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 20088 19496 20116 20266
rect 20640 20244 20668 20538
rect 20824 20534 20852 20703
rect 20812 20528 20864 20534
rect 20812 20470 20864 20476
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 20640 20216 20760 20244
rect 20628 19916 20680 19922
rect 20628 19858 20680 19864
rect 20214 19612 20522 19632
rect 20214 19610 20220 19612
rect 20276 19610 20300 19612
rect 20356 19610 20380 19612
rect 20436 19610 20460 19612
rect 20516 19610 20522 19612
rect 20276 19558 20278 19610
rect 20458 19558 20460 19610
rect 20214 19556 20220 19558
rect 20276 19556 20300 19558
rect 20356 19556 20380 19558
rect 20436 19556 20460 19558
rect 20516 19556 20522 19558
rect 20214 19536 20522 19556
rect 20640 19496 20668 19858
rect 20732 19514 20760 20216
rect 20088 19468 20300 19496
rect 19984 19440 20036 19446
rect 19904 19400 19984 19428
rect 19984 19382 20036 19388
rect 19800 19304 19852 19310
rect 19800 19246 19852 19252
rect 19812 18154 19840 19246
rect 20272 19174 20300 19468
rect 20548 19468 20668 19496
rect 20720 19508 20772 19514
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20352 19304 20404 19310
rect 20350 19272 20352 19281
rect 20404 19272 20406 19281
rect 20350 19207 20406 19216
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20456 18970 20484 19382
rect 20548 19334 20576 19468
rect 20720 19450 20772 19456
rect 20548 19306 20668 19334
rect 20260 18964 20312 18970
rect 20260 18906 20312 18912
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 19892 18896 19944 18902
rect 19892 18838 19944 18844
rect 20272 18850 20300 18906
rect 20548 18850 20576 18906
rect 19800 18148 19852 18154
rect 19800 18090 19852 18096
rect 19904 17785 19932 18838
rect 19984 18828 20036 18834
rect 20272 18822 20576 18850
rect 20036 18788 20208 18816
rect 19984 18770 20036 18776
rect 20180 18714 20208 18788
rect 20352 18760 20404 18766
rect 20180 18708 20352 18714
rect 20180 18702 20404 18708
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20180 18686 20392 18702
rect 20456 18612 20484 18702
rect 20088 18584 20484 18612
rect 19890 17776 19946 17785
rect 19890 17711 19946 17720
rect 19720 17564 19932 17592
rect 19798 17504 19854 17513
rect 19798 17439 19854 17448
rect 19616 17128 19668 17134
rect 19616 17070 19668 17076
rect 19812 17066 19840 17439
rect 19800 17060 19852 17066
rect 19800 17002 19852 17008
rect 19616 16992 19668 16998
rect 19616 16934 19668 16940
rect 19628 16697 19656 16934
rect 19614 16688 19670 16697
rect 19614 16623 19670 16632
rect 19812 16590 19840 17002
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 19708 16448 19760 16454
rect 19706 16416 19708 16425
rect 19800 16448 19852 16454
rect 19760 16416 19762 16425
rect 19800 16390 19852 16396
rect 19706 16351 19762 16360
rect 19706 16144 19762 16153
rect 19706 16079 19762 16088
rect 19720 16046 19748 16079
rect 19708 16040 19760 16046
rect 19708 15982 19760 15988
rect 19708 15496 19760 15502
rect 19708 15438 19760 15444
rect 19522 15056 19578 15065
rect 19522 14991 19578 15000
rect 19720 15008 19748 15438
rect 19812 15201 19840 16390
rect 19904 16114 19932 17564
rect 20088 17513 20116 18584
rect 20214 18524 20522 18544
rect 20214 18522 20220 18524
rect 20276 18522 20300 18524
rect 20356 18522 20380 18524
rect 20436 18522 20460 18524
rect 20516 18522 20522 18524
rect 20276 18470 20278 18522
rect 20458 18470 20460 18522
rect 20214 18468 20220 18470
rect 20276 18468 20300 18470
rect 20356 18468 20380 18470
rect 20436 18468 20460 18470
rect 20516 18468 20522 18470
rect 20214 18448 20522 18468
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 20364 17678 20392 18226
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20074 17504 20130 17513
rect 20074 17439 20130 17448
rect 20214 17436 20522 17456
rect 20214 17434 20220 17436
rect 20276 17434 20300 17436
rect 20356 17434 20380 17436
rect 20436 17434 20460 17436
rect 20516 17434 20522 17436
rect 20276 17382 20278 17434
rect 20458 17382 20460 17434
rect 20214 17380 20220 17382
rect 20276 17380 20300 17382
rect 20356 17380 20380 17382
rect 20436 17380 20460 17382
rect 20516 17380 20522 17382
rect 20074 17368 20130 17377
rect 20214 17360 20522 17380
rect 20640 17320 20668 19306
rect 20720 18692 20772 18698
rect 20720 18634 20772 18640
rect 20732 18154 20760 18634
rect 20720 18148 20772 18154
rect 20720 18090 20772 18096
rect 20718 17912 20774 17921
rect 20718 17847 20720 17856
rect 20772 17847 20774 17856
rect 20720 17818 20772 17824
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20732 17513 20760 17614
rect 20718 17504 20774 17513
rect 20718 17439 20774 17448
rect 20074 17303 20130 17312
rect 19984 17264 20036 17270
rect 19984 17206 20036 17212
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19798 15192 19854 15201
rect 19798 15127 19854 15136
rect 19536 14618 19564 14991
rect 19720 14980 19840 15008
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19616 14544 19668 14550
rect 19616 14486 19668 14492
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 19536 11558 19564 14350
rect 19628 14074 19656 14486
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19628 13258 19656 14010
rect 19616 13252 19668 13258
rect 19616 13194 19668 13200
rect 19708 12912 19760 12918
rect 19708 12854 19760 12860
rect 19720 12442 19748 12854
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19340 11144 19392 11150
rect 19338 11112 19340 11121
rect 19392 11112 19394 11121
rect 19338 11047 19394 11056
rect 19536 9674 19564 11494
rect 19708 11348 19760 11354
rect 19708 11290 19760 11296
rect 19720 10266 19748 11290
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19812 10130 19840 14980
rect 19800 10124 19852 10130
rect 19800 10066 19852 10072
rect 19444 9646 19564 9674
rect 19444 8430 19472 9646
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19904 7857 19932 15846
rect 19996 14414 20024 17206
rect 20088 16697 20116 17303
rect 20548 17292 20668 17320
rect 20260 17196 20312 17202
rect 20260 17138 20312 17144
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20074 16688 20130 16697
rect 20074 16623 20130 16632
rect 20074 16552 20130 16561
rect 20272 16522 20300 17138
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20364 16522 20392 16934
rect 20456 16794 20484 17138
rect 20548 16810 20576 17292
rect 20628 17196 20680 17202
rect 20732 17184 20760 17439
rect 20680 17156 20760 17184
rect 20628 17138 20680 17144
rect 20444 16788 20496 16794
rect 20548 16782 20668 16810
rect 20444 16730 20496 16736
rect 20536 16720 20588 16726
rect 20536 16662 20588 16668
rect 20548 16561 20576 16662
rect 20534 16552 20590 16561
rect 20074 16487 20130 16496
rect 20260 16516 20312 16522
rect 20088 16454 20116 16487
rect 20260 16458 20312 16464
rect 20352 16516 20404 16522
rect 20534 16487 20590 16496
rect 20352 16458 20404 16464
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 20214 16348 20522 16368
rect 20214 16346 20220 16348
rect 20276 16346 20300 16348
rect 20356 16346 20380 16348
rect 20436 16346 20460 16348
rect 20516 16346 20522 16348
rect 20276 16294 20278 16346
rect 20458 16294 20460 16346
rect 20214 16292 20220 16294
rect 20276 16292 20300 16294
rect 20356 16292 20380 16294
rect 20436 16292 20460 16294
rect 20516 16292 20522 16294
rect 20214 16272 20522 16292
rect 20548 16182 20576 16213
rect 20536 16176 20588 16182
rect 20534 16144 20536 16153
rect 20588 16144 20590 16153
rect 20076 16108 20128 16114
rect 20534 16079 20590 16088
rect 20076 16050 20128 16056
rect 20088 15706 20116 16050
rect 20168 16040 20220 16046
rect 20168 15982 20220 15988
rect 20180 15881 20208 15982
rect 20166 15872 20222 15881
rect 20166 15807 20222 15816
rect 20076 15700 20128 15706
rect 20076 15642 20128 15648
rect 20166 15600 20222 15609
rect 20166 15535 20222 15544
rect 20180 15502 20208 15535
rect 20548 15502 20576 16079
rect 20168 15496 20220 15502
rect 20074 15464 20130 15473
rect 20168 15438 20220 15444
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20074 15399 20130 15408
rect 20088 15366 20116 15399
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 20214 15260 20522 15280
rect 20214 15258 20220 15260
rect 20276 15258 20300 15260
rect 20356 15258 20380 15260
rect 20436 15258 20460 15260
rect 20516 15258 20522 15260
rect 20276 15206 20278 15258
rect 20458 15206 20460 15258
rect 20214 15204 20220 15206
rect 20276 15204 20300 15206
rect 20356 15204 20380 15206
rect 20436 15204 20460 15206
rect 20516 15204 20522 15206
rect 20214 15184 20522 15204
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 20088 14929 20116 14962
rect 20260 14952 20312 14958
rect 20074 14920 20130 14929
rect 20260 14894 20312 14900
rect 20074 14855 20130 14864
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 19996 10810 20024 13874
rect 20088 13530 20116 14418
rect 20180 14414 20208 14758
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20272 14260 20300 14894
rect 20640 14822 20668 16782
rect 20720 16720 20772 16726
rect 20720 16662 20772 16668
rect 20732 16114 20760 16662
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20720 15972 20772 15978
rect 20720 15914 20772 15920
rect 20732 15881 20760 15914
rect 20718 15872 20774 15881
rect 20718 15807 20774 15816
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20364 14550 20392 14758
rect 20732 14634 20760 15438
rect 20640 14606 20760 14634
rect 20640 14550 20668 14606
rect 20352 14544 20404 14550
rect 20352 14486 20404 14492
rect 20444 14544 20496 14550
rect 20444 14486 20496 14492
rect 20628 14544 20680 14550
rect 20628 14486 20680 14492
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 20352 14340 20404 14346
rect 20456 14328 20484 14486
rect 20536 14408 20588 14414
rect 20588 14368 20668 14396
rect 20536 14350 20588 14356
rect 20404 14300 20484 14328
rect 20352 14282 20404 14288
rect 20153 14232 20300 14260
rect 20153 14056 20181 14232
rect 20214 14172 20522 14192
rect 20214 14170 20220 14172
rect 20276 14170 20300 14172
rect 20356 14170 20380 14172
rect 20436 14170 20460 14172
rect 20516 14170 20522 14172
rect 20276 14118 20278 14170
rect 20458 14118 20460 14170
rect 20214 14116 20220 14118
rect 20276 14116 20300 14118
rect 20356 14116 20380 14118
rect 20436 14116 20460 14118
rect 20516 14116 20522 14118
rect 20214 14096 20522 14116
rect 20153 14028 20208 14056
rect 20180 13977 20208 14028
rect 20166 13968 20222 13977
rect 20166 13903 20222 13912
rect 20534 13968 20590 13977
rect 20534 13903 20536 13912
rect 20588 13903 20590 13912
rect 20536 13874 20588 13880
rect 20444 13864 20496 13870
rect 20442 13832 20444 13841
rect 20496 13832 20498 13841
rect 20442 13767 20498 13776
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 20088 12986 20116 13466
rect 20214 13084 20522 13104
rect 20214 13082 20220 13084
rect 20276 13082 20300 13084
rect 20356 13082 20380 13084
rect 20436 13082 20460 13084
rect 20516 13082 20522 13084
rect 20276 13030 20278 13082
rect 20458 13030 20460 13082
rect 20214 13028 20220 13030
rect 20276 13028 20300 13030
rect 20356 13028 20380 13030
rect 20436 13028 20460 13030
rect 20516 13028 20522 13030
rect 20214 13008 20522 13028
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 20088 10470 20116 12582
rect 20214 11996 20522 12016
rect 20214 11994 20220 11996
rect 20276 11994 20300 11996
rect 20356 11994 20380 11996
rect 20436 11994 20460 11996
rect 20516 11994 20522 11996
rect 20276 11942 20278 11994
rect 20458 11942 20460 11994
rect 20214 11940 20220 11942
rect 20276 11940 20300 11942
rect 20356 11940 20380 11942
rect 20436 11940 20460 11942
rect 20516 11940 20522 11942
rect 20214 11920 20522 11940
rect 20442 11384 20498 11393
rect 20442 11319 20498 11328
rect 20456 11286 20484 11319
rect 20640 11286 20668 14368
rect 20732 14278 20760 14486
rect 20824 14482 20852 20334
rect 20916 19514 20944 21286
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 21008 19938 21036 20878
rect 21100 20398 21128 22714
rect 21180 21956 21232 21962
rect 21180 21898 21232 21904
rect 21192 21690 21220 21898
rect 21272 21888 21324 21894
rect 21272 21830 21324 21836
rect 21180 21684 21232 21690
rect 21180 21626 21232 21632
rect 21180 21480 21232 21486
rect 21180 21422 21232 21428
rect 21088 20392 21140 20398
rect 21088 20334 21140 20340
rect 21192 20262 21220 21422
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 21178 20088 21234 20097
rect 21178 20023 21234 20032
rect 21192 19990 21220 20023
rect 21180 19984 21232 19990
rect 21008 19910 21128 19938
rect 21180 19926 21232 19932
rect 20996 19780 21048 19786
rect 20996 19722 21048 19728
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 20916 18834 20944 19314
rect 20904 18828 20956 18834
rect 20904 18770 20956 18776
rect 21008 18426 21036 19722
rect 21100 19553 21128 19910
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 21086 19544 21142 19553
rect 21086 19479 21142 19488
rect 21100 18834 21128 19479
rect 21088 18828 21140 18834
rect 21088 18770 21140 18776
rect 21088 18624 21140 18630
rect 21192 18601 21220 19790
rect 21284 19242 21312 21830
rect 21376 20602 21404 23831
rect 21468 22778 21496 25230
rect 21652 24342 21680 25366
rect 21640 24336 21692 24342
rect 21640 24278 21692 24284
rect 21652 23322 21680 24278
rect 21732 23520 21784 23526
rect 21732 23462 21784 23468
rect 21640 23316 21692 23322
rect 21640 23258 21692 23264
rect 21456 22772 21508 22778
rect 21456 22714 21508 22720
rect 21456 22500 21508 22506
rect 21456 22442 21508 22448
rect 21468 20942 21496 22442
rect 21638 21856 21694 21865
rect 21638 21791 21694 21800
rect 21548 21344 21600 21350
rect 21548 21286 21600 21292
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 21456 20596 21508 20602
rect 21456 20538 21508 20544
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21376 19689 21404 20198
rect 21362 19680 21418 19689
rect 21362 19615 21418 19624
rect 21468 19514 21496 20538
rect 21456 19508 21508 19514
rect 21456 19450 21508 19456
rect 21454 19408 21510 19417
rect 21454 19343 21510 19352
rect 21272 19236 21324 19242
rect 21272 19178 21324 19184
rect 21284 18902 21312 19178
rect 21272 18896 21324 18902
rect 21272 18838 21324 18844
rect 21364 18828 21416 18834
rect 21364 18770 21416 18776
rect 21272 18760 21324 18766
rect 21376 18737 21404 18770
rect 21468 18766 21496 19343
rect 21456 18760 21508 18766
rect 21272 18702 21324 18708
rect 21362 18728 21418 18737
rect 21088 18566 21140 18572
rect 21178 18592 21234 18601
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20916 17678 20944 18226
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20916 16794 20944 17614
rect 20996 17604 21048 17610
rect 20996 17546 21048 17552
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 21008 16232 21036 17546
rect 21100 17202 21128 18566
rect 21178 18527 21234 18536
rect 21284 18426 21312 18702
rect 21456 18702 21508 18708
rect 21362 18663 21418 18672
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 21376 17785 21404 18566
rect 21456 18284 21508 18290
rect 21560 18272 21588 21286
rect 21652 20942 21680 21791
rect 21640 20936 21692 20942
rect 21640 20878 21692 20884
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21652 20466 21680 20742
rect 21640 20460 21692 20466
rect 21640 20402 21692 20408
rect 21744 19378 21772 23462
rect 21836 21350 21864 25735
rect 21824 21344 21876 21350
rect 21824 21286 21876 21292
rect 21822 21176 21878 21185
rect 21822 21111 21824 21120
rect 21876 21111 21878 21120
rect 21824 21082 21876 21088
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 21732 19372 21784 19378
rect 21732 19314 21784 19320
rect 21732 18828 21784 18834
rect 21732 18770 21784 18776
rect 21640 18624 21692 18630
rect 21640 18566 21692 18572
rect 21508 18244 21588 18272
rect 21456 18226 21508 18232
rect 21362 17776 21418 17785
rect 21180 17740 21232 17746
rect 21362 17711 21418 17720
rect 21180 17682 21232 17688
rect 21192 17338 21220 17682
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21284 16590 21312 17478
rect 21362 17368 21418 17377
rect 21362 17303 21418 17312
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 21272 16584 21324 16590
rect 21272 16526 21324 16532
rect 21192 16425 21220 16526
rect 21272 16448 21324 16454
rect 21178 16416 21234 16425
rect 21272 16390 21324 16396
rect 21178 16351 21234 16360
rect 21008 16204 21220 16232
rect 21086 16144 21142 16153
rect 21086 16079 21142 16088
rect 21100 16046 21128 16079
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 21192 15858 21220 16204
rect 21008 15830 21220 15858
rect 20902 15600 20958 15609
rect 20902 15535 20904 15544
rect 20956 15535 20958 15544
rect 20904 15506 20956 15512
rect 20904 15360 20956 15366
rect 20902 15328 20904 15337
rect 20956 15328 20958 15337
rect 20902 15263 20958 15272
rect 20902 15192 20958 15201
rect 20902 15127 20904 15136
rect 20956 15127 20958 15136
rect 20904 15098 20956 15104
rect 20902 14920 20958 14929
rect 20902 14855 20958 14864
rect 20916 14657 20944 14855
rect 20902 14648 20958 14657
rect 20902 14583 20958 14592
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 20824 13870 20852 14418
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20916 14113 20944 14350
rect 20902 14104 20958 14113
rect 21008 14074 21036 15830
rect 21284 15706 21312 16390
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 21100 14657 21128 15642
rect 21180 15632 21232 15638
rect 21376 15586 21404 17303
rect 21180 15574 21232 15580
rect 21192 15201 21220 15574
rect 21284 15558 21404 15586
rect 21178 15192 21234 15201
rect 21178 15127 21234 15136
rect 21284 15076 21312 15558
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21192 15048 21312 15076
rect 21086 14648 21142 14657
rect 21086 14583 21142 14592
rect 21086 14376 21142 14385
rect 21086 14311 21142 14320
rect 20902 14039 20958 14048
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20994 13968 21050 13977
rect 20994 13903 20996 13912
rect 21048 13903 21050 13912
rect 20996 13874 21048 13880
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20718 13560 20774 13569
rect 20718 13495 20774 13504
rect 20732 12850 20760 13495
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 20824 13161 20852 13262
rect 20810 13152 20866 13161
rect 20810 13087 20866 13096
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20916 12442 20944 13670
rect 21100 13569 21128 14311
rect 21192 14006 21220 15048
rect 21272 14544 21324 14550
rect 21272 14486 21324 14492
rect 21284 14414 21312 14486
rect 21376 14414 21404 15438
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 21364 14408 21416 14414
rect 21364 14350 21416 14356
rect 21180 14000 21232 14006
rect 21180 13942 21232 13948
rect 21272 13728 21324 13734
rect 21178 13696 21234 13705
rect 21272 13670 21324 13676
rect 21362 13696 21418 13705
rect 21178 13631 21234 13640
rect 21086 13560 21142 13569
rect 21086 13495 21142 13504
rect 20996 13252 21048 13258
rect 20996 13194 21048 13200
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20902 12064 20958 12073
rect 20902 11999 20958 12008
rect 20444 11280 20496 11286
rect 20444 11222 20496 11228
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20916 11150 20944 11999
rect 21008 11762 21036 13194
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 21008 11558 21036 11698
rect 20996 11552 21048 11558
rect 20996 11494 21048 11500
rect 21192 11506 21220 13631
rect 21284 13190 21312 13670
rect 21362 13631 21418 13640
rect 21376 13326 21404 13631
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21272 13184 21324 13190
rect 21272 13126 21324 13132
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20214 10908 20522 10928
rect 20214 10906 20220 10908
rect 20276 10906 20300 10908
rect 20356 10906 20380 10908
rect 20436 10906 20460 10908
rect 20516 10906 20522 10908
rect 20276 10854 20278 10906
rect 20458 10854 20460 10906
rect 20214 10852 20220 10854
rect 20276 10852 20300 10854
rect 20356 10852 20380 10854
rect 20436 10852 20460 10854
rect 20516 10852 20522 10854
rect 20214 10832 20522 10852
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20214 9820 20522 9840
rect 20214 9818 20220 9820
rect 20276 9818 20300 9820
rect 20356 9818 20380 9820
rect 20436 9818 20460 9820
rect 20516 9818 20522 9820
rect 20276 9766 20278 9818
rect 20458 9766 20460 9818
rect 20214 9764 20220 9766
rect 20276 9764 20300 9766
rect 20356 9764 20380 9766
rect 20436 9764 20460 9766
rect 20516 9764 20522 9766
rect 20214 9744 20522 9764
rect 20640 8838 20668 10406
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20214 8732 20522 8752
rect 20214 8730 20220 8732
rect 20276 8730 20300 8732
rect 20356 8730 20380 8732
rect 20436 8730 20460 8732
rect 20516 8730 20522 8732
rect 20276 8678 20278 8730
rect 20458 8678 20460 8730
rect 20214 8676 20220 8678
rect 20276 8676 20300 8678
rect 20356 8676 20380 8678
rect 20436 8676 20460 8678
rect 20516 8676 20522 8678
rect 20214 8656 20522 8676
rect 19890 7848 19946 7857
rect 19890 7783 19946 7792
rect 20214 7644 20522 7664
rect 20214 7642 20220 7644
rect 20276 7642 20300 7644
rect 20356 7642 20380 7644
rect 20436 7642 20460 7644
rect 20516 7642 20522 7644
rect 20276 7590 20278 7642
rect 20458 7590 20460 7642
rect 20214 7588 20220 7590
rect 20276 7588 20300 7590
rect 20356 7588 20380 7590
rect 20436 7588 20460 7590
rect 20516 7588 20522 7590
rect 20214 7568 20522 7588
rect 19168 6886 19288 6914
rect 18432 5370 18460 6886
rect 18420 5364 18472 5370
rect 18420 5306 18472 5312
rect 19260 4078 19288 6886
rect 20214 6556 20522 6576
rect 20214 6554 20220 6556
rect 20276 6554 20300 6556
rect 20356 6554 20380 6556
rect 20436 6554 20460 6556
rect 20516 6554 20522 6556
rect 20276 6502 20278 6554
rect 20458 6502 20460 6554
rect 20214 6500 20220 6502
rect 20276 6500 20300 6502
rect 20356 6500 20380 6502
rect 20436 6500 20460 6502
rect 20516 6500 20522 6502
rect 20214 6480 20522 6500
rect 20214 5468 20522 5488
rect 20214 5466 20220 5468
rect 20276 5466 20300 5468
rect 20356 5466 20380 5468
rect 20436 5466 20460 5468
rect 20516 5466 20522 5468
rect 20276 5414 20278 5466
rect 20458 5414 20460 5466
rect 20214 5412 20220 5414
rect 20276 5412 20300 5414
rect 20356 5412 20380 5414
rect 20436 5412 20460 5414
rect 20516 5412 20522 5414
rect 20214 5392 20522 5412
rect 20214 4380 20522 4400
rect 20214 4378 20220 4380
rect 20276 4378 20300 4380
rect 20356 4378 20380 4380
rect 20436 4378 20460 4380
rect 20516 4378 20522 4380
rect 20276 4326 20278 4378
rect 20458 4326 20460 4378
rect 20214 4324 20220 4326
rect 20276 4324 20300 4326
rect 20356 4324 20380 4326
rect 20436 4324 20460 4326
rect 20516 4324 20522 4326
rect 20214 4304 20522 4324
rect 19248 4072 19300 4078
rect 19248 4014 19300 4020
rect 21008 4010 21036 11494
rect 21192 11478 21312 11506
rect 21178 11384 21234 11393
rect 21178 11319 21180 11328
rect 21232 11319 21234 11328
rect 21180 11290 21232 11296
rect 21180 10804 21232 10810
rect 21180 10746 21232 10752
rect 20996 4004 21048 4010
rect 20996 3946 21048 3952
rect 20214 3292 20522 3312
rect 20214 3290 20220 3292
rect 20276 3290 20300 3292
rect 20356 3290 20380 3292
rect 20436 3290 20460 3292
rect 20516 3290 20522 3292
rect 20276 3238 20278 3290
rect 20458 3238 20460 3290
rect 20214 3236 20220 3238
rect 20276 3236 20300 3238
rect 20356 3236 20380 3238
rect 20436 3236 20460 3238
rect 20516 3236 20522 3238
rect 20214 3216 20522 3236
rect 21192 2961 21220 10746
rect 21284 8974 21312 11478
rect 21376 10810 21404 13262
rect 21364 10804 21416 10810
rect 21364 10746 21416 10752
rect 21468 10713 21496 18226
rect 21652 18086 21680 18566
rect 21744 18358 21772 18770
rect 21836 18630 21864 20198
rect 21928 20097 21956 26930
rect 22836 26920 22888 26926
rect 22836 26862 22888 26868
rect 22006 26752 22062 26761
rect 22006 26687 22062 26696
rect 22020 25770 22048 26687
rect 22008 25764 22060 25770
rect 22008 25706 22060 25712
rect 22098 25120 22154 25129
rect 22098 25055 22154 25064
rect 22008 24268 22060 24274
rect 22008 24210 22060 24216
rect 22020 24070 22048 24210
rect 22008 24064 22060 24070
rect 22008 24006 22060 24012
rect 22020 23662 22048 24006
rect 22008 23656 22060 23662
rect 22008 23598 22060 23604
rect 22008 23316 22060 23322
rect 22008 23258 22060 23264
rect 22020 22438 22048 23258
rect 22008 22432 22060 22438
rect 22006 22400 22008 22409
rect 22060 22400 22062 22409
rect 22006 22335 22062 22344
rect 22112 22030 22140 25055
rect 22192 24812 22244 24818
rect 22192 24754 22244 24760
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22204 21894 22232 24754
rect 22284 24676 22336 24682
rect 22284 24618 22336 24624
rect 22296 24206 22324 24618
rect 22744 24608 22796 24614
rect 22744 24550 22796 24556
rect 22756 24449 22784 24550
rect 22742 24440 22798 24449
rect 22742 24375 22798 24384
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 22848 23662 22876 26862
rect 23204 26512 23256 26518
rect 23204 26454 23256 26460
rect 23020 25764 23072 25770
rect 23020 25706 23072 25712
rect 22928 24200 22980 24206
rect 22928 24142 22980 24148
rect 22836 23656 22888 23662
rect 22836 23598 22888 23604
rect 22560 23180 22612 23186
rect 22560 23122 22612 23128
rect 22376 22976 22428 22982
rect 22376 22918 22428 22924
rect 22388 21978 22416 22918
rect 22296 21950 22416 21978
rect 22192 21888 22244 21894
rect 22098 21856 22154 21865
rect 22192 21830 22244 21836
rect 22098 21791 22154 21800
rect 22112 21078 22140 21791
rect 22190 21584 22246 21593
rect 22296 21554 22324 21950
rect 22376 21888 22428 21894
rect 22376 21830 22428 21836
rect 22190 21519 22246 21528
rect 22284 21548 22336 21554
rect 22100 21072 22152 21078
rect 22100 21014 22152 21020
rect 22098 20496 22154 20505
rect 22098 20431 22154 20440
rect 22008 20256 22060 20262
rect 22008 20198 22060 20204
rect 21914 20088 21970 20097
rect 21914 20023 21970 20032
rect 21928 18834 21956 20023
rect 22020 19922 22048 20198
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 22112 19718 22140 20431
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 22204 19514 22232 21519
rect 22284 21490 22336 21496
rect 22284 21344 22336 21350
rect 22284 21286 22336 21292
rect 22296 20534 22324 21286
rect 22284 20528 22336 20534
rect 22284 20470 22336 20476
rect 22284 20392 22336 20398
rect 22284 20334 22336 20340
rect 22192 19508 22244 19514
rect 22192 19450 22244 19456
rect 22190 19408 22246 19417
rect 22190 19343 22192 19352
rect 22244 19343 22246 19352
rect 22192 19314 22244 19320
rect 22192 19236 22244 19242
rect 22192 19178 22244 19184
rect 22008 18896 22060 18902
rect 22008 18838 22060 18844
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 21824 18624 21876 18630
rect 21824 18566 21876 18572
rect 21732 18352 21784 18358
rect 21732 18294 21784 18300
rect 21640 18080 21692 18086
rect 21640 18022 21692 18028
rect 21744 17882 21772 18294
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 21548 17876 21600 17882
rect 21548 17818 21600 17824
rect 21732 17876 21784 17882
rect 21732 17818 21784 17824
rect 21560 16522 21588 17818
rect 21928 17338 21956 18022
rect 22020 17785 22048 18838
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 22006 17776 22062 17785
rect 22006 17711 22062 17720
rect 21916 17332 21968 17338
rect 21916 17274 21968 17280
rect 22112 17270 22140 17818
rect 22100 17264 22152 17270
rect 22100 17206 22152 17212
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 21640 16992 21692 16998
rect 21640 16934 21692 16940
rect 21652 16658 21680 16934
rect 21730 16688 21786 16697
rect 21640 16652 21692 16658
rect 21730 16623 21732 16632
rect 21640 16594 21692 16600
rect 21784 16623 21786 16632
rect 21732 16594 21784 16600
rect 21548 16516 21600 16522
rect 21548 16458 21600 16464
rect 21638 16280 21694 16289
rect 21638 16215 21694 16224
rect 21546 16144 21602 16153
rect 21652 16114 21680 16215
rect 21546 16079 21602 16088
rect 21640 16108 21692 16114
rect 21560 15570 21588 16079
rect 21640 16050 21692 16056
rect 21732 16108 21784 16114
rect 21836 16096 21864 17138
rect 21914 17096 21970 17105
rect 21914 17031 21916 17040
rect 21968 17031 21970 17040
rect 21916 17002 21968 17008
rect 22204 16794 22232 19178
rect 22296 17377 22324 20334
rect 22388 20074 22416 21830
rect 22572 21010 22600 23122
rect 22744 22976 22796 22982
rect 22744 22918 22796 22924
rect 22756 22817 22784 22918
rect 22742 22808 22798 22817
rect 22742 22743 22798 22752
rect 22756 22234 22784 22743
rect 22836 22568 22888 22574
rect 22836 22510 22888 22516
rect 22848 22438 22876 22510
rect 22836 22432 22888 22438
rect 22834 22400 22836 22409
rect 22888 22400 22890 22409
rect 22834 22335 22890 22344
rect 22744 22228 22796 22234
rect 22744 22170 22796 22176
rect 22940 22030 22968 24142
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22756 21486 22784 21966
rect 22834 21720 22890 21729
rect 22834 21655 22890 21664
rect 22848 21622 22876 21655
rect 22836 21616 22888 21622
rect 22836 21558 22888 21564
rect 22928 21616 22980 21622
rect 22928 21558 22980 21564
rect 22744 21480 22796 21486
rect 22940 21457 22968 21558
rect 22744 21422 22796 21428
rect 22926 21448 22982 21457
rect 22560 21004 22612 21010
rect 22560 20946 22612 20952
rect 22558 20632 22614 20641
rect 22558 20567 22614 20576
rect 22388 20046 22508 20074
rect 22374 19952 22430 19961
rect 22480 19922 22508 20046
rect 22374 19887 22430 19896
rect 22468 19916 22520 19922
rect 22388 19378 22416 19887
rect 22468 19858 22520 19864
rect 22376 19372 22428 19378
rect 22376 19314 22428 19320
rect 22466 19136 22522 19145
rect 22466 19071 22522 19080
rect 22376 18692 22428 18698
rect 22376 18634 22428 18640
rect 22388 18465 22416 18634
rect 22374 18456 22430 18465
rect 22374 18391 22430 18400
rect 22480 18290 22508 19071
rect 22468 18284 22520 18290
rect 22468 18226 22520 18232
rect 22572 18170 22600 20567
rect 22652 19916 22704 19922
rect 22652 19858 22704 19864
rect 22664 19378 22692 19858
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22388 18142 22600 18170
rect 22388 17610 22416 18142
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 22376 17604 22428 17610
rect 22376 17546 22428 17552
rect 22480 17513 22508 17682
rect 22466 17504 22522 17513
rect 22466 17439 22522 17448
rect 22282 17368 22338 17377
rect 22282 17303 22338 17312
rect 22376 17128 22428 17134
rect 22664 17116 22692 19314
rect 22428 17088 22692 17116
rect 22376 17070 22428 17076
rect 22192 16788 22244 16794
rect 22192 16730 22244 16736
rect 22008 16584 22060 16590
rect 22480 16561 22508 17088
rect 22008 16526 22060 16532
rect 22466 16552 22522 16561
rect 21784 16068 21864 16096
rect 21732 16050 21784 16056
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 21548 15564 21600 15570
rect 21548 15506 21600 15512
rect 21546 15328 21602 15337
rect 21546 15263 21602 15272
rect 21560 15094 21588 15263
rect 21548 15088 21600 15094
rect 21548 15030 21600 15036
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 21560 14482 21588 14758
rect 21548 14476 21600 14482
rect 21548 14418 21600 14424
rect 21548 14272 21600 14278
rect 21548 14214 21600 14220
rect 21560 13977 21588 14214
rect 21546 13968 21602 13977
rect 21546 13903 21602 13912
rect 21548 13796 21600 13802
rect 21548 13738 21600 13744
rect 21560 13569 21588 13738
rect 21546 13560 21602 13569
rect 21546 13495 21602 13504
rect 21560 12442 21588 13495
rect 21652 12714 21680 15846
rect 21744 15638 21772 16050
rect 21732 15632 21784 15638
rect 21732 15574 21784 15580
rect 21730 15328 21786 15337
rect 21730 15263 21786 15272
rect 21744 15162 21772 15263
rect 21732 15156 21784 15162
rect 21732 15098 21784 15104
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21732 15020 21784 15026
rect 21732 14962 21784 14968
rect 21744 13462 21772 14962
rect 21836 14890 21864 15098
rect 21824 14884 21876 14890
rect 21824 14826 21876 14832
rect 21916 14884 21968 14890
rect 21916 14826 21968 14832
rect 21824 14476 21876 14482
rect 21824 14418 21876 14424
rect 21732 13456 21784 13462
rect 21732 13398 21784 13404
rect 21640 12708 21692 12714
rect 21640 12650 21692 12656
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21546 11520 21602 11529
rect 21546 11455 21602 11464
rect 21560 11354 21588 11455
rect 21548 11348 21600 11354
rect 21548 11290 21600 11296
rect 21454 10704 21510 10713
rect 21454 10639 21510 10648
rect 21744 9042 21772 13398
rect 21836 12918 21864 14418
rect 21928 14346 21956 14826
rect 21916 14340 21968 14346
rect 21916 14282 21968 14288
rect 22020 14226 22048 16526
rect 22284 16516 22336 16522
rect 22466 16487 22522 16496
rect 22284 16458 22336 16464
rect 22190 16144 22246 16153
rect 22190 16079 22246 16088
rect 22098 15736 22154 15745
rect 22098 15671 22154 15680
rect 22112 15434 22140 15671
rect 22204 15502 22232 16079
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 22100 15428 22152 15434
rect 22100 15370 22152 15376
rect 22296 15162 22324 16458
rect 22560 16448 22612 16454
rect 22560 16390 22612 16396
rect 22468 16040 22520 16046
rect 22468 15982 22520 15988
rect 22376 15972 22428 15978
rect 22376 15914 22428 15920
rect 22284 15156 22336 15162
rect 22284 15098 22336 15104
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 22112 14822 22140 14962
rect 22284 14884 22336 14890
rect 22284 14826 22336 14832
rect 22100 14816 22152 14822
rect 22100 14758 22152 14764
rect 22190 14512 22246 14521
rect 22296 14482 22324 14826
rect 22190 14447 22246 14456
rect 22284 14476 22336 14482
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 22112 14278 22140 14350
rect 21928 14198 22048 14226
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 21928 13190 21956 14198
rect 22006 14104 22062 14113
rect 22006 14039 22062 14048
rect 22020 13802 22048 14039
rect 22008 13796 22060 13802
rect 22008 13738 22060 13744
rect 22006 13560 22062 13569
rect 22006 13495 22008 13504
rect 22060 13495 22062 13504
rect 22008 13466 22060 13472
rect 22008 13388 22060 13394
rect 22008 13330 22060 13336
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 21928 12986 21956 13126
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 21824 12912 21876 12918
rect 21824 12854 21876 12860
rect 21822 12472 21878 12481
rect 21822 12407 21878 12416
rect 21916 12436 21968 12442
rect 21836 12238 21864 12407
rect 21916 12378 21968 12384
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 21928 11529 21956 12378
rect 22020 11830 22048 13330
rect 22112 12374 22140 14214
rect 22204 13938 22232 14447
rect 22284 14418 22336 14424
rect 22192 13932 22244 13938
rect 22244 13892 22324 13920
rect 22192 13874 22244 13880
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22204 13326 22232 13466
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22296 12968 22324 13892
rect 22388 13870 22416 15914
rect 22480 15609 22508 15982
rect 22466 15600 22522 15609
rect 22466 15535 22522 15544
rect 22468 14340 22520 14346
rect 22468 14282 22520 14288
rect 22376 13864 22428 13870
rect 22376 13806 22428 13812
rect 22480 13802 22508 14282
rect 22468 13796 22520 13802
rect 22468 13738 22520 13744
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 22388 13138 22416 13670
rect 22388 13110 22508 13138
rect 22296 12940 22416 12968
rect 22192 12912 22244 12918
rect 22192 12854 22244 12860
rect 22100 12368 22152 12374
rect 22100 12310 22152 12316
rect 22204 11898 22232 12854
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22192 11892 22244 11898
rect 22192 11834 22244 11840
rect 22008 11824 22060 11830
rect 22008 11766 22060 11772
rect 21914 11520 21970 11529
rect 21914 11455 21970 11464
rect 21914 11384 21970 11393
rect 21914 11319 21970 11328
rect 21732 9036 21784 9042
rect 21732 8978 21784 8984
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21178 2952 21234 2961
rect 21178 2887 21234 2896
rect 17960 2576 18012 2582
rect 17960 2518 18012 2524
rect 21928 2417 21956 11319
rect 22296 11082 22324 12786
rect 22388 12374 22416 12940
rect 22480 12481 22508 13110
rect 22466 12472 22522 12481
rect 22466 12407 22522 12416
rect 22376 12368 22428 12374
rect 22376 12310 22428 12316
rect 22388 11762 22416 12310
rect 22480 11898 22508 12407
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22376 11756 22428 11762
rect 22376 11698 22428 11704
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 22572 10305 22600 16390
rect 22756 16130 22784 21422
rect 22926 21383 22982 21392
rect 22928 21344 22980 21350
rect 22928 21286 22980 21292
rect 22940 20874 22968 21286
rect 23032 21010 23060 25706
rect 23112 24608 23164 24614
rect 23112 24550 23164 24556
rect 23124 22030 23152 24550
rect 23216 22098 23244 26454
rect 23388 26444 23440 26450
rect 23388 26386 23440 26392
rect 23400 24410 23428 26386
rect 23952 25430 23980 27882
rect 23940 25424 23992 25430
rect 23940 25366 23992 25372
rect 23848 25220 23900 25226
rect 23848 25162 23900 25168
rect 23388 24404 23440 24410
rect 23388 24346 23440 24352
rect 23572 24336 23624 24342
rect 23572 24278 23624 24284
rect 23584 24070 23612 24278
rect 23664 24132 23716 24138
rect 23664 24074 23716 24080
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23296 23588 23348 23594
rect 23296 23530 23348 23536
rect 23308 23254 23336 23530
rect 23296 23248 23348 23254
rect 23296 23190 23348 23196
rect 23480 23044 23532 23050
rect 23480 22986 23532 22992
rect 23296 22976 23348 22982
rect 23296 22918 23348 22924
rect 23308 22778 23336 22918
rect 23296 22772 23348 22778
rect 23296 22714 23348 22720
rect 23204 22092 23256 22098
rect 23204 22034 23256 22040
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 23124 21457 23152 21966
rect 23308 21962 23336 22714
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23400 22273 23428 22374
rect 23386 22264 23442 22273
rect 23386 22199 23442 22208
rect 23296 21956 23348 21962
rect 23296 21898 23348 21904
rect 23204 21616 23256 21622
rect 23204 21558 23256 21564
rect 23110 21448 23166 21457
rect 23110 21383 23166 21392
rect 23124 21049 23152 21383
rect 23110 21040 23166 21049
rect 23020 21004 23072 21010
rect 23110 20975 23166 20984
rect 23020 20946 23072 20952
rect 22928 20868 22980 20874
rect 22928 20810 22980 20816
rect 22836 20800 22888 20806
rect 22834 20768 22836 20777
rect 22888 20768 22890 20777
rect 22834 20703 22890 20712
rect 23216 20466 23244 21558
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 23204 20460 23256 20466
rect 23204 20402 23256 20408
rect 23020 20324 23072 20330
rect 23020 20266 23072 20272
rect 22928 19848 22980 19854
rect 22928 19790 22980 19796
rect 22940 19378 22968 19790
rect 22928 19372 22980 19378
rect 22928 19314 22980 19320
rect 22940 17746 22968 19314
rect 23032 18601 23060 20266
rect 23400 19530 23428 21490
rect 23492 20641 23520 22986
rect 23584 22574 23612 24006
rect 23572 22568 23624 22574
rect 23572 22510 23624 22516
rect 23572 22228 23624 22234
rect 23572 22170 23624 22176
rect 23584 20942 23612 22170
rect 23572 20936 23624 20942
rect 23572 20878 23624 20884
rect 23478 20632 23534 20641
rect 23478 20567 23534 20576
rect 23676 20398 23704 24074
rect 23860 22642 23888 25162
rect 24124 24676 24176 24682
rect 24124 24618 24176 24624
rect 24136 23798 24164 24618
rect 24124 23792 24176 23798
rect 24124 23734 24176 23740
rect 24124 23112 24176 23118
rect 24124 23054 24176 23060
rect 23940 22976 23992 22982
rect 23940 22918 23992 22924
rect 24032 22976 24084 22982
rect 24032 22918 24084 22924
rect 23848 22636 23900 22642
rect 23848 22578 23900 22584
rect 23756 22568 23808 22574
rect 23756 22510 23808 22516
rect 23768 21128 23796 22510
rect 23952 22030 23980 22918
rect 23940 22024 23992 22030
rect 23940 21966 23992 21972
rect 23952 21350 23980 21966
rect 23940 21344 23992 21350
rect 23940 21286 23992 21292
rect 23768 21100 23980 21128
rect 23754 21040 23810 21049
rect 23754 20975 23756 20984
rect 23808 20975 23810 20984
rect 23756 20946 23808 20952
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23768 20398 23796 20470
rect 23664 20392 23716 20398
rect 23664 20334 23716 20340
rect 23756 20392 23808 20398
rect 23756 20334 23808 20340
rect 23570 20088 23626 20097
rect 23570 20023 23626 20032
rect 23584 19718 23612 20023
rect 23664 19984 23716 19990
rect 23664 19926 23716 19932
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23204 19508 23256 19514
rect 23400 19502 23612 19530
rect 23676 19514 23704 19926
rect 23204 19450 23256 19456
rect 23110 18728 23166 18737
rect 23110 18663 23166 18672
rect 23018 18592 23074 18601
rect 23018 18527 23074 18536
rect 23020 18420 23072 18426
rect 23020 18362 23072 18368
rect 22928 17740 22980 17746
rect 22928 17682 22980 17688
rect 23032 17626 23060 18362
rect 22836 17604 22888 17610
rect 22836 17546 22888 17552
rect 22940 17598 23060 17626
rect 22848 17338 22876 17546
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 22756 16102 22876 16130
rect 22744 16040 22796 16046
rect 22744 15982 22796 15988
rect 22650 15736 22706 15745
rect 22650 15671 22652 15680
rect 22704 15671 22706 15680
rect 22652 15642 22704 15648
rect 22756 15337 22784 15982
rect 22742 15328 22798 15337
rect 22742 15263 22798 15272
rect 22652 15020 22704 15026
rect 22652 14962 22704 14968
rect 22664 12986 22692 14962
rect 22744 14816 22796 14822
rect 22744 14758 22796 14764
rect 22756 13734 22784 14758
rect 22848 14550 22876 16102
rect 22940 15026 22968 17598
rect 23020 17536 23072 17542
rect 23020 17478 23072 17484
rect 23032 17270 23060 17478
rect 23020 17264 23072 17270
rect 23020 17206 23072 17212
rect 22928 15020 22980 15026
rect 22928 14962 22980 14968
rect 22928 14816 22980 14822
rect 22928 14758 22980 14764
rect 22836 14544 22888 14550
rect 22836 14486 22888 14492
rect 22836 13932 22888 13938
rect 22836 13874 22888 13880
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22652 12980 22704 12986
rect 22652 12922 22704 12928
rect 22848 12850 22876 13874
rect 22836 12844 22888 12850
rect 22836 12786 22888 12792
rect 22744 11756 22796 11762
rect 22744 11698 22796 11704
rect 22650 10840 22706 10849
rect 22650 10775 22652 10784
rect 22704 10775 22706 10784
rect 22652 10746 22704 10752
rect 22558 10296 22614 10305
rect 22558 10231 22614 10240
rect 22008 9444 22060 9450
rect 22008 9386 22060 9392
rect 22020 5574 22048 9386
rect 22756 6730 22784 11698
rect 22848 11354 22876 12786
rect 22940 11762 22968 14758
rect 23032 13938 23060 17206
rect 23124 16046 23152 18663
rect 23112 16040 23164 16046
rect 23112 15982 23164 15988
rect 23216 15201 23244 19450
rect 23480 18080 23532 18086
rect 23386 18048 23442 18057
rect 23480 18022 23532 18028
rect 23386 17983 23442 17992
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 23308 15366 23336 17070
rect 23400 16017 23428 17983
rect 23386 16008 23442 16017
rect 23386 15943 23442 15952
rect 23492 15706 23520 18022
rect 23480 15700 23532 15706
rect 23480 15642 23532 15648
rect 23584 15609 23612 19502
rect 23664 19508 23716 19514
rect 23664 19450 23716 19456
rect 23846 19408 23902 19417
rect 23846 19343 23902 19352
rect 23860 18834 23888 19343
rect 23952 18834 23980 21100
rect 24044 20534 24072 22918
rect 24136 22642 24164 23054
rect 24228 22710 24256 28455
rect 24504 27606 24532 29200
rect 29846 27772 30154 27792
rect 29846 27770 29852 27772
rect 29908 27770 29932 27772
rect 29988 27770 30012 27772
rect 30068 27770 30092 27772
rect 30148 27770 30154 27772
rect 29908 27718 29910 27770
rect 30090 27718 30092 27770
rect 29846 27716 29852 27718
rect 29908 27716 29932 27718
rect 29988 27716 30012 27718
rect 30068 27716 30092 27718
rect 30148 27716 30154 27718
rect 29846 27696 30154 27716
rect 30208 27606 30236 29294
rect 32312 28212 32364 28218
rect 32312 28154 32364 28160
rect 30470 27976 30526 27985
rect 30470 27911 30526 27920
rect 30288 27668 30340 27674
rect 30288 27610 30340 27616
rect 24492 27600 24544 27606
rect 24492 27542 24544 27548
rect 30196 27600 30248 27606
rect 30196 27542 30248 27548
rect 28632 27464 28684 27470
rect 28632 27406 28684 27412
rect 28814 27432 28870 27441
rect 25780 27328 25832 27334
rect 25780 27270 25832 27276
rect 26424 27328 26476 27334
rect 26424 27270 26476 27276
rect 28540 27328 28592 27334
rect 28540 27270 28592 27276
rect 25792 27130 25820 27270
rect 25780 27124 25832 27130
rect 25780 27066 25832 27072
rect 25136 26784 25188 26790
rect 25136 26726 25188 26732
rect 25148 26246 25176 26726
rect 24676 26240 24728 26246
rect 24676 26182 24728 26188
rect 25136 26240 25188 26246
rect 25136 26182 25188 26188
rect 25412 26240 25464 26246
rect 25412 26182 25464 26188
rect 24582 26072 24638 26081
rect 24582 26007 24638 26016
rect 24400 25696 24452 25702
rect 24400 25638 24452 25644
rect 24412 25537 24440 25638
rect 24398 25528 24454 25537
rect 24398 25463 24454 25472
rect 24306 24984 24362 24993
rect 24306 24919 24362 24928
rect 24216 22704 24268 22710
rect 24216 22646 24268 22652
rect 24124 22636 24176 22642
rect 24124 22578 24176 22584
rect 24136 22545 24164 22578
rect 24122 22536 24178 22545
rect 24122 22471 24178 22480
rect 24124 22228 24176 22234
rect 24124 22170 24176 22176
rect 24136 21622 24164 22170
rect 24216 22092 24268 22098
rect 24216 22034 24268 22040
rect 24124 21616 24176 21622
rect 24124 21558 24176 21564
rect 24228 21350 24256 22034
rect 24124 21344 24176 21350
rect 24124 21286 24176 21292
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 24032 20528 24084 20534
rect 24032 20470 24084 20476
rect 24044 20398 24072 20429
rect 24032 20392 24084 20398
rect 24136 20346 24164 21286
rect 24320 21185 24348 24919
rect 24400 24608 24452 24614
rect 24400 24550 24452 24556
rect 24412 22681 24440 24550
rect 24596 24070 24624 26007
rect 24688 25974 24716 26182
rect 24676 25968 24728 25974
rect 24676 25910 24728 25916
rect 24860 25696 24912 25702
rect 24860 25638 24912 25644
rect 25044 25696 25096 25702
rect 25044 25638 25096 25644
rect 24584 24064 24636 24070
rect 24584 24006 24636 24012
rect 24492 23112 24544 23118
rect 24596 23089 24624 24006
rect 24872 23662 24900 25638
rect 24952 25152 25004 25158
rect 24952 25094 25004 25100
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 24860 23248 24912 23254
rect 24860 23190 24912 23196
rect 24768 23180 24820 23186
rect 24768 23122 24820 23128
rect 24676 23112 24728 23118
rect 24492 23054 24544 23060
rect 24582 23080 24638 23089
rect 24398 22672 24454 22681
rect 24398 22607 24454 22616
rect 24412 22574 24440 22607
rect 24400 22568 24452 22574
rect 24400 22510 24452 22516
rect 24504 22098 24532 23054
rect 24676 23054 24728 23060
rect 24582 23015 24638 23024
rect 24688 22930 24716 23054
rect 24596 22902 24716 22930
rect 24492 22092 24544 22098
rect 24492 22034 24544 22040
rect 24596 21842 24624 22902
rect 24674 22400 24730 22409
rect 24674 22335 24730 22344
rect 24412 21814 24624 21842
rect 24306 21176 24362 21185
rect 24306 21111 24362 21120
rect 24320 20534 24348 21111
rect 24308 20528 24360 20534
rect 24308 20470 24360 20476
rect 24084 20340 24164 20346
rect 24032 20334 24164 20340
rect 24044 20318 24164 20334
rect 24308 20324 24360 20330
rect 23848 18828 23900 18834
rect 23848 18770 23900 18776
rect 23940 18828 23992 18834
rect 23940 18770 23992 18776
rect 23846 18728 23902 18737
rect 23846 18663 23902 18672
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23676 18329 23704 18362
rect 23662 18320 23718 18329
rect 23860 18290 23888 18663
rect 23662 18255 23718 18264
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 23664 17672 23716 17678
rect 23664 17614 23716 17620
rect 23570 15600 23626 15609
rect 23570 15535 23626 15544
rect 23572 15428 23624 15434
rect 23572 15370 23624 15376
rect 23296 15360 23348 15366
rect 23296 15302 23348 15308
rect 23202 15192 23258 15201
rect 23112 15156 23164 15162
rect 23202 15127 23258 15136
rect 23112 15098 23164 15104
rect 23124 14793 23152 15098
rect 23204 15020 23256 15026
rect 23204 14962 23256 14968
rect 23110 14784 23166 14793
rect 23110 14719 23166 14728
rect 23020 13932 23072 13938
rect 23020 13874 23072 13880
rect 23032 13258 23060 13874
rect 23020 13252 23072 13258
rect 23020 13194 23072 13200
rect 23032 12646 23060 13194
rect 23020 12640 23072 12646
rect 23020 12582 23072 12588
rect 22928 11756 22980 11762
rect 22928 11698 22980 11704
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 23020 11076 23072 11082
rect 23020 11018 23072 11024
rect 23032 7585 23060 11018
rect 23124 10169 23152 14719
rect 23216 14414 23244 14962
rect 23204 14408 23256 14414
rect 23204 14350 23256 14356
rect 23308 14346 23336 15302
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 23388 14952 23440 14958
rect 23386 14920 23388 14929
rect 23440 14920 23442 14929
rect 23386 14855 23442 14864
rect 23386 14784 23442 14793
rect 23386 14719 23442 14728
rect 23400 14414 23428 14719
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 23296 14340 23348 14346
rect 23296 14282 23348 14288
rect 23202 14240 23258 14249
rect 23202 14175 23258 14184
rect 23216 13870 23244 14175
rect 23204 13864 23256 13870
rect 23204 13806 23256 13812
rect 23204 12640 23256 12646
rect 23204 12582 23256 12588
rect 23110 10160 23166 10169
rect 23110 10095 23166 10104
rect 23018 7576 23074 7585
rect 23018 7511 23074 7520
rect 22744 6724 22796 6730
rect 22744 6666 22796 6672
rect 23216 6633 23244 12582
rect 23308 10198 23336 14282
rect 23400 12782 23428 14350
rect 23492 12850 23520 14962
rect 23584 13394 23612 15370
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23480 12844 23532 12850
rect 23480 12786 23532 12792
rect 23388 12776 23440 12782
rect 23676 12730 23704 17614
rect 23940 16652 23992 16658
rect 23940 16594 23992 16600
rect 23756 16584 23808 16590
rect 23754 16552 23756 16561
rect 23808 16552 23810 16561
rect 23754 16487 23810 16496
rect 23952 16454 23980 16594
rect 24044 16561 24072 20318
rect 24308 20266 24360 20272
rect 24124 19848 24176 19854
rect 24124 19790 24176 19796
rect 24030 16552 24086 16561
rect 24030 16487 24086 16496
rect 23848 16448 23900 16454
rect 23848 16390 23900 16396
rect 23940 16448 23992 16454
rect 23940 16390 23992 16396
rect 23860 15162 23888 16390
rect 24032 15700 24084 15706
rect 24032 15642 24084 15648
rect 23848 15156 23900 15162
rect 23848 15098 23900 15104
rect 23940 15088 23992 15094
rect 23754 15056 23810 15065
rect 23940 15030 23992 15036
rect 23754 14991 23756 15000
rect 23808 14991 23810 15000
rect 23756 14962 23808 14968
rect 23846 13968 23902 13977
rect 23952 13938 23980 15030
rect 23846 13903 23848 13912
rect 23900 13903 23902 13912
rect 23940 13932 23992 13938
rect 23848 13874 23900 13880
rect 23940 13874 23992 13880
rect 23860 13410 23888 13874
rect 23860 13382 23980 13410
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 23388 12718 23440 12724
rect 23492 12702 23704 12730
rect 23756 12776 23808 12782
rect 23756 12718 23808 12724
rect 23492 12170 23520 12702
rect 23664 12640 23716 12646
rect 23664 12582 23716 12588
rect 23676 12434 23704 12582
rect 23584 12406 23704 12434
rect 23584 12238 23612 12406
rect 23572 12232 23624 12238
rect 23768 12209 23796 12718
rect 23572 12174 23624 12180
rect 23754 12200 23810 12209
rect 23480 12164 23532 12170
rect 23480 12106 23532 12112
rect 23492 11898 23520 12106
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23584 11218 23612 12174
rect 23754 12135 23810 12144
rect 23664 11824 23716 11830
rect 23662 11792 23664 11801
rect 23716 11792 23718 11801
rect 23662 11727 23718 11736
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 23480 11008 23532 11014
rect 23480 10950 23532 10956
rect 23492 10674 23520 10950
rect 23756 10804 23808 10810
rect 23756 10746 23808 10752
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 23388 10600 23440 10606
rect 23388 10542 23440 10548
rect 23296 10192 23348 10198
rect 23296 10134 23348 10140
rect 23296 8832 23348 8838
rect 23296 8774 23348 8780
rect 23308 8430 23336 8774
rect 23296 8424 23348 8430
rect 23296 8366 23348 8372
rect 23400 7410 23428 10542
rect 23492 10266 23520 10610
rect 23768 10266 23796 10746
rect 23480 10260 23532 10266
rect 23480 10202 23532 10208
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 23492 9382 23520 10202
rect 23860 9586 23888 13262
rect 23952 11354 23980 13382
rect 24044 12646 24072 15642
rect 24136 15638 24164 19790
rect 24216 19712 24268 19718
rect 24216 19654 24268 19660
rect 24228 19378 24256 19654
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 24216 18828 24268 18834
rect 24216 18770 24268 18776
rect 24228 18222 24256 18770
rect 24216 18216 24268 18222
rect 24216 18158 24268 18164
rect 24320 17610 24348 20266
rect 24412 17678 24440 21814
rect 24582 21720 24638 21729
rect 24582 21655 24638 21664
rect 24596 21622 24624 21655
rect 24584 21616 24636 21622
rect 24584 21558 24636 21564
rect 24492 21344 24544 21350
rect 24492 21286 24544 21292
rect 24504 21146 24532 21286
rect 24492 21140 24544 21146
rect 24492 21082 24544 21088
rect 24492 20936 24544 20942
rect 24492 20878 24544 20884
rect 24596 20890 24624 21558
rect 24688 21010 24716 22335
rect 24780 21554 24808 23122
rect 24768 21548 24820 21554
rect 24768 21490 24820 21496
rect 24768 21344 24820 21350
rect 24768 21286 24820 21292
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24504 19378 24532 20878
rect 24596 20862 24716 20890
rect 24582 20632 24638 20641
rect 24582 20567 24638 20576
rect 24596 19990 24624 20567
rect 24584 19984 24636 19990
rect 24584 19926 24636 19932
rect 24492 19372 24544 19378
rect 24492 19314 24544 19320
rect 24492 19236 24544 19242
rect 24492 19178 24544 19184
rect 24504 17921 24532 19178
rect 24688 18766 24716 20862
rect 24780 19854 24808 21286
rect 24872 20942 24900 23190
rect 24964 22642 24992 25094
rect 24952 22636 25004 22642
rect 24952 22578 25004 22584
rect 24964 22545 24992 22578
rect 25056 22574 25084 25638
rect 25148 23798 25176 26182
rect 25424 26042 25452 26182
rect 25412 26036 25464 26042
rect 25412 25978 25464 25984
rect 25424 25702 25452 25978
rect 25412 25696 25464 25702
rect 25412 25638 25464 25644
rect 25792 25498 25820 27066
rect 26436 26489 26464 27270
rect 27528 26920 27580 26926
rect 27526 26888 27528 26897
rect 27580 26888 27582 26897
rect 27448 26846 27526 26874
rect 27344 26784 27396 26790
rect 27344 26726 27396 26732
rect 26422 26480 26478 26489
rect 26422 26415 26478 26424
rect 26792 25900 26844 25906
rect 26792 25842 26844 25848
rect 25780 25492 25832 25498
rect 25780 25434 25832 25440
rect 26424 25492 26476 25498
rect 26424 25434 26476 25440
rect 25228 25424 25280 25430
rect 25228 25366 25280 25372
rect 26240 25424 26292 25430
rect 26240 25366 26292 25372
rect 25240 25265 25268 25366
rect 25780 25356 25832 25362
rect 25780 25298 25832 25304
rect 25226 25256 25282 25265
rect 25226 25191 25282 25200
rect 25504 24948 25556 24954
rect 25504 24890 25556 24896
rect 25516 24750 25544 24890
rect 25504 24744 25556 24750
rect 25504 24686 25556 24692
rect 25688 24744 25740 24750
rect 25688 24686 25740 24692
rect 25320 24676 25372 24682
rect 25320 24618 25372 24624
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 25136 23792 25188 23798
rect 25136 23734 25188 23740
rect 25148 22574 25176 23734
rect 25240 23118 25268 24210
rect 25228 23112 25280 23118
rect 25228 23054 25280 23060
rect 25044 22568 25096 22574
rect 24950 22536 25006 22545
rect 25044 22510 25096 22516
rect 25136 22568 25188 22574
rect 25136 22510 25188 22516
rect 24950 22471 25006 22480
rect 25332 22098 25360 24618
rect 25412 24608 25464 24614
rect 25412 24550 25464 24556
rect 25424 24177 25452 24550
rect 25410 24168 25466 24177
rect 25410 24103 25412 24112
rect 25464 24103 25466 24112
rect 25412 24074 25464 24080
rect 25410 24032 25466 24041
rect 25410 23967 25466 23976
rect 25424 23050 25452 23967
rect 25412 23044 25464 23050
rect 25412 22986 25464 22992
rect 25412 22500 25464 22506
rect 25412 22442 25464 22448
rect 25320 22092 25372 22098
rect 25320 22034 25372 22040
rect 25228 22024 25280 22030
rect 25134 21992 25190 22001
rect 25228 21966 25280 21972
rect 25424 21978 25452 22442
rect 25516 22166 25544 24686
rect 25596 24608 25648 24614
rect 25596 24550 25648 24556
rect 25608 24041 25636 24550
rect 25594 24032 25650 24041
rect 25594 23967 25650 23976
rect 25700 23866 25728 24686
rect 25688 23860 25740 23866
rect 25688 23802 25740 23808
rect 25792 23730 25820 25298
rect 26148 25152 26200 25158
rect 26148 25094 26200 25100
rect 26160 24614 26188 25094
rect 26148 24608 26200 24614
rect 26148 24550 26200 24556
rect 25964 24200 26016 24206
rect 25964 24142 26016 24148
rect 26054 24168 26110 24177
rect 25872 24064 25924 24070
rect 25872 24006 25924 24012
rect 25884 23866 25912 24006
rect 25872 23860 25924 23866
rect 25872 23802 25924 23808
rect 25596 23724 25648 23730
rect 25780 23724 25832 23730
rect 25648 23684 25728 23712
rect 25596 23666 25648 23672
rect 25594 23624 25650 23633
rect 25594 23559 25650 23568
rect 25608 22710 25636 23559
rect 25700 22778 25728 23684
rect 25780 23666 25832 23672
rect 25872 23656 25924 23662
rect 25778 23624 25834 23633
rect 25872 23598 25924 23604
rect 25778 23559 25834 23568
rect 25792 23186 25820 23559
rect 25780 23180 25832 23186
rect 25780 23122 25832 23128
rect 25688 22772 25740 22778
rect 25688 22714 25740 22720
rect 25596 22704 25648 22710
rect 25780 22704 25832 22710
rect 25596 22646 25648 22652
rect 25778 22672 25780 22681
rect 25832 22672 25834 22681
rect 25778 22607 25834 22616
rect 25596 22568 25648 22574
rect 25596 22510 25648 22516
rect 25504 22160 25556 22166
rect 25504 22102 25556 22108
rect 25134 21927 25190 21936
rect 24952 21616 25004 21622
rect 24952 21558 25004 21564
rect 24964 21350 24992 21558
rect 25042 21448 25098 21457
rect 25042 21383 25098 21392
rect 24952 21344 25004 21350
rect 24952 21286 25004 21292
rect 24952 21140 25004 21146
rect 24952 21082 25004 21088
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24872 20097 24900 20878
rect 24964 20330 24992 21082
rect 25056 20448 25084 21383
rect 25148 21146 25176 21927
rect 25136 21140 25188 21146
rect 25136 21082 25188 21088
rect 25240 20602 25268 21966
rect 25424 21950 25544 21978
rect 25412 21888 25464 21894
rect 25412 21830 25464 21836
rect 25424 21554 25452 21830
rect 25412 21548 25464 21554
rect 25412 21490 25464 21496
rect 25320 21072 25372 21078
rect 25320 21014 25372 21020
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 25056 20420 25268 20448
rect 24952 20324 25004 20330
rect 24952 20266 25004 20272
rect 25136 20324 25188 20330
rect 25136 20266 25188 20272
rect 25044 20256 25096 20262
rect 25044 20198 25096 20204
rect 24858 20088 24914 20097
rect 24858 20023 24914 20032
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24872 19689 24900 20023
rect 24858 19680 24914 19689
rect 24858 19615 24914 19624
rect 24950 19272 25006 19281
rect 24950 19207 25006 19216
rect 24858 19000 24914 19009
rect 24858 18935 24914 18944
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 24676 18760 24728 18766
rect 24676 18702 24728 18708
rect 24490 17912 24546 17921
rect 24596 17882 24624 18702
rect 24674 17912 24730 17921
rect 24490 17847 24546 17856
rect 24584 17876 24636 17882
rect 24674 17847 24730 17856
rect 24584 17818 24636 17824
rect 24400 17672 24452 17678
rect 24400 17614 24452 17620
rect 24308 17604 24360 17610
rect 24308 17546 24360 17552
rect 24490 17504 24546 17513
rect 24490 17439 24546 17448
rect 24504 16266 24532 17439
rect 24688 17202 24716 17847
rect 24768 17536 24820 17542
rect 24768 17478 24820 17484
rect 24676 17196 24728 17202
rect 24676 17138 24728 17144
rect 24676 16584 24728 16590
rect 24676 16526 24728 16532
rect 24320 16238 24532 16266
rect 24214 16008 24270 16017
rect 24214 15943 24216 15952
rect 24268 15943 24270 15952
rect 24216 15914 24268 15920
rect 24124 15632 24176 15638
rect 24124 15574 24176 15580
rect 24214 15600 24270 15609
rect 24214 15535 24270 15544
rect 24228 15065 24256 15535
rect 24214 15056 24270 15065
rect 24214 14991 24270 15000
rect 24214 14512 24270 14521
rect 24214 14447 24270 14456
rect 24228 14278 24256 14447
rect 24216 14272 24268 14278
rect 24216 14214 24268 14220
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24136 13190 24164 13874
rect 24124 13184 24176 13190
rect 24228 13161 24256 13874
rect 24124 13126 24176 13132
rect 24214 13152 24270 13161
rect 24136 12968 24164 13126
rect 24214 13087 24270 13096
rect 24136 12940 24256 12968
rect 24124 12844 24176 12850
rect 24124 12786 24176 12792
rect 24032 12640 24084 12646
rect 24032 12582 24084 12588
rect 24136 11694 24164 12786
rect 24228 12306 24256 12940
rect 24320 12646 24348 16238
rect 24492 16176 24544 16182
rect 24492 16118 24544 16124
rect 24400 15020 24452 15026
rect 24400 14962 24452 14968
rect 24308 12640 24360 12646
rect 24308 12582 24360 12588
rect 24216 12300 24268 12306
rect 24216 12242 24268 12248
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24124 11688 24176 11694
rect 24124 11630 24176 11636
rect 23940 11348 23992 11354
rect 23940 11290 23992 11296
rect 24032 11280 24084 11286
rect 24032 11222 24084 11228
rect 24044 11082 24072 11222
rect 24032 11076 24084 11082
rect 24032 11018 24084 11024
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 23570 9480 23626 9489
rect 23570 9415 23572 9424
rect 23624 9415 23626 9424
rect 23572 9386 23624 9392
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 23492 8634 23520 9318
rect 23480 8628 23532 8634
rect 23480 8570 23532 8576
rect 23388 7404 23440 7410
rect 23388 7346 23440 7352
rect 23202 6624 23258 6633
rect 23202 6559 23258 6568
rect 22008 5568 22060 5574
rect 22008 5510 22060 5516
rect 23584 4010 23612 9386
rect 23848 9104 23900 9110
rect 23848 9046 23900 9052
rect 23860 8838 23888 9046
rect 24136 8838 24164 11630
rect 24228 11558 24256 11698
rect 24216 11552 24268 11558
rect 24216 11494 24268 11500
rect 24228 10674 24256 11494
rect 24308 11348 24360 11354
rect 24308 11290 24360 11296
rect 24320 11121 24348 11290
rect 24306 11112 24362 11121
rect 24306 11047 24362 11056
rect 24320 10742 24348 11047
rect 24308 10736 24360 10742
rect 24308 10678 24360 10684
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 24412 10130 24440 14962
rect 24504 14618 24532 16118
rect 24584 15632 24636 15638
rect 24584 15574 24636 15580
rect 24492 14612 24544 14618
rect 24492 14554 24544 14560
rect 24596 14414 24624 15574
rect 24688 15502 24716 16526
rect 24780 15910 24808 17478
rect 24872 16153 24900 18935
rect 24964 18698 24992 19207
rect 24952 18692 25004 18698
rect 24952 18634 25004 18640
rect 24952 18352 25004 18358
rect 24950 18320 24952 18329
rect 25004 18320 25006 18329
rect 24950 18255 25006 18264
rect 25056 18193 25084 20198
rect 25042 18184 25098 18193
rect 25042 18119 25098 18128
rect 25148 17610 25176 20266
rect 25136 17604 25188 17610
rect 25136 17546 25188 17552
rect 25044 17264 25096 17270
rect 24950 17232 25006 17241
rect 25044 17206 25096 17212
rect 24950 17167 25006 17176
rect 24964 16794 24992 17167
rect 24952 16788 25004 16794
rect 24952 16730 25004 16736
rect 24964 16658 24992 16730
rect 24952 16652 25004 16658
rect 24952 16594 25004 16600
rect 24858 16144 24914 16153
rect 24858 16079 24914 16088
rect 24860 15972 24912 15978
rect 24860 15914 24912 15920
rect 24768 15904 24820 15910
rect 24768 15846 24820 15852
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24766 15328 24822 15337
rect 24766 15263 24822 15272
rect 24676 14952 24728 14958
rect 24676 14894 24728 14900
rect 24584 14408 24636 14414
rect 24584 14350 24636 14356
rect 24492 14272 24544 14278
rect 24492 14214 24544 14220
rect 24504 14074 24532 14214
rect 24492 14068 24544 14074
rect 24492 14010 24544 14016
rect 24584 14068 24636 14074
rect 24584 14010 24636 14016
rect 24596 13802 24624 14010
rect 24688 13841 24716 14894
rect 24674 13832 24730 13841
rect 24584 13796 24636 13802
rect 24674 13767 24730 13776
rect 24584 13738 24636 13744
rect 24676 13456 24728 13462
rect 24674 13424 24676 13433
rect 24728 13424 24730 13433
rect 24674 13359 24730 13368
rect 24780 13326 24808 15263
rect 24872 15094 24900 15914
rect 24860 15088 24912 15094
rect 24860 15030 24912 15036
rect 24952 14952 25004 14958
rect 24952 14894 25004 14900
rect 24858 14784 24914 14793
rect 24858 14719 24914 14728
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24584 12980 24636 12986
rect 24584 12922 24636 12928
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24596 12646 24624 12922
rect 24780 12753 24808 12922
rect 24766 12744 24822 12753
rect 24766 12679 24822 12688
rect 24872 12646 24900 14719
rect 24964 13841 24992 14894
rect 25056 14550 25084 17206
rect 25136 16516 25188 16522
rect 25136 16458 25188 16464
rect 25148 15638 25176 16458
rect 25240 16250 25268 20420
rect 25228 16244 25280 16250
rect 25228 16186 25280 16192
rect 25136 15632 25188 15638
rect 25332 15609 25360 21014
rect 25424 21010 25452 21490
rect 25516 21457 25544 21950
rect 25502 21448 25558 21457
rect 25502 21383 25558 21392
rect 25412 21004 25464 21010
rect 25412 20946 25464 20952
rect 25504 20596 25556 20602
rect 25608 20584 25636 22510
rect 25688 22500 25740 22506
rect 25688 22442 25740 22448
rect 25780 22500 25832 22506
rect 25780 22442 25832 22448
rect 25700 21554 25728 22442
rect 25792 22166 25820 22442
rect 25780 22160 25832 22166
rect 25780 22102 25832 22108
rect 25688 21548 25740 21554
rect 25688 21490 25740 21496
rect 25556 20556 25636 20584
rect 25504 20538 25556 20544
rect 25412 19916 25464 19922
rect 25412 19858 25464 19864
rect 25424 19786 25452 19858
rect 25412 19780 25464 19786
rect 25412 19722 25464 19728
rect 25608 19514 25636 20556
rect 25700 20924 25728 21490
rect 25884 21418 25912 23598
rect 25872 21412 25924 21418
rect 25872 21354 25924 21360
rect 25780 20936 25832 20942
rect 25700 20896 25780 20924
rect 25596 19508 25648 19514
rect 25596 19450 25648 19456
rect 25410 19272 25466 19281
rect 25410 19207 25466 19216
rect 25424 18358 25452 19207
rect 25596 18624 25648 18630
rect 25596 18566 25648 18572
rect 25608 18426 25636 18566
rect 25596 18420 25648 18426
rect 25596 18362 25648 18368
rect 25412 18352 25464 18358
rect 25412 18294 25464 18300
rect 25700 17882 25728 20896
rect 25780 20878 25832 20884
rect 25780 20392 25832 20398
rect 25976 20346 26004 24142
rect 26054 24103 26110 24112
rect 26068 23254 26096 24103
rect 26148 24064 26200 24070
rect 26148 24006 26200 24012
rect 26056 23248 26108 23254
rect 26056 23190 26108 23196
rect 26056 21888 26108 21894
rect 26056 21830 26108 21836
rect 26068 21486 26096 21830
rect 26056 21480 26108 21486
rect 26056 21422 26108 21428
rect 26056 20392 26108 20398
rect 25832 20340 26004 20346
rect 25780 20334 26004 20340
rect 25792 20318 26004 20334
rect 25778 20088 25834 20097
rect 25778 20023 25834 20032
rect 25688 17876 25740 17882
rect 25688 17818 25740 17824
rect 25410 17776 25466 17785
rect 25410 17711 25466 17720
rect 25424 15706 25452 17711
rect 25596 16652 25648 16658
rect 25596 16594 25648 16600
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25412 15700 25464 15706
rect 25412 15642 25464 15648
rect 25136 15574 25188 15580
rect 25318 15600 25374 15609
rect 25318 15535 25374 15544
rect 25320 14952 25372 14958
rect 25320 14894 25372 14900
rect 25136 14612 25188 14618
rect 25136 14554 25188 14560
rect 25044 14544 25096 14550
rect 25044 14486 25096 14492
rect 25148 14362 25176 14554
rect 25056 14334 25176 14362
rect 25332 14346 25360 14894
rect 25320 14340 25372 14346
rect 24950 13832 25006 13841
rect 24950 13767 25006 13776
rect 24950 13288 25006 13297
rect 24950 13223 24952 13232
rect 25004 13223 25006 13232
rect 24952 13194 25004 13200
rect 24952 12776 25004 12782
rect 24952 12718 25004 12724
rect 24584 12640 24636 12646
rect 24584 12582 24636 12588
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 24596 12442 24624 12582
rect 24674 12472 24730 12481
rect 24584 12436 24636 12442
rect 24674 12407 24730 12416
rect 24584 12378 24636 12384
rect 24688 12306 24716 12407
rect 24964 12374 24992 12718
rect 24768 12368 24820 12374
rect 24766 12336 24768 12345
rect 24952 12368 25004 12374
rect 24820 12336 24822 12345
rect 24676 12300 24728 12306
rect 24766 12271 24822 12280
rect 24872 12328 24952 12356
rect 24676 12242 24728 12248
rect 24674 12200 24730 12209
rect 24584 12164 24636 12170
rect 24504 12124 24584 12152
rect 24504 10198 24532 12124
rect 24674 12135 24730 12144
rect 24584 12106 24636 12112
rect 24584 11892 24636 11898
rect 24584 11834 24636 11840
rect 24596 11762 24624 11834
rect 24584 11756 24636 11762
rect 24584 11698 24636 11704
rect 24596 10266 24624 11698
rect 24688 11694 24716 12135
rect 24872 11744 24900 12328
rect 24952 12310 25004 12316
rect 25056 11762 25084 14334
rect 25320 14282 25372 14288
rect 25332 14090 25360 14282
rect 25240 14062 25360 14090
rect 25240 14006 25268 14062
rect 25228 14000 25280 14006
rect 25228 13942 25280 13948
rect 25136 13184 25188 13190
rect 25424 13172 25452 15642
rect 25516 13274 25544 16186
rect 25608 13530 25636 16594
rect 25688 15156 25740 15162
rect 25688 15098 25740 15104
rect 25596 13524 25648 13530
rect 25596 13466 25648 13472
rect 25516 13246 25636 13274
rect 25424 13144 25544 13172
rect 25136 13126 25188 13132
rect 25148 12753 25176 13126
rect 25410 13016 25466 13025
rect 25410 12951 25466 12960
rect 25424 12918 25452 12951
rect 25412 12912 25464 12918
rect 25412 12854 25464 12860
rect 25228 12844 25280 12850
rect 25228 12786 25280 12792
rect 25134 12744 25190 12753
rect 25134 12679 25190 12688
rect 25240 12646 25268 12786
rect 25412 12708 25464 12714
rect 25412 12650 25464 12656
rect 25228 12640 25280 12646
rect 25228 12582 25280 12588
rect 25320 12640 25372 12646
rect 25320 12582 25372 12588
rect 25136 12436 25188 12442
rect 25136 12378 25188 12384
rect 25148 11830 25176 12378
rect 25228 12300 25280 12306
rect 25228 12242 25280 12248
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 24780 11716 24900 11744
rect 25044 11756 25096 11762
rect 24676 11688 24728 11694
rect 24676 11630 24728 11636
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24688 10441 24716 11086
rect 24780 10810 24808 11716
rect 25044 11698 25096 11704
rect 25136 11688 25188 11694
rect 25136 11630 25188 11636
rect 24860 11620 24912 11626
rect 24860 11562 24912 11568
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24766 10704 24822 10713
rect 24766 10639 24822 10648
rect 24780 10538 24808 10639
rect 24768 10532 24820 10538
rect 24768 10474 24820 10480
rect 24674 10432 24730 10441
rect 24674 10367 24730 10376
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24492 10192 24544 10198
rect 24492 10134 24544 10140
rect 24400 10124 24452 10130
rect 24400 10066 24452 10072
rect 24688 9722 24716 10367
rect 24676 9716 24728 9722
rect 24676 9658 24728 9664
rect 24872 9636 24900 11562
rect 25042 11384 25098 11393
rect 25042 11319 25098 11328
rect 25056 11150 25084 11319
rect 25044 11144 25096 11150
rect 25044 11086 25096 11092
rect 24950 10704 25006 10713
rect 24950 10639 24952 10648
rect 25004 10639 25006 10648
rect 24952 10610 25004 10616
rect 24780 9608 24900 9636
rect 24780 9450 24808 9608
rect 24768 9444 24820 9450
rect 24768 9386 24820 9392
rect 24400 9376 24452 9382
rect 24400 9318 24452 9324
rect 23848 8832 23900 8838
rect 23848 8774 23900 8780
rect 24124 8832 24176 8838
rect 24124 8774 24176 8780
rect 23860 5545 23888 8774
rect 23846 5536 23902 5545
rect 23846 5471 23902 5480
rect 23572 4004 23624 4010
rect 23572 3946 23624 3952
rect 21914 2408 21970 2417
rect 21914 2343 21970 2352
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 14554 2000 14610 2009
rect 14554 1935 14610 1944
rect 17972 800 18000 2246
rect 20214 2204 20522 2224
rect 20214 2202 20220 2204
rect 20276 2202 20300 2204
rect 20356 2202 20380 2204
rect 20436 2202 20460 2204
rect 20516 2202 20522 2204
rect 20276 2150 20278 2202
rect 20458 2150 20460 2202
rect 20214 2148 20220 2150
rect 20276 2148 20300 2150
rect 20356 2148 20380 2150
rect 20436 2148 20460 2150
rect 20516 2148 20522 2150
rect 20214 2128 20522 2148
rect 24412 2106 24440 9318
rect 24964 8634 24992 10610
rect 25056 9518 25084 11086
rect 25044 9512 25096 9518
rect 25044 9454 25096 9460
rect 25148 9110 25176 11630
rect 25240 10266 25268 12242
rect 25228 10260 25280 10266
rect 25228 10202 25280 10208
rect 25332 10062 25360 12582
rect 25424 11150 25452 12650
rect 25412 11144 25464 11150
rect 25412 11086 25464 11092
rect 25412 10600 25464 10606
rect 25412 10542 25464 10548
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25424 9654 25452 10542
rect 25412 9648 25464 9654
rect 25412 9590 25464 9596
rect 25136 9104 25188 9110
rect 25136 9046 25188 9052
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 25516 8566 25544 13144
rect 25608 12646 25636 13246
rect 25596 12640 25648 12646
rect 25596 12582 25648 12588
rect 25608 12442 25636 12582
rect 25596 12436 25648 12442
rect 25596 12378 25648 12384
rect 25594 11384 25650 11393
rect 25594 11319 25596 11328
rect 25648 11319 25650 11328
rect 25596 11290 25648 11296
rect 25596 11144 25648 11150
rect 25596 11086 25648 11092
rect 25504 8560 25556 8566
rect 25504 8502 25556 8508
rect 25608 8480 25636 11086
rect 25700 8945 25728 15098
rect 25792 14929 25820 20023
rect 25976 19514 26004 20318
rect 26054 20360 26056 20369
rect 26108 20360 26110 20369
rect 26054 20295 26110 20304
rect 25964 19508 26016 19514
rect 25964 19450 26016 19456
rect 26056 19168 26108 19174
rect 26056 19110 26108 19116
rect 26068 18970 26096 19110
rect 26056 18964 26108 18970
rect 26056 18906 26108 18912
rect 26054 18864 26110 18873
rect 26054 18799 26110 18808
rect 25872 18420 25924 18426
rect 25872 18362 25924 18368
rect 25778 14920 25834 14929
rect 25778 14855 25834 14864
rect 25780 13388 25832 13394
rect 25780 13330 25832 13336
rect 25792 11762 25820 13330
rect 25884 12442 25912 18362
rect 26068 17746 26096 18799
rect 26056 17740 26108 17746
rect 26056 17682 26108 17688
rect 26054 17232 26110 17241
rect 26054 17167 26056 17176
rect 26108 17167 26110 17176
rect 26056 17138 26108 17144
rect 25964 16652 26016 16658
rect 25964 16594 26016 16600
rect 25976 15434 26004 16594
rect 26160 16182 26188 24006
rect 26252 22953 26280 25366
rect 26332 24608 26384 24614
rect 26332 24550 26384 24556
rect 26344 23798 26372 24550
rect 26332 23792 26384 23798
rect 26332 23734 26384 23740
rect 26330 23216 26386 23225
rect 26330 23151 26332 23160
rect 26384 23151 26386 23160
rect 26332 23122 26384 23128
rect 26330 23080 26386 23089
rect 26330 23015 26386 23024
rect 26238 22944 26294 22953
rect 26238 22879 26294 22888
rect 26238 22672 26294 22681
rect 26238 22607 26294 22616
rect 26252 22234 26280 22607
rect 26240 22228 26292 22234
rect 26240 22170 26292 22176
rect 26252 22098 26280 22170
rect 26240 22092 26292 22098
rect 26240 22034 26292 22040
rect 26344 22030 26372 23015
rect 26436 22642 26464 25434
rect 26516 24608 26568 24614
rect 26516 24550 26568 24556
rect 26528 23526 26556 24550
rect 26700 24132 26752 24138
rect 26700 24074 26752 24080
rect 26608 23724 26660 23730
rect 26608 23666 26660 23672
rect 26516 23520 26568 23526
rect 26516 23462 26568 23468
rect 26424 22636 26476 22642
rect 26424 22578 26476 22584
rect 26528 22438 26556 23462
rect 26424 22432 26476 22438
rect 26424 22374 26476 22380
rect 26516 22432 26568 22438
rect 26516 22374 26568 22380
rect 26332 22024 26384 22030
rect 26332 21966 26384 21972
rect 26332 21888 26384 21894
rect 26332 21830 26384 21836
rect 26344 21690 26372 21830
rect 26332 21684 26384 21690
rect 26332 21626 26384 21632
rect 26332 21548 26384 21554
rect 26332 21490 26384 21496
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 26252 19446 26280 21286
rect 26344 20942 26372 21490
rect 26332 20936 26384 20942
rect 26332 20878 26384 20884
rect 26240 19440 26292 19446
rect 26240 19382 26292 19388
rect 26240 16992 26292 16998
rect 26240 16934 26292 16940
rect 26148 16176 26200 16182
rect 26148 16118 26200 16124
rect 25964 15428 26016 15434
rect 25964 15370 26016 15376
rect 25976 14346 26004 15370
rect 26148 15360 26200 15366
rect 26148 15302 26200 15308
rect 25964 14340 26016 14346
rect 25964 14282 26016 14288
rect 25976 14074 26004 14282
rect 25964 14068 26016 14074
rect 25964 14010 26016 14016
rect 26056 13728 26108 13734
rect 26056 13670 26108 13676
rect 25964 13184 26016 13190
rect 25964 13126 26016 13132
rect 25976 12714 26004 13126
rect 25964 12708 26016 12714
rect 25964 12650 26016 12656
rect 26068 12594 26096 13670
rect 26160 13326 26188 15302
rect 26252 14958 26280 16934
rect 26436 16114 26464 22374
rect 26516 22228 26568 22234
rect 26516 22170 26568 22176
rect 26528 21894 26556 22170
rect 26620 22166 26648 23666
rect 26712 23497 26740 24074
rect 26698 23488 26754 23497
rect 26698 23423 26754 23432
rect 26700 23112 26752 23118
rect 26700 23054 26752 23060
rect 26712 22545 26740 23054
rect 26698 22536 26754 22545
rect 26698 22471 26754 22480
rect 26608 22160 26660 22166
rect 26608 22102 26660 22108
rect 26804 22094 26832 25842
rect 27252 25764 27304 25770
rect 27252 25706 27304 25712
rect 27160 25696 27212 25702
rect 27160 25638 27212 25644
rect 26884 25288 26936 25294
rect 26884 25230 26936 25236
rect 26896 24721 26924 25230
rect 27172 25158 27200 25638
rect 27264 25265 27292 25706
rect 27250 25256 27306 25265
rect 27250 25191 27306 25200
rect 27160 25152 27212 25158
rect 27160 25094 27212 25100
rect 26882 24712 26938 24721
rect 26882 24647 26938 24656
rect 27172 24410 27200 25094
rect 27160 24404 27212 24410
rect 27160 24346 27212 24352
rect 27252 24404 27304 24410
rect 27252 24346 27304 24352
rect 26976 24132 27028 24138
rect 26976 24074 27028 24080
rect 26884 24064 26936 24070
rect 26882 24032 26884 24041
rect 26936 24032 26938 24041
rect 26882 23967 26938 23976
rect 26882 23080 26938 23089
rect 26882 23015 26884 23024
rect 26936 23015 26938 23024
rect 26884 22986 26936 22992
rect 26882 22944 26938 22953
rect 26882 22879 26938 22888
rect 26896 22710 26924 22879
rect 26884 22704 26936 22710
rect 26884 22646 26936 22652
rect 26988 22234 27016 24074
rect 27172 23712 27200 24346
rect 27264 24206 27292 24346
rect 27356 24313 27384 26726
rect 27448 24585 27476 26846
rect 27526 26823 27582 26832
rect 28356 26784 28408 26790
rect 28356 26726 28408 26732
rect 28368 26382 28396 26726
rect 28446 26616 28502 26625
rect 28446 26551 28502 26560
rect 27712 26376 27764 26382
rect 27618 26344 27674 26353
rect 27712 26318 27764 26324
rect 28356 26376 28408 26382
rect 28356 26318 28408 26324
rect 27618 26279 27674 26288
rect 27528 24812 27580 24818
rect 27528 24754 27580 24760
rect 27434 24576 27490 24585
rect 27434 24511 27490 24520
rect 27436 24336 27488 24342
rect 27342 24304 27398 24313
rect 27436 24278 27488 24284
rect 27342 24239 27398 24248
rect 27356 24206 27384 24239
rect 27252 24200 27304 24206
rect 27252 24142 27304 24148
rect 27344 24200 27396 24206
rect 27344 24142 27396 24148
rect 27356 24041 27384 24142
rect 27342 24032 27398 24041
rect 27342 23967 27398 23976
rect 27342 23896 27398 23905
rect 27342 23831 27398 23840
rect 27252 23724 27304 23730
rect 27172 23684 27252 23712
rect 27252 23666 27304 23672
rect 27158 23624 27214 23633
rect 27158 23559 27160 23568
rect 27212 23559 27214 23568
rect 27160 23530 27212 23536
rect 27264 23508 27292 23666
rect 27356 23662 27384 23831
rect 27344 23656 27396 23662
rect 27344 23598 27396 23604
rect 27344 23520 27396 23526
rect 27264 23480 27344 23508
rect 27344 23462 27396 23468
rect 27066 23352 27122 23361
rect 27066 23287 27122 23296
rect 26976 22228 27028 22234
rect 26976 22170 27028 22176
rect 26804 22066 26924 22094
rect 26608 22024 26660 22030
rect 26608 21966 26660 21972
rect 26516 21888 26568 21894
rect 26516 21830 26568 21836
rect 26516 21616 26568 21622
rect 26516 21558 26568 21564
rect 26424 16108 26476 16114
rect 26424 16050 26476 16056
rect 26424 15564 26476 15570
rect 26424 15506 26476 15512
rect 26330 15192 26386 15201
rect 26330 15127 26386 15136
rect 26240 14952 26292 14958
rect 26240 14894 26292 14900
rect 26238 14104 26294 14113
rect 26238 14039 26294 14048
rect 26252 13841 26280 14039
rect 26238 13832 26294 13841
rect 26238 13767 26294 13776
rect 26148 13320 26200 13326
rect 26148 13262 26200 13268
rect 26240 13252 26292 13258
rect 26240 13194 26292 13200
rect 25976 12566 26096 12594
rect 25872 12436 25924 12442
rect 25872 12378 25924 12384
rect 25976 12306 26004 12566
rect 26054 12472 26110 12481
rect 26054 12407 26110 12416
rect 26068 12374 26096 12407
rect 26056 12368 26108 12374
rect 26056 12310 26108 12316
rect 25964 12300 26016 12306
rect 25964 12242 26016 12248
rect 25872 12232 25924 12238
rect 25872 12174 25924 12180
rect 25780 11756 25832 11762
rect 25780 11698 25832 11704
rect 25792 11014 25820 11698
rect 25884 11354 25912 12174
rect 25964 12096 26016 12102
rect 25964 12038 26016 12044
rect 25872 11348 25924 11354
rect 25872 11290 25924 11296
rect 25780 11008 25832 11014
rect 25780 10950 25832 10956
rect 25792 10674 25820 10950
rect 25780 10668 25832 10674
rect 25780 10610 25832 10616
rect 25792 9178 25820 10610
rect 25872 10260 25924 10266
rect 25872 10202 25924 10208
rect 25884 10062 25912 10202
rect 25872 10056 25924 10062
rect 25872 9998 25924 10004
rect 25976 9654 26004 12038
rect 25964 9648 26016 9654
rect 25964 9590 26016 9596
rect 25780 9172 25832 9178
rect 25780 9114 25832 9120
rect 25686 8936 25742 8945
rect 25686 8871 25742 8880
rect 25780 8492 25832 8498
rect 25608 8452 25780 8480
rect 25780 8434 25832 8440
rect 24582 8120 24638 8129
rect 24582 8055 24638 8064
rect 24766 8120 24822 8129
rect 24766 8055 24768 8064
rect 24596 6866 24624 8055
rect 24820 8055 24822 8064
rect 24768 8026 24820 8032
rect 24584 6860 24636 6866
rect 24584 6802 24636 6808
rect 24780 2774 24808 8026
rect 25504 7744 25556 7750
rect 25504 7686 25556 7692
rect 24858 3360 24914 3369
rect 24858 3295 24914 3304
rect 24596 2746 24808 2774
rect 24596 2553 24624 2746
rect 24582 2544 24638 2553
rect 24872 2514 24900 3295
rect 24582 2479 24638 2488
rect 24860 2508 24912 2514
rect 24860 2450 24912 2456
rect 24400 2100 24452 2106
rect 24400 2042 24452 2048
rect 25516 2038 25544 7686
rect 25792 4185 25820 8434
rect 25962 8120 26018 8129
rect 26068 8090 26096 12310
rect 26252 12073 26280 13194
rect 26344 12306 26372 15127
rect 26436 14550 26464 15506
rect 26424 14544 26476 14550
rect 26424 14486 26476 14492
rect 26422 14104 26478 14113
rect 26422 14039 26478 14048
rect 26436 13870 26464 14039
rect 26424 13864 26476 13870
rect 26424 13806 26476 13812
rect 26422 13016 26478 13025
rect 26422 12951 26424 12960
rect 26476 12951 26478 12960
rect 26424 12922 26476 12928
rect 26424 12368 26476 12374
rect 26424 12310 26476 12316
rect 26332 12300 26384 12306
rect 26332 12242 26384 12248
rect 26238 12064 26294 12073
rect 26238 11999 26294 12008
rect 26238 11928 26294 11937
rect 26436 11898 26464 12310
rect 26238 11863 26294 11872
rect 26424 11892 26476 11898
rect 26148 11756 26200 11762
rect 26148 11698 26200 11704
rect 26160 11393 26188 11698
rect 26252 11558 26280 11863
rect 26424 11834 26476 11840
rect 26332 11824 26384 11830
rect 26332 11766 26384 11772
rect 26344 11558 26372 11766
rect 26424 11620 26476 11626
rect 26424 11562 26476 11568
rect 26240 11552 26292 11558
rect 26240 11494 26292 11500
rect 26332 11552 26384 11558
rect 26332 11494 26384 11500
rect 26146 11384 26202 11393
rect 26146 11319 26202 11328
rect 26332 11212 26384 11218
rect 26332 11154 26384 11160
rect 26148 11076 26200 11082
rect 26148 11018 26200 11024
rect 26160 10674 26188 11018
rect 26148 10668 26200 10674
rect 26148 10610 26200 10616
rect 26160 9722 26188 10610
rect 26344 10470 26372 11154
rect 26436 11121 26464 11562
rect 26422 11112 26478 11121
rect 26422 11047 26478 11056
rect 26332 10464 26384 10470
rect 26332 10406 26384 10412
rect 26238 10296 26294 10305
rect 26238 10231 26240 10240
rect 26292 10231 26294 10240
rect 26240 10202 26292 10208
rect 26148 9716 26200 9722
rect 26148 9658 26200 9664
rect 26240 9580 26292 9586
rect 26240 9522 26292 9528
rect 26252 9432 26280 9522
rect 26332 9512 26384 9518
rect 26332 9454 26384 9460
rect 26160 9404 26280 9432
rect 25962 8055 25964 8064
rect 26016 8055 26018 8064
rect 26056 8084 26108 8090
rect 25964 8026 26016 8032
rect 26056 8026 26108 8032
rect 25872 7540 25924 7546
rect 25872 7482 25924 7488
rect 25778 4176 25834 4185
rect 25778 4111 25834 4120
rect 25884 2514 25912 7482
rect 25976 2774 26004 8026
rect 26160 7750 26188 9404
rect 26344 8634 26372 9454
rect 26424 9444 26476 9450
rect 26424 9386 26476 9392
rect 26436 8906 26464 9386
rect 26528 9178 26556 21558
rect 26620 21010 26648 21966
rect 26896 21894 26924 22066
rect 27080 22001 27108 23287
rect 27252 22772 27304 22778
rect 27252 22714 27304 22720
rect 27264 22642 27292 22714
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 27252 22636 27304 22642
rect 27252 22578 27304 22584
rect 27172 22166 27200 22578
rect 27356 22409 27384 23462
rect 27342 22400 27398 22409
rect 27342 22335 27398 22344
rect 27342 22264 27398 22273
rect 27342 22199 27398 22208
rect 27160 22160 27212 22166
rect 27160 22102 27212 22108
rect 27066 21992 27122 22001
rect 27066 21927 27122 21936
rect 26884 21888 26936 21894
rect 26884 21830 26936 21836
rect 26792 21344 26844 21350
rect 26792 21286 26844 21292
rect 27068 21344 27120 21350
rect 27068 21286 27120 21292
rect 27250 21312 27306 21321
rect 26608 21004 26660 21010
rect 26608 20946 26660 20952
rect 26804 20874 26832 21286
rect 26976 21072 27028 21078
rect 26976 21014 27028 21020
rect 26884 20936 26936 20942
rect 26884 20878 26936 20884
rect 26792 20868 26844 20874
rect 26792 20810 26844 20816
rect 26700 20596 26752 20602
rect 26700 20538 26752 20544
rect 26608 20460 26660 20466
rect 26608 20402 26660 20408
rect 26620 19922 26648 20402
rect 26712 20398 26740 20538
rect 26700 20392 26752 20398
rect 26700 20334 26752 20340
rect 26698 19952 26754 19961
rect 26608 19916 26660 19922
rect 26698 19887 26700 19896
rect 26608 19858 26660 19864
rect 26752 19887 26754 19896
rect 26700 19858 26752 19864
rect 26620 17202 26648 19858
rect 26700 19712 26752 19718
rect 26804 19700 26832 20810
rect 26896 20534 26924 20878
rect 26884 20528 26936 20534
rect 26884 20470 26936 20476
rect 26896 19786 26924 20470
rect 26988 20466 27016 21014
rect 26976 20460 27028 20466
rect 26976 20402 27028 20408
rect 26884 19780 26936 19786
rect 26884 19722 26936 19728
rect 26752 19672 26832 19700
rect 26700 19654 26752 19660
rect 27080 18737 27108 21286
rect 27250 21247 27306 21256
rect 27264 21146 27292 21247
rect 27252 21140 27304 21146
rect 27252 21082 27304 21088
rect 27264 20505 27292 21082
rect 27250 20496 27306 20505
rect 27250 20431 27306 20440
rect 27356 20398 27384 22199
rect 27344 20392 27396 20398
rect 27344 20334 27396 20340
rect 27158 20224 27214 20233
rect 27158 20159 27214 20168
rect 27172 19990 27200 20159
rect 27160 19984 27212 19990
rect 27448 19972 27476 24278
rect 27540 22710 27568 24754
rect 27632 23730 27660 26279
rect 27724 25362 27752 26318
rect 28264 26308 28316 26314
rect 28264 26250 28316 26256
rect 28080 26240 28132 26246
rect 28080 26182 28132 26188
rect 27804 25968 27856 25974
rect 27804 25910 27856 25916
rect 27712 25356 27764 25362
rect 27712 25298 27764 25304
rect 27724 24886 27752 25298
rect 27712 24880 27764 24886
rect 27712 24822 27764 24828
rect 27712 24676 27764 24682
rect 27712 24618 27764 24624
rect 27620 23724 27672 23730
rect 27620 23666 27672 23672
rect 27620 23520 27672 23526
rect 27620 23462 27672 23468
rect 27632 23186 27660 23462
rect 27620 23180 27672 23186
rect 27620 23122 27672 23128
rect 27620 23044 27672 23050
rect 27620 22986 27672 22992
rect 27632 22778 27660 22986
rect 27620 22772 27672 22778
rect 27620 22714 27672 22720
rect 27528 22704 27580 22710
rect 27528 22646 27580 22652
rect 27528 22432 27580 22438
rect 27528 22374 27580 22380
rect 27540 22098 27568 22374
rect 27528 22092 27580 22098
rect 27528 22034 27580 22040
rect 27620 21684 27672 21690
rect 27540 21644 27620 21672
rect 27540 21486 27568 21644
rect 27620 21626 27672 21632
rect 27618 21584 27674 21593
rect 27618 21519 27620 21528
rect 27672 21519 27674 21528
rect 27620 21490 27672 21496
rect 27528 21480 27580 21486
rect 27528 21422 27580 21428
rect 27212 19944 27476 19972
rect 27160 19926 27212 19932
rect 27448 19689 27476 19944
rect 27158 19680 27214 19689
rect 27158 19615 27214 19624
rect 27434 19680 27490 19689
rect 27434 19615 27490 19624
rect 27066 18728 27122 18737
rect 26976 18692 27028 18698
rect 27066 18663 27122 18672
rect 26976 18634 27028 18640
rect 26608 17196 26660 17202
rect 26608 17138 26660 17144
rect 26792 17196 26844 17202
rect 26792 17138 26844 17144
rect 26698 16552 26754 16561
rect 26698 16487 26754 16496
rect 26712 16454 26740 16487
rect 26700 16448 26752 16454
rect 26700 16390 26752 16396
rect 26606 15736 26662 15745
rect 26606 15671 26662 15680
rect 26620 11830 26648 15671
rect 26804 15570 26832 17138
rect 26792 15564 26844 15570
rect 26792 15506 26844 15512
rect 26804 15026 26832 15506
rect 26792 15020 26844 15026
rect 26792 14962 26844 14968
rect 26700 14816 26752 14822
rect 26700 14758 26752 14764
rect 26608 11824 26660 11830
rect 26608 11766 26660 11772
rect 26712 10674 26740 14758
rect 26804 13938 26832 14962
rect 26884 14544 26936 14550
rect 26884 14486 26936 14492
rect 26792 13932 26844 13938
rect 26792 13874 26844 13880
rect 26790 13560 26846 13569
rect 26790 13495 26846 13504
rect 26804 12442 26832 13495
rect 26792 12436 26844 12442
rect 26792 12378 26844 12384
rect 26792 12300 26844 12306
rect 26792 12242 26844 12248
rect 26804 12170 26832 12242
rect 26896 12209 26924 14486
rect 26988 13433 27016 18634
rect 27172 18612 27200 19615
rect 27436 19372 27488 19378
rect 27436 19314 27488 19320
rect 27252 18760 27304 18766
rect 27250 18728 27252 18737
rect 27304 18728 27306 18737
rect 27250 18663 27306 18672
rect 27172 18584 27292 18612
rect 27160 18216 27212 18222
rect 27160 18158 27212 18164
rect 27068 17604 27120 17610
rect 27068 17546 27120 17552
rect 26974 13424 27030 13433
rect 26974 13359 27030 13368
rect 26976 13320 27028 13326
rect 26976 13262 27028 13268
rect 26988 12986 27016 13262
rect 26976 12980 27028 12986
rect 26976 12922 27028 12928
rect 26882 12200 26938 12209
rect 26792 12164 26844 12170
rect 26882 12135 26938 12144
rect 26792 12106 26844 12112
rect 26790 11656 26846 11665
rect 26790 11591 26846 11600
rect 26804 11286 26832 11591
rect 26792 11280 26844 11286
rect 26792 11222 26844 11228
rect 26792 11144 26844 11150
rect 26792 11086 26844 11092
rect 26804 10742 26832 11086
rect 26792 10736 26844 10742
rect 26792 10678 26844 10684
rect 26700 10668 26752 10674
rect 26700 10610 26752 10616
rect 26700 10056 26752 10062
rect 26700 9998 26752 10004
rect 26516 9172 26568 9178
rect 26516 9114 26568 9120
rect 26528 8906 26556 9114
rect 26424 8900 26476 8906
rect 26424 8842 26476 8848
rect 26516 8900 26568 8906
rect 26516 8842 26568 8848
rect 26332 8628 26384 8634
rect 26332 8570 26384 8576
rect 26238 8392 26294 8401
rect 26238 8327 26294 8336
rect 26148 7744 26200 7750
rect 26148 7686 26200 7692
rect 26252 7546 26280 8327
rect 26436 7546 26464 8842
rect 26240 7540 26292 7546
rect 26240 7482 26292 7488
rect 26424 7540 26476 7546
rect 26424 7482 26476 7488
rect 26712 7206 26740 9998
rect 26804 9994 26832 10678
rect 26792 9988 26844 9994
rect 26792 9930 26844 9936
rect 26896 9586 26924 12135
rect 27080 11121 27108 17546
rect 27172 16590 27200 18158
rect 27264 16674 27292 18584
rect 27344 17264 27396 17270
rect 27344 17206 27396 17212
rect 27356 16833 27384 17206
rect 27342 16824 27398 16833
rect 27342 16759 27398 16768
rect 27264 16646 27384 16674
rect 27160 16584 27212 16590
rect 27160 16526 27212 16532
rect 27172 16114 27200 16526
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27158 15872 27214 15881
rect 27158 15807 27214 15816
rect 27172 14278 27200 15807
rect 27252 15496 27304 15502
rect 27252 15438 27304 15444
rect 27160 14272 27212 14278
rect 27160 14214 27212 14220
rect 27160 13932 27212 13938
rect 27160 13874 27212 13880
rect 27172 12238 27200 13874
rect 27160 12232 27212 12238
rect 27160 12174 27212 12180
rect 27066 11112 27122 11121
rect 26976 11076 27028 11082
rect 27066 11047 27122 11056
rect 26976 11018 27028 11024
rect 26988 10577 27016 11018
rect 26974 10568 27030 10577
rect 26974 10503 27030 10512
rect 26884 9580 26936 9586
rect 26884 9522 26936 9528
rect 26988 8974 27016 10503
rect 27172 10452 27200 12174
rect 27264 10606 27292 15438
rect 27356 14550 27384 16646
rect 27344 14544 27396 14550
rect 27344 14486 27396 14492
rect 27342 14240 27398 14249
rect 27342 14175 27398 14184
rect 27356 14006 27384 14175
rect 27344 14000 27396 14006
rect 27344 13942 27396 13948
rect 27344 13524 27396 13530
rect 27344 13466 27396 13472
rect 27356 12986 27384 13466
rect 27344 12980 27396 12986
rect 27344 12922 27396 12928
rect 27344 12776 27396 12782
rect 27344 12718 27396 12724
rect 27356 12345 27384 12718
rect 27342 12336 27398 12345
rect 27342 12271 27398 12280
rect 27342 11384 27398 11393
rect 27342 11319 27344 11328
rect 27396 11319 27398 11328
rect 27344 11290 27396 11296
rect 27252 10600 27304 10606
rect 27252 10542 27304 10548
rect 27344 10464 27396 10470
rect 27172 10424 27344 10452
rect 27344 10406 27396 10412
rect 27356 10146 27384 10406
rect 27448 10266 27476 19314
rect 27528 17536 27580 17542
rect 27528 17478 27580 17484
rect 27540 16726 27568 17478
rect 27724 17338 27752 24618
rect 27816 23662 27844 25910
rect 28092 25702 28120 26182
rect 28080 25696 28132 25702
rect 28080 25638 28132 25644
rect 27896 25152 27948 25158
rect 27896 25094 27948 25100
rect 27804 23656 27856 23662
rect 27804 23598 27856 23604
rect 27816 22574 27844 23598
rect 27804 22568 27856 22574
rect 27804 22510 27856 22516
rect 27816 21690 27844 22510
rect 27908 22234 27936 25094
rect 28092 24274 28120 25638
rect 28172 25288 28224 25294
rect 28172 25230 28224 25236
rect 28080 24268 28132 24274
rect 28080 24210 28132 24216
rect 27986 24168 28042 24177
rect 27986 24103 28042 24112
rect 28000 24070 28028 24103
rect 27988 24064 28040 24070
rect 27988 24006 28040 24012
rect 27986 23488 28042 23497
rect 27986 23423 28042 23432
rect 28000 23322 28028 23423
rect 28184 23361 28212 25230
rect 28276 24138 28304 26250
rect 28368 25974 28396 26318
rect 28356 25968 28408 25974
rect 28356 25910 28408 25916
rect 28460 25242 28488 26551
rect 28552 25770 28580 27270
rect 28644 27062 28672 27406
rect 28814 27367 28870 27376
rect 29644 27396 29696 27402
rect 28632 27056 28684 27062
rect 28632 26998 28684 27004
rect 28540 25764 28592 25770
rect 28540 25706 28592 25712
rect 28368 25214 28488 25242
rect 28264 24132 28316 24138
rect 28264 24074 28316 24080
rect 28262 24032 28318 24041
rect 28262 23967 28318 23976
rect 28276 23526 28304 23967
rect 28264 23520 28316 23526
rect 28264 23462 28316 23468
rect 28170 23352 28226 23361
rect 27988 23316 28040 23322
rect 28170 23287 28226 23296
rect 27988 23258 28040 23264
rect 28184 23118 28212 23287
rect 27988 23112 28040 23118
rect 27986 23080 27988 23089
rect 28172 23112 28224 23118
rect 28040 23080 28042 23089
rect 28368 23089 28396 25214
rect 28448 25152 28500 25158
rect 28446 25120 28448 25129
rect 28500 25120 28502 25129
rect 28446 25055 28502 25064
rect 28448 24880 28500 24886
rect 28448 24822 28500 24828
rect 28172 23054 28224 23060
rect 28354 23080 28410 23089
rect 27986 23015 28042 23024
rect 28354 23015 28410 23024
rect 28080 22976 28132 22982
rect 28264 22976 28316 22982
rect 28080 22918 28132 22924
rect 28184 22936 28264 22964
rect 28092 22817 28120 22918
rect 28078 22808 28134 22817
rect 27988 22772 28040 22778
rect 28078 22743 28134 22752
rect 27988 22714 28040 22720
rect 28000 22438 28028 22714
rect 28184 22692 28212 22936
rect 28264 22918 28316 22924
rect 28092 22664 28212 22692
rect 28092 22545 28120 22664
rect 28264 22636 28316 22642
rect 28264 22578 28316 22584
rect 28078 22536 28134 22545
rect 28078 22471 28134 22480
rect 27988 22432 28040 22438
rect 27988 22374 28040 22380
rect 27986 22264 28042 22273
rect 27896 22228 27948 22234
rect 28276 22234 28304 22578
rect 27986 22199 28042 22208
rect 28264 22228 28316 22234
rect 27896 22170 27948 22176
rect 27894 21720 27950 21729
rect 27804 21684 27856 21690
rect 27894 21655 27896 21664
rect 27804 21626 27856 21632
rect 27948 21655 27950 21664
rect 27896 21626 27948 21632
rect 28000 21622 28028 22199
rect 28264 22170 28316 22176
rect 28078 22128 28134 22137
rect 28078 22063 28134 22072
rect 27988 21616 28040 21622
rect 27988 21558 28040 21564
rect 27988 20052 28040 20058
rect 27988 19994 28040 20000
rect 27896 18624 27948 18630
rect 27896 18566 27948 18572
rect 27908 18086 27936 18566
rect 27896 18080 27948 18086
rect 27896 18022 27948 18028
rect 28000 17746 28028 19994
rect 27988 17740 28040 17746
rect 27988 17682 28040 17688
rect 27712 17332 27764 17338
rect 27712 17274 27764 17280
rect 27804 17264 27856 17270
rect 27804 17206 27856 17212
rect 27528 16720 27580 16726
rect 27528 16662 27580 16668
rect 27816 16658 27844 17206
rect 27804 16652 27856 16658
rect 27856 16612 28028 16640
rect 27804 16594 27856 16600
rect 27526 16280 27582 16289
rect 27526 16215 27528 16224
rect 27580 16215 27582 16224
rect 27528 16186 27580 16192
rect 28000 15434 28028 16612
rect 27988 15428 28040 15434
rect 27988 15370 28040 15376
rect 27528 14816 27580 14822
rect 27528 14758 27580 14764
rect 27540 13705 27568 14758
rect 27618 14648 27674 14657
rect 27618 14583 27674 14592
rect 27526 13696 27582 13705
rect 27526 13631 27582 13640
rect 27526 13288 27582 13297
rect 27526 13223 27582 13232
rect 27540 12170 27568 13223
rect 27528 12164 27580 12170
rect 27528 12106 27580 12112
rect 27528 11348 27580 11354
rect 27528 11290 27580 11296
rect 27436 10260 27488 10266
rect 27436 10202 27488 10208
rect 27356 10118 27476 10146
rect 27252 10056 27304 10062
rect 27252 9998 27304 10004
rect 26976 8968 27028 8974
rect 26976 8910 27028 8916
rect 27068 8968 27120 8974
rect 27068 8910 27120 8916
rect 27080 8634 27108 8910
rect 27068 8628 27120 8634
rect 27068 8570 27120 8576
rect 26792 8424 26844 8430
rect 26792 8366 26844 8372
rect 26700 7200 26752 7206
rect 26700 7142 26752 7148
rect 26804 6662 26832 8366
rect 27264 8090 27292 9998
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 27252 8084 27304 8090
rect 27252 8026 27304 8032
rect 27252 7200 27304 7206
rect 27252 7142 27304 7148
rect 27264 6730 27292 7142
rect 27356 6730 27384 9522
rect 27252 6724 27304 6730
rect 27252 6666 27304 6672
rect 27344 6724 27396 6730
rect 27344 6666 27396 6672
rect 26240 6656 26292 6662
rect 26240 6598 26292 6604
rect 26792 6656 26844 6662
rect 26792 6598 26844 6604
rect 26252 6118 26280 6598
rect 26804 6322 26832 6598
rect 26792 6316 26844 6322
rect 26792 6258 26844 6264
rect 27264 6254 27292 6666
rect 27448 6610 27476 10118
rect 27540 7546 27568 11290
rect 27632 11150 27660 14583
rect 27986 14512 28042 14521
rect 27986 14447 28042 14456
rect 27894 14240 27950 14249
rect 27894 14175 27950 14184
rect 27908 14074 27936 14175
rect 27896 14068 27948 14074
rect 27896 14010 27948 14016
rect 27804 12980 27856 12986
rect 27804 12922 27856 12928
rect 27816 11286 27844 12922
rect 27896 12300 27948 12306
rect 27896 12242 27948 12248
rect 27908 12209 27936 12242
rect 27894 12200 27950 12209
rect 27894 12135 27950 12144
rect 27894 11792 27950 11801
rect 27894 11727 27896 11736
rect 27948 11727 27950 11736
rect 27896 11698 27948 11704
rect 27896 11620 27948 11626
rect 27896 11562 27948 11568
rect 27804 11280 27856 11286
rect 27804 11222 27856 11228
rect 27620 11144 27672 11150
rect 27620 11086 27672 11092
rect 27632 8634 27660 11086
rect 27908 11082 27936 11562
rect 28000 11218 28028 14447
rect 28092 13705 28120 22063
rect 28170 21992 28226 22001
rect 28170 21927 28172 21936
rect 28224 21927 28226 21936
rect 28172 21898 28224 21904
rect 28170 21448 28226 21457
rect 28170 21383 28226 21392
rect 28184 19802 28212 21383
rect 28264 19916 28316 19922
rect 28368 19904 28396 23015
rect 28460 21486 28488 24822
rect 28552 24818 28580 25706
rect 28644 25294 28672 26998
rect 28828 26450 28856 27367
rect 29644 27338 29696 27344
rect 29460 26784 29512 26790
rect 29460 26726 29512 26732
rect 29550 26752 29606 26761
rect 28816 26444 28868 26450
rect 28816 26386 28868 26392
rect 28724 25764 28776 25770
rect 28724 25706 28776 25712
rect 28736 25430 28764 25706
rect 28724 25424 28776 25430
rect 28724 25366 28776 25372
rect 28828 25362 28856 26386
rect 29092 26240 29144 26246
rect 28998 26208 29054 26217
rect 29092 26182 29144 26188
rect 28998 26143 29054 26152
rect 29012 25809 29040 26143
rect 28998 25800 29054 25809
rect 28998 25735 29054 25744
rect 28908 25696 28960 25702
rect 28906 25664 28908 25673
rect 28960 25664 28962 25673
rect 28906 25599 28962 25608
rect 28906 25392 28962 25401
rect 28816 25356 28868 25362
rect 28906 25327 28962 25336
rect 29000 25356 29052 25362
rect 28816 25298 28868 25304
rect 28632 25288 28684 25294
rect 28632 25230 28684 25236
rect 28540 24812 28592 24818
rect 28540 24754 28592 24760
rect 28552 24070 28580 24754
rect 28540 24064 28592 24070
rect 28540 24006 28592 24012
rect 28448 21480 28500 21486
rect 28448 21422 28500 21428
rect 28552 21321 28580 24006
rect 28644 22545 28672 25230
rect 28724 24268 28776 24274
rect 28724 24210 28776 24216
rect 28736 24177 28764 24210
rect 28722 24168 28778 24177
rect 28722 24103 28778 24112
rect 28816 24064 28868 24070
rect 28816 24006 28868 24012
rect 28828 23866 28856 24006
rect 28816 23860 28868 23866
rect 28816 23802 28868 23808
rect 28920 23798 28948 25327
rect 29000 25298 29052 25304
rect 28908 23792 28960 23798
rect 28908 23734 28960 23740
rect 28724 23588 28776 23594
rect 28724 23530 28776 23536
rect 28630 22536 28686 22545
rect 28630 22471 28686 22480
rect 28632 22432 28684 22438
rect 28632 22374 28684 22380
rect 28538 21312 28594 21321
rect 28538 21247 28594 21256
rect 28644 21162 28672 22374
rect 28460 21134 28672 21162
rect 28460 20806 28488 21134
rect 28632 21004 28684 21010
rect 28552 20964 28632 20992
rect 28448 20800 28500 20806
rect 28448 20742 28500 20748
rect 28316 19876 28396 19904
rect 28264 19858 28316 19864
rect 28184 19774 28304 19802
rect 28170 19408 28226 19417
rect 28170 19343 28226 19352
rect 28078 13696 28134 13705
rect 28078 13631 28134 13640
rect 28080 13524 28132 13530
rect 28080 13466 28132 13472
rect 27988 11212 28040 11218
rect 27988 11154 28040 11160
rect 27896 11076 27948 11082
rect 27896 11018 27948 11024
rect 27710 10976 27766 10985
rect 27710 10911 27766 10920
rect 27724 10606 27752 10911
rect 27712 10600 27764 10606
rect 27712 10542 27764 10548
rect 27802 10432 27858 10441
rect 27802 10367 27858 10376
rect 27816 10198 27844 10367
rect 27712 10192 27764 10198
rect 27712 10134 27764 10140
rect 27804 10192 27856 10198
rect 27804 10134 27856 10140
rect 27724 9722 27752 10134
rect 27804 9988 27856 9994
rect 27908 9976 27936 11018
rect 27986 10840 28042 10849
rect 27986 10775 28042 10784
rect 28000 10538 28028 10775
rect 27988 10532 28040 10538
rect 27988 10474 28040 10480
rect 27986 10296 28042 10305
rect 27986 10231 28042 10240
rect 27856 9948 27936 9976
rect 27804 9930 27856 9936
rect 27712 9716 27764 9722
rect 27712 9658 27764 9664
rect 27710 9616 27766 9625
rect 27710 9551 27766 9560
rect 27724 9450 27752 9551
rect 27816 9518 27844 9930
rect 28000 9722 28028 10231
rect 28092 10130 28120 13466
rect 28184 13258 28212 19343
rect 28276 18193 28304 19774
rect 28552 19281 28580 20964
rect 28632 20946 28684 20952
rect 28736 19990 28764 23530
rect 28906 23488 28962 23497
rect 28906 23423 28962 23432
rect 28814 23352 28870 23361
rect 28920 23322 28948 23423
rect 28814 23287 28870 23296
rect 28908 23316 28960 23322
rect 28724 19984 28776 19990
rect 28630 19952 28686 19961
rect 28724 19926 28776 19932
rect 28630 19887 28686 19896
rect 28644 19854 28672 19887
rect 28632 19848 28684 19854
rect 28632 19790 28684 19796
rect 28538 19272 28594 19281
rect 28538 19207 28594 19216
rect 28262 18184 28318 18193
rect 28318 18142 28396 18170
rect 28262 18119 28318 18128
rect 28264 14340 28316 14346
rect 28264 14282 28316 14288
rect 28276 14249 28304 14282
rect 28262 14240 28318 14249
rect 28262 14175 28318 14184
rect 28262 13832 28318 13841
rect 28262 13767 28318 13776
rect 28276 13394 28304 13767
rect 28368 13530 28396 18142
rect 28630 18048 28686 18057
rect 28630 17983 28686 17992
rect 28540 17876 28592 17882
rect 28540 17818 28592 17824
rect 28552 17134 28580 17818
rect 28644 17338 28672 17983
rect 28722 17776 28778 17785
rect 28722 17711 28778 17720
rect 28632 17332 28684 17338
rect 28632 17274 28684 17280
rect 28540 17128 28592 17134
rect 28540 17070 28592 17076
rect 28538 16552 28594 16561
rect 28736 16522 28764 17711
rect 28538 16487 28594 16496
rect 28724 16516 28776 16522
rect 28552 15570 28580 16487
rect 28724 16458 28776 16464
rect 28828 16402 28856 23287
rect 28908 23258 28960 23264
rect 28908 23180 28960 23186
rect 28908 23122 28960 23128
rect 28920 22545 28948 23122
rect 28906 22536 28962 22545
rect 28906 22471 28962 22480
rect 28906 22400 28962 22409
rect 28906 22335 28962 22344
rect 28920 22030 28948 22335
rect 28908 22024 28960 22030
rect 28908 21966 28960 21972
rect 29012 21672 29040 25298
rect 29104 24070 29132 26182
rect 29274 25936 29330 25945
rect 29274 25871 29330 25880
rect 29368 25900 29420 25906
rect 29182 25800 29238 25809
rect 29182 25735 29238 25744
rect 29196 25226 29224 25735
rect 29184 25220 29236 25226
rect 29184 25162 29236 25168
rect 29184 24744 29236 24750
rect 29184 24686 29236 24692
rect 29092 24064 29144 24070
rect 29092 24006 29144 24012
rect 29092 23860 29144 23866
rect 29092 23802 29144 23808
rect 28920 21644 29040 21672
rect 28920 21434 28948 21644
rect 28920 21406 29040 21434
rect 28906 21312 28962 21321
rect 28906 21247 28962 21256
rect 28920 17882 28948 21247
rect 29012 20058 29040 21406
rect 29000 20052 29052 20058
rect 29000 19994 29052 20000
rect 29000 19236 29052 19242
rect 29000 19178 29052 19184
rect 29012 18970 29040 19178
rect 29000 18964 29052 18970
rect 29000 18906 29052 18912
rect 29104 18358 29132 23802
rect 29196 23662 29224 24686
rect 29184 23656 29236 23662
rect 29184 23598 29236 23604
rect 29184 23180 29236 23186
rect 29184 23122 29236 23128
rect 29196 22710 29224 23122
rect 29288 23118 29316 25871
rect 29368 25842 29420 25848
rect 29276 23112 29328 23118
rect 29276 23054 29328 23060
rect 29184 22704 29236 22710
rect 29184 22646 29236 22652
rect 29196 22438 29224 22646
rect 29184 22432 29236 22438
rect 29184 22374 29236 22380
rect 29274 22400 29330 22409
rect 29274 22335 29330 22344
rect 29184 22092 29236 22098
rect 29184 22034 29236 22040
rect 29196 21418 29224 22034
rect 29184 21412 29236 21418
rect 29184 21354 29236 21360
rect 29288 21010 29316 22335
rect 29276 21004 29328 21010
rect 29276 20946 29328 20952
rect 29184 20936 29236 20942
rect 29182 20904 29184 20913
rect 29236 20904 29238 20913
rect 29182 20839 29238 20848
rect 29276 20868 29328 20874
rect 29276 20810 29328 20816
rect 29184 20596 29236 20602
rect 29184 20538 29236 20544
rect 29196 19417 29224 20538
rect 29288 19553 29316 20810
rect 29380 19802 29408 25842
rect 29472 25786 29500 26726
rect 29550 26687 29606 26696
rect 29564 26518 29592 26687
rect 29552 26512 29604 26518
rect 29552 26454 29604 26460
rect 29656 25838 29684 27338
rect 29734 27024 29790 27033
rect 29734 26959 29790 26968
rect 29748 26489 29776 26959
rect 30196 26852 30248 26858
rect 30196 26794 30248 26800
rect 29846 26684 30154 26704
rect 29846 26682 29852 26684
rect 29908 26682 29932 26684
rect 29988 26682 30012 26684
rect 30068 26682 30092 26684
rect 30148 26682 30154 26684
rect 29908 26630 29910 26682
rect 30090 26630 30092 26682
rect 29846 26628 29852 26630
rect 29908 26628 29932 26630
rect 29988 26628 30012 26630
rect 30068 26628 30092 26630
rect 30148 26628 30154 26630
rect 29846 26608 30154 26628
rect 29734 26480 29790 26489
rect 29734 26415 29790 26424
rect 29748 26382 29776 26415
rect 29736 26376 29788 26382
rect 29736 26318 29788 26324
rect 29920 25968 29972 25974
rect 29734 25936 29790 25945
rect 29920 25910 29972 25916
rect 29734 25871 29790 25880
rect 29644 25832 29696 25838
rect 29472 25758 29592 25786
rect 29644 25774 29696 25780
rect 29460 25696 29512 25702
rect 29460 25638 29512 25644
rect 29472 20534 29500 25638
rect 29564 24256 29592 25758
rect 29748 25378 29776 25871
rect 29932 25770 29960 25910
rect 29920 25764 29972 25770
rect 29920 25706 29972 25712
rect 29846 25596 30154 25616
rect 29846 25594 29852 25596
rect 29908 25594 29932 25596
rect 29988 25594 30012 25596
rect 30068 25594 30092 25596
rect 30148 25594 30154 25596
rect 29908 25542 29910 25594
rect 30090 25542 30092 25594
rect 29846 25540 29852 25542
rect 29908 25540 29932 25542
rect 29988 25540 30012 25542
rect 30068 25540 30092 25542
rect 30148 25540 30154 25542
rect 29846 25520 30154 25540
rect 29656 25350 29776 25378
rect 29656 24750 29684 25350
rect 29736 25220 29788 25226
rect 29736 25162 29788 25168
rect 29748 24993 29776 25162
rect 29734 24984 29790 24993
rect 29734 24919 29790 24928
rect 29920 24812 29972 24818
rect 29748 24772 29920 24800
rect 29644 24744 29696 24750
rect 29644 24686 29696 24692
rect 29644 24268 29696 24274
rect 29564 24228 29644 24256
rect 29644 24210 29696 24216
rect 29656 23769 29684 24210
rect 29642 23760 29698 23769
rect 29552 23724 29604 23730
rect 29642 23695 29698 23704
rect 29552 23666 29604 23672
rect 29564 23322 29592 23666
rect 29552 23316 29604 23322
rect 29552 23258 29604 23264
rect 29644 23248 29696 23254
rect 29644 23190 29696 23196
rect 29552 23112 29604 23118
rect 29552 23054 29604 23060
rect 29564 22098 29592 23054
rect 29552 22092 29604 22098
rect 29552 22034 29604 22040
rect 29552 21888 29604 21894
rect 29552 21830 29604 21836
rect 29564 21690 29592 21830
rect 29552 21684 29604 21690
rect 29552 21626 29604 21632
rect 29552 21480 29604 21486
rect 29552 21422 29604 21428
rect 29564 21078 29592 21422
rect 29552 21072 29604 21078
rect 29552 21014 29604 21020
rect 29656 20874 29684 23190
rect 29748 22234 29776 24772
rect 29920 24754 29972 24760
rect 29846 24508 30154 24528
rect 29846 24506 29852 24508
rect 29908 24506 29932 24508
rect 29988 24506 30012 24508
rect 30068 24506 30092 24508
rect 30148 24506 30154 24508
rect 29908 24454 29910 24506
rect 30090 24454 30092 24506
rect 29846 24452 29852 24454
rect 29908 24452 29932 24454
rect 29988 24452 30012 24454
rect 30068 24452 30092 24454
rect 30148 24452 30154 24454
rect 29846 24432 30154 24452
rect 30104 24064 30156 24070
rect 30104 24006 30156 24012
rect 30116 23769 30144 24006
rect 30102 23760 30158 23769
rect 30102 23695 30158 23704
rect 30012 23656 30064 23662
rect 30010 23624 30012 23633
rect 30064 23624 30066 23633
rect 30208 23610 30236 26794
rect 30300 25294 30328 27610
rect 30380 27464 30432 27470
rect 30380 27406 30432 27412
rect 30392 25922 30420 27406
rect 30484 26586 30512 27911
rect 31942 27840 31998 27849
rect 31942 27775 31998 27784
rect 30748 27600 30800 27606
rect 30748 27542 30800 27548
rect 30564 26784 30616 26790
rect 30564 26726 30616 26732
rect 30472 26580 30524 26586
rect 30472 26522 30524 26528
rect 30470 26072 30526 26081
rect 30470 26007 30472 26016
rect 30524 26007 30526 26016
rect 30472 25978 30524 25984
rect 30392 25894 30512 25922
rect 30380 25764 30432 25770
rect 30380 25706 30432 25712
rect 30392 25673 30420 25706
rect 30378 25664 30434 25673
rect 30378 25599 30434 25608
rect 30392 25401 30420 25599
rect 30378 25392 30434 25401
rect 30378 25327 30434 25336
rect 30288 25288 30340 25294
rect 30288 25230 30340 25236
rect 30380 24200 30432 24206
rect 30378 24168 30380 24177
rect 30432 24168 30434 24177
rect 30378 24103 30434 24112
rect 30484 23882 30512 25894
rect 30576 25294 30604 26726
rect 30760 26450 30788 27542
rect 31576 27328 31628 27334
rect 31576 27270 31628 27276
rect 30840 26784 30892 26790
rect 30838 26752 30840 26761
rect 31484 26784 31536 26790
rect 30892 26752 30894 26761
rect 31484 26726 31536 26732
rect 30838 26687 30894 26696
rect 31206 26616 31262 26625
rect 31206 26551 31208 26560
rect 31260 26551 31262 26560
rect 31208 26522 31260 26528
rect 30748 26444 30800 26450
rect 30748 26386 30800 26392
rect 31208 26376 31260 26382
rect 31496 26353 31524 26726
rect 31208 26318 31260 26324
rect 31482 26344 31538 26353
rect 31022 26208 31078 26217
rect 31022 26143 31078 26152
rect 30932 25832 30984 25838
rect 30932 25774 30984 25780
rect 30840 25696 30892 25702
rect 30840 25638 30892 25644
rect 30564 25288 30616 25294
rect 30562 25256 30564 25265
rect 30616 25256 30618 25265
rect 30562 25191 30618 25200
rect 30656 24812 30708 24818
rect 30656 24754 30708 24760
rect 30564 24744 30616 24750
rect 30564 24686 30616 24692
rect 30576 24342 30604 24686
rect 30564 24336 30616 24342
rect 30564 24278 30616 24284
rect 30668 24256 30696 24754
rect 30668 24228 30788 24256
rect 30300 23854 30512 23882
rect 30300 23798 30328 23854
rect 30288 23792 30340 23798
rect 30288 23734 30340 23740
rect 30208 23582 30328 23610
rect 30010 23559 30066 23568
rect 30196 23520 30248 23526
rect 30196 23462 30248 23468
rect 29846 23420 30154 23440
rect 29846 23418 29852 23420
rect 29908 23418 29932 23420
rect 29988 23418 30012 23420
rect 30068 23418 30092 23420
rect 30148 23418 30154 23420
rect 29908 23366 29910 23418
rect 30090 23366 30092 23418
rect 29846 23364 29852 23366
rect 29908 23364 29932 23366
rect 29988 23364 30012 23366
rect 30068 23364 30092 23366
rect 30148 23364 30154 23366
rect 29846 23344 30154 23364
rect 30208 23322 30236 23462
rect 30196 23316 30248 23322
rect 30196 23258 30248 23264
rect 30300 23202 30328 23582
rect 30208 23174 30328 23202
rect 30104 23044 30156 23050
rect 30104 22986 30156 22992
rect 30116 22681 30144 22986
rect 30102 22672 30158 22681
rect 30102 22607 30158 22616
rect 29846 22332 30154 22352
rect 29846 22330 29852 22332
rect 29908 22330 29932 22332
rect 29988 22330 30012 22332
rect 30068 22330 30092 22332
rect 30148 22330 30154 22332
rect 29908 22278 29910 22330
rect 30090 22278 30092 22330
rect 29846 22276 29852 22278
rect 29908 22276 29932 22278
rect 29988 22276 30012 22278
rect 30068 22276 30092 22278
rect 30148 22276 30154 22278
rect 29846 22256 30154 22276
rect 29736 22228 29788 22234
rect 29736 22170 29788 22176
rect 29644 20868 29696 20874
rect 29644 20810 29696 20816
rect 29550 20768 29606 20777
rect 29550 20703 29606 20712
rect 29460 20528 29512 20534
rect 29460 20470 29512 20476
rect 29380 19774 29500 19802
rect 29368 19712 29420 19718
rect 29368 19654 29420 19660
rect 29274 19544 29330 19553
rect 29274 19479 29330 19488
rect 29182 19408 29238 19417
rect 29182 19343 29238 19352
rect 29276 19372 29328 19378
rect 29276 19314 29328 19320
rect 29288 19258 29316 19314
rect 29196 19230 29316 19258
rect 29092 18352 29144 18358
rect 29092 18294 29144 18300
rect 28908 17876 28960 17882
rect 28908 17818 28960 17824
rect 28908 17332 28960 17338
rect 28908 17274 28960 17280
rect 28920 17066 28948 17274
rect 28908 17060 28960 17066
rect 28908 17002 28960 17008
rect 29092 16788 29144 16794
rect 29092 16730 29144 16736
rect 29000 16720 29052 16726
rect 28998 16688 29000 16697
rect 29052 16688 29054 16697
rect 29104 16658 29132 16730
rect 29196 16726 29224 19230
rect 29276 19168 29328 19174
rect 29276 19110 29328 19116
rect 29288 18057 29316 19110
rect 29380 19009 29408 19654
rect 29472 19378 29500 19774
rect 29460 19372 29512 19378
rect 29460 19314 29512 19320
rect 29460 19168 29512 19174
rect 29460 19110 29512 19116
rect 29366 19000 29422 19009
rect 29366 18935 29422 18944
rect 29472 18766 29500 19110
rect 29460 18760 29512 18766
rect 29460 18702 29512 18708
rect 29472 18222 29500 18702
rect 29368 18216 29420 18222
rect 29368 18158 29420 18164
rect 29460 18216 29512 18222
rect 29460 18158 29512 18164
rect 29274 18048 29330 18057
rect 29274 17983 29330 17992
rect 29276 16992 29328 16998
rect 29276 16934 29328 16940
rect 29288 16794 29316 16934
rect 29276 16788 29328 16794
rect 29276 16730 29328 16736
rect 29184 16720 29236 16726
rect 29184 16662 29236 16668
rect 28998 16623 29054 16632
rect 29092 16652 29144 16658
rect 29092 16594 29144 16600
rect 29276 16516 29328 16522
rect 29276 16458 29328 16464
rect 29182 16416 29238 16425
rect 28828 16374 28994 16402
rect 28966 16266 28994 16374
rect 29182 16351 29238 16360
rect 28966 16238 29132 16266
rect 28724 15904 28776 15910
rect 28724 15846 28776 15852
rect 28540 15564 28592 15570
rect 28540 15506 28592 15512
rect 28448 15360 28500 15366
rect 28736 15337 28764 15846
rect 28814 15736 28870 15745
rect 28814 15671 28870 15680
rect 28448 15302 28500 15308
rect 28722 15328 28778 15337
rect 28356 13524 28408 13530
rect 28356 13466 28408 13472
rect 28264 13388 28316 13394
rect 28264 13330 28316 13336
rect 28172 13252 28224 13258
rect 28172 13194 28224 13200
rect 28354 13152 28410 13161
rect 28354 13087 28410 13096
rect 28262 12608 28318 12617
rect 28262 12543 28318 12552
rect 28276 12170 28304 12543
rect 28264 12164 28316 12170
rect 28264 12106 28316 12112
rect 28264 11756 28316 11762
rect 28264 11698 28316 11704
rect 28172 11552 28224 11558
rect 28172 11494 28224 11500
rect 28080 10124 28132 10130
rect 28080 10066 28132 10072
rect 27896 9716 27948 9722
rect 27896 9658 27948 9664
rect 27988 9716 28040 9722
rect 27988 9658 28040 9664
rect 27804 9512 27856 9518
rect 27804 9454 27856 9460
rect 27712 9444 27764 9450
rect 27712 9386 27764 9392
rect 27710 9208 27766 9217
rect 27710 9143 27712 9152
rect 27764 9143 27766 9152
rect 27712 9114 27764 9120
rect 27712 9036 27764 9042
rect 27712 8978 27764 8984
rect 27724 8634 27752 8978
rect 27620 8628 27672 8634
rect 27620 8570 27672 8576
rect 27712 8628 27764 8634
rect 27712 8570 27764 8576
rect 27816 8022 27844 9454
rect 27804 8016 27856 8022
rect 27804 7958 27856 7964
rect 27528 7540 27580 7546
rect 27528 7482 27580 7488
rect 27908 7313 27936 9658
rect 28000 8634 28028 9658
rect 28092 9450 28120 10066
rect 28184 10062 28212 11494
rect 28172 10056 28224 10062
rect 28172 9998 28224 10004
rect 28080 9444 28132 9450
rect 28080 9386 28132 9392
rect 28092 9042 28120 9386
rect 28080 9036 28132 9042
rect 28080 8978 28132 8984
rect 27988 8628 28040 8634
rect 27988 8570 28040 8576
rect 27894 7304 27950 7313
rect 27894 7239 27950 7248
rect 27356 6582 27476 6610
rect 27252 6248 27304 6254
rect 27252 6190 27304 6196
rect 27356 6118 27384 6582
rect 28000 6390 28028 8570
rect 28092 8090 28120 8978
rect 28184 8634 28212 9998
rect 28276 9042 28304 11698
rect 28368 11626 28396 13087
rect 28356 11620 28408 11626
rect 28356 11562 28408 11568
rect 28356 10532 28408 10538
rect 28356 10474 28408 10480
rect 28368 9586 28396 10474
rect 28460 10266 28488 15302
rect 28722 15263 28778 15272
rect 28540 15088 28592 15094
rect 28540 15030 28592 15036
rect 28552 14929 28580 15030
rect 28538 14920 28594 14929
rect 28538 14855 28594 14864
rect 28538 14648 28594 14657
rect 28538 14583 28594 14592
rect 28552 14074 28580 14583
rect 28632 14340 28684 14346
rect 28632 14282 28684 14288
rect 28540 14068 28592 14074
rect 28540 14010 28592 14016
rect 28448 10260 28500 10266
rect 28448 10202 28500 10208
rect 28552 10130 28580 14010
rect 28644 10282 28672 14282
rect 28724 13252 28776 13258
rect 28724 13194 28776 13200
rect 28736 13025 28764 13194
rect 28722 13016 28778 13025
rect 28722 12951 28778 12960
rect 28724 11892 28776 11898
rect 28724 11834 28776 11840
rect 28736 11801 28764 11834
rect 28722 11792 28778 11801
rect 28722 11727 28778 11736
rect 28828 11529 28856 15671
rect 28998 15192 29054 15201
rect 28998 15127 29054 15136
rect 29012 15094 29040 15127
rect 29000 15088 29052 15094
rect 29000 15030 29052 15036
rect 28906 13696 28962 13705
rect 28906 13631 28962 13640
rect 28920 12782 28948 13631
rect 29000 13320 29052 13326
rect 29000 13262 29052 13268
rect 28908 12776 28960 12782
rect 28908 12718 28960 12724
rect 28906 12064 28962 12073
rect 28906 11999 28962 12008
rect 28920 11762 28948 11999
rect 28908 11756 28960 11762
rect 28908 11698 28960 11704
rect 28908 11620 28960 11626
rect 28908 11562 28960 11568
rect 28814 11520 28870 11529
rect 28814 11455 28870 11464
rect 28724 11144 28776 11150
rect 28724 11086 28776 11092
rect 28736 10441 28764 11086
rect 28722 10432 28778 10441
rect 28722 10367 28778 10376
rect 28644 10254 28764 10282
rect 28540 10124 28592 10130
rect 28540 10066 28592 10072
rect 28538 10024 28594 10033
rect 28448 9988 28500 9994
rect 28538 9959 28594 9968
rect 28448 9930 28500 9936
rect 28460 9722 28488 9930
rect 28448 9716 28500 9722
rect 28552 9704 28580 9959
rect 28632 9716 28684 9722
rect 28552 9676 28632 9704
rect 28448 9658 28500 9664
rect 28632 9658 28684 9664
rect 28460 9625 28488 9658
rect 28446 9616 28502 9625
rect 28356 9580 28408 9586
rect 28736 9568 28764 10254
rect 28446 9551 28502 9560
rect 28356 9522 28408 9528
rect 28644 9540 28764 9568
rect 28264 9036 28316 9042
rect 28264 8978 28316 8984
rect 28172 8628 28224 8634
rect 28172 8570 28224 8576
rect 28080 8084 28132 8090
rect 28080 8026 28132 8032
rect 28368 6798 28396 9522
rect 28448 9376 28500 9382
rect 28448 9318 28500 9324
rect 28460 9110 28488 9318
rect 28644 9178 28672 9540
rect 28722 9480 28778 9489
rect 28722 9415 28778 9424
rect 28632 9172 28684 9178
rect 28632 9114 28684 9120
rect 28448 9104 28500 9110
rect 28448 9046 28500 9052
rect 28538 9072 28594 9081
rect 28632 9036 28684 9042
rect 28594 9016 28632 9024
rect 28538 9007 28632 9016
rect 28552 8996 28632 9007
rect 28552 7546 28580 8996
rect 28632 8978 28684 8984
rect 28736 8974 28764 9415
rect 28724 8968 28776 8974
rect 28724 8910 28776 8916
rect 28722 8664 28778 8673
rect 28722 8599 28724 8608
rect 28644 8566 28672 8597
rect 28776 8599 28778 8608
rect 28724 8570 28776 8576
rect 28632 8560 28684 8566
rect 28630 8528 28632 8537
rect 28684 8528 28686 8537
rect 28828 8498 28856 11455
rect 28920 10305 28948 11562
rect 28906 10296 28962 10305
rect 28906 10231 28962 10240
rect 28908 10124 28960 10130
rect 28908 10066 28960 10072
rect 28630 8463 28686 8472
rect 28816 8492 28868 8498
rect 28540 7540 28592 7546
rect 28540 7482 28592 7488
rect 28356 6792 28408 6798
rect 28356 6734 28408 6740
rect 28644 6730 28672 8463
rect 28816 8434 28868 8440
rect 28632 6724 28684 6730
rect 28632 6666 28684 6672
rect 28446 6488 28502 6497
rect 28446 6423 28502 6432
rect 27988 6384 28040 6390
rect 27988 6326 28040 6332
rect 26240 6112 26292 6118
rect 26240 6054 26292 6060
rect 27344 6112 27396 6118
rect 27344 6054 27396 6060
rect 27356 5234 27384 6054
rect 28460 5914 28488 6423
rect 28828 5914 28856 8434
rect 28920 7546 28948 10066
rect 28908 7540 28960 7546
rect 28908 7482 28960 7488
rect 29012 7478 29040 13262
rect 29104 12986 29132 16238
rect 29196 14006 29224 16351
rect 29184 14000 29236 14006
rect 29184 13942 29236 13948
rect 29288 13569 29316 16458
rect 29274 13560 29330 13569
rect 29274 13495 29330 13504
rect 29276 13456 29328 13462
rect 29182 13424 29238 13433
rect 29276 13398 29328 13404
rect 29182 13359 29238 13368
rect 29092 12980 29144 12986
rect 29092 12922 29144 12928
rect 29090 12744 29146 12753
rect 29090 12679 29092 12688
rect 29144 12679 29146 12688
rect 29092 12650 29144 12656
rect 29092 12164 29144 12170
rect 29092 12106 29144 12112
rect 29104 7721 29132 12106
rect 29196 11762 29224 13359
rect 29288 12288 29316 13398
rect 29380 12442 29408 18158
rect 29472 17678 29500 18158
rect 29460 17672 29512 17678
rect 29460 17614 29512 17620
rect 29472 17320 29500 17614
rect 29564 17610 29592 20703
rect 29552 17604 29604 17610
rect 29552 17546 29604 17552
rect 29552 17332 29604 17338
rect 29472 17292 29552 17320
rect 29552 17274 29604 17280
rect 29460 16992 29512 16998
rect 29460 16934 29512 16940
rect 29472 16182 29500 16934
rect 29564 16590 29592 17274
rect 29552 16584 29604 16590
rect 29552 16526 29604 16532
rect 29460 16176 29512 16182
rect 29460 16118 29512 16124
rect 29656 15960 29684 20810
rect 29748 19854 29776 22170
rect 30208 21690 30236 23174
rect 30484 22438 30512 23854
rect 30760 23798 30788 24228
rect 30852 23905 30880 25638
rect 30838 23896 30894 23905
rect 30838 23831 30894 23840
rect 30748 23792 30800 23798
rect 30800 23752 30880 23780
rect 30748 23734 30800 23740
rect 30656 23656 30708 23662
rect 30656 23598 30708 23604
rect 30472 22432 30524 22438
rect 30472 22374 30524 22380
rect 30484 22250 30512 22374
rect 30300 22222 30512 22250
rect 30196 21684 30248 21690
rect 30196 21626 30248 21632
rect 30300 21298 30328 22222
rect 30380 22092 30432 22098
rect 30380 22034 30432 22040
rect 30392 21622 30420 22034
rect 30472 21684 30524 21690
rect 30472 21626 30524 21632
rect 30380 21616 30432 21622
rect 30380 21558 30432 21564
rect 30300 21270 30420 21298
rect 29846 21244 30154 21264
rect 29846 21242 29852 21244
rect 29908 21242 29932 21244
rect 29988 21242 30012 21244
rect 30068 21242 30092 21244
rect 30148 21242 30154 21244
rect 29908 21190 29910 21242
rect 30090 21190 30092 21242
rect 29846 21188 29852 21190
rect 29908 21188 29932 21190
rect 29988 21188 30012 21190
rect 30068 21188 30092 21190
rect 30148 21188 30154 21190
rect 29846 21168 30154 21188
rect 30286 21176 30342 21185
rect 30286 21111 30342 21120
rect 30012 21004 30064 21010
rect 30300 20992 30328 21111
rect 30064 20964 30328 20992
rect 30012 20946 30064 20952
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 29918 20904 29974 20913
rect 29840 20369 29868 20878
rect 30392 20890 30420 21270
rect 30484 21010 30512 21626
rect 30562 21312 30618 21321
rect 30562 21247 30618 21256
rect 30576 21146 30604 21247
rect 30564 21140 30616 21146
rect 30564 21082 30616 21088
rect 30472 21004 30524 21010
rect 30472 20946 30524 20952
rect 29918 20839 29974 20848
rect 30300 20862 30420 20890
rect 29932 20806 29960 20839
rect 29920 20800 29972 20806
rect 29920 20742 29972 20748
rect 29826 20360 29882 20369
rect 29826 20295 29882 20304
rect 29846 20156 30154 20176
rect 29846 20154 29852 20156
rect 29908 20154 29932 20156
rect 29988 20154 30012 20156
rect 30068 20154 30092 20156
rect 30148 20154 30154 20156
rect 29908 20102 29910 20154
rect 30090 20102 30092 20154
rect 29846 20100 29852 20102
rect 29908 20100 29932 20102
rect 29988 20100 30012 20102
rect 30068 20100 30092 20102
rect 30148 20100 30154 20102
rect 29846 20080 30154 20100
rect 29736 19848 29788 19854
rect 29736 19790 29788 19796
rect 29748 19446 29776 19790
rect 30196 19712 30248 19718
rect 30196 19654 30248 19660
rect 30208 19514 30236 19654
rect 30196 19508 30248 19514
rect 30196 19450 30248 19456
rect 29736 19440 29788 19446
rect 29736 19382 29788 19388
rect 29846 19068 30154 19088
rect 29846 19066 29852 19068
rect 29908 19066 29932 19068
rect 29988 19066 30012 19068
rect 30068 19066 30092 19068
rect 30148 19066 30154 19068
rect 29908 19014 29910 19066
rect 30090 19014 30092 19066
rect 29846 19012 29852 19014
rect 29908 19012 29932 19014
rect 29988 19012 30012 19014
rect 30068 19012 30092 19014
rect 30148 19012 30154 19014
rect 29846 18992 30154 19012
rect 30208 18986 30236 19450
rect 30300 19174 30328 20862
rect 30380 20800 30432 20806
rect 30378 20768 30380 20777
rect 30432 20768 30434 20777
rect 30378 20703 30434 20712
rect 30484 20233 30512 20946
rect 30470 20224 30526 20233
rect 30470 20159 30526 20168
rect 30564 19916 30616 19922
rect 30564 19858 30616 19864
rect 30288 19168 30340 19174
rect 30288 19110 30340 19116
rect 30380 19168 30432 19174
rect 30380 19110 30432 19116
rect 30392 18986 30420 19110
rect 30208 18958 30420 18986
rect 29826 18864 29882 18873
rect 30378 18864 30434 18873
rect 29826 18799 29882 18808
rect 30300 18808 30378 18816
rect 30300 18799 30434 18808
rect 29736 18692 29788 18698
rect 29736 18634 29788 18640
rect 29472 15932 29684 15960
rect 29368 12436 29420 12442
rect 29368 12378 29420 12384
rect 29368 12300 29420 12306
rect 29288 12260 29368 12288
rect 29368 12242 29420 12248
rect 29184 11756 29236 11762
rect 29184 11698 29236 11704
rect 29090 7712 29146 7721
rect 29090 7647 29146 7656
rect 29196 7546 29224 11698
rect 29276 11552 29328 11558
rect 29274 11520 29276 11529
rect 29328 11520 29330 11529
rect 29274 11455 29330 11464
rect 29274 11384 29330 11393
rect 29274 11319 29330 11328
rect 29288 11150 29316 11319
rect 29276 11144 29328 11150
rect 29276 11086 29328 11092
rect 29288 9674 29316 11086
rect 29380 10169 29408 12242
rect 29366 10160 29422 10169
rect 29366 10095 29422 10104
rect 29288 9646 29408 9674
rect 29276 9580 29328 9586
rect 29276 9522 29328 9528
rect 29184 7540 29236 7546
rect 29184 7482 29236 7488
rect 29000 7472 29052 7478
rect 29000 7414 29052 7420
rect 29288 6798 29316 9522
rect 29380 9178 29408 9646
rect 29472 9586 29500 15932
rect 29550 15872 29606 15881
rect 29550 15807 29606 15816
rect 29564 15638 29592 15807
rect 29552 15632 29604 15638
rect 29552 15574 29604 15580
rect 29552 15428 29604 15434
rect 29552 15370 29604 15376
rect 29564 15094 29592 15370
rect 29644 15360 29696 15366
rect 29644 15302 29696 15308
rect 29552 15088 29604 15094
rect 29552 15030 29604 15036
rect 29552 14884 29604 14890
rect 29552 14826 29604 14832
rect 29564 14793 29592 14826
rect 29550 14784 29606 14793
rect 29550 14719 29606 14728
rect 29656 14618 29684 15302
rect 29644 14612 29696 14618
rect 29644 14554 29696 14560
rect 29552 14408 29604 14414
rect 29552 14350 29604 14356
rect 29642 14376 29698 14385
rect 29564 13462 29592 14350
rect 29642 14311 29698 14320
rect 29656 14074 29684 14311
rect 29644 14068 29696 14074
rect 29644 14010 29696 14016
rect 29644 13864 29696 13870
rect 29644 13806 29696 13812
rect 29552 13456 29604 13462
rect 29552 13398 29604 13404
rect 29552 12776 29604 12782
rect 29552 12718 29604 12724
rect 29564 12617 29592 12718
rect 29550 12608 29606 12617
rect 29550 12543 29606 12552
rect 29552 12232 29604 12238
rect 29552 12174 29604 12180
rect 29564 10470 29592 12174
rect 29552 10464 29604 10470
rect 29552 10406 29604 10412
rect 29564 10130 29592 10406
rect 29552 10124 29604 10130
rect 29552 10066 29604 10072
rect 29550 9888 29606 9897
rect 29550 9823 29606 9832
rect 29460 9580 29512 9586
rect 29460 9522 29512 9528
rect 29460 9376 29512 9382
rect 29460 9318 29512 9324
rect 29368 9172 29420 9178
rect 29368 9114 29420 9120
rect 29368 8832 29420 8838
rect 29368 8774 29420 8780
rect 29380 8566 29408 8774
rect 29368 8560 29420 8566
rect 29368 8502 29420 8508
rect 29368 8424 29420 8430
rect 29368 8366 29420 8372
rect 29380 6866 29408 8366
rect 29368 6860 29420 6866
rect 29368 6802 29420 6808
rect 28908 6792 28960 6798
rect 28908 6734 28960 6740
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 28920 6390 28948 6734
rect 29380 6458 29408 6802
rect 29472 6497 29500 9318
rect 29458 6488 29514 6497
rect 29368 6452 29420 6458
rect 29458 6423 29514 6432
rect 29368 6394 29420 6400
rect 28908 6384 28960 6390
rect 28908 6326 28960 6332
rect 28448 5908 28500 5914
rect 28448 5850 28500 5856
rect 28816 5908 28868 5914
rect 28816 5850 28868 5856
rect 27344 5228 27396 5234
rect 27344 5170 27396 5176
rect 25976 2746 26096 2774
rect 25872 2508 25924 2514
rect 25872 2450 25924 2456
rect 25504 2032 25556 2038
rect 25504 1974 25556 1980
rect 26068 1970 26096 2746
rect 26056 1964 26108 1970
rect 26056 1906 26108 1912
rect 28460 1601 28488 5850
rect 29458 5400 29514 5409
rect 29458 5335 29460 5344
rect 29512 5335 29514 5344
rect 29460 5306 29512 5312
rect 29564 4826 29592 9823
rect 29656 8537 29684 13806
rect 29642 8528 29698 8537
rect 29642 8463 29698 8472
rect 29748 8430 29776 18634
rect 29840 18630 29868 18799
rect 30300 18788 30420 18799
rect 29828 18624 29880 18630
rect 29828 18566 29880 18572
rect 29846 17980 30154 18000
rect 29846 17978 29852 17980
rect 29908 17978 29932 17980
rect 29988 17978 30012 17980
rect 30068 17978 30092 17980
rect 30148 17978 30154 17980
rect 29908 17926 29910 17978
rect 30090 17926 30092 17978
rect 29846 17924 29852 17926
rect 29908 17924 29932 17926
rect 29988 17924 30012 17926
rect 30068 17924 30092 17926
rect 30148 17924 30154 17926
rect 29846 17904 30154 17924
rect 29846 16892 30154 16912
rect 29846 16890 29852 16892
rect 29908 16890 29932 16892
rect 29988 16890 30012 16892
rect 30068 16890 30092 16892
rect 30148 16890 30154 16892
rect 29908 16838 29910 16890
rect 30090 16838 30092 16890
rect 29846 16836 29852 16838
rect 29908 16836 29932 16838
rect 29988 16836 30012 16838
rect 30068 16836 30092 16838
rect 30148 16836 30154 16838
rect 29846 16816 30154 16836
rect 29920 16720 29972 16726
rect 29920 16662 29972 16668
rect 29932 16182 29960 16662
rect 29920 16176 29972 16182
rect 29920 16118 29972 16124
rect 30196 16108 30248 16114
rect 30196 16050 30248 16056
rect 29846 15804 30154 15824
rect 29846 15802 29852 15804
rect 29908 15802 29932 15804
rect 29988 15802 30012 15804
rect 30068 15802 30092 15804
rect 30148 15802 30154 15804
rect 29908 15750 29910 15802
rect 30090 15750 30092 15802
rect 29846 15748 29852 15750
rect 29908 15748 29932 15750
rect 29988 15748 30012 15750
rect 30068 15748 30092 15750
rect 30148 15748 30154 15750
rect 29846 15728 30154 15748
rect 30208 15366 30236 16050
rect 30300 15910 30328 18788
rect 30380 18624 30432 18630
rect 30380 18566 30432 18572
rect 30392 18426 30420 18566
rect 30380 18420 30432 18426
rect 30380 18362 30432 18368
rect 30380 18216 30432 18222
rect 30380 18158 30432 18164
rect 30288 15904 30340 15910
rect 30288 15846 30340 15852
rect 30288 15428 30340 15434
rect 30288 15370 30340 15376
rect 30196 15360 30248 15366
rect 30196 15302 30248 15308
rect 29846 14716 30154 14736
rect 29846 14714 29852 14716
rect 29908 14714 29932 14716
rect 29988 14714 30012 14716
rect 30068 14714 30092 14716
rect 30148 14714 30154 14716
rect 29908 14662 29910 14714
rect 30090 14662 30092 14714
rect 29846 14660 29852 14662
rect 29908 14660 29932 14662
rect 29988 14660 30012 14662
rect 30068 14660 30092 14662
rect 30148 14660 30154 14662
rect 29846 14640 30154 14660
rect 29828 14544 29880 14550
rect 29828 14486 29880 14492
rect 29840 13870 29868 14486
rect 29920 14408 29972 14414
rect 29920 14350 29972 14356
rect 29932 13870 29960 14350
rect 29828 13864 29880 13870
rect 29828 13806 29880 13812
rect 29920 13864 29972 13870
rect 29920 13806 29972 13812
rect 29846 13628 30154 13648
rect 29846 13626 29852 13628
rect 29908 13626 29932 13628
rect 29988 13626 30012 13628
rect 30068 13626 30092 13628
rect 30148 13626 30154 13628
rect 29908 13574 29910 13626
rect 30090 13574 30092 13626
rect 29846 13572 29852 13574
rect 29908 13572 29932 13574
rect 29988 13572 30012 13574
rect 30068 13572 30092 13574
rect 30148 13572 30154 13574
rect 29846 13552 30154 13572
rect 30196 13524 30248 13530
rect 30196 13466 30248 13472
rect 29826 13424 29882 13433
rect 29826 13359 29882 13368
rect 29840 13326 29868 13359
rect 29828 13320 29880 13326
rect 29828 13262 29880 13268
rect 29840 13161 29868 13262
rect 29826 13152 29882 13161
rect 29826 13087 29882 13096
rect 29846 12540 30154 12560
rect 29846 12538 29852 12540
rect 29908 12538 29932 12540
rect 29988 12538 30012 12540
rect 30068 12538 30092 12540
rect 30148 12538 30154 12540
rect 29908 12486 29910 12538
rect 30090 12486 30092 12538
rect 29846 12484 29852 12486
rect 29908 12484 29932 12486
rect 29988 12484 30012 12486
rect 30068 12484 30092 12486
rect 30148 12484 30154 12486
rect 29846 12464 30154 12484
rect 30208 12102 30236 13466
rect 30300 12782 30328 15370
rect 30392 14958 30420 18158
rect 30470 17504 30526 17513
rect 30470 17439 30526 17448
rect 30484 16697 30512 17439
rect 30470 16688 30526 16697
rect 30470 16623 30526 16632
rect 30470 16416 30526 16425
rect 30470 16351 30526 16360
rect 30484 15609 30512 16351
rect 30470 15600 30526 15609
rect 30470 15535 30526 15544
rect 30380 14952 30432 14958
rect 30380 14894 30432 14900
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 30288 12776 30340 12782
rect 30288 12718 30340 12724
rect 30392 12617 30420 14214
rect 30378 12608 30434 12617
rect 30378 12543 30434 12552
rect 30196 12096 30248 12102
rect 30196 12038 30248 12044
rect 30286 11792 30342 11801
rect 30286 11727 30342 11736
rect 30196 11688 30248 11694
rect 30196 11630 30248 11636
rect 29846 11452 30154 11472
rect 29846 11450 29852 11452
rect 29908 11450 29932 11452
rect 29988 11450 30012 11452
rect 30068 11450 30092 11452
rect 30148 11450 30154 11452
rect 29908 11398 29910 11450
rect 30090 11398 30092 11450
rect 29846 11396 29852 11398
rect 29908 11396 29932 11398
rect 29988 11396 30012 11398
rect 30068 11396 30092 11398
rect 30148 11396 30154 11398
rect 29846 11376 30154 11396
rect 29846 10364 30154 10384
rect 29846 10362 29852 10364
rect 29908 10362 29932 10364
rect 29988 10362 30012 10364
rect 30068 10362 30092 10364
rect 30148 10362 30154 10364
rect 29908 10310 29910 10362
rect 30090 10310 30092 10362
rect 29846 10308 29852 10310
rect 29908 10308 29932 10310
rect 29988 10308 30012 10310
rect 30068 10308 30092 10310
rect 30148 10308 30154 10310
rect 29846 10288 30154 10308
rect 30208 10169 30236 11630
rect 30300 11218 30328 11727
rect 30288 11212 30340 11218
rect 30288 11154 30340 11160
rect 30380 11008 30432 11014
rect 30380 10950 30432 10956
rect 30288 10668 30340 10674
rect 30288 10610 30340 10616
rect 29918 10160 29974 10169
rect 30194 10160 30250 10169
rect 29918 10095 29974 10104
rect 30012 10124 30064 10130
rect 29828 9580 29880 9586
rect 29828 9522 29880 9528
rect 29840 9450 29868 9522
rect 29828 9444 29880 9450
rect 29828 9386 29880 9392
rect 29932 9364 29960 10095
rect 30012 10066 30064 10072
rect 30104 10124 30156 10130
rect 30194 10095 30250 10104
rect 30104 10066 30156 10072
rect 30024 9897 30052 10066
rect 30116 9994 30144 10066
rect 30104 9988 30156 9994
rect 30104 9930 30156 9936
rect 30010 9888 30066 9897
rect 30010 9823 30066 9832
rect 30300 9704 30328 10610
rect 30392 10538 30420 10950
rect 30380 10532 30432 10538
rect 30380 10474 30432 10480
rect 30300 9676 30420 9704
rect 30102 9616 30158 9625
rect 30102 9551 30104 9560
rect 30156 9551 30158 9560
rect 30104 9522 30156 9528
rect 30116 9432 30144 9522
rect 30116 9404 30328 9432
rect 29932 9336 30236 9364
rect 29846 9276 30154 9296
rect 29846 9274 29852 9276
rect 29908 9274 29932 9276
rect 29988 9274 30012 9276
rect 30068 9274 30092 9276
rect 30148 9274 30154 9276
rect 29908 9222 29910 9274
rect 30090 9222 30092 9274
rect 29846 9220 29852 9222
rect 29908 9220 29932 9222
rect 29988 9220 30012 9222
rect 30068 9220 30092 9222
rect 30148 9220 30154 9222
rect 29846 9200 30154 9220
rect 30208 9160 30236 9336
rect 29840 9132 30236 9160
rect 29736 8424 29788 8430
rect 29642 8392 29698 8401
rect 29736 8366 29788 8372
rect 29642 8327 29698 8336
rect 29656 8090 29684 8327
rect 29840 8276 29868 9132
rect 29918 9072 29974 9081
rect 29918 9007 29974 9016
rect 30104 9036 30156 9042
rect 29932 8838 29960 9007
rect 30104 8978 30156 8984
rect 30012 8900 30064 8906
rect 30012 8842 30064 8848
rect 29920 8832 29972 8838
rect 29920 8774 29972 8780
rect 29918 8664 29974 8673
rect 29918 8599 29974 8608
rect 29932 8430 29960 8599
rect 30024 8566 30052 8842
rect 30116 8566 30144 8978
rect 30012 8560 30064 8566
rect 30012 8502 30064 8508
rect 30104 8560 30156 8566
rect 30104 8502 30156 8508
rect 30194 8528 30250 8537
rect 30194 8463 30196 8472
rect 30248 8463 30250 8472
rect 30196 8434 30248 8440
rect 29920 8424 29972 8430
rect 29920 8366 29972 8372
rect 29748 8248 29868 8276
rect 29644 8084 29696 8090
rect 29644 8026 29696 8032
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 29656 6390 29684 7346
rect 29748 6866 29776 8248
rect 29846 8188 30154 8208
rect 29846 8186 29852 8188
rect 29908 8186 29932 8188
rect 29988 8186 30012 8188
rect 30068 8186 30092 8188
rect 30148 8186 30154 8188
rect 29908 8134 29910 8186
rect 30090 8134 30092 8186
rect 29846 8132 29852 8134
rect 29908 8132 29932 8134
rect 29988 8132 30012 8134
rect 30068 8132 30092 8134
rect 30148 8132 30154 8134
rect 29846 8112 30154 8132
rect 29846 7100 30154 7120
rect 29846 7098 29852 7100
rect 29908 7098 29932 7100
rect 29988 7098 30012 7100
rect 30068 7098 30092 7100
rect 30148 7098 30154 7100
rect 29908 7046 29910 7098
rect 30090 7046 30092 7098
rect 29846 7044 29852 7046
rect 29908 7044 29932 7046
rect 29988 7044 30012 7046
rect 30068 7044 30092 7046
rect 30148 7044 30154 7046
rect 29846 7024 30154 7044
rect 29736 6860 29788 6866
rect 29736 6802 29788 6808
rect 30208 6458 30236 8434
rect 30300 7750 30328 9404
rect 30288 7744 30340 7750
rect 30288 7686 30340 7692
rect 30300 7585 30328 7686
rect 30286 7576 30342 7585
rect 30286 7511 30342 7520
rect 30288 7404 30340 7410
rect 30288 7346 30340 7352
rect 30196 6452 30248 6458
rect 30196 6394 30248 6400
rect 29644 6384 29696 6390
rect 29644 6326 29696 6332
rect 29656 5914 29684 6326
rect 29846 6012 30154 6032
rect 29846 6010 29852 6012
rect 29908 6010 29932 6012
rect 29988 6010 30012 6012
rect 30068 6010 30092 6012
rect 30148 6010 30154 6012
rect 29908 5958 29910 6010
rect 30090 5958 30092 6010
rect 29846 5956 29852 5958
rect 29908 5956 29932 5958
rect 29988 5956 30012 5958
rect 30068 5956 30092 5958
rect 30148 5956 30154 5958
rect 29846 5936 30154 5956
rect 30300 5914 30328 7346
rect 29644 5908 29696 5914
rect 29644 5850 29696 5856
rect 30288 5908 30340 5914
rect 30288 5850 30340 5856
rect 30392 5370 30420 9676
rect 30484 9178 30512 15535
rect 30576 15162 30604 19858
rect 30668 19334 30696 23598
rect 30748 23044 30800 23050
rect 30748 22986 30800 22992
rect 30760 20641 30788 22986
rect 30852 22778 30880 23752
rect 30840 22772 30892 22778
rect 30840 22714 30892 22720
rect 30852 21690 30880 22714
rect 30840 21684 30892 21690
rect 30840 21626 30892 21632
rect 30746 20632 30802 20641
rect 30746 20567 30802 20576
rect 30840 20528 30892 20534
rect 30840 20470 30892 20476
rect 30746 20360 30802 20369
rect 30746 20295 30802 20304
rect 30760 20262 30788 20295
rect 30748 20256 30800 20262
rect 30748 20198 30800 20204
rect 30852 19718 30880 20470
rect 30944 20262 30972 25774
rect 31036 22273 31064 26143
rect 31116 25152 31168 25158
rect 31116 25094 31168 25100
rect 31022 22264 31078 22273
rect 31022 22199 31078 22208
rect 30932 20256 30984 20262
rect 30932 20198 30984 20204
rect 30840 19712 30892 19718
rect 30840 19654 30892 19660
rect 30668 19306 30788 19334
rect 30760 18136 30788 19306
rect 30852 18680 30880 19654
rect 30944 19310 30972 20198
rect 30932 19304 30984 19310
rect 30932 19246 30984 19252
rect 31024 18692 31076 18698
rect 30852 18652 31024 18680
rect 31024 18634 31076 18640
rect 31036 18290 31064 18634
rect 31128 18340 31156 25094
rect 31220 23497 31248 26318
rect 31482 26279 31538 26288
rect 31484 26240 31536 26246
rect 31588 26217 31616 27270
rect 31668 26784 31720 26790
rect 31668 26726 31720 26732
rect 31484 26182 31536 26188
rect 31574 26208 31630 26217
rect 31392 25832 31444 25838
rect 31392 25774 31444 25780
rect 31496 25786 31524 26182
rect 31574 26143 31630 26152
rect 31588 25906 31616 26143
rect 31576 25900 31628 25906
rect 31576 25842 31628 25848
rect 31404 24698 31432 25774
rect 31496 25758 31616 25786
rect 31588 25498 31616 25758
rect 31576 25492 31628 25498
rect 31576 25434 31628 25440
rect 31588 25294 31616 25434
rect 31576 25288 31628 25294
rect 31482 25256 31538 25265
rect 31576 25230 31628 25236
rect 31482 25191 31484 25200
rect 31536 25191 31538 25200
rect 31484 25162 31536 25168
rect 31576 24812 31628 24818
rect 31680 24800 31708 26726
rect 31956 26382 31984 27775
rect 32218 27432 32274 27441
rect 32128 27396 32180 27402
rect 32218 27367 32274 27376
rect 32128 27338 32180 27344
rect 32036 26988 32088 26994
rect 32036 26930 32088 26936
rect 31944 26376 31996 26382
rect 31944 26318 31996 26324
rect 31852 26308 31904 26314
rect 31852 26250 31904 26256
rect 31760 25696 31812 25702
rect 31760 25638 31812 25644
rect 31772 24954 31800 25638
rect 31760 24948 31812 24954
rect 31760 24890 31812 24896
rect 31628 24772 31708 24800
rect 31576 24754 31628 24760
rect 31404 24670 31616 24698
rect 31300 24608 31352 24614
rect 31484 24608 31536 24614
rect 31352 24568 31432 24596
rect 31300 24550 31352 24556
rect 31298 24168 31354 24177
rect 31298 24103 31354 24112
rect 31206 23488 31262 23497
rect 31206 23423 31262 23432
rect 31208 22432 31260 22438
rect 31208 22374 31260 22380
rect 31220 22166 31248 22374
rect 31208 22160 31260 22166
rect 31208 22102 31260 22108
rect 31206 19544 31262 19553
rect 31206 19479 31262 19488
rect 31220 18902 31248 19479
rect 31208 18896 31260 18902
rect 31208 18838 31260 18844
rect 31208 18760 31260 18766
rect 31208 18702 31260 18708
rect 31128 18312 31174 18340
rect 31024 18284 31076 18290
rect 31024 18226 31076 18232
rect 31146 18204 31174 18312
rect 31220 18222 31248 18702
rect 31128 18176 31174 18204
rect 31208 18216 31260 18222
rect 30760 18108 31064 18136
rect 30838 18048 30894 18057
rect 30838 17983 30894 17992
rect 30656 17876 30708 17882
rect 30656 17818 30708 17824
rect 30668 17513 30696 17818
rect 30852 17542 30880 17983
rect 30840 17536 30892 17542
rect 30654 17504 30710 17513
rect 30840 17478 30892 17484
rect 30932 17536 30984 17542
rect 30932 17478 30984 17484
rect 30654 17439 30710 17448
rect 30656 17264 30708 17270
rect 30944 17252 30972 17478
rect 30708 17224 30972 17252
rect 30656 17206 30708 17212
rect 30654 16824 30710 16833
rect 30654 16759 30710 16768
rect 30668 15745 30696 16759
rect 30748 16176 30800 16182
rect 30748 16118 30800 16124
rect 30654 15736 30710 15745
rect 30654 15671 30710 15680
rect 30656 15360 30708 15366
rect 30656 15302 30708 15308
rect 30564 15156 30616 15162
rect 30564 15098 30616 15104
rect 30576 13870 30604 15098
rect 30668 14793 30696 15302
rect 30654 14784 30710 14793
rect 30654 14719 30710 14728
rect 30760 14634 30788 16118
rect 30852 16046 30880 17224
rect 30930 16824 30986 16833
rect 30930 16759 30986 16768
rect 30840 16040 30892 16046
rect 30840 15982 30892 15988
rect 30840 15904 30892 15910
rect 30840 15846 30892 15852
rect 30852 15366 30880 15846
rect 30840 15360 30892 15366
rect 30840 15302 30892 15308
rect 30840 15088 30892 15094
rect 30840 15030 30892 15036
rect 30668 14606 30788 14634
rect 30668 14414 30696 14606
rect 30746 14512 30802 14521
rect 30746 14447 30748 14456
rect 30800 14447 30802 14456
rect 30748 14418 30800 14424
rect 30656 14408 30708 14414
rect 30656 14350 30708 14356
rect 30656 14272 30708 14278
rect 30656 14214 30708 14220
rect 30564 13864 30616 13870
rect 30564 13806 30616 13812
rect 30562 11792 30618 11801
rect 30562 11727 30618 11736
rect 30576 11014 30604 11727
rect 30564 11008 30616 11014
rect 30564 10950 30616 10956
rect 30562 10704 30618 10713
rect 30562 10639 30618 10648
rect 30576 10130 30604 10639
rect 30564 10124 30616 10130
rect 30564 10066 30616 10072
rect 30564 9716 30616 9722
rect 30564 9658 30616 9664
rect 30576 9625 30604 9658
rect 30562 9616 30618 9625
rect 30562 9551 30618 9560
rect 30668 9450 30696 14214
rect 30748 13728 30800 13734
rect 30748 13670 30800 13676
rect 30760 13410 30788 13670
rect 30852 13512 30880 15030
rect 30944 13734 30972 16759
rect 31036 15162 31064 18108
rect 31024 15156 31076 15162
rect 31024 15098 31076 15104
rect 31022 15056 31078 15065
rect 31022 14991 31078 15000
rect 30932 13728 30984 13734
rect 30932 13670 30984 13676
rect 30852 13484 30972 13512
rect 30760 13382 30880 13410
rect 30746 12472 30802 12481
rect 30746 12407 30802 12416
rect 30760 11393 30788 12407
rect 30746 11384 30802 11393
rect 30746 11319 30802 11328
rect 30746 9888 30802 9897
rect 30746 9823 30802 9832
rect 30656 9444 30708 9450
rect 30656 9386 30708 9392
rect 30472 9172 30524 9178
rect 30472 9114 30524 9120
rect 30484 8106 30512 9114
rect 30656 9036 30708 9042
rect 30656 8978 30708 8984
rect 30564 8968 30616 8974
rect 30562 8936 30564 8945
rect 30616 8936 30618 8945
rect 30562 8871 30618 8880
rect 30576 8673 30604 8871
rect 30562 8664 30618 8673
rect 30562 8599 30618 8608
rect 30484 8078 30604 8106
rect 30472 8016 30524 8022
rect 30472 7958 30524 7964
rect 30484 7857 30512 7958
rect 30470 7848 30526 7857
rect 30470 7783 30526 7792
rect 30472 7744 30524 7750
rect 30472 7686 30524 7692
rect 30484 7274 30512 7686
rect 30472 7268 30524 7274
rect 30472 7210 30524 7216
rect 30484 5914 30512 7210
rect 30576 6458 30604 8078
rect 30668 7993 30696 8978
rect 30654 7984 30710 7993
rect 30654 7919 30710 7928
rect 30656 7812 30708 7818
rect 30656 7754 30708 7760
rect 30564 6452 30616 6458
rect 30564 6394 30616 6400
rect 30668 6186 30696 7754
rect 30760 7546 30788 9823
rect 30852 8294 30880 13382
rect 30944 11937 30972 13484
rect 31036 13433 31064 14991
rect 31128 14482 31156 18176
rect 31208 18158 31260 18164
rect 31220 16833 31248 18158
rect 31206 16824 31262 16833
rect 31206 16759 31262 16768
rect 31208 16584 31260 16590
rect 31208 16526 31260 16532
rect 31220 16114 31248 16526
rect 31208 16108 31260 16114
rect 31208 16050 31260 16056
rect 31116 14476 31168 14482
rect 31116 14418 31168 14424
rect 31114 13832 31170 13841
rect 31114 13767 31170 13776
rect 31128 13462 31156 13767
rect 31220 13530 31248 16050
rect 31208 13524 31260 13530
rect 31208 13466 31260 13472
rect 31116 13456 31168 13462
rect 31022 13424 31078 13433
rect 31116 13398 31168 13404
rect 31022 13359 31078 13368
rect 31208 13320 31260 13326
rect 31208 13262 31260 13268
rect 31116 12980 31168 12986
rect 31116 12922 31168 12928
rect 31128 12374 31156 12922
rect 31220 12850 31248 13262
rect 31312 12986 31340 24103
rect 31404 23186 31432 24568
rect 31484 24550 31536 24556
rect 31496 24138 31524 24550
rect 31484 24132 31536 24138
rect 31484 24074 31536 24080
rect 31392 23180 31444 23186
rect 31392 23122 31444 23128
rect 31404 22506 31432 23122
rect 31482 22808 31538 22817
rect 31482 22743 31538 22752
rect 31392 22500 31444 22506
rect 31392 22442 31444 22448
rect 31496 22094 31524 22743
rect 31588 22438 31616 24670
rect 31576 22432 31628 22438
rect 31576 22374 31628 22380
rect 31588 22234 31616 22374
rect 31576 22228 31628 22234
rect 31576 22170 31628 22176
rect 31404 22066 31524 22094
rect 31404 20346 31432 22066
rect 31576 21616 31628 21622
rect 31576 21558 31628 21564
rect 31588 21146 31616 21558
rect 31576 21140 31628 21146
rect 31576 21082 31628 21088
rect 31484 20528 31536 20534
rect 31588 20516 31616 21082
rect 31536 20488 31616 20516
rect 31484 20470 31536 20476
rect 31680 20466 31708 24772
rect 31864 24750 31892 26250
rect 32048 25294 32076 26930
rect 32036 25288 32088 25294
rect 31956 25248 32036 25276
rect 31956 25129 31984 25248
rect 32036 25230 32088 25236
rect 32036 25152 32088 25158
rect 31942 25120 31998 25129
rect 32036 25094 32088 25100
rect 31942 25055 31998 25064
rect 32048 24750 32076 25094
rect 32140 24818 32168 27338
rect 32232 25226 32260 27367
rect 32324 26994 32352 28154
rect 32864 28076 32916 28082
rect 32864 28018 32916 28024
rect 32876 27334 32904 28018
rect 34058 27704 34114 27713
rect 34058 27639 34114 27648
rect 33508 27532 33560 27538
rect 33508 27474 33560 27480
rect 32864 27328 32916 27334
rect 32864 27270 32916 27276
rect 33140 27328 33192 27334
rect 33140 27270 33192 27276
rect 32312 26988 32364 26994
rect 32312 26930 32364 26936
rect 32324 25702 32352 26930
rect 32588 26784 32640 26790
rect 32588 26726 32640 26732
rect 32496 26376 32548 26382
rect 32494 26344 32496 26353
rect 32548 26344 32550 26353
rect 32494 26279 32550 26288
rect 32600 26228 32628 26726
rect 32508 26200 32628 26228
rect 32680 26240 32732 26246
rect 32508 26042 32536 26200
rect 32680 26182 32732 26188
rect 32496 26036 32548 26042
rect 32496 25978 32548 25984
rect 32312 25696 32364 25702
rect 32312 25638 32364 25644
rect 32404 25696 32456 25702
rect 32404 25638 32456 25644
rect 32220 25220 32272 25226
rect 32220 25162 32272 25168
rect 32310 25120 32366 25129
rect 32310 25055 32366 25064
rect 32324 24954 32352 25055
rect 32220 24948 32272 24954
rect 32220 24890 32272 24896
rect 32312 24948 32364 24954
rect 32312 24890 32364 24896
rect 32232 24818 32260 24890
rect 32128 24812 32180 24818
rect 32128 24754 32180 24760
rect 32220 24812 32272 24818
rect 32220 24754 32272 24760
rect 31852 24744 31904 24750
rect 31852 24686 31904 24692
rect 32036 24744 32088 24750
rect 32036 24686 32088 24692
rect 31760 24676 31812 24682
rect 31760 24618 31812 24624
rect 31772 23089 31800 24618
rect 31864 23254 31892 24686
rect 32036 24608 32088 24614
rect 32140 24596 32168 24754
rect 32310 24712 32366 24721
rect 32310 24647 32366 24656
rect 32140 24568 32260 24596
rect 32036 24550 32088 24556
rect 32048 24138 32076 24550
rect 32126 24168 32182 24177
rect 32036 24132 32088 24138
rect 32126 24103 32182 24112
rect 32036 24074 32088 24080
rect 32140 24070 32168 24103
rect 32128 24064 32180 24070
rect 32128 24006 32180 24012
rect 32034 23760 32090 23769
rect 32034 23695 32090 23704
rect 31944 23588 31996 23594
rect 31944 23530 31996 23536
rect 31956 23322 31984 23530
rect 31944 23316 31996 23322
rect 31944 23258 31996 23264
rect 31852 23248 31904 23254
rect 31852 23190 31904 23196
rect 31758 23080 31814 23089
rect 31758 23015 31814 23024
rect 31852 22568 31904 22574
rect 31852 22510 31904 22516
rect 31864 21418 31892 22510
rect 31944 21888 31996 21894
rect 31944 21830 31996 21836
rect 31956 21729 31984 21830
rect 31942 21720 31998 21729
rect 31942 21655 31998 21664
rect 31852 21412 31904 21418
rect 31852 21354 31904 21360
rect 32048 21026 32076 23695
rect 32128 23316 32180 23322
rect 32128 23258 32180 23264
rect 32140 22982 32168 23258
rect 32128 22976 32180 22982
rect 32128 22918 32180 22924
rect 32126 22808 32182 22817
rect 32126 22743 32182 22752
rect 32140 21128 32168 22743
rect 32232 21321 32260 24568
rect 32324 24206 32352 24647
rect 32416 24614 32444 25638
rect 32404 24608 32456 24614
rect 32404 24550 32456 24556
rect 32508 24426 32536 25978
rect 32588 25764 32640 25770
rect 32588 25706 32640 25712
rect 32600 25158 32628 25706
rect 32588 25152 32640 25158
rect 32588 25094 32640 25100
rect 32600 24954 32628 25094
rect 32588 24948 32640 24954
rect 32588 24890 32640 24896
rect 32692 24818 32720 26182
rect 32680 24812 32732 24818
rect 32680 24754 32732 24760
rect 32416 24398 32536 24426
rect 32312 24200 32364 24206
rect 32312 24142 32364 24148
rect 32416 22817 32444 24398
rect 32588 24268 32640 24274
rect 32588 24210 32640 24216
rect 32402 22808 32458 22817
rect 32402 22743 32458 22752
rect 32404 22500 32456 22506
rect 32404 22442 32456 22448
rect 32312 22024 32364 22030
rect 32312 21966 32364 21972
rect 32218 21312 32274 21321
rect 32218 21247 32274 21256
rect 32140 21100 32260 21128
rect 31956 20998 32076 21026
rect 32128 21004 32180 21010
rect 31668 20460 31720 20466
rect 31668 20402 31720 20408
rect 31404 20318 31616 20346
rect 31484 20256 31536 20262
rect 31484 20198 31536 20204
rect 31392 18284 31444 18290
rect 31392 18226 31444 18232
rect 31404 17542 31432 18226
rect 31392 17536 31444 17542
rect 31392 17478 31444 17484
rect 31496 17270 31524 20198
rect 31588 19378 31616 20318
rect 31576 19372 31628 19378
rect 31576 19314 31628 19320
rect 31588 17882 31616 19314
rect 31680 19258 31708 20402
rect 31852 19712 31904 19718
rect 31852 19654 31904 19660
rect 31680 19230 31800 19258
rect 31772 18834 31800 19230
rect 31760 18828 31812 18834
rect 31760 18770 31812 18776
rect 31772 17882 31800 18770
rect 31576 17876 31628 17882
rect 31576 17818 31628 17824
rect 31760 17876 31812 17882
rect 31760 17818 31812 17824
rect 31588 17762 31616 17818
rect 31588 17734 31800 17762
rect 31668 17672 31720 17678
rect 31668 17614 31720 17620
rect 31680 17338 31708 17614
rect 31668 17332 31720 17338
rect 31668 17274 31720 17280
rect 31484 17264 31536 17270
rect 31772 17218 31800 17734
rect 31864 17610 31892 19654
rect 31852 17604 31904 17610
rect 31852 17546 31904 17552
rect 31850 17504 31906 17513
rect 31850 17439 31906 17448
rect 31864 17338 31892 17439
rect 31852 17332 31904 17338
rect 31852 17274 31904 17280
rect 31484 17206 31536 17212
rect 31588 17190 31800 17218
rect 31390 17096 31446 17105
rect 31390 17031 31392 17040
rect 31444 17031 31446 17040
rect 31392 17002 31444 17008
rect 31392 16788 31444 16794
rect 31392 16730 31444 16736
rect 31300 12980 31352 12986
rect 31300 12922 31352 12928
rect 31208 12844 31260 12850
rect 31208 12786 31260 12792
rect 31312 12753 31340 12922
rect 31298 12744 31354 12753
rect 31298 12679 31354 12688
rect 31404 12628 31432 16730
rect 31484 16516 31536 16522
rect 31484 16458 31536 16464
rect 31496 16266 31524 16458
rect 31588 16425 31616 17190
rect 31668 17128 31720 17134
rect 31668 17070 31720 17076
rect 31760 17128 31812 17134
rect 31760 17070 31812 17076
rect 31850 17096 31906 17105
rect 31574 16416 31630 16425
rect 31574 16351 31630 16360
rect 31496 16250 31616 16266
rect 31496 16244 31628 16250
rect 31496 16238 31576 16244
rect 31576 16186 31628 16192
rect 31588 16046 31616 16186
rect 31576 16040 31628 16046
rect 31576 15982 31628 15988
rect 31588 15722 31616 15982
rect 31496 15694 31616 15722
rect 31496 15366 31524 15694
rect 31576 15428 31628 15434
rect 31576 15370 31628 15376
rect 31484 15360 31536 15366
rect 31588 15337 31616 15370
rect 31484 15302 31536 15308
rect 31574 15328 31630 15337
rect 31496 14006 31524 15302
rect 31574 15263 31630 15272
rect 31576 15156 31628 15162
rect 31576 15098 31628 15104
rect 31484 14000 31536 14006
rect 31484 13942 31536 13948
rect 31220 12600 31432 12628
rect 31116 12368 31168 12374
rect 31116 12310 31168 12316
rect 31220 12220 31248 12600
rect 31300 12368 31352 12374
rect 31484 12368 31536 12374
rect 31300 12310 31352 12316
rect 31482 12336 31484 12345
rect 31536 12336 31538 12345
rect 31128 12192 31248 12220
rect 31022 12064 31078 12073
rect 31022 11999 31078 12008
rect 30930 11928 30986 11937
rect 30930 11863 30986 11872
rect 30930 11656 30986 11665
rect 30930 11591 30986 11600
rect 30944 9110 30972 11591
rect 31036 11150 31064 11999
rect 31024 11144 31076 11150
rect 31024 11086 31076 11092
rect 31024 9920 31076 9926
rect 31024 9862 31076 9868
rect 31036 9722 31064 9862
rect 31024 9716 31076 9722
rect 31024 9658 31076 9664
rect 31128 9586 31156 12192
rect 31208 11076 31260 11082
rect 31208 11018 31260 11024
rect 31116 9580 31168 9586
rect 31116 9522 31168 9528
rect 31024 9512 31076 9518
rect 31024 9454 31076 9460
rect 30932 9104 30984 9110
rect 30932 9046 30984 9052
rect 30932 8492 30984 8498
rect 31036 8480 31064 9454
rect 30984 8452 31064 8480
rect 30932 8434 30984 8440
rect 30944 8294 30972 8434
rect 30840 8288 30892 8294
rect 30944 8266 31064 8294
rect 30840 8230 30892 8236
rect 30748 7540 30800 7546
rect 30748 7482 30800 7488
rect 30852 7002 30880 8230
rect 30932 7880 30984 7886
rect 30930 7848 30932 7857
rect 30984 7848 30986 7857
rect 31036 7818 31064 8266
rect 31128 8090 31156 9522
rect 31116 8084 31168 8090
rect 31116 8026 31168 8032
rect 31116 7880 31168 7886
rect 31116 7822 31168 7828
rect 30930 7783 30986 7792
rect 31024 7812 31076 7818
rect 31024 7754 31076 7760
rect 31022 7576 31078 7585
rect 31022 7511 31024 7520
rect 31076 7511 31078 7520
rect 31024 7482 31076 7488
rect 31128 7449 31156 7822
rect 31114 7440 31170 7449
rect 31114 7375 31170 7384
rect 30840 6996 30892 7002
rect 30840 6938 30892 6944
rect 30656 6180 30708 6186
rect 30656 6122 30708 6128
rect 31128 5914 31156 7375
rect 30472 5908 30524 5914
rect 30472 5850 30524 5856
rect 31116 5908 31168 5914
rect 31116 5850 31168 5856
rect 31128 5681 31156 5850
rect 31114 5672 31170 5681
rect 31114 5607 31170 5616
rect 30380 5364 30432 5370
rect 30380 5306 30432 5312
rect 30564 5364 30616 5370
rect 30564 5306 30616 5312
rect 29846 4924 30154 4944
rect 29846 4922 29852 4924
rect 29908 4922 29932 4924
rect 29988 4922 30012 4924
rect 30068 4922 30092 4924
rect 30148 4922 30154 4924
rect 29908 4870 29910 4922
rect 30090 4870 30092 4922
rect 29846 4868 29852 4870
rect 29908 4868 29932 4870
rect 29988 4868 30012 4870
rect 30068 4868 30092 4870
rect 30148 4868 30154 4870
rect 29846 4848 30154 4868
rect 29552 4820 29604 4826
rect 29552 4762 29604 4768
rect 29846 3836 30154 3856
rect 29846 3834 29852 3836
rect 29908 3834 29932 3836
rect 29988 3834 30012 3836
rect 30068 3834 30092 3836
rect 30148 3834 30154 3836
rect 29908 3782 29910 3834
rect 30090 3782 30092 3834
rect 29846 3780 29852 3782
rect 29908 3780 29932 3782
rect 29988 3780 30012 3782
rect 30068 3780 30092 3782
rect 30148 3780 30154 3782
rect 29846 3760 30154 3780
rect 29846 2748 30154 2768
rect 29846 2746 29852 2748
rect 29908 2746 29932 2748
rect 29988 2746 30012 2748
rect 30068 2746 30092 2748
rect 30148 2746 30154 2748
rect 29908 2694 29910 2746
rect 30090 2694 30092 2746
rect 29846 2692 29852 2694
rect 29908 2692 29932 2694
rect 29988 2692 30012 2694
rect 30068 2692 30092 2694
rect 30148 2692 30154 2694
rect 29846 2672 30154 2692
rect 30576 2650 30604 5306
rect 30564 2644 30616 2650
rect 30564 2586 30616 2592
rect 29920 2440 29972 2446
rect 29920 2382 29972 2388
rect 28446 1592 28502 1601
rect 28446 1527 28502 1536
rect 29932 800 29960 2382
rect 31220 2310 31248 11018
rect 31312 10742 31340 12310
rect 31482 12271 31538 12280
rect 31392 11824 31444 11830
rect 31392 11766 31444 11772
rect 31404 11529 31432 11766
rect 31588 11642 31616 15098
rect 31680 15094 31708 17070
rect 31772 16726 31800 17070
rect 31850 17031 31906 17040
rect 31864 16998 31892 17031
rect 31852 16992 31904 16998
rect 31852 16934 31904 16940
rect 31760 16720 31812 16726
rect 31760 16662 31812 16668
rect 31772 15178 31800 16662
rect 31852 16652 31904 16658
rect 31852 16594 31904 16600
rect 31864 15337 31892 16594
rect 31956 15434 31984 20998
rect 32128 20946 32180 20952
rect 32140 20602 32168 20946
rect 32128 20596 32180 20602
rect 32128 20538 32180 20544
rect 32232 19417 32260 21100
rect 32324 20777 32352 21966
rect 32416 21146 32444 22442
rect 32600 22001 32628 24210
rect 32586 21992 32642 22001
rect 32586 21927 32642 21936
rect 32692 21894 32720 24754
rect 32772 24404 32824 24410
rect 32772 24346 32824 24352
rect 32784 23798 32812 24346
rect 32876 24138 32904 27270
rect 33152 27062 33180 27270
rect 33048 27056 33100 27062
rect 33048 26998 33100 27004
rect 33140 27056 33192 27062
rect 33140 26998 33192 27004
rect 33060 26858 33088 26998
rect 33232 26920 33284 26926
rect 33232 26862 33284 26868
rect 33048 26852 33100 26858
rect 33048 26794 33100 26800
rect 32956 25832 33008 25838
rect 32956 25774 33008 25780
rect 32968 24274 32996 25774
rect 33060 25498 33088 26794
rect 33244 26382 33272 26862
rect 33324 26784 33376 26790
rect 33324 26726 33376 26732
rect 33232 26376 33284 26382
rect 33232 26318 33284 26324
rect 33140 26308 33192 26314
rect 33140 26250 33192 26256
rect 33048 25492 33100 25498
rect 33048 25434 33100 25440
rect 33048 25288 33100 25294
rect 33048 25230 33100 25236
rect 32956 24268 33008 24274
rect 32956 24210 33008 24216
rect 32864 24132 32916 24138
rect 32864 24074 32916 24080
rect 32968 23905 32996 24210
rect 32954 23896 33010 23905
rect 32954 23831 33010 23840
rect 32772 23792 32824 23798
rect 32772 23734 32824 23740
rect 33060 23730 33088 25230
rect 33152 24698 33180 26250
rect 33232 25152 33284 25158
rect 33232 25094 33284 25100
rect 33244 24886 33272 25094
rect 33232 24880 33284 24886
rect 33232 24822 33284 24828
rect 33152 24670 33272 24698
rect 33140 24608 33192 24614
rect 33140 24550 33192 24556
rect 33048 23724 33100 23730
rect 33048 23666 33100 23672
rect 32864 23656 32916 23662
rect 32864 23598 32916 23604
rect 32876 22778 32904 23598
rect 33152 23497 33180 24550
rect 33138 23488 33194 23497
rect 33138 23423 33194 23432
rect 32772 22772 32824 22778
rect 32772 22714 32824 22720
rect 32864 22772 32916 22778
rect 32864 22714 32916 22720
rect 32680 21888 32732 21894
rect 32680 21830 32732 21836
rect 32496 21480 32548 21486
rect 32548 21440 32628 21468
rect 32496 21422 32548 21428
rect 32494 21312 32550 21321
rect 32494 21247 32550 21256
rect 32404 21140 32456 21146
rect 32404 21082 32456 21088
rect 32404 20868 32456 20874
rect 32404 20810 32456 20816
rect 32310 20768 32366 20777
rect 32310 20703 32366 20712
rect 32416 20448 32444 20810
rect 32324 20420 32444 20448
rect 32324 19786 32352 20420
rect 32312 19780 32364 19786
rect 32312 19722 32364 19728
rect 32218 19408 32274 19417
rect 32218 19343 32274 19352
rect 32324 19310 32352 19722
rect 32312 19304 32364 19310
rect 32312 19246 32364 19252
rect 32404 18692 32456 18698
rect 32404 18634 32456 18640
rect 32128 18624 32180 18630
rect 32128 18566 32180 18572
rect 32036 18148 32088 18154
rect 32036 18090 32088 18096
rect 31944 15428 31996 15434
rect 31944 15370 31996 15376
rect 31850 15328 31906 15337
rect 31850 15263 31906 15272
rect 31772 15162 31892 15178
rect 31772 15156 31904 15162
rect 31772 15150 31852 15156
rect 31852 15098 31904 15104
rect 31668 15088 31720 15094
rect 31668 15030 31720 15036
rect 31760 14544 31812 14550
rect 31760 14486 31812 14492
rect 31666 14104 31722 14113
rect 31666 14039 31722 14048
rect 31680 13938 31708 14039
rect 31668 13932 31720 13938
rect 31668 13874 31720 13880
rect 31668 12844 31720 12850
rect 31668 12786 31720 12792
rect 31680 12306 31708 12786
rect 31668 12300 31720 12306
rect 31668 12242 31720 12248
rect 31668 12164 31720 12170
rect 31668 12106 31720 12112
rect 31496 11614 31616 11642
rect 31390 11520 31446 11529
rect 31390 11455 31446 11464
rect 31392 11212 31444 11218
rect 31392 11154 31444 11160
rect 31404 10742 31432 11154
rect 31496 10826 31524 11614
rect 31576 11552 31628 11558
rect 31680 11540 31708 12106
rect 31772 11665 31800 14486
rect 31864 13870 31892 15098
rect 32048 14890 32076 18090
rect 32140 15026 32168 18566
rect 32312 18216 32364 18222
rect 32312 18158 32364 18164
rect 32324 16572 32352 18158
rect 32232 16544 32352 16572
rect 32128 15020 32180 15026
rect 32128 14962 32180 14968
rect 32036 14884 32088 14890
rect 32036 14826 32088 14832
rect 31852 13864 31904 13870
rect 31852 13806 31904 13812
rect 31864 13444 31892 13806
rect 31944 13728 31996 13734
rect 31944 13670 31996 13676
rect 32036 13728 32088 13734
rect 32036 13670 32088 13676
rect 31956 13569 31984 13670
rect 31942 13560 31998 13569
rect 32048 13530 32076 13670
rect 31942 13495 31998 13504
rect 32036 13524 32088 13530
rect 32036 13466 32088 13472
rect 31864 13416 31984 13444
rect 31852 13320 31904 13326
rect 31852 13262 31904 13268
rect 31758 11656 31814 11665
rect 31758 11591 31814 11600
rect 31680 11512 31800 11540
rect 31576 11494 31628 11500
rect 31588 11121 31616 11494
rect 31668 11212 31720 11218
rect 31668 11154 31720 11160
rect 31574 11112 31630 11121
rect 31574 11047 31630 11056
rect 31680 11014 31708 11154
rect 31772 11082 31800 11512
rect 31760 11076 31812 11082
rect 31760 11018 31812 11024
rect 31668 11008 31720 11014
rect 31668 10950 31720 10956
rect 31496 10798 31708 10826
rect 31300 10736 31352 10742
rect 31300 10678 31352 10684
rect 31392 10736 31444 10742
rect 31392 10678 31444 10684
rect 31496 10674 31524 10798
rect 31484 10668 31536 10674
rect 31484 10610 31536 10616
rect 31680 10062 31708 10798
rect 31668 10056 31720 10062
rect 31668 9998 31720 10004
rect 31576 9920 31628 9926
rect 31576 9862 31628 9868
rect 31300 9444 31352 9450
rect 31300 9386 31352 9392
rect 31484 9444 31536 9450
rect 31484 9386 31536 9392
rect 31312 8566 31340 9386
rect 31496 9353 31524 9386
rect 31482 9344 31538 9353
rect 31482 9279 31538 9288
rect 31588 9178 31616 9862
rect 31576 9172 31628 9178
rect 31576 9114 31628 9120
rect 31680 9110 31708 9998
rect 31772 9994 31800 11018
rect 31760 9988 31812 9994
rect 31760 9930 31812 9936
rect 31864 9897 31892 13262
rect 31956 12238 31984 13416
rect 32140 12458 32168 14962
rect 32232 12646 32260 16544
rect 32312 15632 32364 15638
rect 32312 15574 32364 15580
rect 32324 15502 32352 15574
rect 32312 15496 32364 15502
rect 32312 15438 32364 15444
rect 32312 15360 32364 15366
rect 32312 15302 32364 15308
rect 32220 12640 32272 12646
rect 32220 12582 32272 12588
rect 32324 12481 32352 15302
rect 32416 14278 32444 18634
rect 32508 18154 32536 21247
rect 32496 18148 32548 18154
rect 32496 18090 32548 18096
rect 32494 17640 32550 17649
rect 32494 17575 32550 17584
rect 32508 17542 32536 17575
rect 32496 17536 32548 17542
rect 32496 17478 32548 17484
rect 32496 16516 32548 16522
rect 32496 16458 32548 16464
rect 32508 15473 32536 16458
rect 32494 15464 32550 15473
rect 32600 15434 32628 21440
rect 32678 20088 32734 20097
rect 32678 20023 32734 20032
rect 32692 19922 32720 20023
rect 32680 19916 32732 19922
rect 32680 19858 32732 19864
rect 32784 18222 32812 22714
rect 32876 22574 32904 22714
rect 32956 22704 33008 22710
rect 32956 22646 33008 22652
rect 32864 22568 32916 22574
rect 32864 22510 32916 22516
rect 32968 21622 32996 22646
rect 33140 22568 33192 22574
rect 33140 22510 33192 22516
rect 33152 22409 33180 22510
rect 33138 22400 33194 22409
rect 33138 22335 33194 22344
rect 33138 22128 33194 22137
rect 33138 22063 33194 22072
rect 33152 21894 33180 22063
rect 33140 21888 33192 21894
rect 33140 21830 33192 21836
rect 33046 21720 33102 21729
rect 33046 21655 33102 21664
rect 32956 21616 33008 21622
rect 32956 21558 33008 21564
rect 32968 20942 32996 21558
rect 33060 21486 33088 21655
rect 33048 21480 33100 21486
rect 33048 21422 33100 21428
rect 32956 20936 33008 20942
rect 32956 20878 33008 20884
rect 32968 20602 32996 20878
rect 32956 20596 33008 20602
rect 32956 20538 33008 20544
rect 32954 20224 33010 20233
rect 32954 20159 33010 20168
rect 32772 18216 32824 18222
rect 32772 18158 32824 18164
rect 32680 18148 32732 18154
rect 32680 18090 32732 18096
rect 32494 15399 32550 15408
rect 32588 15428 32640 15434
rect 32588 15370 32640 15376
rect 32692 15042 32720 18090
rect 32784 17649 32812 18158
rect 32862 17776 32918 17785
rect 32862 17711 32918 17720
rect 32770 17640 32826 17649
rect 32770 17575 32826 17584
rect 32772 16992 32824 16998
rect 32772 16934 32824 16940
rect 32784 15638 32812 16934
rect 32772 15632 32824 15638
rect 32772 15574 32824 15580
rect 32600 15014 32720 15042
rect 32600 14618 32628 15014
rect 32680 14952 32732 14958
rect 32680 14894 32732 14900
rect 32588 14612 32640 14618
rect 32588 14554 32640 14560
rect 32404 14272 32456 14278
rect 32404 14214 32456 14220
rect 32404 12912 32456 12918
rect 32402 12880 32404 12889
rect 32456 12880 32458 12889
rect 32402 12815 32458 12824
rect 32692 12594 32720 14894
rect 32508 12566 32720 12594
rect 32310 12472 32366 12481
rect 32140 12430 32260 12458
rect 31944 12232 31996 12238
rect 31944 12174 31996 12180
rect 31956 11762 31984 12174
rect 31944 11756 31996 11762
rect 31944 11698 31996 11704
rect 31942 11248 31998 11257
rect 31942 11183 31998 11192
rect 31956 10690 31984 11183
rect 31956 10662 32168 10690
rect 32036 10600 32088 10606
rect 32036 10542 32088 10548
rect 31944 10464 31996 10470
rect 31944 10406 31996 10412
rect 31956 10130 31984 10406
rect 31944 10124 31996 10130
rect 31944 10066 31996 10072
rect 31942 10024 31998 10033
rect 31942 9959 31998 9968
rect 31850 9888 31906 9897
rect 31850 9823 31906 9832
rect 31852 9716 31904 9722
rect 31852 9658 31904 9664
rect 31864 9217 31892 9658
rect 31956 9654 31984 9959
rect 31944 9648 31996 9654
rect 31944 9590 31996 9596
rect 31850 9208 31906 9217
rect 31850 9143 31906 9152
rect 31668 9104 31720 9110
rect 31668 9046 31720 9052
rect 31392 8832 31444 8838
rect 31390 8800 31392 8809
rect 31444 8800 31446 8809
rect 31390 8735 31446 8744
rect 31300 8560 31352 8566
rect 31300 8502 31352 8508
rect 31300 8288 31352 8294
rect 31300 8230 31352 8236
rect 31312 7002 31340 8230
rect 31404 7721 31432 8735
rect 31576 8356 31628 8362
rect 31576 8298 31628 8304
rect 31588 8129 31616 8298
rect 31680 8265 31708 9046
rect 31864 8786 31892 9143
rect 32048 8974 32076 10542
rect 32140 9897 32168 10662
rect 32126 9888 32182 9897
rect 32126 9823 32182 9832
rect 32126 9752 32182 9761
rect 32126 9687 32182 9696
rect 32036 8968 32088 8974
rect 32036 8910 32088 8916
rect 31864 8758 32076 8786
rect 31850 8664 31906 8673
rect 31850 8599 31906 8608
rect 31760 8492 31812 8498
rect 31760 8434 31812 8440
rect 31772 8276 31800 8434
rect 31666 8256 31722 8265
rect 31666 8191 31722 8200
rect 31764 8248 31800 8276
rect 31864 8276 31892 8599
rect 32048 8362 32076 8758
rect 32140 8498 32168 9687
rect 32232 8634 32260 12430
rect 32310 12407 32366 12416
rect 32404 12436 32456 12442
rect 32404 12378 32456 12384
rect 32312 12164 32364 12170
rect 32312 12106 32364 12112
rect 32324 11121 32352 12106
rect 32310 11112 32366 11121
rect 32310 11047 32366 11056
rect 32416 10146 32444 12378
rect 32508 10674 32536 12566
rect 32586 12472 32642 12481
rect 32586 12407 32642 12416
rect 32496 10668 32548 10674
rect 32496 10610 32548 10616
rect 32324 10118 32444 10146
rect 32324 9674 32352 10118
rect 32404 10056 32456 10062
rect 32508 10044 32536 10610
rect 32456 10016 32536 10044
rect 32404 9998 32456 10004
rect 32494 9888 32550 9897
rect 32494 9823 32550 9832
rect 32324 9646 32444 9674
rect 32508 9654 32536 9823
rect 32416 9586 32444 9646
rect 32496 9648 32548 9654
rect 32496 9590 32548 9596
rect 32404 9580 32456 9586
rect 32404 9522 32456 9528
rect 32312 9376 32364 9382
rect 32312 9318 32364 9324
rect 32324 9058 32352 9318
rect 32324 9042 32444 9058
rect 32324 9036 32456 9042
rect 32324 9030 32404 9036
rect 32220 8628 32272 8634
rect 32220 8570 32272 8576
rect 32128 8492 32180 8498
rect 32128 8434 32180 8440
rect 32036 8356 32088 8362
rect 32036 8298 32088 8304
rect 31944 8288 31996 8294
rect 31864 8248 31944 8276
rect 31574 8120 31630 8129
rect 31764 8106 31792 8248
rect 31944 8230 31996 8236
rect 32034 8120 32090 8129
rect 31764 8078 31800 8106
rect 31574 8055 31630 8064
rect 31390 7712 31446 7721
rect 31390 7647 31446 7656
rect 31772 7546 31800 8078
rect 32034 8055 32090 8064
rect 31760 7540 31812 7546
rect 31760 7482 31812 7488
rect 31300 6996 31352 7002
rect 31300 6938 31352 6944
rect 32048 6730 32076 8055
rect 31944 6724 31996 6730
rect 31944 6666 31996 6672
rect 32036 6724 32088 6730
rect 32036 6666 32088 6672
rect 31956 6186 31984 6666
rect 32140 6458 32168 8434
rect 32218 8120 32274 8129
rect 32218 8055 32220 8064
rect 32272 8055 32274 8064
rect 32220 8026 32272 8032
rect 32324 7750 32352 9030
rect 32404 8978 32456 8984
rect 32600 8634 32628 12407
rect 32680 12164 32732 12170
rect 32680 12106 32732 12112
rect 32692 11830 32720 12106
rect 32680 11824 32732 11830
rect 32680 11766 32732 11772
rect 32692 10441 32720 11766
rect 32784 11286 32812 15574
rect 32876 15094 32904 17711
rect 32968 16998 32996 20159
rect 33046 19816 33102 19825
rect 33046 19751 33102 19760
rect 33060 18086 33088 19751
rect 33048 18080 33100 18086
rect 33048 18022 33100 18028
rect 33048 17604 33100 17610
rect 33048 17546 33100 17552
rect 33060 17270 33088 17546
rect 33048 17264 33100 17270
rect 33048 17206 33100 17212
rect 32956 16992 33008 16998
rect 32956 16934 33008 16940
rect 32956 16516 33008 16522
rect 33060 16504 33088 17206
rect 33152 16794 33180 21830
rect 33244 20913 33272 24670
rect 33336 24206 33364 26726
rect 33520 26042 33548 27474
rect 34072 27130 34100 27639
rect 34150 27432 34206 27441
rect 34150 27367 34152 27376
rect 34204 27367 34206 27376
rect 34152 27338 34204 27344
rect 34060 27124 34112 27130
rect 33888 27084 34060 27112
rect 33784 26308 33836 26314
rect 33784 26250 33836 26256
rect 33508 26036 33560 26042
rect 33508 25978 33560 25984
rect 33520 25294 33548 25978
rect 33692 25900 33744 25906
rect 33692 25842 33744 25848
rect 33704 25809 33732 25842
rect 33690 25800 33746 25809
rect 33690 25735 33746 25744
rect 33600 25696 33652 25702
rect 33600 25638 33652 25644
rect 33508 25288 33560 25294
rect 33428 25248 33508 25276
rect 33428 24256 33456 25248
rect 33508 25230 33560 25236
rect 33506 24576 33562 24585
rect 33506 24511 33562 24520
rect 33520 24410 33548 24511
rect 33508 24404 33560 24410
rect 33508 24346 33560 24352
rect 33428 24228 33548 24256
rect 33324 24200 33376 24206
rect 33324 24142 33376 24148
rect 33416 24132 33468 24138
rect 33416 24074 33468 24080
rect 33322 23624 33378 23633
rect 33322 23559 33378 23568
rect 33230 20904 33286 20913
rect 33230 20839 33286 20848
rect 33336 19922 33364 23559
rect 33428 20346 33456 24074
rect 33520 22930 33548 24228
rect 33612 23050 33640 25638
rect 33692 24200 33744 24206
rect 33692 24142 33744 24148
rect 33704 24018 33732 24142
rect 33796 24138 33824 26250
rect 33888 24342 33916 27084
rect 34060 27066 34112 27072
rect 33968 26444 34020 26450
rect 33968 26386 34020 26392
rect 34244 26444 34296 26450
rect 34244 26386 34296 26392
rect 33980 26081 34008 26386
rect 34150 26344 34206 26353
rect 34060 26308 34112 26314
rect 34150 26279 34206 26288
rect 34060 26250 34112 26256
rect 33966 26072 34022 26081
rect 33966 26007 34022 26016
rect 33968 24812 34020 24818
rect 33968 24754 34020 24760
rect 33876 24336 33928 24342
rect 33876 24278 33928 24284
rect 33876 24200 33928 24206
rect 33874 24168 33876 24177
rect 33928 24168 33930 24177
rect 33784 24132 33836 24138
rect 33874 24103 33930 24112
rect 33784 24074 33836 24080
rect 33704 23990 33824 24018
rect 33600 23044 33652 23050
rect 33600 22986 33652 22992
rect 33692 23044 33744 23050
rect 33692 22986 33744 22992
rect 33520 22902 33640 22930
rect 33506 22808 33562 22817
rect 33506 22743 33562 22752
rect 33520 21962 33548 22743
rect 33612 22556 33640 22902
rect 33704 22710 33732 22986
rect 33692 22704 33744 22710
rect 33692 22646 33744 22652
rect 33612 22528 33732 22556
rect 33704 22030 33732 22528
rect 33692 22024 33744 22030
rect 33690 21992 33692 22001
rect 33744 21992 33746 22001
rect 33508 21956 33560 21962
rect 33690 21927 33746 21936
rect 33508 21898 33560 21904
rect 33600 21344 33652 21350
rect 33600 21286 33652 21292
rect 33612 20534 33640 21286
rect 33600 20528 33652 20534
rect 33600 20470 33652 20476
rect 33428 20318 33548 20346
rect 33414 20224 33470 20233
rect 33414 20159 33470 20168
rect 33324 19916 33376 19922
rect 33324 19858 33376 19864
rect 33322 19680 33378 19689
rect 33428 19666 33456 20159
rect 33378 19638 33456 19666
rect 33322 19615 33378 19624
rect 33232 17332 33284 17338
rect 33232 17274 33284 17280
rect 33140 16788 33192 16794
rect 33140 16730 33192 16736
rect 33008 16476 33088 16504
rect 32956 16458 33008 16464
rect 32968 16250 32996 16458
rect 32956 16244 33008 16250
rect 32956 16186 33008 16192
rect 33048 15428 33100 15434
rect 33048 15370 33100 15376
rect 33140 15428 33192 15434
rect 33140 15370 33192 15376
rect 32864 15088 32916 15094
rect 32864 15030 32916 15036
rect 32864 14000 32916 14006
rect 32864 13942 32916 13948
rect 32876 12889 32904 13942
rect 32956 13728 33008 13734
rect 32956 13670 33008 13676
rect 32862 12880 32918 12889
rect 32862 12815 32918 12824
rect 32876 11830 32904 12815
rect 32864 11824 32916 11830
rect 32864 11766 32916 11772
rect 32862 11520 32918 11529
rect 32862 11455 32918 11464
rect 32772 11280 32824 11286
rect 32772 11222 32824 11228
rect 32678 10432 32734 10441
rect 32678 10367 32734 10376
rect 32692 10062 32720 10367
rect 32680 10056 32732 10062
rect 32680 9998 32732 10004
rect 32680 9444 32732 9450
rect 32680 9386 32732 9392
rect 32692 8838 32720 9386
rect 32876 9042 32904 11455
rect 32968 9178 32996 13670
rect 33060 12186 33088 15370
rect 33152 14414 33180 15370
rect 33140 14408 33192 14414
rect 33140 14350 33192 14356
rect 33060 12158 33180 12186
rect 33048 12096 33100 12102
rect 33048 12038 33100 12044
rect 33060 10713 33088 12038
rect 33152 11558 33180 12158
rect 33140 11552 33192 11558
rect 33140 11494 33192 11500
rect 33152 11082 33180 11494
rect 33140 11076 33192 11082
rect 33140 11018 33192 11024
rect 33244 10962 33272 17274
rect 33336 11014 33364 19615
rect 33416 19304 33468 19310
rect 33416 19246 33468 19252
rect 33428 18222 33456 19246
rect 33416 18216 33468 18222
rect 33416 18158 33468 18164
rect 33428 18086 33456 18158
rect 33416 18080 33468 18086
rect 33416 18022 33468 18028
rect 33520 16232 33548 20318
rect 33796 19961 33824 23990
rect 33980 23746 34008 24754
rect 34072 24177 34100 26250
rect 34164 24342 34192 26279
rect 34256 24562 34284 26386
rect 34428 25900 34480 25906
rect 34428 25842 34480 25848
rect 34336 25696 34388 25702
rect 34336 25638 34388 25644
rect 34348 24993 34376 25638
rect 34334 24984 34390 24993
rect 34334 24919 34390 24928
rect 34440 24682 34468 25842
rect 34624 25498 34652 29543
rect 34704 25696 34756 25702
rect 34704 25638 34756 25644
rect 34612 25492 34664 25498
rect 34612 25434 34664 25440
rect 34612 24812 34664 24818
rect 34612 24754 34664 24760
rect 34428 24676 34480 24682
rect 34428 24618 34480 24624
rect 34256 24534 34376 24562
rect 34152 24336 34204 24342
rect 34152 24278 34204 24284
rect 34244 24336 34296 24342
rect 34244 24278 34296 24284
rect 34058 24168 34114 24177
rect 34058 24103 34060 24112
rect 34112 24103 34114 24112
rect 34060 24074 34112 24080
rect 34256 24018 34284 24278
rect 33888 23730 34008 23746
rect 33876 23724 34008 23730
rect 33928 23718 34008 23724
rect 34072 23990 34284 24018
rect 33876 23666 33928 23672
rect 33888 23361 33916 23666
rect 33968 23656 34020 23662
rect 33968 23598 34020 23604
rect 33874 23352 33930 23361
rect 33874 23287 33930 23296
rect 33876 22568 33928 22574
rect 33876 22510 33928 22516
rect 33888 22234 33916 22510
rect 33876 22228 33928 22234
rect 33876 22170 33928 22176
rect 33782 19952 33838 19961
rect 33888 19922 33916 22170
rect 33980 21962 34008 23598
rect 34072 23118 34100 23990
rect 34244 23588 34296 23594
rect 34244 23530 34296 23536
rect 34152 23248 34204 23254
rect 34152 23190 34204 23196
rect 34060 23112 34112 23118
rect 34060 23054 34112 23060
rect 33968 21956 34020 21962
rect 33968 21898 34020 21904
rect 34072 21554 34100 23054
rect 34060 21548 34112 21554
rect 34060 21490 34112 21496
rect 34060 21004 34112 21010
rect 34060 20946 34112 20952
rect 33782 19887 33838 19896
rect 33876 19916 33928 19922
rect 33876 19858 33928 19864
rect 33692 19848 33744 19854
rect 33692 19790 33744 19796
rect 33598 19408 33654 19417
rect 33598 19343 33654 19352
rect 33428 16204 33548 16232
rect 33428 14822 33456 16204
rect 33508 16108 33560 16114
rect 33508 16050 33560 16056
rect 33416 14816 33468 14822
rect 33416 14758 33468 14764
rect 33520 13530 33548 16050
rect 33612 13870 33640 19343
rect 33704 18970 33732 19790
rect 33692 18964 33744 18970
rect 33692 18906 33744 18912
rect 33968 18692 34020 18698
rect 33968 18634 34020 18640
rect 33784 18420 33836 18426
rect 33784 18362 33836 18368
rect 33796 18222 33824 18362
rect 33784 18216 33836 18222
rect 33784 18158 33836 18164
rect 33874 18184 33930 18193
rect 33874 18119 33930 18128
rect 33692 17808 33744 17814
rect 33692 17750 33744 17756
rect 33704 15978 33732 17750
rect 33784 16788 33836 16794
rect 33784 16730 33836 16736
rect 33796 16114 33824 16730
rect 33888 16726 33916 18119
rect 33980 18086 34008 18634
rect 33968 18080 34020 18086
rect 33968 18022 34020 18028
rect 33980 17066 34008 18022
rect 33968 17060 34020 17066
rect 33968 17002 34020 17008
rect 33876 16720 33928 16726
rect 33876 16662 33928 16668
rect 33876 16448 33928 16454
rect 33874 16416 33876 16425
rect 33928 16416 33930 16425
rect 33874 16351 33930 16360
rect 33784 16108 33836 16114
rect 33784 16050 33836 16056
rect 33980 16046 34008 17002
rect 33876 16040 33928 16046
rect 33876 15982 33928 15988
rect 33968 16040 34020 16046
rect 33968 15982 34020 15988
rect 33692 15972 33744 15978
rect 33692 15914 33744 15920
rect 33692 14884 33744 14890
rect 33692 14826 33744 14832
rect 33600 13864 33652 13870
rect 33600 13806 33652 13812
rect 33508 13524 33560 13530
rect 33508 13466 33560 13472
rect 33416 12640 33468 12646
rect 33416 12582 33468 12588
rect 33152 10934 33272 10962
rect 33324 11008 33376 11014
rect 33324 10950 33376 10956
rect 33046 10704 33102 10713
rect 33046 10639 33102 10648
rect 33152 10606 33180 10934
rect 33324 10736 33376 10742
rect 33324 10678 33376 10684
rect 33140 10600 33192 10606
rect 33140 10542 33192 10548
rect 33336 10452 33364 10678
rect 33428 10470 33456 12582
rect 33520 11937 33548 13466
rect 33704 13410 33732 14826
rect 33888 14618 33916 15982
rect 33980 15434 34008 15982
rect 33968 15428 34020 15434
rect 33968 15370 34020 15376
rect 33876 14612 33928 14618
rect 33876 14554 33928 14560
rect 33968 14408 34020 14414
rect 33968 14350 34020 14356
rect 33784 14272 33836 14278
rect 33784 14214 33836 14220
rect 33796 13530 33824 14214
rect 33784 13524 33836 13530
rect 33784 13466 33836 13472
rect 33704 13382 33824 13410
rect 33600 12776 33652 12782
rect 33600 12718 33652 12724
rect 33612 12374 33640 12718
rect 33692 12708 33744 12714
rect 33692 12650 33744 12656
rect 33600 12368 33652 12374
rect 33600 12310 33652 12316
rect 33506 11928 33562 11937
rect 33506 11863 33562 11872
rect 33508 11076 33560 11082
rect 33508 11018 33560 11024
rect 33244 10424 33364 10452
rect 33416 10464 33468 10470
rect 33244 9994 33272 10424
rect 33416 10406 33468 10412
rect 33324 10124 33376 10130
rect 33324 10066 33376 10072
rect 33232 9988 33284 9994
rect 33232 9930 33284 9936
rect 33140 9716 33192 9722
rect 33140 9658 33192 9664
rect 33048 9648 33100 9654
rect 33046 9616 33048 9625
rect 33100 9616 33102 9625
rect 33046 9551 33102 9560
rect 32956 9172 33008 9178
rect 32956 9114 33008 9120
rect 32864 9036 32916 9042
rect 32864 8978 32916 8984
rect 33048 9036 33100 9042
rect 33048 8978 33100 8984
rect 32680 8832 32732 8838
rect 32680 8774 32732 8780
rect 32692 8634 32720 8774
rect 32588 8628 32640 8634
rect 32588 8570 32640 8576
rect 32680 8628 32732 8634
rect 32680 8570 32732 8576
rect 32956 8560 33008 8566
rect 32862 8528 32918 8537
rect 32956 8502 33008 8508
rect 32862 8463 32864 8472
rect 32916 8463 32918 8472
rect 32864 8434 32916 8440
rect 32680 8288 32732 8294
rect 32586 8256 32642 8265
rect 32680 8230 32732 8236
rect 32586 8191 32642 8200
rect 32312 7744 32364 7750
rect 32312 7686 32364 7692
rect 32600 7478 32628 8191
rect 32692 7546 32720 8230
rect 32968 8090 32996 8502
rect 33060 8498 33088 8978
rect 33048 8492 33100 8498
rect 33048 8434 33100 8440
rect 33048 8356 33100 8362
rect 33048 8298 33100 8304
rect 33060 8265 33088 8298
rect 33046 8256 33102 8265
rect 33046 8191 33102 8200
rect 32956 8084 33008 8090
rect 32956 8026 33008 8032
rect 33152 7954 33180 9658
rect 33336 9178 33364 10066
rect 33324 9172 33376 9178
rect 33324 9114 33376 9120
rect 33416 8628 33468 8634
rect 33416 8570 33468 8576
rect 33140 7948 33192 7954
rect 33140 7890 33192 7896
rect 32864 7880 32916 7886
rect 32864 7822 32916 7828
rect 32680 7540 32732 7546
rect 32680 7482 32732 7488
rect 32588 7472 32640 7478
rect 32588 7414 32640 7420
rect 32600 7002 32628 7414
rect 32772 7404 32824 7410
rect 32876 7392 32904 7822
rect 32824 7364 32904 7392
rect 32772 7346 32824 7352
rect 32588 6996 32640 7002
rect 32588 6938 32640 6944
rect 32784 6458 32812 7346
rect 33428 6662 33456 8570
rect 33416 6656 33468 6662
rect 33416 6598 33468 6604
rect 32128 6452 32180 6458
rect 32128 6394 32180 6400
rect 32772 6452 32824 6458
rect 32772 6394 32824 6400
rect 31944 6180 31996 6186
rect 31944 6122 31996 6128
rect 32220 5908 32272 5914
rect 32220 5850 32272 5856
rect 32232 5302 32260 5850
rect 32784 5778 32812 6394
rect 32862 5944 32918 5953
rect 32862 5879 32918 5888
rect 32876 5846 32904 5879
rect 33520 5846 33548 11018
rect 33704 10742 33732 12650
rect 33796 11558 33824 13382
rect 33876 12368 33928 12374
rect 33876 12310 33928 12316
rect 33784 11552 33836 11558
rect 33784 11494 33836 11500
rect 33782 11248 33838 11257
rect 33782 11183 33838 11192
rect 33796 11150 33824 11183
rect 33784 11144 33836 11150
rect 33784 11086 33836 11092
rect 33692 10736 33744 10742
rect 33692 10678 33744 10684
rect 33782 10704 33838 10713
rect 33782 10639 33838 10648
rect 33796 10538 33824 10639
rect 33692 10532 33744 10538
rect 33692 10474 33744 10480
rect 33784 10532 33836 10538
rect 33784 10474 33836 10480
rect 33704 10441 33732 10474
rect 33690 10432 33746 10441
rect 33690 10367 33746 10376
rect 33888 10282 33916 12310
rect 33980 12238 34008 14350
rect 34072 13326 34100 20946
rect 34164 20806 34192 23190
rect 34256 23050 34284 23530
rect 34348 23474 34376 24534
rect 34440 24274 34468 24618
rect 34520 24608 34572 24614
rect 34520 24550 34572 24556
rect 34428 24268 34480 24274
rect 34428 24210 34480 24216
rect 34426 23896 34482 23905
rect 34426 23831 34482 23840
rect 34440 23594 34468 23831
rect 34428 23588 34480 23594
rect 34428 23530 34480 23536
rect 34348 23446 34468 23474
rect 34336 23316 34388 23322
rect 34336 23258 34388 23264
rect 34244 23044 34296 23050
rect 34244 22986 34296 22992
rect 34242 22944 34298 22953
rect 34242 22879 34298 22888
rect 34256 21690 34284 22879
rect 34348 22030 34376 23258
rect 34336 22024 34388 22030
rect 34336 21966 34388 21972
rect 34244 21684 34296 21690
rect 34244 21626 34296 21632
rect 34256 20924 34284 21626
rect 34348 21078 34376 21966
rect 34336 21072 34388 21078
rect 34336 21014 34388 21020
rect 34440 21010 34468 23446
rect 34532 22982 34560 24550
rect 34520 22976 34572 22982
rect 34520 22918 34572 22924
rect 34520 22160 34572 22166
rect 34520 22102 34572 22108
rect 34428 21004 34480 21010
rect 34428 20946 34480 20952
rect 34532 20942 34560 22102
rect 34624 21622 34652 24754
rect 34716 24410 34744 25638
rect 34992 25498 35020 29679
rect 35346 29322 35402 30000
rect 39118 29880 39174 29889
rect 39118 29815 39174 29824
rect 35346 29294 35664 29322
rect 35346 29200 35402 29294
rect 35636 27606 35664 29294
rect 38200 28144 38252 28150
rect 37830 28112 37886 28121
rect 38200 28086 38252 28092
rect 37830 28047 37886 28056
rect 37464 28008 37516 28014
rect 37464 27950 37516 27956
rect 37372 27872 37424 27878
rect 37372 27814 37424 27820
rect 35348 27600 35400 27606
rect 35348 27542 35400 27548
rect 35624 27600 35676 27606
rect 35624 27542 35676 27548
rect 35070 25936 35126 25945
rect 35070 25871 35126 25880
rect 34796 25492 34848 25498
rect 34796 25434 34848 25440
rect 34980 25492 35032 25498
rect 34980 25434 35032 25440
rect 34704 24404 34756 24410
rect 34704 24346 34756 24352
rect 34808 23848 34836 25434
rect 35084 24721 35112 25871
rect 35256 25832 35308 25838
rect 35256 25774 35308 25780
rect 35164 24812 35216 24818
rect 35164 24754 35216 24760
rect 35070 24712 35126 24721
rect 35070 24647 35126 24656
rect 34888 24200 34940 24206
rect 34888 24142 34940 24148
rect 34716 23820 34836 23848
rect 34716 22982 34744 23820
rect 34796 23724 34848 23730
rect 34796 23666 34848 23672
rect 34704 22976 34756 22982
rect 34704 22918 34756 22924
rect 34704 22568 34756 22574
rect 34704 22510 34756 22516
rect 34612 21616 34664 21622
rect 34612 21558 34664 21564
rect 34520 20936 34572 20942
rect 34256 20896 34376 20924
rect 34152 20800 34204 20806
rect 34152 20742 34204 20748
rect 34242 20768 34298 20777
rect 34164 20466 34192 20742
rect 34242 20703 34298 20712
rect 34152 20460 34204 20466
rect 34152 20402 34204 20408
rect 34152 19168 34204 19174
rect 34152 19110 34204 19116
rect 34164 16998 34192 19110
rect 34152 16992 34204 16998
rect 34150 16960 34152 16969
rect 34204 16960 34206 16969
rect 34150 16895 34206 16904
rect 34150 16824 34206 16833
rect 34150 16759 34206 16768
rect 34164 16182 34192 16759
rect 34152 16176 34204 16182
rect 34152 16118 34204 16124
rect 34152 15972 34204 15978
rect 34152 15914 34204 15920
rect 34164 14958 34192 15914
rect 34152 14952 34204 14958
rect 34152 14894 34204 14900
rect 34152 14340 34204 14346
rect 34152 14282 34204 14288
rect 34164 13938 34192 14282
rect 34152 13932 34204 13938
rect 34152 13874 34204 13880
rect 34150 13696 34206 13705
rect 34150 13631 34206 13640
rect 34060 13320 34112 13326
rect 34060 13262 34112 13268
rect 34072 12782 34100 13262
rect 34164 12850 34192 13631
rect 34256 13258 34284 20703
rect 34348 20618 34376 20896
rect 34520 20878 34572 20884
rect 34716 20754 34744 22510
rect 34624 20726 34744 20754
rect 34348 20590 34560 20618
rect 34532 20398 34560 20590
rect 34336 20392 34388 20398
rect 34336 20334 34388 20340
rect 34520 20392 34572 20398
rect 34520 20334 34572 20340
rect 34348 18329 34376 20334
rect 34532 19378 34560 20334
rect 34624 19446 34652 20726
rect 34808 20618 34836 23666
rect 34900 23118 34928 24142
rect 34978 24032 35034 24041
rect 34978 23967 35034 23976
rect 34888 23112 34940 23118
rect 34888 23054 34940 23060
rect 34888 22976 34940 22982
rect 34888 22918 34940 22924
rect 34716 20590 34836 20618
rect 34612 19440 34664 19446
rect 34612 19382 34664 19388
rect 34520 19372 34572 19378
rect 34520 19314 34572 19320
rect 34716 19334 34744 20590
rect 34900 19786 34928 22918
rect 34992 19922 35020 23967
rect 35070 23896 35126 23905
rect 35070 23831 35126 23840
rect 35084 23730 35112 23831
rect 35072 23724 35124 23730
rect 35072 23666 35124 23672
rect 35072 23180 35124 23186
rect 35072 23122 35124 23128
rect 35084 23089 35112 23122
rect 35070 23080 35126 23089
rect 35070 23015 35126 23024
rect 35072 22228 35124 22234
rect 35072 22170 35124 22176
rect 35084 21865 35112 22170
rect 35176 21894 35204 24754
rect 35268 23186 35296 25774
rect 35360 23746 35388 27542
rect 37096 26920 37148 26926
rect 37096 26862 37148 26868
rect 35716 26784 35768 26790
rect 35716 26726 35768 26732
rect 35900 26784 35952 26790
rect 35900 26726 35952 26732
rect 35440 26512 35492 26518
rect 35440 26454 35492 26460
rect 35452 23866 35480 26454
rect 35728 26382 35756 26726
rect 35808 26512 35860 26518
rect 35806 26480 35808 26489
rect 35860 26480 35862 26489
rect 35806 26415 35862 26424
rect 35716 26376 35768 26382
rect 35912 26330 35940 26726
rect 36912 26580 36964 26586
rect 36912 26522 36964 26528
rect 35716 26318 35768 26324
rect 35820 26302 35940 26330
rect 36924 26314 36952 26522
rect 36176 26308 36228 26314
rect 35820 26246 35848 26302
rect 36176 26250 36228 26256
rect 36912 26308 36964 26314
rect 36912 26250 36964 26256
rect 35624 26240 35676 26246
rect 35624 26182 35676 26188
rect 35808 26240 35860 26246
rect 35808 26182 35860 26188
rect 35530 25800 35586 25809
rect 35530 25735 35532 25744
rect 35584 25735 35586 25744
rect 35532 25706 35584 25712
rect 35636 25430 35664 26182
rect 35716 25764 35768 25770
rect 35716 25706 35768 25712
rect 35532 25424 35584 25430
rect 35532 25366 35584 25372
rect 35624 25424 35676 25430
rect 35624 25366 35676 25372
rect 35544 24206 35572 25366
rect 35636 25294 35664 25366
rect 35728 25294 35756 25706
rect 35624 25288 35676 25294
rect 35624 25230 35676 25236
rect 35716 25288 35768 25294
rect 35716 25230 35768 25236
rect 35636 25158 35664 25230
rect 35624 25152 35676 25158
rect 35728 25129 35756 25230
rect 35900 25152 35952 25158
rect 35624 25094 35676 25100
rect 35714 25120 35770 25129
rect 35900 25094 35952 25100
rect 35714 25055 35770 25064
rect 35622 24984 35678 24993
rect 35622 24919 35678 24928
rect 35636 24818 35664 24919
rect 35624 24812 35676 24818
rect 35624 24754 35676 24760
rect 35532 24200 35584 24206
rect 35532 24142 35584 24148
rect 35624 24132 35676 24138
rect 35624 24074 35676 24080
rect 35532 24064 35584 24070
rect 35530 24032 35532 24041
rect 35584 24032 35586 24041
rect 35530 23967 35586 23976
rect 35440 23860 35492 23866
rect 35440 23802 35492 23808
rect 35360 23718 35572 23746
rect 35256 23180 35308 23186
rect 35256 23122 35308 23128
rect 35346 22672 35402 22681
rect 35346 22607 35402 22616
rect 35360 22137 35388 22607
rect 35346 22128 35402 22137
rect 35346 22063 35402 22072
rect 35164 21888 35216 21894
rect 35070 21856 35126 21865
rect 35164 21830 35216 21836
rect 35070 21791 35126 21800
rect 35072 21480 35124 21486
rect 35072 21422 35124 21428
rect 34980 19916 35032 19922
rect 34980 19858 35032 19864
rect 34888 19780 34940 19786
rect 34888 19722 34940 19728
rect 34716 19306 34836 19334
rect 34612 19168 34664 19174
rect 34612 19110 34664 19116
rect 34428 18896 34480 18902
rect 34428 18838 34480 18844
rect 34440 18737 34468 18838
rect 34624 18834 34652 19110
rect 34612 18828 34664 18834
rect 34612 18770 34664 18776
rect 34704 18760 34756 18766
rect 34426 18728 34482 18737
rect 34704 18702 34756 18708
rect 34426 18663 34482 18672
rect 34716 18630 34744 18702
rect 34704 18624 34756 18630
rect 34704 18566 34756 18572
rect 34716 18465 34744 18566
rect 34702 18456 34758 18465
rect 34702 18391 34758 18400
rect 34334 18320 34390 18329
rect 34334 18255 34390 18264
rect 34704 18216 34756 18222
rect 34334 18184 34390 18193
rect 34704 18158 34756 18164
rect 34334 18119 34390 18128
rect 34348 17134 34376 18119
rect 34716 17610 34744 18158
rect 34808 18057 34836 19306
rect 34794 18048 34850 18057
rect 34794 17983 34850 17992
rect 34704 17604 34756 17610
rect 34704 17546 34756 17552
rect 34808 17320 34836 17983
rect 34900 17542 34928 19722
rect 35084 18630 35112 21422
rect 35348 20528 35400 20534
rect 35348 20470 35400 20476
rect 35164 20392 35216 20398
rect 35164 20334 35216 20340
rect 35176 20262 35204 20334
rect 35164 20256 35216 20262
rect 35164 20198 35216 20204
rect 35162 19952 35218 19961
rect 35162 19887 35218 19896
rect 35072 18624 35124 18630
rect 35072 18566 35124 18572
rect 35070 18456 35126 18465
rect 35070 18391 35126 18400
rect 35084 18222 35112 18391
rect 35072 18216 35124 18222
rect 35072 18158 35124 18164
rect 35072 17604 35124 17610
rect 35072 17546 35124 17552
rect 34888 17536 34940 17542
rect 34888 17478 34940 17484
rect 34808 17292 35020 17320
rect 34336 17128 34388 17134
rect 34888 17128 34940 17134
rect 34336 17070 34388 17076
rect 34702 17096 34758 17105
rect 34348 16833 34376 17070
rect 34888 17070 34940 17076
rect 34702 17031 34758 17040
rect 34334 16824 34390 16833
rect 34334 16759 34390 16768
rect 34716 16658 34744 17031
rect 34704 16652 34756 16658
rect 34704 16594 34756 16600
rect 34520 16516 34572 16522
rect 34520 16458 34572 16464
rect 34336 16448 34388 16454
rect 34336 16390 34388 16396
rect 34244 13252 34296 13258
rect 34244 13194 34296 13200
rect 34152 12844 34204 12850
rect 34152 12786 34204 12792
rect 34060 12776 34112 12782
rect 34060 12718 34112 12724
rect 34072 12646 34100 12718
rect 34060 12640 34112 12646
rect 34060 12582 34112 12588
rect 33968 12232 34020 12238
rect 33968 12174 34020 12180
rect 34244 12232 34296 12238
rect 34244 12174 34296 12180
rect 34060 11756 34112 11762
rect 34060 11698 34112 11704
rect 33968 11552 34020 11558
rect 33968 11494 34020 11500
rect 33980 11150 34008 11494
rect 34072 11218 34100 11698
rect 34256 11218 34284 12174
rect 34348 11694 34376 16390
rect 34426 15464 34482 15473
rect 34426 15399 34482 15408
rect 34440 15162 34468 15399
rect 34428 15156 34480 15162
rect 34428 15098 34480 15104
rect 34532 14550 34560 16458
rect 34612 16244 34664 16250
rect 34612 16186 34664 16192
rect 34624 15502 34652 16186
rect 34612 15496 34664 15502
rect 34612 15438 34664 15444
rect 34612 15360 34664 15366
rect 34612 15302 34664 15308
rect 34520 14544 34572 14550
rect 34520 14486 34572 14492
rect 34520 14408 34572 14414
rect 34518 14376 34520 14385
rect 34572 14376 34574 14385
rect 34518 14311 34574 14320
rect 34428 12912 34480 12918
rect 34428 12854 34480 12860
rect 34336 11688 34388 11694
rect 34336 11630 34388 11636
rect 34060 11212 34112 11218
rect 34060 11154 34112 11160
rect 34244 11212 34296 11218
rect 34244 11154 34296 11160
rect 33968 11144 34020 11150
rect 33968 11086 34020 11092
rect 33968 11008 34020 11014
rect 33968 10950 34020 10956
rect 33980 10470 34008 10950
rect 33968 10464 34020 10470
rect 33968 10406 34020 10412
rect 33704 10254 33916 10282
rect 33704 8974 33732 10254
rect 33784 9920 33836 9926
rect 33784 9862 33836 9868
rect 33876 9920 33928 9926
rect 33876 9862 33928 9868
rect 33692 8968 33744 8974
rect 33692 8910 33744 8916
rect 33600 8084 33652 8090
rect 33600 8026 33652 8032
rect 33612 7993 33640 8026
rect 33598 7984 33654 7993
rect 33796 7954 33824 9862
rect 33888 9761 33916 9862
rect 33874 9752 33930 9761
rect 33874 9687 33930 9696
rect 33598 7919 33654 7928
rect 33784 7948 33836 7954
rect 33784 7890 33836 7896
rect 33796 6798 33824 7890
rect 33888 7546 33916 9687
rect 33980 8634 34008 10406
rect 34072 9994 34100 11154
rect 34152 11008 34204 11014
rect 34152 10950 34204 10956
rect 34164 10674 34192 10950
rect 34152 10668 34204 10674
rect 34152 10610 34204 10616
rect 34244 10668 34296 10674
rect 34244 10610 34296 10616
rect 34152 10532 34204 10538
rect 34152 10474 34204 10480
rect 34164 10282 34192 10474
rect 34256 10441 34284 10610
rect 34242 10432 34298 10441
rect 34242 10367 34298 10376
rect 34164 10254 34284 10282
rect 34152 10192 34204 10198
rect 34152 10134 34204 10140
rect 34164 10033 34192 10134
rect 34256 10130 34284 10254
rect 34244 10124 34296 10130
rect 34244 10066 34296 10072
rect 34150 10024 34206 10033
rect 34060 9988 34112 9994
rect 34150 9959 34206 9968
rect 34060 9930 34112 9936
rect 34164 9926 34192 9959
rect 34152 9920 34204 9926
rect 34072 9868 34152 9874
rect 34072 9862 34204 9868
rect 34072 9846 34192 9862
rect 33968 8628 34020 8634
rect 33968 8570 34020 8576
rect 33968 7880 34020 7886
rect 33966 7848 33968 7857
rect 34020 7848 34022 7857
rect 33966 7783 34022 7792
rect 33876 7540 33928 7546
rect 33876 7482 33928 7488
rect 34072 6866 34100 9846
rect 34164 9797 34192 9846
rect 34152 9648 34204 9654
rect 34152 9590 34204 9596
rect 34164 8673 34192 9590
rect 34244 9580 34296 9586
rect 34244 9522 34296 9528
rect 34256 9450 34284 9522
rect 34244 9444 34296 9450
rect 34244 9386 34296 9392
rect 34348 9042 34376 11630
rect 34440 10130 34468 12854
rect 34624 12434 34652 15302
rect 34716 15201 34744 16594
rect 34796 16040 34848 16046
rect 34796 15982 34848 15988
rect 34702 15192 34758 15201
rect 34702 15127 34758 15136
rect 34704 14952 34756 14958
rect 34704 14894 34756 14900
rect 34716 13841 34744 14894
rect 34702 13832 34758 13841
rect 34702 13767 34758 13776
rect 34702 13560 34758 13569
rect 34702 13495 34758 13504
rect 34532 12406 34652 12434
rect 34532 11014 34560 12406
rect 34716 11762 34744 13495
rect 34704 11756 34756 11762
rect 34704 11698 34756 11704
rect 34808 11540 34836 15982
rect 34624 11512 34836 11540
rect 34520 11008 34572 11014
rect 34520 10950 34572 10956
rect 34624 10849 34652 11512
rect 34794 11384 34850 11393
rect 34794 11319 34796 11328
rect 34848 11319 34850 11328
rect 34796 11290 34848 11296
rect 34796 11212 34848 11218
rect 34796 11154 34848 11160
rect 34704 11144 34756 11150
rect 34704 11086 34756 11092
rect 34610 10840 34666 10849
rect 34520 10804 34572 10810
rect 34610 10775 34666 10784
rect 34520 10746 34572 10752
rect 34428 10124 34480 10130
rect 34428 10066 34480 10072
rect 34532 10062 34560 10746
rect 34612 10464 34664 10470
rect 34612 10406 34664 10412
rect 34624 10146 34652 10406
rect 34716 10266 34744 11086
rect 34808 11014 34836 11154
rect 34796 11008 34848 11014
rect 34796 10950 34848 10956
rect 34796 10668 34848 10674
rect 34796 10610 34848 10616
rect 34704 10260 34756 10266
rect 34704 10202 34756 10208
rect 34808 10198 34836 10610
rect 34796 10192 34848 10198
rect 34624 10118 34744 10146
rect 34796 10134 34848 10140
rect 34520 10056 34572 10062
rect 34520 9998 34572 10004
rect 34612 9988 34664 9994
rect 34612 9930 34664 9936
rect 34520 9920 34572 9926
rect 34520 9862 34572 9868
rect 34532 9761 34560 9862
rect 34518 9752 34574 9761
rect 34518 9687 34574 9696
rect 34426 9616 34482 9625
rect 34426 9551 34428 9560
rect 34480 9551 34482 9560
rect 34428 9522 34480 9528
rect 34440 9178 34468 9522
rect 34520 9376 34572 9382
rect 34520 9318 34572 9324
rect 34428 9172 34480 9178
rect 34428 9114 34480 9120
rect 34336 9036 34388 9042
rect 34336 8978 34388 8984
rect 34244 8968 34296 8974
rect 34244 8910 34296 8916
rect 34150 8664 34206 8673
rect 34150 8599 34152 8608
rect 34204 8599 34206 8608
rect 34152 8570 34204 8576
rect 34256 6866 34284 8910
rect 34428 8900 34480 8906
rect 34428 8842 34480 8848
rect 34440 7206 34468 8842
rect 34532 7313 34560 9318
rect 34624 8634 34652 9930
rect 34716 9897 34744 10118
rect 34900 10033 34928 17070
rect 34992 14521 35020 17292
rect 35084 16658 35112 17546
rect 35072 16652 35124 16658
rect 35072 16594 35124 16600
rect 35084 16046 35112 16594
rect 35072 16040 35124 16046
rect 35072 15982 35124 15988
rect 34978 14512 35034 14521
rect 34978 14447 35034 14456
rect 34980 14340 35032 14346
rect 34980 14282 35032 14288
rect 34886 10024 34942 10033
rect 34886 9959 34942 9968
rect 34702 9888 34758 9897
rect 34702 9823 34758 9832
rect 34716 8906 34744 9823
rect 34992 9738 35020 14282
rect 35084 14090 35112 15982
rect 35176 14226 35204 19887
rect 35360 19768 35388 20470
rect 35440 19780 35492 19786
rect 35360 19740 35440 19768
rect 35440 19722 35492 19728
rect 35440 19440 35492 19446
rect 35440 19382 35492 19388
rect 35452 18698 35480 19382
rect 35256 18692 35308 18698
rect 35256 18634 35308 18640
rect 35440 18692 35492 18698
rect 35440 18634 35492 18640
rect 35268 16522 35296 18634
rect 35440 16720 35492 16726
rect 35440 16662 35492 16668
rect 35256 16516 35308 16522
rect 35256 16458 35308 16464
rect 35268 16250 35296 16458
rect 35256 16244 35308 16250
rect 35256 16186 35308 16192
rect 35348 16244 35400 16250
rect 35348 16186 35400 16192
rect 35268 15094 35296 16186
rect 35360 15910 35388 16186
rect 35348 15904 35400 15910
rect 35348 15846 35400 15852
rect 35256 15088 35308 15094
rect 35256 15030 35308 15036
rect 35452 14521 35480 16662
rect 35438 14512 35494 14521
rect 35438 14447 35494 14456
rect 35176 14198 35296 14226
rect 35084 14062 35204 14090
rect 35072 14000 35124 14006
rect 35072 13942 35124 13948
rect 34808 9710 35020 9738
rect 35084 9722 35112 13942
rect 35176 13326 35204 14062
rect 35268 13569 35296 14198
rect 35348 13864 35400 13870
rect 35348 13806 35400 13812
rect 35254 13560 35310 13569
rect 35254 13495 35310 13504
rect 35164 13320 35216 13326
rect 35164 13262 35216 13268
rect 35176 12850 35204 13262
rect 35254 12880 35310 12889
rect 35164 12844 35216 12850
rect 35254 12815 35256 12824
rect 35164 12786 35216 12792
rect 35308 12815 35310 12824
rect 35256 12786 35308 12792
rect 35256 12708 35308 12714
rect 35256 12650 35308 12656
rect 35268 12617 35296 12650
rect 35254 12608 35310 12617
rect 35254 12543 35310 12552
rect 35256 12232 35308 12238
rect 35256 12174 35308 12180
rect 35162 11248 35218 11257
rect 35162 11183 35164 11192
rect 35216 11183 35218 11192
rect 35164 11154 35216 11160
rect 35268 11150 35296 12174
rect 35256 11144 35308 11150
rect 35256 11086 35308 11092
rect 35164 10736 35216 10742
rect 35164 10678 35216 10684
rect 35176 10470 35204 10678
rect 35164 10464 35216 10470
rect 35164 10406 35216 10412
rect 35254 10432 35310 10441
rect 35254 10367 35310 10376
rect 35072 9716 35124 9722
rect 34704 8900 34756 8906
rect 34704 8842 34756 8848
rect 34612 8628 34664 8634
rect 34612 8570 34664 8576
rect 34716 7818 34744 8842
rect 34808 8129 34836 9710
rect 35072 9658 35124 9664
rect 35164 9716 35216 9722
rect 35164 9658 35216 9664
rect 34886 9616 34942 9625
rect 35176 9602 35204 9658
rect 34886 9551 34942 9560
rect 34980 9580 35032 9586
rect 34900 9353 34928 9551
rect 34980 9522 35032 9528
rect 35084 9574 35204 9602
rect 34886 9344 34942 9353
rect 34886 9279 34942 9288
rect 34992 8537 35020 9522
rect 35084 9217 35112 9574
rect 35162 9480 35218 9489
rect 35162 9415 35218 9424
rect 35176 9382 35204 9415
rect 35164 9376 35216 9382
rect 35164 9318 35216 9324
rect 35070 9208 35126 9217
rect 35268 9178 35296 10367
rect 35360 9654 35388 13806
rect 35440 13252 35492 13258
rect 35440 13194 35492 13200
rect 35452 12646 35480 13194
rect 35440 12640 35492 12646
rect 35440 12582 35492 12588
rect 35544 12238 35572 23718
rect 35636 21622 35664 24074
rect 35728 23730 35756 25055
rect 35808 24812 35860 24818
rect 35808 24754 35860 24760
rect 35716 23724 35768 23730
rect 35716 23666 35768 23672
rect 35728 23633 35756 23666
rect 35714 23624 35770 23633
rect 35714 23559 35770 23568
rect 35624 21616 35676 21622
rect 35820 21593 35848 24754
rect 35912 23866 35940 25094
rect 36188 24857 36216 26250
rect 36636 25900 36688 25906
rect 36636 25842 36688 25848
rect 36452 25696 36504 25702
rect 36452 25638 36504 25644
rect 36360 25220 36412 25226
rect 36360 25162 36412 25168
rect 36174 24848 36230 24857
rect 36174 24783 36176 24792
rect 36228 24783 36230 24792
rect 36176 24754 36228 24760
rect 35992 24744 36044 24750
rect 35990 24712 35992 24721
rect 36044 24712 36046 24721
rect 35990 24647 36046 24656
rect 36176 24676 36228 24682
rect 36176 24618 36228 24624
rect 36084 24608 36136 24614
rect 36084 24550 36136 24556
rect 35992 24064 36044 24070
rect 35992 24006 36044 24012
rect 35900 23860 35952 23866
rect 35900 23802 35952 23808
rect 35912 23662 35940 23802
rect 35900 23656 35952 23662
rect 35900 23598 35952 23604
rect 35898 23488 35954 23497
rect 35898 23423 35954 23432
rect 35912 23066 35940 23423
rect 36004 23186 36032 24006
rect 35992 23180 36044 23186
rect 35992 23122 36044 23128
rect 35912 23038 36032 23066
rect 35898 22808 35954 22817
rect 35898 22743 35954 22752
rect 35912 22642 35940 22743
rect 35900 22636 35952 22642
rect 35900 22578 35952 22584
rect 35912 22234 35940 22578
rect 36004 22438 36032 23038
rect 35992 22432 36044 22438
rect 35992 22374 36044 22380
rect 35900 22228 35952 22234
rect 35900 22170 35952 22176
rect 36004 22001 36032 22374
rect 36096 22098 36124 24550
rect 36188 24206 36216 24618
rect 36268 24404 36320 24410
rect 36268 24346 36320 24352
rect 36280 24206 36308 24346
rect 36176 24200 36228 24206
rect 36176 24142 36228 24148
rect 36268 24200 36320 24206
rect 36268 24142 36320 24148
rect 36188 23769 36216 24142
rect 36268 24064 36320 24070
rect 36268 24006 36320 24012
rect 36174 23760 36230 23769
rect 36174 23695 36230 23704
rect 36176 23656 36228 23662
rect 36176 23598 36228 23604
rect 36188 22642 36216 23598
rect 36176 22636 36228 22642
rect 36176 22578 36228 22584
rect 36174 22264 36230 22273
rect 36174 22199 36176 22208
rect 36228 22199 36230 22208
rect 36176 22170 36228 22176
rect 36084 22092 36136 22098
rect 36084 22034 36136 22040
rect 35990 21992 36046 22001
rect 35990 21927 36046 21936
rect 36084 21956 36136 21962
rect 36084 21898 36136 21904
rect 35624 21558 35676 21564
rect 35806 21584 35862 21593
rect 35806 21519 35862 21528
rect 36096 21418 36124 21898
rect 35624 21412 35676 21418
rect 35624 21354 35676 21360
rect 36084 21412 36136 21418
rect 36084 21354 36136 21360
rect 35636 20233 35664 21354
rect 35808 21344 35860 21350
rect 35808 21286 35860 21292
rect 35716 20868 35768 20874
rect 35716 20810 35768 20816
rect 35728 20602 35756 20810
rect 35716 20596 35768 20602
rect 35716 20538 35768 20544
rect 35622 20224 35678 20233
rect 35622 20159 35678 20168
rect 35714 19544 35770 19553
rect 35714 19479 35770 19488
rect 35728 17105 35756 19479
rect 35820 19310 35848 21286
rect 36084 20460 36136 20466
rect 36084 20402 36136 20408
rect 36096 20058 36124 20402
rect 36084 20052 36136 20058
rect 36084 19994 36136 20000
rect 35898 19544 35954 19553
rect 35898 19479 35954 19488
rect 35912 19446 35940 19479
rect 35900 19440 35952 19446
rect 35900 19382 35952 19388
rect 35808 19304 35860 19310
rect 35808 19246 35860 19252
rect 35912 19122 35940 19382
rect 35820 19094 35940 19122
rect 35820 18630 35848 19094
rect 36280 18698 36308 24006
rect 36372 18834 36400 25162
rect 36464 24750 36492 25638
rect 36544 25152 36596 25158
rect 36544 25094 36596 25100
rect 36452 24744 36504 24750
rect 36452 24686 36504 24692
rect 36464 23798 36492 24686
rect 36452 23792 36504 23798
rect 36452 23734 36504 23740
rect 36556 23526 36584 25094
rect 36452 23520 36504 23526
rect 36544 23520 36596 23526
rect 36452 23462 36504 23468
rect 36542 23488 36544 23497
rect 36596 23488 36598 23497
rect 36464 22098 36492 23462
rect 36542 23423 36598 23432
rect 36648 23186 36676 25842
rect 36728 24812 36780 24818
rect 36728 24754 36780 24760
rect 36740 23594 36768 24754
rect 36910 24440 36966 24449
rect 36910 24375 36966 24384
rect 36820 24336 36872 24342
rect 36820 24278 36872 24284
rect 36832 23633 36860 24278
rect 36924 24070 36952 24375
rect 36912 24064 36964 24070
rect 36912 24006 36964 24012
rect 37002 24032 37058 24041
rect 36924 23662 36952 24006
rect 37002 23967 37058 23976
rect 37016 23866 37044 23967
rect 37004 23860 37056 23866
rect 37004 23802 37056 23808
rect 36912 23656 36964 23662
rect 36818 23624 36874 23633
rect 36728 23588 36780 23594
rect 36912 23598 36964 23604
rect 36818 23559 36874 23568
rect 36728 23530 36780 23536
rect 37108 23361 37136 26862
rect 37280 26036 37332 26042
rect 37280 25978 37332 25984
rect 37188 25356 37240 25362
rect 37188 25298 37240 25304
rect 37200 23730 37228 25298
rect 37292 25294 37320 25978
rect 37384 25498 37412 27814
rect 37372 25492 37424 25498
rect 37372 25434 37424 25440
rect 37280 25288 37332 25294
rect 37280 25230 37332 25236
rect 37280 24608 37332 24614
rect 37280 24550 37332 24556
rect 37292 23905 37320 24550
rect 37372 24200 37424 24206
rect 37372 24142 37424 24148
rect 37278 23896 37334 23905
rect 37278 23831 37334 23840
rect 37384 23730 37412 24142
rect 37188 23724 37240 23730
rect 37188 23666 37240 23672
rect 37372 23724 37424 23730
rect 37372 23666 37424 23672
rect 37476 23610 37504 27950
rect 37556 26784 37608 26790
rect 37556 26726 37608 26732
rect 37568 26450 37596 26726
rect 37556 26444 37608 26450
rect 37556 26386 37608 26392
rect 37740 25968 37792 25974
rect 37740 25910 37792 25916
rect 37646 25664 37702 25673
rect 37646 25599 37702 25608
rect 37556 25492 37608 25498
rect 37556 25434 37608 25440
rect 37292 23582 37504 23610
rect 36910 23352 36966 23361
rect 37094 23352 37150 23361
rect 36910 23287 36966 23296
rect 37016 23310 37094 23338
rect 36636 23180 36688 23186
rect 36636 23122 36688 23128
rect 36820 22976 36872 22982
rect 36820 22918 36872 22924
rect 36726 22672 36782 22681
rect 36556 22616 36726 22624
rect 36556 22596 36728 22616
rect 36452 22092 36504 22098
rect 36452 22034 36504 22040
rect 36556 21536 36584 22596
rect 36780 22607 36782 22616
rect 36728 22578 36780 22584
rect 36832 22574 36860 22918
rect 36820 22568 36872 22574
rect 36820 22510 36872 22516
rect 36728 22432 36780 22438
rect 36728 22374 36780 22380
rect 36740 22273 36768 22374
rect 36726 22264 36782 22273
rect 36636 22228 36688 22234
rect 36726 22199 36782 22208
rect 36636 22170 36688 22176
rect 36648 21554 36676 22170
rect 36924 22094 36952 23287
rect 37016 22506 37044 23310
rect 37094 23287 37150 23296
rect 37096 23044 37148 23050
rect 37096 22986 37148 22992
rect 37108 22778 37136 22986
rect 37188 22976 37240 22982
rect 37188 22918 37240 22924
rect 37096 22772 37148 22778
rect 37096 22714 37148 22720
rect 37004 22500 37056 22506
rect 37004 22442 37056 22448
rect 36832 22066 36952 22094
rect 36832 21570 36860 22066
rect 37200 22012 37228 22918
rect 37292 22778 37320 23582
rect 37372 23112 37424 23118
rect 37372 23054 37424 23060
rect 37464 23112 37516 23118
rect 37464 23054 37516 23060
rect 37280 22772 37332 22778
rect 37280 22714 37332 22720
rect 37384 22030 37412 23054
rect 37476 22094 37504 23054
rect 37568 22438 37596 25434
rect 37660 22438 37688 25599
rect 37556 22432 37608 22438
rect 37556 22374 37608 22380
rect 37648 22432 37700 22438
rect 37648 22374 37700 22380
rect 37476 22066 37688 22094
rect 37108 21984 37228 22012
rect 37372 22024 37424 22030
rect 37004 21888 37056 21894
rect 37004 21830 37056 21836
rect 36464 21508 36584 21536
rect 36636 21548 36688 21554
rect 36464 20534 36492 21508
rect 36636 21490 36688 21496
rect 36740 21542 36860 21570
rect 36912 21548 36964 21554
rect 36648 21434 36676 21490
rect 36556 21406 36676 21434
rect 36556 20806 36584 21406
rect 36636 21344 36688 21350
rect 36636 21286 36688 21292
rect 36544 20800 36596 20806
rect 36648 20777 36676 21286
rect 36544 20742 36596 20748
rect 36634 20768 36690 20777
rect 36452 20528 36504 20534
rect 36452 20470 36504 20476
rect 36452 19712 36504 19718
rect 36452 19654 36504 19660
rect 36360 18828 36412 18834
rect 36360 18770 36412 18776
rect 36268 18692 36320 18698
rect 36268 18634 36320 18640
rect 35808 18624 35860 18630
rect 35808 18566 35860 18572
rect 36174 18592 36230 18601
rect 36174 18527 36230 18536
rect 35900 17808 35952 17814
rect 35900 17750 35952 17756
rect 35714 17096 35770 17105
rect 35714 17031 35770 17040
rect 35808 17060 35860 17066
rect 35808 17002 35860 17008
rect 35820 16697 35848 17002
rect 35806 16688 35862 16697
rect 35806 16623 35862 16632
rect 35912 15688 35940 17750
rect 35992 17740 36044 17746
rect 35992 17682 36044 17688
rect 35636 15660 35940 15688
rect 35636 12753 35664 15660
rect 35806 15600 35862 15609
rect 35806 15535 35862 15544
rect 35820 15178 35848 15535
rect 35716 15156 35768 15162
rect 35820 15150 35940 15178
rect 35716 15098 35768 15104
rect 35728 15065 35756 15098
rect 35714 15056 35770 15065
rect 35714 14991 35770 15000
rect 35716 13320 35768 13326
rect 35716 13262 35768 13268
rect 35808 13320 35860 13326
rect 35808 13262 35860 13268
rect 35728 12850 35756 13262
rect 35716 12844 35768 12850
rect 35716 12786 35768 12792
rect 35820 12782 35848 13262
rect 35808 12776 35860 12782
rect 35622 12744 35678 12753
rect 35808 12718 35860 12724
rect 35622 12679 35678 12688
rect 35912 12646 35940 15150
rect 36004 14249 36032 17682
rect 36188 15434 36216 18527
rect 36268 18216 36320 18222
rect 36268 18158 36320 18164
rect 36280 17649 36308 18158
rect 36464 17864 36492 19654
rect 36556 19310 36584 20742
rect 36634 20703 36690 20712
rect 36636 20392 36688 20398
rect 36636 20334 36688 20340
rect 36648 19514 36676 20334
rect 36636 19508 36688 19514
rect 36636 19450 36688 19456
rect 36544 19304 36596 19310
rect 36544 19246 36596 19252
rect 36740 19174 36768 21542
rect 36912 21490 36964 21496
rect 36924 21321 36952 21490
rect 36910 21312 36966 21321
rect 36910 21247 36966 21256
rect 37016 21010 37044 21830
rect 37004 21004 37056 21010
rect 37004 20946 37056 20952
rect 36912 20868 36964 20874
rect 36912 20810 36964 20816
rect 36544 19168 36596 19174
rect 36544 19110 36596 19116
rect 36728 19168 36780 19174
rect 36728 19110 36780 19116
rect 36556 18902 36584 19110
rect 36544 18896 36596 18902
rect 36544 18838 36596 18844
rect 36726 18184 36782 18193
rect 36726 18119 36782 18128
rect 36372 17836 36492 17864
rect 36266 17640 36322 17649
rect 36266 17575 36322 17584
rect 36280 15745 36308 17575
rect 36266 15736 36322 15745
rect 36266 15671 36322 15680
rect 36176 15428 36228 15434
rect 36176 15370 36228 15376
rect 36188 15065 36216 15370
rect 36174 15056 36230 15065
rect 36174 14991 36230 15000
rect 36176 14816 36228 14822
rect 36174 14784 36176 14793
rect 36228 14784 36230 14793
rect 36174 14719 36230 14728
rect 36372 14634 36400 17836
rect 36740 17814 36768 18119
rect 36728 17808 36780 17814
rect 36728 17750 36780 17756
rect 36820 17740 36872 17746
rect 36820 17682 36872 17688
rect 36832 17649 36860 17682
rect 36818 17640 36874 17649
rect 36818 17575 36874 17584
rect 36728 17332 36780 17338
rect 36728 17274 36780 17280
rect 36452 16584 36504 16590
rect 36452 16526 36504 16532
rect 36464 15502 36492 16526
rect 36544 15564 36596 15570
rect 36544 15506 36596 15512
rect 36452 15496 36504 15502
rect 36450 15464 36452 15473
rect 36504 15464 36506 15473
rect 36450 15399 36506 15408
rect 36556 15094 36584 15506
rect 36544 15088 36596 15094
rect 36544 15030 36596 15036
rect 36188 14606 36400 14634
rect 36450 14648 36506 14657
rect 36084 14408 36136 14414
rect 36084 14350 36136 14356
rect 35990 14240 36046 14249
rect 35990 14175 36046 14184
rect 35990 13832 36046 13841
rect 35990 13767 35992 13776
rect 36044 13767 36046 13776
rect 35992 13738 36044 13744
rect 35990 13016 36046 13025
rect 35990 12951 36046 12960
rect 36004 12714 36032 12951
rect 35992 12708 36044 12714
rect 35992 12650 36044 12656
rect 35900 12640 35952 12646
rect 35622 12608 35678 12617
rect 35900 12582 35952 12588
rect 35622 12543 35678 12552
rect 35636 12374 35664 12543
rect 36096 12434 36124 14350
rect 36188 13274 36216 14606
rect 36450 14583 36506 14592
rect 36464 14550 36492 14583
rect 36452 14544 36504 14550
rect 36452 14486 36504 14492
rect 36360 14476 36412 14482
rect 36360 14418 36412 14424
rect 36268 13864 36320 13870
rect 36268 13806 36320 13812
rect 36280 13394 36308 13806
rect 36268 13388 36320 13394
rect 36268 13330 36320 13336
rect 36188 13246 36308 13274
rect 36176 12980 36228 12986
rect 36176 12922 36228 12928
rect 35912 12406 36124 12434
rect 35624 12368 35676 12374
rect 35624 12310 35676 12316
rect 35806 12336 35862 12345
rect 35806 12271 35862 12280
rect 35532 12232 35584 12238
rect 35532 12174 35584 12180
rect 35624 12096 35676 12102
rect 35624 12038 35676 12044
rect 35636 11762 35664 12038
rect 35714 11792 35770 11801
rect 35624 11756 35676 11762
rect 35820 11762 35848 12271
rect 35714 11727 35770 11736
rect 35808 11756 35860 11762
rect 35624 11698 35676 11704
rect 35636 11665 35664 11698
rect 35728 11694 35756 11727
rect 35808 11698 35860 11704
rect 35716 11688 35768 11694
rect 35622 11656 35678 11665
rect 35716 11630 35768 11636
rect 35622 11591 35678 11600
rect 35728 11370 35756 11630
rect 35806 11520 35862 11529
rect 35806 11455 35862 11464
rect 35636 11342 35756 11370
rect 35636 11218 35664 11342
rect 35716 11280 35768 11286
rect 35716 11222 35768 11228
rect 35624 11212 35676 11218
rect 35624 11154 35676 11160
rect 35728 11150 35756 11222
rect 35440 11144 35492 11150
rect 35440 11086 35492 11092
rect 35716 11144 35768 11150
rect 35716 11086 35768 11092
rect 35452 10418 35480 11086
rect 35624 11076 35676 11082
rect 35624 11018 35676 11024
rect 35636 10985 35664 11018
rect 35820 11014 35848 11455
rect 35716 11008 35768 11014
rect 35622 10976 35678 10985
rect 35716 10950 35768 10956
rect 35808 11008 35860 11014
rect 35808 10950 35860 10956
rect 35622 10911 35678 10920
rect 35728 10656 35756 10950
rect 35808 10668 35860 10674
rect 35728 10628 35808 10656
rect 35808 10610 35860 10616
rect 35530 10568 35586 10577
rect 35530 10503 35532 10512
rect 35584 10503 35586 10512
rect 35532 10474 35584 10480
rect 35716 10464 35768 10470
rect 35452 10390 35572 10418
rect 35716 10406 35768 10412
rect 35440 10056 35492 10062
rect 35440 9998 35492 10004
rect 35348 9648 35400 9654
rect 35348 9590 35400 9596
rect 35070 9143 35126 9152
rect 35256 9172 35308 9178
rect 35256 9114 35308 9120
rect 35256 9036 35308 9042
rect 35256 8978 35308 8984
rect 34978 8528 35034 8537
rect 35268 8498 35296 8978
rect 34978 8463 35034 8472
rect 35256 8492 35308 8498
rect 34794 8120 34850 8129
rect 34794 8055 34850 8064
rect 34992 8022 35020 8463
rect 35256 8434 35308 8440
rect 34980 8016 35032 8022
rect 34980 7958 35032 7964
rect 34704 7812 34756 7818
rect 34704 7754 34756 7760
rect 34992 7546 35020 7958
rect 35268 7818 35296 8434
rect 35256 7812 35308 7818
rect 35256 7754 35308 7760
rect 35348 7812 35400 7818
rect 35348 7754 35400 7760
rect 34980 7540 35032 7546
rect 34980 7482 35032 7488
rect 34518 7304 34574 7313
rect 35268 7274 35296 7754
rect 34518 7239 34574 7248
rect 35256 7268 35308 7274
rect 35256 7210 35308 7216
rect 35360 7206 35388 7754
rect 34428 7200 34480 7206
rect 34428 7142 34480 7148
rect 35348 7200 35400 7206
rect 35348 7142 35400 7148
rect 34060 6860 34112 6866
rect 34060 6802 34112 6808
rect 34244 6860 34296 6866
rect 34244 6802 34296 6808
rect 33784 6792 33836 6798
rect 33784 6734 33836 6740
rect 34256 6390 34284 6802
rect 34440 6798 34468 7142
rect 34428 6792 34480 6798
rect 34428 6734 34480 6740
rect 35360 6662 35388 7142
rect 35348 6656 35400 6662
rect 35452 6633 35480 9998
rect 35544 9042 35572 10390
rect 35728 10266 35756 10406
rect 35716 10260 35768 10266
rect 35716 10202 35768 10208
rect 35624 10056 35676 10062
rect 35624 9998 35676 10004
rect 35532 9036 35584 9042
rect 35532 8978 35584 8984
rect 35636 8430 35664 9998
rect 35728 8566 35756 10202
rect 35820 9926 35848 10610
rect 35808 9920 35860 9926
rect 35808 9862 35860 9868
rect 35716 8560 35768 8566
rect 35716 8502 35768 8508
rect 35624 8424 35676 8430
rect 35624 8366 35676 8372
rect 35912 7585 35940 12406
rect 36084 12164 36136 12170
rect 36084 12106 36136 12112
rect 36096 11778 36124 12106
rect 36188 11898 36216 12922
rect 36280 12850 36308 13246
rect 36268 12844 36320 12850
rect 36268 12786 36320 12792
rect 36266 12744 36322 12753
rect 36266 12679 36322 12688
rect 36280 12442 36308 12679
rect 36268 12436 36320 12442
rect 36268 12378 36320 12384
rect 36176 11892 36228 11898
rect 36176 11834 36228 11840
rect 36096 11750 36216 11778
rect 36084 11212 36136 11218
rect 36084 11154 36136 11160
rect 35992 11008 36044 11014
rect 35992 10950 36044 10956
rect 36004 10713 36032 10950
rect 35990 10704 36046 10713
rect 35990 10639 36046 10648
rect 36096 10033 36124 11154
rect 36082 10024 36138 10033
rect 36082 9959 36138 9968
rect 36188 8809 36216 11750
rect 36280 10962 36308 12378
rect 36372 11150 36400 14418
rect 36556 13938 36584 15030
rect 36636 14816 36688 14822
rect 36636 14758 36688 14764
rect 36648 14249 36676 14758
rect 36634 14240 36690 14249
rect 36634 14175 36690 14184
rect 36648 14074 36676 14175
rect 36636 14068 36688 14074
rect 36636 14010 36688 14016
rect 36544 13932 36596 13938
rect 36544 13874 36596 13880
rect 36452 13796 36504 13802
rect 36452 13738 36504 13744
rect 36464 11354 36492 13738
rect 36452 11348 36504 11354
rect 36452 11290 36504 11296
rect 36360 11144 36412 11150
rect 36412 11104 36492 11132
rect 36360 11086 36412 11092
rect 36280 10934 36400 10962
rect 36266 10840 36322 10849
rect 36266 10775 36268 10784
rect 36320 10775 36322 10784
rect 36268 10746 36320 10752
rect 36268 10668 36320 10674
rect 36268 10610 36320 10616
rect 36280 9518 36308 10610
rect 36268 9512 36320 9518
rect 36268 9454 36320 9460
rect 36280 9178 36308 9454
rect 36268 9172 36320 9178
rect 36268 9114 36320 9120
rect 36372 8906 36400 10934
rect 36464 10810 36492 11104
rect 36452 10804 36504 10810
rect 36452 10746 36504 10752
rect 36556 10198 36584 13874
rect 36740 13802 36768 17274
rect 36818 15872 36874 15881
rect 36818 15807 36874 15816
rect 36832 15570 36860 15807
rect 36820 15564 36872 15570
rect 36820 15506 36872 15512
rect 36820 14952 36872 14958
rect 36820 14894 36872 14900
rect 36832 14414 36860 14894
rect 36820 14408 36872 14414
rect 36820 14350 36872 14356
rect 36832 13870 36860 14350
rect 36924 14074 36952 20810
rect 37004 20528 37056 20534
rect 37004 20470 37056 20476
rect 37016 19666 37044 20470
rect 37108 19786 37136 21984
rect 37372 21966 37424 21972
rect 37556 22024 37608 22030
rect 37556 21966 37608 21972
rect 37188 21888 37240 21894
rect 37188 21830 37240 21836
rect 37280 21888 37332 21894
rect 37280 21830 37332 21836
rect 37200 20913 37228 21830
rect 37186 20904 37242 20913
rect 37186 20839 37242 20848
rect 37292 20330 37320 21830
rect 37568 21690 37596 21966
rect 37660 21690 37688 22066
rect 37556 21684 37608 21690
rect 37556 21626 37608 21632
rect 37648 21684 37700 21690
rect 37648 21626 37700 21632
rect 37464 21480 37516 21486
rect 37464 21422 37516 21428
rect 37280 20324 37332 20330
rect 37280 20266 37332 20272
rect 37476 19786 37504 21422
rect 37568 20058 37596 21626
rect 37646 20496 37702 20505
rect 37646 20431 37648 20440
rect 37700 20431 37702 20440
rect 37648 20402 37700 20408
rect 37556 20052 37608 20058
rect 37556 19994 37608 20000
rect 37096 19780 37148 19786
rect 37096 19722 37148 19728
rect 37464 19780 37516 19786
rect 37464 19722 37516 19728
rect 37556 19712 37608 19718
rect 37462 19680 37518 19689
rect 37016 19638 37136 19666
rect 37002 19272 37058 19281
rect 37002 19207 37058 19216
rect 37016 17746 37044 19207
rect 37004 17740 37056 17746
rect 37004 17682 37056 17688
rect 37108 14498 37136 19638
rect 37556 19654 37608 19660
rect 37462 19615 37518 19624
rect 37278 19272 37334 19281
rect 37476 19258 37504 19615
rect 37568 19446 37596 19654
rect 37556 19440 37608 19446
rect 37556 19382 37608 19388
rect 37476 19230 37596 19258
rect 37278 19207 37334 19216
rect 37292 17746 37320 19207
rect 37462 18592 37518 18601
rect 37462 18527 37518 18536
rect 37476 18358 37504 18527
rect 37464 18352 37516 18358
rect 37464 18294 37516 18300
rect 37462 18048 37518 18057
rect 37462 17983 37518 17992
rect 37280 17740 37332 17746
rect 37280 17682 37332 17688
rect 37372 17740 37424 17746
rect 37372 17682 37424 17688
rect 37384 17610 37412 17682
rect 37372 17604 37424 17610
rect 37372 17546 37424 17552
rect 37370 16688 37426 16697
rect 37280 16652 37332 16658
rect 37370 16623 37426 16632
rect 37280 16594 37332 16600
rect 37292 16561 37320 16594
rect 37278 16552 37334 16561
rect 37278 16487 37334 16496
rect 37280 15428 37332 15434
rect 37016 14470 37136 14498
rect 37200 15388 37280 15416
rect 36912 14068 36964 14074
rect 36912 14010 36964 14016
rect 36820 13864 36872 13870
rect 36820 13806 36872 13812
rect 36728 13796 36780 13802
rect 36728 13738 36780 13744
rect 37016 13716 37044 14470
rect 37096 14408 37148 14414
rect 37096 14350 37148 14356
rect 37108 13938 37136 14350
rect 37096 13932 37148 13938
rect 37096 13874 37148 13880
rect 36832 13688 37044 13716
rect 36726 13424 36782 13433
rect 36726 13359 36782 13368
rect 36740 12918 36768 13359
rect 36728 12912 36780 12918
rect 36728 12854 36780 12860
rect 36728 12776 36780 12782
rect 36726 12744 36728 12753
rect 36780 12744 36782 12753
rect 36726 12679 36782 12688
rect 36726 12472 36782 12481
rect 36832 12458 36860 13688
rect 37108 13326 37136 13874
rect 37096 13320 37148 13326
rect 37096 13262 37148 13268
rect 36912 12980 36964 12986
rect 36912 12922 36964 12928
rect 36924 12481 36952 12922
rect 37004 12844 37056 12850
rect 37004 12786 37056 12792
rect 36782 12442 36860 12458
rect 36910 12472 36966 12481
rect 36782 12436 36872 12442
rect 36782 12430 36820 12436
rect 36726 12407 36782 12416
rect 36910 12407 36966 12416
rect 36820 12378 36872 12384
rect 36832 12345 36860 12378
rect 37016 12374 37044 12786
rect 37096 12640 37148 12646
rect 37096 12582 37148 12588
rect 37108 12442 37136 12582
rect 37096 12436 37148 12442
rect 37096 12378 37148 12384
rect 37004 12368 37056 12374
rect 36818 12336 36874 12345
rect 37004 12310 37056 12316
rect 36818 12271 36874 12280
rect 36636 12096 36688 12102
rect 36636 12038 36688 12044
rect 36544 10192 36596 10198
rect 36544 10134 36596 10140
rect 36360 8900 36412 8906
rect 36360 8842 36412 8848
rect 36174 8800 36230 8809
rect 36174 8735 36230 8744
rect 36084 8560 36136 8566
rect 36084 8502 36136 8508
rect 35898 7576 35954 7585
rect 36096 7546 36124 8502
rect 36360 7744 36412 7750
rect 36360 7686 36412 7692
rect 35898 7511 35954 7520
rect 36084 7540 36136 7546
rect 36084 7482 36136 7488
rect 35900 7268 35952 7274
rect 35900 7210 35952 7216
rect 35912 6662 35940 7210
rect 35900 6656 35952 6662
rect 35348 6598 35400 6604
rect 35438 6624 35494 6633
rect 34244 6384 34296 6390
rect 34244 6326 34296 6332
rect 35360 6322 35388 6598
rect 35900 6598 35952 6604
rect 35438 6559 35494 6568
rect 35348 6316 35400 6322
rect 35348 6258 35400 6264
rect 35912 5846 35940 6598
rect 36096 6458 36124 7482
rect 36084 6452 36136 6458
rect 36084 6394 36136 6400
rect 36372 5914 36400 7686
rect 36648 6254 36676 12038
rect 36820 11824 36872 11830
rect 37200 11778 37228 15388
rect 37280 15370 37332 15376
rect 37384 15162 37412 16623
rect 37476 16425 37504 17983
rect 37568 17270 37596 19230
rect 37648 18352 37700 18358
rect 37752 18340 37780 25910
rect 37844 23118 37872 28047
rect 38108 25152 38160 25158
rect 38108 25094 38160 25100
rect 38120 24993 38148 25094
rect 38106 24984 38162 24993
rect 38106 24919 38162 24928
rect 38108 24132 38160 24138
rect 38108 24074 38160 24080
rect 38120 23730 38148 24074
rect 38108 23724 38160 23730
rect 38108 23666 38160 23672
rect 38016 23520 38068 23526
rect 38016 23462 38068 23468
rect 37832 23112 37884 23118
rect 37832 23054 37884 23060
rect 37924 22432 37976 22438
rect 37924 22374 37976 22380
rect 37936 22030 37964 22374
rect 37924 22024 37976 22030
rect 37924 21966 37976 21972
rect 37832 21956 37884 21962
rect 37832 21898 37884 21904
rect 37700 18312 37780 18340
rect 37648 18294 37700 18300
rect 37844 17338 37872 21898
rect 38028 21078 38056 23462
rect 38212 22642 38240 28086
rect 38384 26240 38436 26246
rect 38384 26182 38436 26188
rect 38396 26042 38424 26182
rect 38384 26036 38436 26042
rect 38384 25978 38436 25984
rect 38292 25696 38344 25702
rect 38292 25638 38344 25644
rect 38304 25430 38332 25638
rect 38292 25424 38344 25430
rect 38292 25366 38344 25372
rect 38304 24206 38332 25366
rect 38752 25152 38804 25158
rect 38752 25094 38804 25100
rect 38660 24880 38712 24886
rect 38660 24822 38712 24828
rect 38568 24608 38620 24614
rect 38568 24550 38620 24556
rect 38384 24404 38436 24410
rect 38384 24346 38436 24352
rect 38292 24200 38344 24206
rect 38292 24142 38344 24148
rect 38200 22636 38252 22642
rect 38200 22578 38252 22584
rect 38108 22568 38160 22574
rect 38108 22510 38160 22516
rect 38120 22098 38148 22510
rect 38200 22500 38252 22506
rect 38200 22442 38252 22448
rect 38108 22092 38160 22098
rect 38108 22034 38160 22040
rect 38106 21584 38162 21593
rect 38106 21519 38162 21528
rect 38016 21072 38068 21078
rect 38016 21014 38068 21020
rect 37924 20460 37976 20466
rect 37924 20402 37976 20408
rect 37936 20369 37964 20402
rect 37922 20360 37978 20369
rect 37922 20295 37978 20304
rect 37924 20052 37976 20058
rect 37924 19994 37976 20000
rect 37832 17332 37884 17338
rect 37832 17274 37884 17280
rect 37556 17264 37608 17270
rect 37556 17206 37608 17212
rect 37648 17264 37700 17270
rect 37936 17218 37964 19994
rect 38120 18601 38148 21519
rect 38212 20534 38240 22442
rect 38200 20528 38252 20534
rect 38200 20470 38252 20476
rect 38304 19514 38332 24142
rect 38396 24070 38424 24346
rect 38580 24313 38608 24550
rect 38566 24304 38622 24313
rect 38566 24239 38622 24248
rect 38384 24064 38436 24070
rect 38384 24006 38436 24012
rect 38384 23044 38436 23050
rect 38384 22986 38436 22992
rect 38396 20942 38424 22986
rect 38474 22944 38530 22953
rect 38474 22879 38530 22888
rect 38488 22098 38516 22879
rect 38580 22642 38608 24239
rect 38672 22953 38700 24822
rect 38764 24138 38792 25094
rect 39132 24274 39160 29815
rect 40774 29322 40830 30000
rect 46294 29322 46350 30000
rect 51722 29322 51778 30000
rect 40774 29294 40908 29322
rect 40774 29200 40830 29294
rect 39856 27668 39908 27674
rect 39856 27610 39908 27616
rect 39478 27228 39786 27248
rect 39478 27226 39484 27228
rect 39540 27226 39564 27228
rect 39620 27226 39644 27228
rect 39700 27226 39724 27228
rect 39780 27226 39786 27228
rect 39540 27174 39542 27226
rect 39722 27174 39724 27226
rect 39478 27172 39484 27174
rect 39540 27172 39564 27174
rect 39620 27172 39644 27174
rect 39700 27172 39724 27174
rect 39780 27172 39786 27174
rect 39478 27152 39786 27172
rect 39478 26140 39786 26160
rect 39478 26138 39484 26140
rect 39540 26138 39564 26140
rect 39620 26138 39644 26140
rect 39700 26138 39724 26140
rect 39780 26138 39786 26140
rect 39540 26086 39542 26138
rect 39722 26086 39724 26138
rect 39478 26084 39484 26086
rect 39540 26084 39564 26086
rect 39620 26084 39644 26086
rect 39700 26084 39724 26086
rect 39780 26084 39786 26086
rect 39478 26064 39786 26084
rect 39212 25832 39264 25838
rect 39212 25774 39264 25780
rect 39120 24268 39172 24274
rect 39120 24210 39172 24216
rect 38752 24132 38804 24138
rect 38752 24074 38804 24080
rect 38844 24064 38896 24070
rect 38844 24006 38896 24012
rect 38856 23769 38884 24006
rect 38842 23760 38898 23769
rect 38842 23695 38898 23704
rect 38936 23588 38988 23594
rect 38936 23530 38988 23536
rect 38750 23216 38806 23225
rect 38750 23151 38752 23160
rect 38804 23151 38806 23160
rect 38752 23122 38804 23128
rect 38658 22944 38714 22953
rect 38658 22879 38714 22888
rect 38764 22794 38792 23122
rect 38844 22976 38896 22982
rect 38844 22918 38896 22924
rect 38672 22766 38792 22794
rect 38568 22636 38620 22642
rect 38568 22578 38620 22584
rect 38568 22160 38620 22166
rect 38568 22102 38620 22108
rect 38476 22092 38528 22098
rect 38476 22034 38528 22040
rect 38580 21049 38608 22102
rect 38566 21040 38622 21049
rect 38566 20975 38622 20984
rect 38384 20936 38436 20942
rect 38384 20878 38436 20884
rect 38672 20058 38700 22766
rect 38752 22432 38804 22438
rect 38752 22374 38804 22380
rect 38764 20942 38792 22374
rect 38856 22137 38884 22918
rect 38842 22128 38898 22137
rect 38842 22063 38898 22072
rect 38856 21554 38884 22063
rect 38844 21548 38896 21554
rect 38844 21490 38896 21496
rect 38844 21412 38896 21418
rect 38844 21354 38896 21360
rect 38752 20936 38804 20942
rect 38752 20878 38804 20884
rect 38752 20800 38804 20806
rect 38752 20742 38804 20748
rect 38660 20052 38712 20058
rect 38660 19994 38712 20000
rect 38764 19854 38792 20742
rect 38856 20330 38884 21354
rect 38948 20398 38976 23530
rect 39028 23520 39080 23526
rect 39028 23462 39080 23468
rect 39040 22817 39068 23462
rect 39026 22808 39082 22817
rect 39026 22743 39082 22752
rect 38936 20392 38988 20398
rect 38936 20334 38988 20340
rect 38844 20324 38896 20330
rect 38844 20266 38896 20272
rect 38752 19848 38804 19854
rect 38752 19790 38804 19796
rect 38936 19848 38988 19854
rect 38936 19790 38988 19796
rect 38844 19780 38896 19786
rect 38844 19722 38896 19728
rect 38292 19508 38344 19514
rect 38292 19450 38344 19456
rect 38750 19408 38806 19417
rect 38750 19343 38806 19352
rect 38658 19272 38714 19281
rect 38658 19207 38714 19216
rect 38568 18828 38620 18834
rect 38568 18770 38620 18776
rect 38476 18760 38528 18766
rect 38476 18702 38528 18708
rect 38200 18692 38252 18698
rect 38200 18634 38252 18640
rect 38106 18592 38162 18601
rect 38106 18527 38162 18536
rect 38212 17377 38240 18634
rect 38488 18465 38516 18702
rect 38474 18456 38530 18465
rect 38474 18391 38530 18400
rect 38580 18154 38608 18770
rect 38672 18290 38700 19207
rect 38764 18902 38792 19343
rect 38752 18896 38804 18902
rect 38752 18838 38804 18844
rect 38856 18578 38884 19722
rect 38764 18550 38884 18578
rect 38660 18284 38712 18290
rect 38660 18226 38712 18232
rect 38568 18148 38620 18154
rect 38568 18090 38620 18096
rect 38198 17368 38254 17377
rect 38198 17303 38254 17312
rect 37648 17206 37700 17212
rect 37556 17128 37608 17134
rect 37556 17070 37608 17076
rect 37462 16416 37518 16425
rect 37462 16351 37518 16360
rect 37464 16176 37516 16182
rect 37462 16144 37464 16153
rect 37516 16144 37518 16153
rect 37462 16079 37518 16088
rect 37372 15156 37424 15162
rect 37372 15098 37424 15104
rect 37372 14340 37424 14346
rect 37372 14282 37424 14288
rect 37384 13326 37412 14282
rect 37372 13320 37424 13326
rect 37278 13288 37334 13297
rect 37372 13262 37424 13268
rect 37278 13223 37334 13232
rect 37292 12986 37320 13223
rect 37280 12980 37332 12986
rect 37280 12922 37332 12928
rect 37384 12889 37412 13262
rect 37370 12880 37426 12889
rect 37370 12815 37426 12824
rect 37464 12776 37516 12782
rect 37464 12718 37516 12724
rect 37280 12708 37332 12714
rect 37280 12650 37332 12656
rect 37292 12209 37320 12650
rect 37278 12200 37334 12209
rect 37278 12135 37334 12144
rect 36820 11766 36872 11772
rect 36728 11756 36780 11762
rect 36728 11698 36780 11704
rect 36740 11354 36768 11698
rect 36728 11348 36780 11354
rect 36728 11290 36780 11296
rect 36832 11257 36860 11766
rect 37108 11750 37228 11778
rect 37372 11824 37424 11830
rect 37372 11766 37424 11772
rect 36912 11620 36964 11626
rect 36912 11562 36964 11568
rect 36818 11248 36874 11257
rect 36818 11183 36874 11192
rect 36832 9110 36860 11183
rect 36924 11082 36952 11562
rect 37004 11280 37056 11286
rect 37004 11222 37056 11228
rect 36912 11076 36964 11082
rect 36912 11018 36964 11024
rect 37016 10742 37044 11222
rect 37004 10736 37056 10742
rect 37004 10678 37056 10684
rect 37004 9580 37056 9586
rect 37004 9522 37056 9528
rect 36912 9444 36964 9450
rect 36912 9386 36964 9392
rect 36820 9104 36872 9110
rect 36820 9046 36872 9052
rect 36924 7750 36952 9386
rect 37016 9382 37044 9522
rect 37004 9376 37056 9382
rect 37004 9318 37056 9324
rect 37016 8809 37044 9318
rect 37002 8800 37058 8809
rect 37002 8735 37058 8744
rect 37108 8265 37136 11750
rect 37384 10742 37412 11766
rect 37280 10736 37332 10742
rect 37280 10678 37332 10684
rect 37372 10736 37424 10742
rect 37372 10678 37424 10684
rect 37292 10470 37320 10678
rect 37280 10464 37332 10470
rect 37280 10406 37332 10412
rect 37188 9920 37240 9926
rect 37188 9862 37240 9868
rect 37200 9654 37228 9862
rect 37188 9648 37240 9654
rect 37188 9590 37240 9596
rect 37200 8294 37228 9590
rect 37292 8634 37320 10406
rect 37476 8974 37504 12718
rect 37568 12374 37596 17070
rect 37660 16794 37688 17206
rect 37844 17190 37964 17218
rect 38106 17232 38162 17241
rect 37648 16788 37700 16794
rect 37648 16730 37700 16736
rect 37648 16652 37700 16658
rect 37648 16594 37700 16600
rect 37660 15609 37688 16594
rect 37646 15600 37702 15609
rect 37646 15535 37702 15544
rect 37648 15020 37700 15026
rect 37648 14962 37700 14968
rect 37660 14414 37688 14962
rect 37648 14408 37700 14414
rect 37648 14350 37700 14356
rect 37648 13728 37700 13734
rect 37648 13670 37700 13676
rect 37660 13258 37688 13670
rect 37648 13252 37700 13258
rect 37648 13194 37700 13200
rect 37660 12434 37688 13194
rect 37844 12753 37872 17190
rect 38106 17167 38162 17176
rect 38120 17066 38148 17167
rect 38108 17060 38160 17066
rect 38108 17002 38160 17008
rect 38292 16992 38344 16998
rect 38290 16960 38292 16969
rect 38660 16992 38712 16998
rect 38344 16960 38346 16969
rect 38660 16934 38712 16940
rect 38290 16895 38346 16904
rect 38014 16824 38070 16833
rect 38014 16759 38070 16768
rect 37924 14816 37976 14822
rect 37924 14758 37976 14764
rect 37936 14550 37964 14758
rect 37924 14544 37976 14550
rect 37924 14486 37976 14492
rect 37924 14340 37976 14346
rect 37924 14282 37976 14288
rect 37936 13938 37964 14282
rect 37924 13932 37976 13938
rect 37924 13874 37976 13880
rect 38028 13462 38056 16759
rect 38672 16250 38700 16934
rect 38764 16289 38792 18550
rect 38844 18420 38896 18426
rect 38844 18362 38896 18368
rect 38856 16794 38884 18362
rect 38948 17814 38976 19790
rect 39040 18426 39068 22743
rect 39132 22030 39160 24210
rect 39120 22024 39172 22030
rect 39120 21966 39172 21972
rect 39120 21480 39172 21486
rect 39120 21422 39172 21428
rect 39132 21146 39160 21422
rect 39120 21140 39172 21146
rect 39120 21082 39172 21088
rect 39120 20800 39172 20806
rect 39118 20768 39120 20777
rect 39172 20768 39174 20777
rect 39118 20703 39174 20712
rect 39120 20596 39172 20602
rect 39120 20538 39172 20544
rect 39132 18766 39160 20538
rect 39224 20398 39252 25774
rect 39478 25052 39786 25072
rect 39478 25050 39484 25052
rect 39540 25050 39564 25052
rect 39620 25050 39644 25052
rect 39700 25050 39724 25052
rect 39780 25050 39786 25052
rect 39540 24998 39542 25050
rect 39722 24998 39724 25050
rect 39478 24996 39484 24998
rect 39540 24996 39564 24998
rect 39620 24996 39644 24998
rect 39700 24996 39724 24998
rect 39780 24996 39786 24998
rect 39478 24976 39786 24996
rect 39488 24608 39540 24614
rect 39486 24576 39488 24585
rect 39540 24576 39542 24585
rect 39486 24511 39542 24520
rect 39304 24404 39356 24410
rect 39304 24346 39356 24352
rect 39316 22166 39344 24346
rect 39478 23964 39786 23984
rect 39478 23962 39484 23964
rect 39540 23962 39564 23964
rect 39620 23962 39644 23964
rect 39700 23962 39724 23964
rect 39780 23962 39786 23964
rect 39540 23910 39542 23962
rect 39722 23910 39724 23962
rect 39478 23908 39484 23910
rect 39540 23908 39564 23910
rect 39620 23908 39644 23910
rect 39700 23908 39724 23910
rect 39780 23908 39786 23910
rect 39478 23888 39786 23908
rect 39396 23520 39448 23526
rect 39396 23462 39448 23468
rect 39408 23225 39436 23462
rect 39394 23216 39450 23225
rect 39394 23151 39450 23160
rect 39408 22778 39436 23151
rect 39478 22876 39786 22896
rect 39478 22874 39484 22876
rect 39540 22874 39564 22876
rect 39620 22874 39644 22876
rect 39700 22874 39724 22876
rect 39780 22874 39786 22876
rect 39540 22822 39542 22874
rect 39722 22822 39724 22874
rect 39478 22820 39484 22822
rect 39540 22820 39564 22822
rect 39620 22820 39644 22822
rect 39700 22820 39724 22822
rect 39780 22820 39786 22822
rect 39478 22800 39786 22820
rect 39396 22772 39448 22778
rect 39868 22760 39896 27610
rect 40880 27470 40908 29294
rect 46294 29294 46428 29322
rect 41510 29200 41566 29209
rect 46294 29200 46350 29294
rect 41510 29135 41566 29144
rect 41420 28144 41472 28150
rect 41420 28086 41472 28092
rect 40868 27464 40920 27470
rect 40868 27406 40920 27412
rect 41052 27328 41104 27334
rect 41052 27270 41104 27276
rect 40960 26308 41012 26314
rect 40960 26250 41012 26256
rect 40592 26036 40644 26042
rect 40592 25978 40644 25984
rect 40604 24818 40632 25978
rect 40866 25256 40922 25265
rect 40866 25191 40922 25200
rect 40592 24812 40644 24818
rect 40592 24754 40644 24760
rect 40604 24410 40632 24754
rect 40592 24404 40644 24410
rect 40592 24346 40644 24352
rect 40604 23866 40632 24346
rect 40776 24200 40828 24206
rect 40776 24142 40828 24148
rect 40224 23860 40276 23866
rect 40224 23802 40276 23808
rect 40592 23860 40644 23866
rect 40592 23802 40644 23808
rect 39396 22714 39448 22720
rect 39776 22732 39896 22760
rect 39578 22536 39634 22545
rect 39578 22471 39580 22480
rect 39632 22471 39634 22480
rect 39580 22442 39632 22448
rect 39304 22160 39356 22166
rect 39304 22102 39356 22108
rect 39776 22094 39804 22732
rect 39856 22432 39908 22438
rect 39856 22374 39908 22380
rect 39868 22166 39896 22374
rect 40236 22166 40264 23802
rect 40500 23724 40552 23730
rect 40500 23666 40552 23672
rect 40512 23361 40540 23666
rect 40498 23352 40554 23361
rect 40604 23322 40632 23802
rect 40788 23730 40816 24142
rect 40776 23724 40828 23730
rect 40776 23666 40828 23672
rect 40684 23656 40736 23662
rect 40684 23598 40736 23604
rect 40774 23624 40830 23633
rect 40498 23287 40554 23296
rect 40592 23316 40644 23322
rect 40408 22976 40460 22982
rect 40408 22918 40460 22924
rect 40420 22681 40448 22918
rect 40406 22672 40462 22681
rect 40406 22607 40462 22616
rect 39856 22160 39908 22166
rect 40040 22160 40092 22166
rect 39856 22102 39908 22108
rect 40038 22128 40040 22137
rect 40224 22160 40276 22166
rect 40092 22128 40094 22137
rect 39408 22066 39804 22094
rect 40224 22102 40276 22108
rect 39304 21888 39356 21894
rect 39304 21830 39356 21836
rect 39316 21049 39344 21830
rect 39302 21040 39358 21049
rect 39302 20975 39358 20984
rect 39212 20392 39264 20398
rect 39212 20334 39264 20340
rect 39304 20256 39356 20262
rect 39304 20198 39356 20204
rect 39212 19984 39264 19990
rect 39210 19952 39212 19961
rect 39264 19952 39266 19961
rect 39210 19887 39266 19896
rect 39224 18834 39252 19887
rect 39316 19514 39344 20198
rect 39408 20058 39436 22066
rect 40038 22063 40094 22072
rect 40132 22024 40184 22030
rect 39854 21992 39910 22001
rect 40132 21966 40184 21972
rect 39854 21927 39910 21936
rect 39478 21788 39786 21808
rect 39478 21786 39484 21788
rect 39540 21786 39564 21788
rect 39620 21786 39644 21788
rect 39700 21786 39724 21788
rect 39780 21786 39786 21788
rect 39540 21734 39542 21786
rect 39722 21734 39724 21786
rect 39478 21732 39484 21734
rect 39540 21732 39564 21734
rect 39620 21732 39644 21734
rect 39700 21732 39724 21734
rect 39780 21732 39786 21734
rect 39478 21712 39786 21732
rect 39868 21690 39896 21927
rect 39856 21684 39908 21690
rect 39856 21626 39908 21632
rect 40040 21684 40092 21690
rect 40040 21626 40092 21632
rect 40052 21570 40080 21626
rect 39868 21542 40080 21570
rect 39868 21418 39896 21542
rect 40040 21480 40092 21486
rect 40040 21422 40092 21428
rect 39856 21412 39908 21418
rect 39856 21354 39908 21360
rect 39948 21412 40000 21418
rect 39948 21354 40000 21360
rect 39488 21344 39540 21350
rect 39488 21286 39540 21292
rect 39500 20942 39528 21286
rect 39960 21146 39988 21354
rect 39948 21140 40000 21146
rect 39868 21100 39948 21128
rect 39488 20936 39540 20942
rect 39488 20878 39540 20884
rect 39478 20700 39786 20720
rect 39478 20698 39484 20700
rect 39540 20698 39564 20700
rect 39620 20698 39644 20700
rect 39700 20698 39724 20700
rect 39780 20698 39786 20700
rect 39540 20646 39542 20698
rect 39722 20646 39724 20698
rect 39478 20644 39484 20646
rect 39540 20644 39564 20646
rect 39620 20644 39644 20646
rect 39700 20644 39724 20646
rect 39780 20644 39786 20646
rect 39478 20624 39786 20644
rect 39762 20088 39818 20097
rect 39396 20052 39448 20058
rect 39762 20023 39818 20032
rect 39396 19994 39448 20000
rect 39776 19854 39804 20023
rect 39764 19848 39816 19854
rect 39764 19790 39816 19796
rect 39478 19612 39786 19632
rect 39478 19610 39484 19612
rect 39540 19610 39564 19612
rect 39620 19610 39644 19612
rect 39700 19610 39724 19612
rect 39780 19610 39786 19612
rect 39540 19558 39542 19610
rect 39722 19558 39724 19610
rect 39478 19556 39484 19558
rect 39540 19556 39564 19558
rect 39620 19556 39644 19558
rect 39700 19556 39724 19558
rect 39780 19556 39786 19558
rect 39478 19536 39786 19556
rect 39304 19508 39356 19514
rect 39304 19450 39356 19456
rect 39316 19378 39344 19450
rect 39304 19372 39356 19378
rect 39304 19314 39356 19320
rect 39488 19304 39540 19310
rect 39488 19246 39540 19252
rect 39580 19304 39632 19310
rect 39580 19246 39632 19252
rect 39396 19168 39448 19174
rect 39396 19110 39448 19116
rect 39212 18828 39264 18834
rect 39212 18770 39264 18776
rect 39120 18760 39172 18766
rect 39120 18702 39172 18708
rect 39212 18624 39264 18630
rect 39212 18566 39264 18572
rect 39028 18420 39080 18426
rect 39028 18362 39080 18368
rect 39224 18358 39252 18566
rect 39304 18420 39356 18426
rect 39304 18362 39356 18368
rect 39212 18352 39264 18358
rect 39316 18329 39344 18362
rect 39212 18294 39264 18300
rect 39302 18320 39358 18329
rect 39302 18255 39358 18264
rect 39302 18184 39358 18193
rect 39408 18170 39436 19110
rect 39500 18873 39528 19246
rect 39592 18902 39620 19246
rect 39580 18896 39632 18902
rect 39486 18864 39542 18873
rect 39580 18838 39632 18844
rect 39486 18799 39542 18808
rect 39478 18524 39786 18544
rect 39478 18522 39484 18524
rect 39540 18522 39564 18524
rect 39620 18522 39644 18524
rect 39700 18522 39724 18524
rect 39780 18522 39786 18524
rect 39540 18470 39542 18522
rect 39722 18470 39724 18522
rect 39478 18468 39484 18470
rect 39540 18468 39564 18470
rect 39620 18468 39644 18470
rect 39700 18468 39724 18470
rect 39780 18468 39786 18470
rect 39478 18448 39786 18468
rect 39868 18408 39896 21100
rect 39948 21082 40000 21088
rect 39948 20868 40000 20874
rect 39948 20810 40000 20816
rect 39960 20534 39988 20810
rect 39948 20528 40000 20534
rect 39948 20470 40000 20476
rect 39948 20324 40000 20330
rect 39948 20266 40000 20272
rect 39960 19718 39988 20266
rect 40052 19990 40080 21422
rect 40144 20262 40172 21966
rect 40236 21622 40264 22102
rect 40408 21888 40460 21894
rect 40408 21830 40460 21836
rect 40224 21616 40276 21622
rect 40224 21558 40276 21564
rect 40316 21548 40368 21554
rect 40316 21490 40368 21496
rect 40328 21078 40356 21490
rect 40316 21072 40368 21078
rect 40316 21014 40368 21020
rect 40328 20466 40356 21014
rect 40420 20505 40448 21830
rect 40512 21486 40540 23287
rect 40592 23258 40644 23264
rect 40592 21548 40644 21554
rect 40592 21490 40644 21496
rect 40500 21480 40552 21486
rect 40604 21457 40632 21490
rect 40500 21422 40552 21428
rect 40590 21448 40646 21457
rect 40590 21383 40646 21392
rect 40500 21344 40552 21350
rect 40500 21286 40552 21292
rect 40512 21185 40540 21286
rect 40498 21176 40554 21185
rect 40498 21111 40554 21120
rect 40592 21140 40644 21146
rect 40592 21082 40644 21088
rect 40406 20496 40462 20505
rect 40316 20460 40368 20466
rect 40406 20431 40462 20440
rect 40316 20402 40368 20408
rect 40224 20392 40276 20398
rect 40224 20334 40276 20340
rect 40132 20256 40184 20262
rect 40132 20198 40184 20204
rect 40040 19984 40092 19990
rect 40040 19926 40092 19932
rect 40040 19848 40092 19854
rect 40040 19790 40092 19796
rect 40130 19816 40186 19825
rect 39948 19712 40000 19718
rect 40052 19689 40080 19790
rect 40130 19751 40186 19760
rect 39948 19654 40000 19660
rect 40038 19680 40094 19689
rect 40038 19615 40094 19624
rect 40052 19530 40080 19615
rect 39776 18380 39896 18408
rect 39960 19502 40080 19530
rect 39408 18142 39528 18170
rect 39302 18119 39358 18128
rect 39316 17814 39344 18119
rect 39500 18086 39528 18142
rect 39396 18080 39448 18086
rect 39396 18022 39448 18028
rect 39488 18080 39540 18086
rect 39488 18022 39540 18028
rect 38936 17808 38988 17814
rect 38936 17750 38988 17756
rect 39304 17808 39356 17814
rect 39304 17750 39356 17756
rect 38844 16788 38896 16794
rect 38844 16730 38896 16736
rect 38948 16726 38976 17750
rect 39028 17536 39080 17542
rect 39028 17478 39080 17484
rect 39040 17134 39068 17478
rect 39028 17128 39080 17134
rect 39304 17128 39356 17134
rect 39028 17070 39080 17076
rect 39118 17096 39174 17105
rect 39304 17070 39356 17076
rect 39118 17031 39174 17040
rect 38936 16720 38988 16726
rect 38936 16662 38988 16668
rect 38750 16280 38806 16289
rect 38660 16244 38712 16250
rect 38750 16215 38806 16224
rect 38660 16186 38712 16192
rect 38752 16040 38804 16046
rect 38752 15982 38804 15988
rect 38384 15564 38436 15570
rect 38384 15506 38436 15512
rect 38200 15156 38252 15162
rect 38200 15098 38252 15104
rect 38212 15026 38240 15098
rect 38200 15020 38252 15026
rect 38200 14962 38252 14968
rect 38108 14816 38160 14822
rect 38108 14758 38160 14764
rect 38120 14346 38148 14758
rect 38212 14414 38240 14962
rect 38200 14408 38252 14414
rect 38200 14350 38252 14356
rect 38108 14340 38160 14346
rect 38108 14282 38160 14288
rect 38120 13734 38148 14282
rect 38108 13728 38160 13734
rect 38108 13670 38160 13676
rect 38290 13560 38346 13569
rect 38290 13495 38346 13504
rect 38016 13456 38068 13462
rect 38016 13398 38068 13404
rect 38304 13394 38332 13495
rect 38108 13388 38160 13394
rect 38292 13388 38344 13394
rect 38160 13348 38240 13376
rect 38108 13330 38160 13336
rect 37924 13320 37976 13326
rect 37924 13262 37976 13268
rect 37830 12744 37886 12753
rect 37830 12679 37886 12688
rect 37660 12406 37780 12434
rect 37556 12368 37608 12374
rect 37556 12310 37608 12316
rect 37556 12096 37608 12102
rect 37556 12038 37608 12044
rect 37464 8968 37516 8974
rect 37464 8910 37516 8916
rect 37370 8664 37426 8673
rect 37280 8628 37332 8634
rect 37370 8599 37372 8608
rect 37280 8570 37332 8576
rect 37424 8599 37426 8608
rect 37372 8570 37424 8576
rect 37188 8288 37240 8294
rect 37094 8256 37150 8265
rect 37188 8230 37240 8236
rect 37094 8191 37150 8200
rect 36912 7744 36964 7750
rect 36912 7686 36964 7692
rect 36924 7274 36952 7686
rect 37200 7342 37228 8230
rect 37568 7886 37596 12038
rect 37648 11552 37700 11558
rect 37646 11520 37648 11529
rect 37700 11520 37702 11529
rect 37646 11455 37702 11464
rect 37648 11076 37700 11082
rect 37648 11018 37700 11024
rect 37660 10130 37688 11018
rect 37648 10124 37700 10130
rect 37648 10066 37700 10072
rect 37648 9104 37700 9110
rect 37648 9046 37700 9052
rect 37556 7880 37608 7886
rect 37556 7822 37608 7828
rect 37660 7410 37688 9046
rect 37648 7404 37700 7410
rect 37648 7346 37700 7352
rect 37188 7336 37240 7342
rect 37188 7278 37240 7284
rect 36912 7268 36964 7274
rect 36912 7210 36964 7216
rect 36636 6248 36688 6254
rect 36636 6190 36688 6196
rect 36360 5908 36412 5914
rect 36360 5850 36412 5856
rect 32864 5840 32916 5846
rect 32864 5782 32916 5788
rect 33508 5840 33560 5846
rect 33508 5782 33560 5788
rect 35900 5840 35952 5846
rect 35900 5782 35952 5788
rect 32772 5772 32824 5778
rect 32772 5714 32824 5720
rect 37200 5642 37228 7278
rect 37188 5636 37240 5642
rect 37188 5578 37240 5584
rect 37752 5522 37780 12406
rect 37844 11354 37872 12679
rect 37832 11348 37884 11354
rect 37832 11290 37884 11296
rect 37832 11144 37884 11150
rect 37832 11086 37884 11092
rect 37844 10985 37872 11086
rect 37830 10976 37886 10985
rect 37830 10911 37886 10920
rect 37936 10470 37964 13262
rect 38016 12844 38068 12850
rect 38016 12786 38068 12792
rect 38028 12753 38056 12786
rect 38014 12744 38070 12753
rect 38014 12679 38070 12688
rect 38028 12306 38056 12679
rect 38016 12300 38068 12306
rect 38016 12242 38068 12248
rect 38108 12232 38160 12238
rect 38108 12174 38160 12180
rect 38016 12164 38068 12170
rect 38016 12106 38068 12112
rect 38028 11898 38056 12106
rect 38016 11892 38068 11898
rect 38016 11834 38068 11840
rect 38016 11688 38068 11694
rect 38016 11630 38068 11636
rect 37924 10464 37976 10470
rect 37924 10406 37976 10412
rect 37832 10056 37884 10062
rect 37830 10024 37832 10033
rect 37884 10024 37886 10033
rect 37830 9959 37886 9968
rect 38028 9382 38056 11630
rect 38120 11529 38148 12174
rect 38212 11762 38240 13348
rect 38292 13330 38344 13336
rect 38200 11756 38252 11762
rect 38200 11698 38252 11704
rect 38106 11520 38162 11529
rect 38106 11455 38162 11464
rect 38016 9376 38068 9382
rect 38016 9318 38068 9324
rect 37832 8900 37884 8906
rect 37832 8842 37884 8848
rect 37844 8294 37872 8842
rect 37832 8288 37884 8294
rect 37832 8230 37884 8236
rect 37844 7818 37872 8230
rect 37832 7812 37884 7818
rect 37832 7754 37884 7760
rect 37752 5494 37872 5522
rect 32220 5296 32272 5302
rect 32220 5238 32272 5244
rect 37278 5128 37334 5137
rect 37278 5063 37280 5072
rect 37332 5063 37334 5072
rect 37280 5034 37332 5040
rect 37844 3534 37872 5494
rect 37832 3528 37884 3534
rect 37832 3470 37884 3476
rect 37738 3360 37794 3369
rect 37738 3295 37794 3304
rect 37752 3058 37780 3295
rect 37740 3052 37792 3058
rect 37740 2994 37792 3000
rect 37752 2446 37780 2994
rect 37740 2440 37792 2446
rect 37740 2382 37792 2388
rect 37844 2378 37872 3470
rect 37924 2916 37976 2922
rect 37924 2858 37976 2864
rect 37936 2378 37964 2858
rect 37832 2372 37884 2378
rect 37832 2314 37884 2320
rect 37924 2372 37976 2378
rect 37924 2314 37976 2320
rect 31208 2304 31260 2310
rect 31208 2246 31260 2252
rect 38028 1737 38056 9318
rect 38120 8362 38148 11455
rect 38304 10266 38332 13330
rect 38396 13326 38424 15506
rect 38764 15473 38792 15982
rect 38948 15502 38976 16662
rect 39026 16280 39082 16289
rect 39026 16215 39082 16224
rect 39040 16114 39068 16215
rect 39028 16108 39080 16114
rect 39028 16050 39080 16056
rect 39028 15904 39080 15910
rect 39028 15846 39080 15852
rect 38936 15496 38988 15502
rect 38750 15464 38806 15473
rect 38936 15438 38988 15444
rect 38750 15399 38806 15408
rect 38844 15428 38896 15434
rect 38844 15370 38896 15376
rect 38856 14822 38884 15370
rect 38844 14816 38896 14822
rect 38844 14758 38896 14764
rect 38568 14476 38620 14482
rect 38568 14418 38620 14424
rect 38474 14104 38530 14113
rect 38474 14039 38530 14048
rect 38488 13462 38516 14039
rect 38476 13456 38528 13462
rect 38476 13398 38528 13404
rect 38384 13320 38436 13326
rect 38384 13262 38436 13268
rect 38476 12980 38528 12986
rect 38476 12922 38528 12928
rect 38384 11688 38436 11694
rect 38384 11630 38436 11636
rect 38396 10742 38424 11630
rect 38384 10736 38436 10742
rect 38384 10678 38436 10684
rect 38292 10260 38344 10266
rect 38292 10202 38344 10208
rect 38488 9518 38516 12922
rect 38580 12850 38608 14418
rect 38752 14340 38804 14346
rect 38672 14300 38752 14328
rect 38672 14249 38700 14300
rect 38752 14282 38804 14288
rect 38658 14240 38714 14249
rect 38658 14175 38714 14184
rect 38842 14240 38898 14249
rect 38842 14175 38898 14184
rect 38660 14000 38712 14006
rect 38660 13942 38712 13948
rect 38672 13841 38700 13942
rect 38658 13832 38714 13841
rect 38658 13767 38714 13776
rect 38660 13388 38712 13394
rect 38660 13330 38712 13336
rect 38568 12844 38620 12850
rect 38568 12786 38620 12792
rect 38672 12434 38700 13330
rect 38856 13258 38884 14175
rect 38844 13252 38896 13258
rect 38844 13194 38896 13200
rect 38936 13184 38988 13190
rect 38936 13126 38988 13132
rect 38750 12880 38806 12889
rect 38948 12850 38976 13126
rect 38750 12815 38806 12824
rect 38936 12844 38988 12850
rect 38764 12442 38792 12815
rect 38936 12786 38988 12792
rect 38844 12776 38896 12782
rect 38844 12718 38896 12724
rect 38934 12744 38990 12753
rect 38580 12406 38700 12434
rect 38752 12436 38804 12442
rect 38580 12084 38608 12406
rect 38752 12378 38804 12384
rect 38658 12336 38714 12345
rect 38658 12271 38714 12280
rect 38672 12238 38700 12271
rect 38660 12232 38712 12238
rect 38660 12174 38712 12180
rect 38752 12096 38804 12102
rect 38580 12056 38700 12084
rect 38568 11620 38620 11626
rect 38568 11562 38620 11568
rect 38580 10962 38608 11562
rect 38672 11121 38700 12056
rect 38752 12038 38804 12044
rect 38764 11898 38792 12038
rect 38752 11892 38804 11898
rect 38752 11834 38804 11840
rect 38752 11756 38804 11762
rect 38752 11698 38804 11704
rect 38658 11112 38714 11121
rect 38658 11047 38714 11056
rect 38580 10934 38700 10962
rect 38568 10736 38620 10742
rect 38568 10678 38620 10684
rect 38580 10130 38608 10678
rect 38568 10124 38620 10130
rect 38568 10066 38620 10072
rect 38476 9512 38528 9518
rect 38476 9454 38528 9460
rect 38580 9110 38608 10066
rect 38672 9382 38700 10934
rect 38660 9376 38712 9382
rect 38660 9318 38712 9324
rect 38672 9178 38700 9318
rect 38660 9172 38712 9178
rect 38660 9114 38712 9120
rect 38568 9104 38620 9110
rect 38568 9046 38620 9052
rect 38764 8566 38792 11698
rect 38856 11626 38884 12718
rect 38934 12679 38936 12688
rect 38988 12679 38990 12688
rect 38936 12650 38988 12656
rect 38948 12102 38976 12650
rect 38936 12096 38988 12102
rect 38936 12038 38988 12044
rect 38844 11620 38896 11626
rect 38844 11562 38896 11568
rect 38842 11384 38898 11393
rect 38842 11319 38844 11328
rect 38896 11319 38898 11328
rect 38844 11290 38896 11296
rect 38934 10160 38990 10169
rect 38934 10095 38936 10104
rect 38988 10095 38990 10104
rect 38936 10066 38988 10072
rect 39040 10010 39068 15846
rect 39132 13938 39160 17031
rect 39212 16584 39264 16590
rect 39212 16526 39264 16532
rect 39224 14074 39252 16526
rect 39316 16130 39344 17070
rect 39408 16250 39436 18022
rect 39776 17882 39804 18380
rect 39764 17876 39816 17882
rect 39764 17818 39816 17824
rect 39960 17592 39988 19502
rect 40144 19378 40172 19751
rect 40132 19372 40184 19378
rect 40132 19314 40184 19320
rect 40130 18592 40186 18601
rect 40130 18527 40186 18536
rect 40144 18426 40172 18527
rect 40132 18420 40184 18426
rect 40132 18362 40184 18368
rect 40236 18170 40264 20334
rect 40500 20324 40552 20330
rect 40500 20266 40552 20272
rect 40408 19440 40460 19446
rect 40408 19382 40460 19388
rect 40420 18698 40448 19382
rect 40408 18692 40460 18698
rect 40408 18634 40460 18640
rect 40316 18624 40368 18630
rect 40316 18566 40368 18572
rect 39868 17564 39988 17592
rect 40052 18142 40264 18170
rect 39478 17436 39786 17456
rect 39478 17434 39484 17436
rect 39540 17434 39564 17436
rect 39620 17434 39644 17436
rect 39700 17434 39724 17436
rect 39780 17434 39786 17436
rect 39540 17382 39542 17434
rect 39722 17382 39724 17434
rect 39478 17380 39484 17382
rect 39540 17380 39564 17382
rect 39620 17380 39644 17382
rect 39700 17380 39724 17382
rect 39780 17380 39786 17382
rect 39478 17360 39786 17380
rect 39868 16454 39896 17564
rect 39946 17504 40002 17513
rect 39946 17439 40002 17448
rect 39960 17270 39988 17439
rect 39948 17264 40000 17270
rect 39948 17206 40000 17212
rect 39856 16448 39908 16454
rect 39856 16390 39908 16396
rect 39478 16348 39786 16368
rect 39478 16346 39484 16348
rect 39540 16346 39564 16348
rect 39620 16346 39644 16348
rect 39700 16346 39724 16348
rect 39780 16346 39786 16348
rect 39540 16294 39542 16346
rect 39722 16294 39724 16346
rect 39478 16292 39484 16294
rect 39540 16292 39564 16294
rect 39620 16292 39644 16294
rect 39700 16292 39724 16294
rect 39780 16292 39786 16294
rect 39478 16272 39786 16292
rect 39396 16244 39448 16250
rect 39396 16186 39448 16192
rect 39316 16102 39436 16130
rect 39408 15502 39436 16102
rect 39856 16108 39908 16114
rect 39856 16050 39908 16056
rect 39868 15638 39896 16050
rect 39856 15632 39908 15638
rect 39856 15574 39908 15580
rect 39396 15496 39448 15502
rect 39396 15438 39448 15444
rect 39304 15360 39356 15366
rect 39304 15302 39356 15308
rect 39212 14068 39264 14074
rect 39212 14010 39264 14016
rect 39210 13968 39266 13977
rect 39120 13932 39172 13938
rect 39210 13903 39266 13912
rect 39120 13874 39172 13880
rect 39224 13870 39252 13903
rect 39212 13864 39264 13870
rect 39212 13806 39264 13812
rect 39212 13728 39264 13734
rect 39212 13670 39264 13676
rect 39120 13184 39172 13190
rect 39120 13126 39172 13132
rect 38856 9982 39068 10010
rect 38752 8560 38804 8566
rect 38752 8502 38804 8508
rect 38108 8356 38160 8362
rect 38108 8298 38160 8304
rect 38856 8090 38884 9982
rect 38936 9920 38988 9926
rect 38936 9862 38988 9868
rect 38948 9382 38976 9862
rect 38936 9376 38988 9382
rect 38936 9318 38988 9324
rect 38948 8906 38976 9318
rect 38936 8900 38988 8906
rect 38936 8842 38988 8848
rect 38844 8084 38896 8090
rect 38844 8026 38896 8032
rect 39132 6186 39160 13126
rect 39224 12850 39252 13670
rect 39316 12986 39344 15302
rect 39408 15026 39436 15438
rect 39948 15428 40000 15434
rect 39948 15370 40000 15376
rect 39478 15260 39786 15280
rect 39478 15258 39484 15260
rect 39540 15258 39564 15260
rect 39620 15258 39644 15260
rect 39700 15258 39724 15260
rect 39780 15258 39786 15260
rect 39540 15206 39542 15258
rect 39722 15206 39724 15258
rect 39478 15204 39484 15206
rect 39540 15204 39564 15206
rect 39620 15204 39644 15206
rect 39700 15204 39724 15206
rect 39780 15204 39786 15206
rect 39478 15184 39786 15204
rect 39960 15026 39988 15370
rect 39396 15020 39448 15026
rect 39396 14962 39448 14968
rect 39948 15020 40000 15026
rect 39948 14962 40000 14968
rect 39854 14920 39910 14929
rect 40052 14906 40080 18142
rect 40132 16108 40184 16114
rect 40132 16050 40184 16056
rect 40144 16017 40172 16050
rect 40130 16008 40186 16017
rect 40130 15943 40186 15952
rect 40224 15972 40276 15978
rect 40224 15914 40276 15920
rect 40236 15881 40264 15914
rect 40222 15872 40278 15881
rect 40222 15807 40278 15816
rect 40224 15020 40276 15026
rect 40224 14962 40276 14968
rect 39854 14855 39910 14864
rect 39960 14878 40080 14906
rect 39762 14784 39818 14793
rect 39762 14719 39818 14728
rect 39776 14521 39804 14719
rect 39762 14512 39818 14521
rect 39396 14476 39448 14482
rect 39762 14447 39818 14456
rect 39396 14418 39448 14424
rect 39408 14056 39436 14418
rect 39764 14408 39816 14414
rect 39762 14376 39764 14385
rect 39816 14376 39818 14385
rect 39762 14311 39818 14320
rect 39478 14172 39786 14192
rect 39478 14170 39484 14172
rect 39540 14170 39564 14172
rect 39620 14170 39644 14172
rect 39700 14170 39724 14172
rect 39780 14170 39786 14172
rect 39540 14118 39542 14170
rect 39722 14118 39724 14170
rect 39478 14116 39484 14118
rect 39540 14116 39564 14118
rect 39620 14116 39644 14118
rect 39700 14116 39724 14118
rect 39780 14116 39786 14118
rect 39478 14096 39786 14116
rect 39408 14028 39620 14056
rect 39488 13932 39540 13938
rect 39488 13874 39540 13880
rect 39396 13864 39448 13870
rect 39396 13806 39448 13812
rect 39304 12980 39356 12986
rect 39304 12922 39356 12928
rect 39212 12844 39264 12850
rect 39212 12786 39264 12792
rect 39302 12744 39358 12753
rect 39302 12679 39358 12688
rect 39316 12481 39344 12679
rect 39302 12472 39358 12481
rect 39302 12407 39358 12416
rect 39316 11898 39344 12407
rect 39304 11892 39356 11898
rect 39304 11834 39356 11840
rect 39408 11218 39436 13806
rect 39500 13258 39528 13874
rect 39592 13734 39620 14028
rect 39580 13728 39632 13734
rect 39580 13670 39632 13676
rect 39488 13252 39540 13258
rect 39488 13194 39540 13200
rect 39478 13084 39786 13104
rect 39478 13082 39484 13084
rect 39540 13082 39564 13084
rect 39620 13082 39644 13084
rect 39700 13082 39724 13084
rect 39780 13082 39786 13084
rect 39540 13030 39542 13082
rect 39722 13030 39724 13082
rect 39478 13028 39484 13030
rect 39540 13028 39564 13030
rect 39620 13028 39644 13030
rect 39700 13028 39724 13030
rect 39780 13028 39786 13030
rect 39478 13008 39786 13028
rect 39868 12986 39896 14855
rect 39856 12980 39908 12986
rect 39856 12922 39908 12928
rect 39488 12708 39540 12714
rect 39488 12650 39540 12656
rect 39500 12481 39528 12650
rect 39486 12472 39542 12481
rect 39486 12407 39542 12416
rect 39960 12374 39988 14878
rect 40040 14816 40092 14822
rect 40040 14758 40092 14764
rect 40052 13705 40080 14758
rect 40236 14618 40264 14962
rect 40224 14612 40276 14618
rect 40224 14554 40276 14560
rect 40132 14544 40184 14550
rect 40132 14486 40184 14492
rect 40144 14249 40172 14486
rect 40130 14240 40186 14249
rect 40130 14175 40186 14184
rect 40130 14104 40186 14113
rect 40130 14039 40132 14048
rect 40184 14039 40186 14048
rect 40132 14010 40184 14016
rect 40130 13968 40186 13977
rect 40130 13903 40132 13912
rect 40184 13903 40186 13912
rect 40132 13874 40184 13880
rect 40236 13802 40264 14554
rect 40224 13796 40276 13802
rect 40224 13738 40276 13744
rect 40132 13728 40184 13734
rect 40038 13696 40094 13705
rect 40132 13670 40184 13676
rect 40038 13631 40094 13640
rect 40040 13320 40092 13326
rect 40040 13262 40092 13268
rect 40052 12918 40080 13262
rect 40040 12912 40092 12918
rect 40038 12880 40040 12889
rect 40092 12880 40094 12889
rect 40038 12815 40094 12824
rect 39948 12368 40000 12374
rect 39948 12310 40000 12316
rect 39856 12232 39908 12238
rect 39856 12174 39908 12180
rect 39478 11996 39786 12016
rect 39478 11994 39484 11996
rect 39540 11994 39564 11996
rect 39620 11994 39644 11996
rect 39700 11994 39724 11996
rect 39780 11994 39786 11996
rect 39540 11942 39542 11994
rect 39722 11942 39724 11994
rect 39478 11940 39484 11942
rect 39540 11940 39564 11942
rect 39620 11940 39644 11942
rect 39700 11940 39724 11942
rect 39780 11940 39786 11942
rect 39478 11920 39786 11940
rect 39868 11354 39896 12174
rect 39856 11348 39908 11354
rect 39856 11290 39908 11296
rect 39396 11212 39448 11218
rect 39396 11154 39448 11160
rect 39478 10908 39786 10928
rect 39478 10906 39484 10908
rect 39540 10906 39564 10908
rect 39620 10906 39644 10908
rect 39700 10906 39724 10908
rect 39780 10906 39786 10908
rect 39540 10854 39542 10906
rect 39722 10854 39724 10906
rect 39478 10852 39484 10854
rect 39540 10852 39564 10854
rect 39620 10852 39644 10854
rect 39700 10852 39724 10854
rect 39780 10852 39786 10854
rect 39478 10832 39786 10852
rect 40052 10266 40080 12815
rect 40040 10260 40092 10266
rect 40040 10202 40092 10208
rect 40052 10062 40080 10202
rect 40040 10056 40092 10062
rect 40040 9998 40092 10004
rect 39478 9820 39786 9840
rect 39478 9818 39484 9820
rect 39540 9818 39564 9820
rect 39620 9818 39644 9820
rect 39700 9818 39724 9820
rect 39780 9818 39786 9820
rect 39540 9766 39542 9818
rect 39722 9766 39724 9818
rect 39478 9764 39484 9766
rect 39540 9764 39564 9766
rect 39620 9764 39644 9766
rect 39700 9764 39724 9766
rect 39780 9764 39786 9766
rect 39478 9744 39786 9764
rect 39478 8732 39786 8752
rect 39478 8730 39484 8732
rect 39540 8730 39564 8732
rect 39620 8730 39644 8732
rect 39700 8730 39724 8732
rect 39780 8730 39786 8732
rect 39540 8678 39542 8730
rect 39722 8678 39724 8730
rect 39478 8676 39484 8678
rect 39540 8676 39564 8678
rect 39620 8676 39644 8678
rect 39700 8676 39724 8678
rect 39780 8676 39786 8678
rect 39478 8656 39786 8676
rect 39478 7644 39786 7664
rect 39478 7642 39484 7644
rect 39540 7642 39564 7644
rect 39620 7642 39644 7644
rect 39700 7642 39724 7644
rect 39780 7642 39786 7644
rect 39540 7590 39542 7642
rect 39722 7590 39724 7642
rect 39478 7588 39484 7590
rect 39540 7588 39564 7590
rect 39620 7588 39644 7590
rect 39700 7588 39724 7590
rect 39780 7588 39786 7590
rect 39478 7568 39786 7588
rect 40144 6769 40172 13670
rect 40224 13184 40276 13190
rect 40224 13126 40276 13132
rect 40236 8634 40264 13126
rect 40328 11898 40356 18566
rect 40406 18456 40462 18465
rect 40406 18391 40462 18400
rect 40420 14822 40448 18391
rect 40408 14816 40460 14822
rect 40408 14758 40460 14764
rect 40408 14408 40460 14414
rect 40408 14350 40460 14356
rect 40420 12850 40448 14350
rect 40408 12844 40460 12850
rect 40408 12786 40460 12792
rect 40420 12617 40448 12786
rect 40512 12753 40540 20266
rect 40604 18834 40632 21082
rect 40696 20262 40724 23598
rect 40774 23559 40830 23568
rect 40788 21146 40816 23559
rect 40776 21140 40828 21146
rect 40776 21082 40828 21088
rect 40880 20890 40908 25191
rect 40788 20862 40908 20890
rect 40684 20256 40736 20262
rect 40684 20198 40736 20204
rect 40788 20058 40816 20862
rect 40972 20398 41000 26250
rect 41064 23254 41092 27270
rect 41236 23588 41288 23594
rect 41236 23530 41288 23536
rect 41052 23248 41104 23254
rect 41052 23190 41104 23196
rect 41248 22642 41276 23530
rect 41328 22976 41380 22982
rect 41328 22918 41380 22924
rect 41236 22636 41288 22642
rect 41236 22578 41288 22584
rect 41144 21956 41196 21962
rect 41144 21898 41196 21904
rect 41052 21480 41104 21486
rect 41052 21422 41104 21428
rect 40960 20392 41012 20398
rect 40960 20334 41012 20340
rect 40776 20052 40828 20058
rect 40776 19994 40828 20000
rect 40868 19984 40920 19990
rect 41064 19938 41092 21422
rect 41156 20330 41184 21898
rect 41248 20788 41276 22578
rect 41340 22438 41368 22918
rect 41432 22778 41460 28086
rect 41420 22772 41472 22778
rect 41420 22714 41472 22720
rect 41328 22432 41380 22438
rect 41328 22374 41380 22380
rect 41524 22001 41552 29135
rect 44362 29064 44418 29073
rect 44362 28999 44418 29008
rect 44272 27940 44324 27946
rect 44272 27882 44324 27888
rect 43350 27704 43406 27713
rect 43350 27639 43406 27648
rect 41604 26852 41656 26858
rect 41604 26794 41656 26800
rect 41616 23526 41644 26794
rect 43166 25936 43222 25945
rect 43166 25871 43222 25880
rect 42892 24880 42944 24886
rect 42892 24822 42944 24828
rect 41696 24336 41748 24342
rect 41696 24278 41748 24284
rect 41604 23520 41656 23526
rect 41604 23462 41656 23468
rect 41708 22250 41736 24278
rect 42708 24064 42760 24070
rect 42708 24006 42760 24012
rect 42064 23792 42116 23798
rect 42064 23734 42116 23740
rect 41788 23520 41840 23526
rect 41788 23462 41840 23468
rect 41616 22222 41736 22250
rect 41510 21992 41566 22001
rect 41510 21927 41566 21936
rect 41328 21888 41380 21894
rect 41328 21830 41380 21836
rect 41340 20942 41368 21830
rect 41512 21480 41564 21486
rect 41512 21422 41564 21428
rect 41524 20942 41552 21422
rect 41328 20936 41380 20942
rect 41328 20878 41380 20884
rect 41512 20936 41564 20942
rect 41512 20878 41564 20884
rect 41248 20760 41368 20788
rect 41144 20324 41196 20330
rect 41144 20266 41196 20272
rect 40868 19926 40920 19932
rect 40880 19446 40908 19926
rect 40972 19910 41092 19938
rect 40972 19530 41000 19910
rect 41052 19848 41104 19854
rect 41050 19816 41052 19825
rect 41104 19816 41106 19825
rect 41050 19751 41106 19760
rect 41144 19780 41196 19786
rect 41144 19722 41196 19728
rect 40972 19502 41092 19530
rect 40868 19440 40920 19446
rect 40868 19382 40920 19388
rect 40958 19408 41014 19417
rect 40958 19343 41014 19352
rect 40972 19174 41000 19343
rect 40960 19168 41012 19174
rect 40960 19110 41012 19116
rect 40592 18828 40644 18834
rect 40592 18770 40644 18776
rect 40958 18184 41014 18193
rect 40958 18119 41014 18128
rect 40972 17746 41000 18119
rect 40960 17740 41012 17746
rect 40960 17682 41012 17688
rect 40592 17604 40644 17610
rect 40592 17546 40644 17552
rect 40604 17270 40632 17546
rect 40592 17264 40644 17270
rect 40592 17206 40644 17212
rect 40604 16522 40632 17206
rect 40592 16516 40644 16522
rect 40592 16458 40644 16464
rect 40604 15502 40632 16458
rect 41064 16250 41092 19502
rect 41156 19242 41184 19722
rect 41236 19440 41288 19446
rect 41236 19382 41288 19388
rect 41144 19236 41196 19242
rect 41144 19178 41196 19184
rect 41248 18766 41276 19382
rect 41236 18760 41288 18766
rect 41236 18702 41288 18708
rect 41340 18465 41368 20760
rect 41616 20346 41644 22222
rect 41696 22092 41748 22098
rect 41696 22034 41748 22040
rect 41708 20806 41736 22034
rect 41696 20800 41748 20806
rect 41696 20742 41748 20748
rect 41432 20318 41644 20346
rect 41326 18456 41382 18465
rect 41326 18391 41382 18400
rect 41432 18306 41460 20318
rect 41604 20256 41656 20262
rect 41604 20198 41656 20204
rect 41616 19417 41644 20198
rect 41602 19408 41658 19417
rect 41602 19343 41658 19352
rect 41602 18592 41658 18601
rect 41602 18527 41658 18536
rect 41616 18426 41644 18527
rect 41604 18420 41656 18426
rect 41604 18362 41656 18368
rect 41340 18290 41460 18306
rect 41328 18284 41460 18290
rect 41380 18278 41460 18284
rect 41510 18320 41566 18329
rect 41510 18255 41566 18264
rect 41328 18226 41380 18232
rect 41328 18080 41380 18086
rect 41420 18080 41472 18086
rect 41328 18022 41380 18028
rect 41418 18048 41420 18057
rect 41472 18048 41474 18057
rect 41340 17898 41368 18022
rect 41418 17983 41474 17992
rect 41340 17870 41460 17898
rect 41328 17604 41380 17610
rect 41328 17546 41380 17552
rect 41142 17368 41198 17377
rect 41236 17332 41288 17338
rect 41198 17312 41236 17320
rect 41142 17303 41236 17312
rect 41156 17292 41236 17303
rect 41052 16244 41104 16250
rect 41052 16186 41104 16192
rect 40960 16040 41012 16046
rect 40960 15982 41012 15988
rect 40972 15910 41000 15982
rect 40960 15904 41012 15910
rect 40960 15846 41012 15852
rect 40972 15745 41000 15846
rect 40958 15736 41014 15745
rect 41064 15706 41092 16186
rect 40958 15671 41014 15680
rect 41052 15700 41104 15706
rect 41052 15642 41104 15648
rect 40592 15496 40644 15502
rect 40592 15438 40644 15444
rect 40866 15464 40922 15473
rect 40604 15162 40632 15438
rect 41156 15434 41184 17292
rect 41236 17274 41288 17280
rect 41340 17241 41368 17546
rect 41326 17232 41382 17241
rect 41326 17167 41382 17176
rect 41432 16522 41460 17870
rect 41524 17649 41552 18255
rect 41708 18057 41736 20742
rect 41800 20058 41828 23462
rect 41970 23080 42026 23089
rect 41970 23015 42026 23024
rect 41878 22264 41934 22273
rect 41878 22199 41934 22208
rect 41788 20052 41840 20058
rect 41788 19994 41840 20000
rect 41892 19242 41920 22199
rect 41880 19236 41932 19242
rect 41880 19178 41932 19184
rect 41788 19168 41840 19174
rect 41788 19110 41840 19116
rect 41694 18048 41750 18057
rect 41694 17983 41750 17992
rect 41800 17796 41828 19110
rect 41984 18970 42012 23015
rect 42076 21894 42104 23734
rect 42340 22976 42392 22982
rect 42340 22918 42392 22924
rect 42616 22976 42668 22982
rect 42616 22918 42668 22924
rect 42064 21888 42116 21894
rect 42064 21830 42116 21836
rect 42154 21584 42210 21593
rect 42154 21519 42210 21528
rect 42062 21176 42118 21185
rect 42168 21146 42196 21519
rect 42062 21111 42064 21120
rect 42116 21111 42118 21120
rect 42156 21140 42208 21146
rect 42064 21082 42116 21088
rect 42156 21082 42208 21088
rect 42064 20460 42116 20466
rect 42064 20402 42116 20408
rect 41972 18964 42024 18970
rect 41972 18906 42024 18912
rect 42076 18329 42104 20402
rect 42168 19854 42196 21082
rect 42246 21040 42302 21049
rect 42246 20975 42302 20984
rect 42156 19848 42208 19854
rect 42156 19790 42208 19796
rect 42062 18320 42118 18329
rect 41880 18284 41932 18290
rect 42062 18255 42118 18264
rect 41880 18226 41932 18232
rect 41616 17768 41828 17796
rect 41510 17640 41566 17649
rect 41510 17575 41566 17584
rect 41512 16992 41564 16998
rect 41512 16934 41564 16940
rect 41420 16516 41472 16522
rect 41420 16458 41472 16464
rect 41524 16402 41552 16934
rect 41616 16810 41644 17768
rect 41800 17678 41828 17709
rect 41788 17672 41840 17678
rect 41786 17640 41788 17649
rect 41840 17640 41842 17649
rect 41892 17610 41920 18226
rect 42064 18216 42116 18222
rect 42064 18158 42116 18164
rect 42076 17626 42104 18158
rect 42260 17814 42288 20975
rect 42248 17808 42300 17814
rect 42248 17750 42300 17756
rect 41786 17575 41842 17584
rect 41880 17604 41932 17610
rect 41696 17536 41748 17542
rect 41696 17478 41748 17484
rect 41708 17105 41736 17478
rect 41800 17270 41828 17575
rect 41880 17546 41932 17552
rect 41984 17598 42104 17626
rect 41788 17264 41840 17270
rect 41788 17206 41840 17212
rect 41694 17096 41750 17105
rect 41694 17031 41750 17040
rect 41616 16782 41736 16810
rect 41604 16720 41656 16726
rect 41604 16662 41656 16668
rect 41432 16374 41552 16402
rect 40866 15399 40922 15408
rect 41144 15428 41196 15434
rect 40592 15156 40644 15162
rect 40592 15098 40644 15104
rect 40604 14958 40632 15098
rect 40880 14958 40908 15399
rect 41144 15370 41196 15376
rect 41052 15020 41104 15026
rect 41052 14962 41104 14968
rect 40592 14952 40644 14958
rect 40868 14952 40920 14958
rect 40592 14894 40644 14900
rect 40866 14920 40868 14929
rect 40920 14920 40922 14929
rect 40776 14884 40828 14890
rect 40866 14855 40922 14864
rect 40776 14826 40828 14832
rect 40684 14816 40736 14822
rect 40684 14758 40736 14764
rect 40592 14612 40644 14618
rect 40592 14554 40644 14560
rect 40498 12744 40554 12753
rect 40498 12679 40554 12688
rect 40406 12608 40462 12617
rect 40406 12543 40462 12552
rect 40604 12442 40632 14554
rect 40696 13977 40724 14758
rect 40788 14346 40816 14826
rect 40880 14618 40908 14855
rect 40958 14784 41014 14793
rect 40958 14719 41014 14728
rect 40868 14612 40920 14618
rect 40868 14554 40920 14560
rect 40972 14550 41000 14719
rect 41064 14618 41092 14962
rect 41052 14612 41104 14618
rect 41052 14554 41104 14560
rect 40960 14544 41012 14550
rect 41156 14498 41184 15370
rect 41328 14612 41380 14618
rect 41328 14554 41380 14560
rect 40960 14486 41012 14492
rect 40868 14476 40920 14482
rect 40868 14418 40920 14424
rect 41064 14470 41184 14498
rect 41234 14512 41290 14521
rect 40776 14340 40828 14346
rect 40776 14282 40828 14288
rect 40682 13968 40738 13977
rect 40788 13938 40816 14282
rect 40682 13903 40738 13912
rect 40776 13932 40828 13938
rect 40776 13874 40828 13880
rect 40776 13796 40828 13802
rect 40776 13738 40828 13744
rect 40592 12436 40644 12442
rect 40592 12378 40644 12384
rect 40408 12368 40460 12374
rect 40406 12336 40408 12345
rect 40460 12336 40462 12345
rect 40406 12271 40462 12280
rect 40788 11898 40816 13738
rect 40880 12714 40908 14418
rect 40960 14408 41012 14414
rect 40960 14350 41012 14356
rect 40868 12708 40920 12714
rect 40868 12650 40920 12656
rect 40868 12096 40920 12102
rect 40972 12084 41000 14350
rect 40920 12056 41000 12084
rect 40868 12038 40920 12044
rect 40316 11892 40368 11898
rect 40316 11834 40368 11840
rect 40776 11892 40828 11898
rect 40776 11834 40828 11840
rect 40328 11801 40356 11834
rect 40314 11792 40370 11801
rect 40314 11727 40370 11736
rect 40498 11792 40554 11801
rect 40498 11727 40554 11736
rect 40512 11529 40540 11727
rect 40498 11520 40554 11529
rect 40498 11455 40554 11464
rect 40880 9722 40908 12038
rect 41064 11914 41092 14470
rect 41234 14447 41290 14456
rect 41144 13932 41196 13938
rect 41144 13874 41196 13880
rect 40972 11886 41092 11914
rect 40972 10130 41000 11886
rect 41052 11756 41104 11762
rect 41052 11698 41104 11704
rect 41064 10266 41092 11698
rect 41156 10742 41184 13874
rect 41248 13530 41276 14447
rect 41340 13841 41368 14554
rect 41432 14006 41460 16374
rect 41512 15700 41564 15706
rect 41512 15642 41564 15648
rect 41524 14618 41552 15642
rect 41512 14612 41564 14618
rect 41512 14554 41564 14560
rect 41512 14272 41564 14278
rect 41512 14214 41564 14220
rect 41524 14006 41552 14214
rect 41420 14000 41472 14006
rect 41420 13942 41472 13948
rect 41512 14000 41564 14006
rect 41512 13942 41564 13948
rect 41512 13864 41564 13870
rect 41326 13832 41382 13841
rect 41512 13806 41564 13812
rect 41326 13767 41382 13776
rect 41236 13524 41288 13530
rect 41288 13484 41460 13512
rect 41236 13466 41288 13472
rect 41236 13252 41288 13258
rect 41236 13194 41288 13200
rect 41328 13252 41380 13258
rect 41328 13194 41380 13200
rect 41248 12714 41276 13194
rect 41340 12918 41368 13194
rect 41432 13190 41460 13484
rect 41420 13184 41472 13190
rect 41420 13126 41472 13132
rect 41432 12986 41460 13126
rect 41420 12980 41472 12986
rect 41420 12922 41472 12928
rect 41328 12912 41380 12918
rect 41328 12854 41380 12860
rect 41236 12708 41288 12714
rect 41236 12650 41288 12656
rect 41418 12064 41474 12073
rect 41418 11999 41474 12008
rect 41432 11898 41460 11999
rect 41420 11892 41472 11898
rect 41420 11834 41472 11840
rect 41524 11370 41552 13806
rect 41616 13326 41644 16662
rect 41708 15570 41736 16782
rect 41800 16590 41828 17206
rect 41892 16998 41920 17546
rect 41880 16992 41932 16998
rect 41880 16934 41932 16940
rect 41984 16810 42012 17598
rect 42064 17536 42116 17542
rect 42064 17478 42116 17484
rect 41892 16782 42012 16810
rect 41788 16584 41840 16590
rect 41788 16526 41840 16532
rect 41892 15910 41920 16782
rect 42076 16697 42104 17478
rect 42246 17368 42302 17377
rect 42246 17303 42302 17312
rect 42156 17196 42208 17202
rect 42156 17138 42208 17144
rect 42062 16688 42118 16697
rect 41972 16652 42024 16658
rect 42062 16623 42118 16632
rect 41972 16594 42024 16600
rect 41984 16289 42012 16594
rect 42168 16538 42196 17138
rect 42260 16658 42288 17303
rect 42248 16652 42300 16658
rect 42248 16594 42300 16600
rect 42076 16510 42196 16538
rect 41970 16280 42026 16289
rect 41970 16215 42026 16224
rect 41880 15904 41932 15910
rect 41880 15846 41932 15852
rect 41696 15564 41748 15570
rect 41696 15506 41748 15512
rect 41708 15076 41736 15506
rect 41892 15366 41920 15846
rect 41972 15496 42024 15502
rect 41972 15438 42024 15444
rect 41880 15360 41932 15366
rect 41880 15302 41932 15308
rect 41788 15088 41840 15094
rect 41708 15048 41788 15076
rect 41708 14414 41736 15048
rect 41788 15030 41840 15036
rect 41788 14952 41840 14958
rect 41840 14900 41920 14906
rect 41788 14894 41920 14900
rect 41800 14878 41920 14894
rect 41788 14816 41840 14822
rect 41788 14758 41840 14764
rect 41696 14408 41748 14414
rect 41696 14350 41748 14356
rect 41708 13870 41736 14350
rect 41696 13864 41748 13870
rect 41696 13806 41748 13812
rect 41696 13728 41748 13734
rect 41696 13670 41748 13676
rect 41604 13320 41656 13326
rect 41604 13262 41656 13268
rect 41604 13184 41656 13190
rect 41708 13172 41736 13670
rect 41656 13144 41736 13172
rect 41604 13126 41656 13132
rect 41236 11348 41288 11354
rect 41236 11290 41288 11296
rect 41432 11342 41552 11370
rect 41248 10810 41276 11290
rect 41236 10804 41288 10810
rect 41236 10746 41288 10752
rect 41144 10736 41196 10742
rect 41144 10678 41196 10684
rect 41432 10305 41460 11342
rect 41512 11212 41564 11218
rect 41512 11154 41564 11160
rect 41418 10296 41474 10305
rect 41052 10260 41104 10266
rect 41418 10231 41474 10240
rect 41052 10202 41104 10208
rect 40960 10124 41012 10130
rect 40960 10066 41012 10072
rect 40868 9716 40920 9722
rect 40868 9658 40920 9664
rect 41524 9625 41552 11154
rect 41510 9616 41566 9625
rect 41510 9551 41566 9560
rect 40224 8628 40276 8634
rect 40224 8570 40276 8576
rect 41616 7449 41644 13126
rect 41696 10804 41748 10810
rect 41696 10746 41748 10752
rect 41708 9518 41736 10746
rect 41696 9512 41748 9518
rect 41696 9454 41748 9460
rect 41602 7440 41658 7449
rect 41602 7375 41658 7384
rect 40130 6760 40186 6769
rect 40130 6695 40186 6704
rect 39478 6556 39786 6576
rect 39478 6554 39484 6556
rect 39540 6554 39564 6556
rect 39620 6554 39644 6556
rect 39700 6554 39724 6556
rect 39780 6554 39786 6556
rect 39540 6502 39542 6554
rect 39722 6502 39724 6554
rect 39478 6500 39484 6502
rect 39540 6500 39564 6502
rect 39620 6500 39644 6502
rect 39700 6500 39724 6502
rect 39780 6500 39786 6502
rect 39478 6480 39786 6500
rect 39120 6180 39172 6186
rect 39120 6122 39172 6128
rect 39478 5468 39786 5488
rect 39478 5466 39484 5468
rect 39540 5466 39564 5468
rect 39620 5466 39644 5468
rect 39700 5466 39724 5468
rect 39780 5466 39786 5468
rect 39540 5414 39542 5466
rect 39722 5414 39724 5466
rect 39478 5412 39484 5414
rect 39540 5412 39564 5414
rect 39620 5412 39644 5414
rect 39700 5412 39724 5414
rect 39780 5412 39786 5414
rect 39478 5392 39786 5412
rect 41708 4554 41736 9454
rect 41800 5370 41828 14758
rect 41892 6730 41920 14878
rect 41984 13734 42012 15438
rect 41972 13728 42024 13734
rect 41972 13670 42024 13676
rect 42076 12434 42104 16510
rect 42248 16108 42300 16114
rect 42248 16050 42300 16056
rect 42156 14952 42208 14958
rect 42156 14894 42208 14900
rect 41984 12406 42104 12434
rect 41984 10198 42012 12406
rect 42064 12096 42116 12102
rect 42064 12038 42116 12044
rect 42076 11801 42104 12038
rect 42062 11792 42118 11801
rect 42062 11727 42118 11736
rect 42168 11694 42196 14894
rect 42260 14414 42288 16050
rect 42352 15638 42380 22918
rect 42628 22234 42656 22918
rect 42616 22228 42668 22234
rect 42616 22170 42668 22176
rect 42720 21894 42748 24006
rect 42800 22500 42852 22506
rect 42800 22442 42852 22448
rect 42432 21888 42484 21894
rect 42432 21830 42484 21836
rect 42708 21888 42760 21894
rect 42708 21830 42760 21836
rect 42444 18426 42472 21830
rect 42524 21344 42576 21350
rect 42524 21286 42576 21292
rect 42536 20534 42564 21286
rect 42524 20528 42576 20534
rect 42524 20470 42576 20476
rect 42616 20460 42668 20466
rect 42616 20402 42668 20408
rect 42524 20256 42576 20262
rect 42628 20233 42656 20402
rect 42524 20198 42576 20204
rect 42614 20224 42670 20233
rect 42536 19825 42564 20198
rect 42614 20159 42670 20168
rect 42522 19816 42578 19825
rect 42522 19751 42578 19760
rect 42706 19408 42762 19417
rect 42812 19378 42840 22442
rect 42706 19343 42708 19352
rect 42760 19343 42762 19352
rect 42800 19372 42852 19378
rect 42708 19314 42760 19320
rect 42800 19314 42852 19320
rect 42800 19236 42852 19242
rect 42800 19178 42852 19184
rect 42524 18896 42576 18902
rect 42524 18838 42576 18844
rect 42432 18420 42484 18426
rect 42432 18362 42484 18368
rect 42430 18048 42486 18057
rect 42430 17983 42486 17992
rect 42444 17542 42472 17983
rect 42432 17536 42484 17542
rect 42432 17478 42484 17484
rect 42536 16046 42564 18838
rect 42812 18737 42840 19178
rect 42798 18728 42854 18737
rect 42904 18698 42932 24822
rect 42984 23316 43036 23322
rect 42984 23258 43036 23264
rect 42996 22778 43024 23258
rect 42984 22772 43036 22778
rect 42984 22714 43036 22720
rect 42996 22234 43024 22714
rect 42984 22228 43036 22234
rect 42984 22170 43036 22176
rect 42984 20868 43036 20874
rect 42984 20810 43036 20816
rect 42996 19854 43024 20810
rect 43076 20800 43128 20806
rect 43076 20742 43128 20748
rect 42984 19848 43036 19854
rect 42984 19790 43036 19796
rect 42984 19372 43036 19378
rect 42984 19314 43036 19320
rect 42996 19174 43024 19314
rect 42984 19168 43036 19174
rect 42984 19110 43036 19116
rect 43088 18834 43116 20742
rect 43180 20602 43208 25871
rect 43260 21888 43312 21894
rect 43260 21830 43312 21836
rect 43272 20874 43300 21830
rect 43260 20868 43312 20874
rect 43260 20810 43312 20816
rect 43168 20596 43220 20602
rect 43168 20538 43220 20544
rect 43272 20466 43300 20810
rect 43260 20460 43312 20466
rect 43260 20402 43312 20408
rect 43166 20360 43222 20369
rect 43166 20295 43222 20304
rect 43180 19378 43208 20295
rect 43272 19961 43300 20402
rect 43258 19952 43314 19961
rect 43258 19887 43314 19896
rect 43168 19372 43220 19378
rect 43168 19314 43220 19320
rect 43260 19372 43312 19378
rect 43260 19314 43312 19320
rect 43272 19145 43300 19314
rect 43258 19136 43314 19145
rect 43258 19071 43314 19080
rect 43076 18828 43128 18834
rect 43076 18770 43128 18776
rect 42798 18663 42854 18672
rect 42892 18692 42944 18698
rect 42812 18290 42840 18663
rect 42892 18634 42944 18640
rect 42800 18284 42852 18290
rect 42800 18226 42852 18232
rect 42904 18222 42932 18634
rect 43088 18630 43116 18770
rect 43260 18760 43312 18766
rect 43260 18702 43312 18708
rect 42984 18624 43036 18630
rect 42984 18566 43036 18572
rect 43076 18624 43128 18630
rect 43272 18601 43300 18702
rect 43076 18566 43128 18572
rect 43258 18592 43314 18601
rect 42708 18216 42760 18222
rect 42708 18158 42760 18164
rect 42892 18216 42944 18222
rect 42892 18158 42944 18164
rect 42720 18086 42748 18158
rect 42708 18080 42760 18086
rect 42708 18022 42760 18028
rect 42706 17912 42762 17921
rect 42706 17847 42762 17856
rect 42616 17740 42668 17746
rect 42616 17682 42668 17688
rect 42628 17066 42656 17682
rect 42720 17338 42748 17847
rect 42800 17536 42852 17542
rect 42800 17478 42852 17484
rect 42708 17332 42760 17338
rect 42708 17274 42760 17280
rect 42812 17105 42840 17478
rect 42996 17105 43024 18566
rect 43258 18527 43314 18536
rect 43168 18284 43220 18290
rect 43168 18226 43220 18232
rect 43074 17776 43130 17785
rect 43074 17711 43130 17720
rect 42798 17096 42854 17105
rect 42616 17060 42668 17066
rect 42798 17031 42854 17040
rect 42982 17096 43038 17105
rect 42982 17031 43038 17040
rect 42616 17002 42668 17008
rect 42890 16960 42946 16969
rect 42890 16895 42946 16904
rect 42708 16584 42760 16590
rect 42708 16526 42760 16532
rect 42524 16040 42576 16046
rect 42524 15982 42576 15988
rect 42432 15904 42484 15910
rect 42432 15846 42484 15852
rect 42340 15632 42392 15638
rect 42340 15574 42392 15580
rect 42340 15360 42392 15366
rect 42444 15337 42472 15846
rect 42536 15706 42564 15982
rect 42524 15700 42576 15706
rect 42524 15642 42576 15648
rect 42616 15632 42668 15638
rect 42616 15574 42668 15580
rect 42524 15428 42576 15434
rect 42524 15370 42576 15376
rect 42340 15302 42392 15308
rect 42430 15328 42486 15337
rect 42248 14408 42300 14414
rect 42248 14350 42300 14356
rect 42352 14362 42380 15302
rect 42430 15263 42486 15272
rect 42536 14958 42564 15370
rect 42524 14952 42576 14958
rect 42524 14894 42576 14900
rect 42352 14334 42472 14362
rect 42340 14272 42392 14278
rect 42340 14214 42392 14220
rect 42352 13841 42380 14214
rect 42338 13832 42394 13841
rect 42338 13767 42394 13776
rect 42444 13138 42472 14334
rect 42524 13728 42576 13734
rect 42524 13670 42576 13676
rect 42352 13110 42472 13138
rect 42352 12986 42380 13110
rect 42340 12980 42392 12986
rect 42340 12922 42392 12928
rect 42432 12980 42484 12986
rect 42432 12922 42484 12928
rect 42444 12714 42472 12922
rect 42536 12850 42564 13670
rect 42628 13530 42656 15574
rect 42720 13938 42748 16526
rect 42904 16114 42932 16895
rect 43088 16726 43116 17711
rect 43076 16720 43128 16726
rect 43076 16662 43128 16668
rect 42800 16108 42852 16114
rect 42800 16050 42852 16056
rect 42892 16108 42944 16114
rect 42892 16050 42944 16056
rect 42812 14006 42840 16050
rect 42904 15201 42932 16050
rect 43180 15978 43208 18226
rect 43258 18184 43314 18193
rect 43258 18119 43314 18128
rect 43272 17814 43300 18119
rect 43260 17808 43312 17814
rect 43260 17750 43312 17756
rect 43260 17060 43312 17066
rect 43260 17002 43312 17008
rect 43168 15972 43220 15978
rect 43168 15914 43220 15920
rect 43168 15496 43220 15502
rect 43168 15438 43220 15444
rect 42984 15360 43036 15366
rect 42984 15302 43036 15308
rect 42890 15192 42946 15201
rect 42890 15127 42946 15136
rect 42892 14816 42944 14822
rect 42996 14804 43024 15302
rect 42944 14776 43024 14804
rect 43076 14816 43128 14822
rect 42892 14758 42944 14764
rect 43076 14758 43128 14764
rect 42800 14000 42852 14006
rect 42800 13942 42852 13948
rect 42708 13932 42760 13938
rect 42708 13874 42760 13880
rect 42616 13524 42668 13530
rect 42616 13466 42668 13472
rect 42524 12844 42576 12850
rect 42524 12786 42576 12792
rect 42432 12708 42484 12714
rect 42432 12650 42484 12656
rect 42156 11688 42208 11694
rect 42156 11630 42208 11636
rect 42536 11082 42564 12786
rect 42628 11626 42656 13466
rect 42812 13394 42840 13942
rect 42800 13388 42852 13394
rect 42800 13330 42852 13336
rect 42904 13190 42932 14758
rect 42984 14544 43036 14550
rect 42984 14486 43036 14492
rect 42996 14074 43024 14486
rect 42984 14068 43036 14074
rect 42984 14010 43036 14016
rect 42892 13184 42944 13190
rect 42892 13126 42944 13132
rect 42708 11892 42760 11898
rect 42708 11834 42760 11840
rect 42616 11620 42668 11626
rect 42616 11562 42668 11568
rect 42720 11354 42748 11834
rect 42708 11348 42760 11354
rect 42708 11290 42760 11296
rect 42524 11076 42576 11082
rect 42524 11018 42576 11024
rect 41972 10192 42024 10198
rect 41972 10134 42024 10140
rect 43088 8022 43116 14758
rect 43180 11393 43208 15438
rect 43166 11384 43222 11393
rect 43166 11319 43222 11328
rect 43272 9586 43300 17002
rect 43364 15706 43392 27639
rect 44180 27056 44232 27062
rect 44180 26998 44232 27004
rect 43442 26480 43498 26489
rect 43442 26415 43498 26424
rect 43536 26444 43588 26450
rect 43456 16114 43484 26415
rect 43536 26386 43588 26392
rect 43548 22506 43576 26386
rect 43904 22704 43956 22710
rect 43904 22646 43956 22652
rect 43536 22500 43588 22506
rect 43536 22442 43588 22448
rect 43916 22166 43944 22646
rect 43904 22160 43956 22166
rect 43904 22102 43956 22108
rect 44088 22092 44140 22098
rect 44088 22034 44140 22040
rect 44100 21690 44128 22034
rect 44088 21684 44140 21690
rect 44088 21626 44140 21632
rect 44100 21146 44128 21626
rect 44088 21140 44140 21146
rect 44088 21082 44140 21088
rect 43720 21004 43772 21010
rect 43720 20946 43772 20952
rect 43534 20904 43590 20913
rect 43534 20839 43590 20848
rect 43444 16108 43496 16114
rect 43444 16050 43496 16056
rect 43444 15972 43496 15978
rect 43444 15914 43496 15920
rect 43456 15706 43484 15914
rect 43352 15700 43404 15706
rect 43352 15642 43404 15648
rect 43444 15700 43496 15706
rect 43444 15642 43496 15648
rect 43352 15428 43404 15434
rect 43352 15370 43404 15376
rect 43364 13326 43392 15370
rect 43548 15162 43576 20839
rect 43628 19168 43680 19174
rect 43628 19110 43680 19116
rect 43640 18902 43668 19110
rect 43628 18896 43680 18902
rect 43628 18838 43680 18844
rect 43732 18766 43760 20946
rect 43812 19848 43864 19854
rect 43812 19790 43864 19796
rect 43824 19378 43852 19790
rect 44088 19712 44140 19718
rect 44088 19654 44140 19660
rect 44100 19446 44128 19654
rect 44088 19440 44140 19446
rect 44088 19382 44140 19388
rect 43812 19372 43864 19378
rect 43812 19314 43864 19320
rect 43902 19000 43958 19009
rect 43902 18935 43958 18944
rect 43720 18760 43772 18766
rect 43720 18702 43772 18708
rect 43628 18624 43680 18630
rect 43628 18566 43680 18572
rect 43812 18624 43864 18630
rect 43812 18566 43864 18572
rect 43640 16046 43668 18566
rect 43824 18358 43852 18566
rect 43812 18352 43864 18358
rect 43812 18294 43864 18300
rect 43916 18222 43944 18935
rect 43994 18456 44050 18465
rect 43994 18391 44050 18400
rect 43904 18216 43956 18222
rect 43904 18158 43956 18164
rect 44008 17134 44036 18391
rect 44100 17678 44128 19382
rect 44192 18426 44220 26998
rect 44180 18420 44232 18426
rect 44180 18362 44232 18368
rect 44284 17882 44312 27882
rect 44180 17876 44232 17882
rect 44180 17818 44232 17824
rect 44272 17876 44324 17882
rect 44272 17818 44324 17824
rect 44088 17672 44140 17678
rect 44088 17614 44140 17620
rect 44192 17270 44220 17818
rect 44180 17264 44232 17270
rect 44180 17206 44232 17212
rect 43996 17128 44048 17134
rect 43996 17070 44048 17076
rect 44180 17128 44232 17134
rect 44180 17070 44232 17076
rect 44192 16833 44220 17070
rect 44178 16824 44234 16833
rect 44178 16759 44234 16768
rect 44272 16788 44324 16794
rect 44272 16730 44324 16736
rect 43904 16448 43956 16454
rect 43904 16390 43956 16396
rect 43628 16040 43680 16046
rect 43628 15982 43680 15988
rect 43812 16040 43864 16046
rect 43812 15982 43864 15988
rect 43640 15366 43668 15982
rect 43720 15972 43772 15978
rect 43720 15914 43772 15920
rect 43732 15502 43760 15914
rect 43720 15496 43772 15502
rect 43720 15438 43772 15444
rect 43628 15360 43680 15366
rect 43628 15302 43680 15308
rect 43640 15162 43668 15302
rect 43536 15156 43588 15162
rect 43536 15098 43588 15104
rect 43628 15156 43680 15162
rect 43628 15098 43680 15104
rect 43536 13864 43588 13870
rect 43536 13806 43588 13812
rect 43548 13530 43576 13806
rect 43536 13524 43588 13530
rect 43536 13466 43588 13472
rect 43352 13320 43404 13326
rect 43350 13288 43352 13297
rect 43404 13288 43406 13297
rect 43350 13223 43406 13232
rect 43548 12374 43576 13466
rect 43732 12782 43760 15438
rect 43824 13870 43852 15982
rect 43812 13864 43864 13870
rect 43812 13806 43864 13812
rect 43720 12776 43772 12782
rect 43720 12718 43772 12724
rect 43536 12368 43588 12374
rect 43536 12310 43588 12316
rect 43548 11762 43576 12310
rect 43720 12096 43772 12102
rect 43720 12038 43772 12044
rect 43536 11756 43588 11762
rect 43536 11698 43588 11704
rect 43548 10810 43576 11698
rect 43732 11665 43760 12038
rect 43718 11656 43774 11665
rect 43718 11591 43774 11600
rect 43536 10804 43588 10810
rect 43536 10746 43588 10752
rect 43260 9580 43312 9586
rect 43260 9522 43312 9528
rect 43824 9042 43852 13806
rect 43916 11830 43944 16390
rect 43996 15904 44048 15910
rect 43996 15846 44048 15852
rect 44180 15904 44232 15910
rect 44180 15846 44232 15852
rect 44008 15473 44036 15846
rect 44192 15609 44220 15846
rect 44178 15600 44234 15609
rect 44178 15535 44234 15544
rect 43994 15464 44050 15473
rect 43994 15399 44050 15408
rect 43996 15360 44048 15366
rect 43994 15328 43996 15337
rect 44048 15328 44050 15337
rect 43994 15263 44050 15272
rect 44178 15192 44234 15201
rect 44178 15127 44180 15136
rect 44232 15127 44234 15136
rect 44180 15098 44232 15104
rect 44088 15088 44140 15094
rect 44088 15030 44140 15036
rect 44100 14822 44128 15030
rect 44180 14952 44232 14958
rect 44284 14929 44312 16730
rect 44376 16114 44404 28999
rect 44638 28928 44694 28937
rect 44638 28863 44694 28872
rect 44454 25800 44510 25809
rect 44454 25735 44510 25744
rect 44468 18834 44496 25735
rect 44548 24676 44600 24682
rect 44548 24618 44600 24624
rect 44560 21350 44588 24618
rect 44652 22094 44680 28863
rect 46400 27470 46428 29294
rect 51722 29294 52040 29322
rect 51722 29200 51778 29294
rect 49110 27772 49418 27792
rect 49110 27770 49116 27772
rect 49172 27770 49196 27772
rect 49252 27770 49276 27772
rect 49332 27770 49356 27772
rect 49412 27770 49418 27772
rect 49172 27718 49174 27770
rect 49354 27718 49356 27770
rect 49110 27716 49116 27718
rect 49172 27716 49196 27718
rect 49252 27716 49276 27718
rect 49332 27716 49356 27718
rect 49412 27716 49418 27718
rect 49110 27696 49418 27716
rect 52012 27606 52040 29294
rect 57150 29200 57206 30000
rect 57242 29200 57298 29209
rect 52000 27600 52052 27606
rect 52000 27542 52052 27548
rect 46388 27464 46440 27470
rect 46388 27406 46440 27412
rect 46480 27464 46532 27470
rect 52460 27464 52512 27470
rect 46480 27406 46532 27412
rect 52458 27432 52460 27441
rect 52512 27432 52514 27441
rect 46296 27328 46348 27334
rect 46296 27270 46348 27276
rect 45008 26512 45060 26518
rect 45008 26454 45060 26460
rect 44652 22066 44772 22094
rect 44548 21344 44600 21350
rect 44548 21286 44600 21292
rect 44548 19712 44600 19718
rect 44548 19654 44600 19660
rect 44560 19417 44588 19654
rect 44546 19408 44602 19417
rect 44546 19343 44602 19352
rect 44640 19372 44692 19378
rect 44640 19314 44692 19320
rect 44456 18828 44508 18834
rect 44456 18770 44508 18776
rect 44548 18624 44600 18630
rect 44548 18566 44600 18572
rect 44456 18420 44508 18426
rect 44456 18362 44508 18368
rect 44364 16108 44416 16114
rect 44364 16050 44416 16056
rect 44180 14894 44232 14900
rect 44270 14920 44326 14929
rect 44088 14816 44140 14822
rect 44088 14758 44140 14764
rect 44192 13938 44220 14894
rect 44270 14855 44326 14864
rect 44376 14618 44404 16050
rect 44468 15638 44496 18362
rect 44560 17678 44588 18566
rect 44652 17746 44680 19314
rect 44640 17740 44692 17746
rect 44640 17682 44692 17688
rect 44548 17672 44600 17678
rect 44744 17626 44772 22066
rect 44824 21344 44876 21350
rect 44824 21286 44876 21292
rect 44914 21312 44970 21321
rect 44836 20806 44864 21286
rect 44914 21247 44970 21256
rect 44824 20800 44876 20806
rect 44824 20742 44876 20748
rect 44824 20256 44876 20262
rect 44824 20198 44876 20204
rect 44836 20058 44864 20198
rect 44824 20052 44876 20058
rect 44824 19994 44876 20000
rect 44928 18358 44956 21247
rect 45020 18426 45048 26454
rect 45560 26376 45612 26382
rect 45560 26318 45612 26324
rect 45190 23216 45246 23225
rect 45190 23151 45246 23160
rect 45204 22094 45232 23151
rect 45468 22568 45520 22574
rect 45468 22510 45520 22516
rect 45376 22432 45428 22438
rect 45376 22374 45428 22380
rect 45204 22066 45324 22094
rect 45192 18624 45244 18630
rect 45192 18566 45244 18572
rect 45008 18420 45060 18426
rect 45008 18362 45060 18368
rect 45100 18420 45152 18426
rect 45100 18362 45152 18368
rect 44916 18352 44968 18358
rect 45112 18306 45140 18362
rect 44916 18294 44968 18300
rect 44824 17740 44876 17746
rect 44824 17682 44876 17688
rect 44548 17614 44600 17620
rect 44652 17598 44772 17626
rect 44652 16810 44680 17598
rect 44652 16782 44772 16810
rect 44640 16720 44692 16726
rect 44640 16662 44692 16668
rect 44548 16584 44600 16590
rect 44548 16526 44600 16532
rect 44560 16250 44588 16526
rect 44548 16244 44600 16250
rect 44548 16186 44600 16192
rect 44548 15904 44600 15910
rect 44548 15846 44600 15852
rect 44456 15632 44508 15638
rect 44456 15574 44508 15580
rect 44364 14612 44416 14618
rect 44364 14554 44416 14560
rect 44468 14074 44496 15574
rect 44272 14068 44324 14074
rect 44272 14010 44324 14016
rect 44456 14068 44508 14074
rect 44456 14010 44508 14016
rect 44180 13932 44232 13938
rect 44180 13874 44232 13880
rect 43904 11824 43956 11830
rect 43904 11766 43956 11772
rect 43812 9036 43864 9042
rect 43812 8978 43864 8984
rect 43076 8016 43128 8022
rect 43076 7958 43128 7964
rect 44284 7954 44312 14010
rect 44364 12708 44416 12714
rect 44364 12650 44416 12656
rect 44376 12481 44404 12650
rect 44362 12472 44418 12481
rect 44362 12407 44418 12416
rect 44364 12096 44416 12102
rect 44364 12038 44416 12044
rect 44376 11898 44404 12038
rect 44364 11892 44416 11898
rect 44364 11834 44416 11840
rect 44560 10713 44588 15846
rect 44652 14958 44680 16662
rect 44744 16425 44772 16782
rect 44730 16416 44786 16425
rect 44730 16351 44786 16360
rect 44732 16244 44784 16250
rect 44732 16186 44784 16192
rect 44640 14952 44692 14958
rect 44640 14894 44692 14900
rect 44640 14340 44692 14346
rect 44640 14282 44692 14288
rect 44652 12646 44680 14282
rect 44744 12986 44772 16186
rect 44836 14657 44864 17682
rect 44928 16998 44956 18294
rect 45020 18290 45140 18306
rect 45008 18284 45140 18290
rect 45060 18278 45140 18284
rect 45008 18226 45060 18232
rect 45098 17912 45154 17921
rect 45098 17847 45100 17856
rect 45152 17847 45154 17856
rect 45100 17818 45152 17824
rect 45204 17762 45232 18566
rect 45112 17734 45232 17762
rect 45112 17134 45140 17734
rect 45296 17202 45324 22066
rect 45388 20602 45416 22374
rect 45376 20596 45428 20602
rect 45376 20538 45428 20544
rect 45284 17196 45336 17202
rect 45284 17138 45336 17144
rect 45100 17128 45152 17134
rect 45100 17070 45152 17076
rect 44916 16992 44968 16998
rect 44916 16934 44968 16940
rect 45006 16688 45062 16697
rect 45006 16623 45008 16632
rect 45060 16623 45062 16632
rect 45008 16594 45060 16600
rect 45008 16448 45060 16454
rect 45008 16390 45060 16396
rect 44916 15904 44968 15910
rect 44916 15846 44968 15852
rect 44928 15337 44956 15846
rect 44914 15328 44970 15337
rect 44914 15263 44970 15272
rect 44822 14648 44878 14657
rect 44822 14583 44878 14592
rect 45020 13802 45048 16390
rect 45008 13796 45060 13802
rect 45008 13738 45060 13744
rect 44732 12980 44784 12986
rect 44732 12922 44784 12928
rect 44640 12640 44692 12646
rect 44640 12582 44692 12588
rect 44652 11694 44680 12582
rect 44640 11688 44692 11694
rect 44640 11630 44692 11636
rect 44546 10704 44602 10713
rect 44546 10639 44602 10648
rect 44272 7948 44324 7954
rect 44272 7890 44324 7896
rect 41880 6724 41932 6730
rect 41880 6666 41932 6672
rect 41788 5364 41840 5370
rect 41788 5306 41840 5312
rect 41696 4548 41748 4554
rect 41696 4490 41748 4496
rect 39478 4380 39786 4400
rect 39478 4378 39484 4380
rect 39540 4378 39564 4380
rect 39620 4378 39644 4380
rect 39700 4378 39724 4380
rect 39780 4378 39786 4380
rect 39540 4326 39542 4378
rect 39722 4326 39724 4378
rect 39478 4324 39484 4326
rect 39540 4324 39564 4326
rect 39620 4324 39644 4326
rect 39700 4324 39724 4326
rect 39780 4324 39786 4326
rect 39478 4304 39786 4324
rect 45112 4078 45140 17070
rect 45192 16992 45244 16998
rect 45192 16934 45244 16940
rect 45204 16833 45232 16934
rect 45190 16824 45246 16833
rect 45296 16794 45324 17138
rect 45374 17096 45430 17105
rect 45374 17031 45430 17040
rect 45190 16759 45246 16768
rect 45284 16788 45336 16794
rect 45284 16730 45336 16736
rect 45192 15700 45244 15706
rect 45192 15642 45244 15648
rect 45204 14618 45232 15642
rect 45282 14920 45338 14929
rect 45282 14855 45284 14864
rect 45336 14855 45338 14864
rect 45284 14826 45336 14832
rect 45192 14612 45244 14618
rect 45192 14554 45244 14560
rect 45296 14074 45324 14826
rect 45284 14068 45336 14074
rect 45284 14010 45336 14016
rect 45192 12640 45244 12646
rect 45192 12582 45244 12588
rect 45204 12209 45232 12582
rect 45190 12200 45246 12209
rect 45190 12135 45246 12144
rect 45100 4072 45152 4078
rect 45100 4014 45152 4020
rect 42432 3664 42484 3670
rect 42432 3606 42484 3612
rect 39478 3292 39786 3312
rect 39478 3290 39484 3292
rect 39540 3290 39564 3292
rect 39620 3290 39644 3292
rect 39700 3290 39724 3292
rect 39780 3290 39786 3292
rect 39540 3238 39542 3290
rect 39722 3238 39724 3290
rect 39478 3236 39484 3238
rect 39540 3236 39564 3238
rect 39620 3236 39644 3238
rect 39700 3236 39724 3238
rect 39780 3236 39786 3238
rect 39478 3216 39786 3236
rect 42444 2446 42472 3606
rect 42432 2440 42484 2446
rect 42432 2382 42484 2388
rect 41972 2304 42024 2310
rect 41972 2246 42024 2252
rect 39478 2204 39786 2224
rect 39478 2202 39484 2204
rect 39540 2202 39564 2204
rect 39620 2202 39644 2204
rect 39700 2202 39724 2204
rect 39780 2202 39786 2204
rect 39540 2150 39542 2202
rect 39722 2150 39724 2202
rect 39478 2148 39484 2150
rect 39540 2148 39564 2150
rect 39620 2148 39644 2150
rect 39700 2148 39724 2150
rect 39780 2148 39786 2150
rect 39478 2128 39786 2148
rect 38014 1728 38070 1737
rect 38014 1663 38070 1672
rect 41984 800 42012 2246
rect 45388 2106 45416 17031
rect 45376 2100 45428 2106
rect 45376 2042 45428 2048
rect 45480 2038 45508 22510
rect 45572 19718 45600 26318
rect 46308 24585 46336 27270
rect 46492 26042 46520 27406
rect 52458 27367 52514 27376
rect 57164 27130 57192 29200
rect 57242 29135 57298 29144
rect 57256 27470 57284 29135
rect 57244 27464 57296 27470
rect 57244 27406 57296 27412
rect 58070 27432 58126 27441
rect 57152 27124 57204 27130
rect 57152 27066 57204 27072
rect 57256 27062 57284 27406
rect 57888 27396 57940 27402
rect 58070 27367 58072 27376
rect 57888 27338 57940 27344
rect 58124 27367 58126 27376
rect 58072 27338 58124 27344
rect 57244 27056 57296 27062
rect 57900 27033 57928 27338
rect 57244 26998 57296 27004
rect 57886 27024 57942 27033
rect 56600 26988 56652 26994
rect 57886 26959 57942 26968
rect 56600 26930 56652 26936
rect 49110 26684 49418 26704
rect 49110 26682 49116 26684
rect 49172 26682 49196 26684
rect 49252 26682 49276 26684
rect 49332 26682 49356 26684
rect 49412 26682 49418 26684
rect 49172 26630 49174 26682
rect 49354 26630 49356 26682
rect 49110 26628 49116 26630
rect 49172 26628 49196 26630
rect 49252 26628 49276 26630
rect 49332 26628 49356 26630
rect 49412 26628 49418 26630
rect 49110 26608 49418 26628
rect 46572 26580 46624 26586
rect 46572 26522 46624 26528
rect 46480 26036 46532 26042
rect 46480 25978 46532 25984
rect 46294 24576 46350 24585
rect 46294 24511 46350 24520
rect 46204 21344 46256 21350
rect 46204 21286 46256 21292
rect 46216 20806 46244 21286
rect 46020 20800 46072 20806
rect 46020 20742 46072 20748
rect 46204 20800 46256 20806
rect 46204 20742 46256 20748
rect 46032 20262 46060 20742
rect 46020 20256 46072 20262
rect 46020 20198 46072 20204
rect 45560 19712 45612 19718
rect 45560 19654 45612 19660
rect 45652 18624 45704 18630
rect 45650 18592 45652 18601
rect 45704 18592 45706 18601
rect 45650 18527 45706 18536
rect 45560 18420 45612 18426
rect 45560 18362 45612 18368
rect 45572 18154 45600 18362
rect 45560 18148 45612 18154
rect 45560 18090 45612 18096
rect 46032 17649 46060 20198
rect 46216 19854 46244 20742
rect 46204 19848 46256 19854
rect 46204 19790 46256 19796
rect 46308 19718 46336 24511
rect 46480 21140 46532 21146
rect 46480 21082 46532 21088
rect 46492 20602 46520 21082
rect 46480 20596 46532 20602
rect 46480 20538 46532 20544
rect 46492 20058 46520 20538
rect 46480 20052 46532 20058
rect 46480 19994 46532 20000
rect 46112 19712 46164 19718
rect 46112 19654 46164 19660
rect 46296 19712 46348 19718
rect 46296 19654 46348 19660
rect 46124 19156 46152 19654
rect 46204 19168 46256 19174
rect 46124 19128 46204 19156
rect 46204 19110 46256 19116
rect 46110 18456 46166 18465
rect 46110 18391 46112 18400
rect 46164 18391 46166 18400
rect 46112 18362 46164 18368
rect 46216 18290 46244 19110
rect 46308 18698 46336 19654
rect 46480 19508 46532 19514
rect 46480 19450 46532 19456
rect 46296 18692 46348 18698
rect 46296 18634 46348 18640
rect 46204 18284 46256 18290
rect 46204 18226 46256 18232
rect 46018 17640 46074 17649
rect 46018 17575 46074 17584
rect 46032 17270 46060 17575
rect 46020 17264 46072 17270
rect 46020 17206 46072 17212
rect 46204 17196 46256 17202
rect 46204 17138 46256 17144
rect 45652 16992 45704 16998
rect 45652 16934 45704 16940
rect 45558 15872 45614 15881
rect 45558 15807 45614 15816
rect 45572 15706 45600 15807
rect 45560 15700 45612 15706
rect 45560 15642 45612 15648
rect 45560 14272 45612 14278
rect 45560 14214 45612 14220
rect 45572 13734 45600 14214
rect 45560 13728 45612 13734
rect 45560 13670 45612 13676
rect 45572 13462 45600 13670
rect 45560 13456 45612 13462
rect 45560 13398 45612 13404
rect 45560 12096 45612 12102
rect 45560 12038 45612 12044
rect 45572 8838 45600 12038
rect 45560 8832 45612 8838
rect 45560 8774 45612 8780
rect 45664 6798 45692 16934
rect 45744 16788 45796 16794
rect 45744 16730 45796 16736
rect 45756 16028 45784 16730
rect 45836 16448 45888 16454
rect 45836 16390 45888 16396
rect 45848 16182 45876 16390
rect 45836 16176 45888 16182
rect 45836 16118 45888 16124
rect 45756 16000 45876 16028
rect 45744 15904 45796 15910
rect 45744 15846 45796 15852
rect 45756 14006 45784 15846
rect 45744 14000 45796 14006
rect 45744 13942 45796 13948
rect 45848 10577 45876 16000
rect 46020 15904 46072 15910
rect 46018 15872 46020 15881
rect 46072 15872 46074 15881
rect 46018 15807 46074 15816
rect 46216 14550 46244 17138
rect 46204 14544 46256 14550
rect 46204 14486 46256 14492
rect 45928 14272 45980 14278
rect 45928 14214 45980 14220
rect 45940 12442 45968 14214
rect 46112 13524 46164 13530
rect 46112 13466 46164 13472
rect 45928 12436 45980 12442
rect 45928 12378 45980 12384
rect 46124 12102 46152 13466
rect 46216 13394 46244 14486
rect 46204 13388 46256 13394
rect 46204 13330 46256 13336
rect 46112 12096 46164 12102
rect 46112 12038 46164 12044
rect 46308 11150 46336 18634
rect 46492 17882 46520 19450
rect 46584 18442 46612 26522
rect 56612 25702 56640 26930
rect 58084 26586 58112 27338
rect 58072 26580 58124 26586
rect 58072 26522 58124 26528
rect 58164 25900 58216 25906
rect 58164 25842 58216 25848
rect 57888 25764 57940 25770
rect 57888 25706 57940 25712
rect 56600 25696 56652 25702
rect 56600 25638 56652 25644
rect 49110 25596 49418 25616
rect 49110 25594 49116 25596
rect 49172 25594 49196 25596
rect 49252 25594 49276 25596
rect 49332 25594 49356 25596
rect 49412 25594 49418 25596
rect 49172 25542 49174 25594
rect 49354 25542 49356 25594
rect 49110 25540 49116 25542
rect 49172 25540 49196 25542
rect 49252 25540 49276 25542
rect 49332 25540 49356 25542
rect 49412 25540 49418 25542
rect 49110 25520 49418 25540
rect 46940 25492 46992 25498
rect 46940 25434 46992 25440
rect 46664 20052 46716 20058
rect 46664 19994 46716 20000
rect 46676 19514 46704 19994
rect 46952 19922 46980 25434
rect 49110 24508 49418 24528
rect 49110 24506 49116 24508
rect 49172 24506 49196 24508
rect 49252 24506 49276 24508
rect 49332 24506 49356 24508
rect 49412 24506 49418 24508
rect 49172 24454 49174 24506
rect 49354 24454 49356 24506
rect 49110 24452 49116 24454
rect 49172 24452 49196 24454
rect 49252 24452 49276 24454
rect 49332 24452 49356 24454
rect 49412 24452 49418 24454
rect 49110 24432 49418 24452
rect 49700 24132 49752 24138
rect 49700 24074 49752 24080
rect 49712 23730 49740 24074
rect 49700 23724 49752 23730
rect 49700 23666 49752 23672
rect 49110 23420 49418 23440
rect 49110 23418 49116 23420
rect 49172 23418 49196 23420
rect 49252 23418 49276 23420
rect 49332 23418 49356 23420
rect 49412 23418 49418 23420
rect 49172 23366 49174 23418
rect 49354 23366 49356 23418
rect 49110 23364 49116 23366
rect 49172 23364 49196 23366
rect 49252 23364 49276 23366
rect 49332 23364 49356 23366
rect 49412 23364 49418 23366
rect 49110 23344 49418 23364
rect 48778 22536 48834 22545
rect 48778 22471 48834 22480
rect 48688 22160 48740 22166
rect 48688 22102 48740 22108
rect 47860 21956 47912 21962
rect 47860 21898 47912 21904
rect 47872 20942 47900 21898
rect 47860 20936 47912 20942
rect 47860 20878 47912 20884
rect 46940 19916 46992 19922
rect 46940 19858 46992 19864
rect 46664 19508 46716 19514
rect 46664 19450 46716 19456
rect 46676 18902 46704 19450
rect 46664 18896 46716 18902
rect 46664 18838 46716 18844
rect 46584 18414 46704 18442
rect 46952 18426 46980 19858
rect 47768 19712 47820 19718
rect 47766 19680 47768 19689
rect 47820 19680 47822 19689
rect 47766 19615 47822 19624
rect 47872 18902 47900 20878
rect 48502 19816 48558 19825
rect 48502 19751 48558 19760
rect 47860 18896 47912 18902
rect 47860 18838 47912 18844
rect 48410 18592 48466 18601
rect 48410 18527 48466 18536
rect 46572 18284 46624 18290
rect 46572 18226 46624 18232
rect 46480 17876 46532 17882
rect 46480 17818 46532 17824
rect 46480 17672 46532 17678
rect 46584 17626 46612 18226
rect 46676 17678 46704 18414
rect 46940 18420 46992 18426
rect 46940 18362 46992 18368
rect 48318 18320 48374 18329
rect 48318 18255 48320 18264
rect 48372 18255 48374 18264
rect 48320 18226 48372 18232
rect 48228 17740 48280 17746
rect 48228 17682 48280 17688
rect 46532 17620 46612 17626
rect 46480 17614 46612 17620
rect 46664 17672 46716 17678
rect 46664 17614 46716 17620
rect 46492 17598 46612 17614
rect 46480 16992 46532 16998
rect 46480 16934 46532 16940
rect 46492 16697 46520 16934
rect 46478 16688 46534 16697
rect 46478 16623 46534 16632
rect 46388 16040 46440 16046
rect 46388 15982 46440 15988
rect 46400 15366 46428 15982
rect 46388 15360 46440 15366
rect 46388 15302 46440 15308
rect 46400 15162 46428 15302
rect 46388 15156 46440 15162
rect 46388 15098 46440 15104
rect 46480 15156 46532 15162
rect 46480 15098 46532 15104
rect 46492 14006 46520 15098
rect 46584 14414 46612 17598
rect 46676 15094 46704 17614
rect 48240 17542 48268 17682
rect 47032 17536 47084 17542
rect 48228 17536 48280 17542
rect 47032 17478 47084 17484
rect 47122 17504 47178 17513
rect 47044 17338 47072 17478
rect 47122 17439 47178 17448
rect 48134 17504 48190 17513
rect 48228 17478 48280 17484
rect 48134 17439 48190 17448
rect 47032 17332 47084 17338
rect 47032 17274 47084 17280
rect 47030 16824 47086 16833
rect 47030 16759 47086 16768
rect 46664 15088 46716 15094
rect 46940 15088 46992 15094
rect 46664 15030 46716 15036
rect 46938 15056 46940 15065
rect 46992 15056 46994 15065
rect 46938 14991 46994 15000
rect 46572 14408 46624 14414
rect 46572 14350 46624 14356
rect 46480 14000 46532 14006
rect 46480 13942 46532 13948
rect 46492 13530 46520 13942
rect 46480 13524 46532 13530
rect 46480 13466 46532 13472
rect 47044 12434 47072 16759
rect 46952 12406 47072 12434
rect 46296 11144 46348 11150
rect 46296 11086 46348 11092
rect 45834 10568 45890 10577
rect 45834 10503 45890 10512
rect 46204 8832 46256 8838
rect 46204 8774 46256 8780
rect 45652 6792 45704 6798
rect 45652 6734 45704 6740
rect 46216 2378 46244 8774
rect 46952 2582 46980 12406
rect 47136 11778 47164 17439
rect 48148 17338 48176 17439
rect 48136 17332 48188 17338
rect 48136 17274 48188 17280
rect 47584 16584 47636 16590
rect 47584 16526 47636 16532
rect 47306 16280 47362 16289
rect 47596 16250 47624 16526
rect 48134 16280 48190 16289
rect 47306 16215 47362 16224
rect 47584 16244 47636 16250
rect 47214 15600 47270 15609
rect 47214 15535 47270 15544
rect 47044 11750 47164 11778
rect 47044 4049 47072 11750
rect 47228 11642 47256 15535
rect 47136 11614 47256 11642
rect 47136 4146 47164 11614
rect 47320 6914 47348 16215
rect 48134 16215 48190 16224
rect 47584 16186 47636 16192
rect 48148 16182 48176 16215
rect 48136 16176 48188 16182
rect 48136 16118 48188 16124
rect 47584 15700 47636 15706
rect 47584 15642 47636 15648
rect 47596 15162 47624 15642
rect 47584 15156 47636 15162
rect 47584 15098 47636 15104
rect 48136 14816 48188 14822
rect 48136 14758 48188 14764
rect 48148 14346 48176 14758
rect 48136 14340 48188 14346
rect 48136 14282 48188 14288
rect 48240 12434 48268 17478
rect 48318 16416 48374 16425
rect 48318 16351 48374 16360
rect 48332 16114 48360 16351
rect 48320 16108 48372 16114
rect 48320 16050 48372 16056
rect 48320 15360 48372 15366
rect 48320 15302 48372 15308
rect 48332 14482 48360 15302
rect 48320 14476 48372 14482
rect 48320 14418 48372 14424
rect 47228 6886 47348 6914
rect 48148 12406 48268 12434
rect 47124 4140 47176 4146
rect 47124 4082 47176 4088
rect 47030 4040 47086 4049
rect 47030 3975 47086 3984
rect 47228 3641 47256 6886
rect 48148 6225 48176 12406
rect 48134 6216 48190 6225
rect 48134 6151 48190 6160
rect 47214 3632 47270 3641
rect 47214 3567 47270 3576
rect 46940 2576 46992 2582
rect 46940 2518 46992 2524
rect 46204 2372 46256 2378
rect 46204 2314 46256 2320
rect 45468 2032 45520 2038
rect 45468 1974 45520 1980
rect 48424 1970 48452 18527
rect 48516 4010 48544 19751
rect 48700 19310 48728 22102
rect 48688 19304 48740 19310
rect 48688 19246 48740 19252
rect 48688 18828 48740 18834
rect 48688 18770 48740 18776
rect 48700 18426 48728 18770
rect 48688 18420 48740 18426
rect 48688 18362 48740 18368
rect 48700 17882 48728 18362
rect 48688 17876 48740 17882
rect 48688 17818 48740 17824
rect 48596 17264 48648 17270
rect 48596 17206 48648 17212
rect 48608 16454 48636 17206
rect 48700 16794 48728 17818
rect 48688 16788 48740 16794
rect 48688 16730 48740 16736
rect 48596 16448 48648 16454
rect 48596 16390 48648 16396
rect 48608 15366 48636 16390
rect 48700 16250 48728 16730
rect 48688 16244 48740 16250
rect 48688 16186 48740 16192
rect 48700 15706 48728 16186
rect 48688 15700 48740 15706
rect 48688 15642 48740 15648
rect 48596 15360 48648 15366
rect 48596 15302 48648 15308
rect 48504 4004 48556 4010
rect 48504 3946 48556 3952
rect 48792 2514 48820 22471
rect 49110 22332 49418 22352
rect 49110 22330 49116 22332
rect 49172 22330 49196 22332
rect 49252 22330 49276 22332
rect 49332 22330 49356 22332
rect 49412 22330 49418 22332
rect 49172 22278 49174 22330
rect 49354 22278 49356 22330
rect 49110 22276 49116 22278
rect 49172 22276 49196 22278
rect 49252 22276 49276 22278
rect 49332 22276 49356 22278
rect 49412 22276 49418 22278
rect 49110 22256 49418 22276
rect 49110 21244 49418 21264
rect 49110 21242 49116 21244
rect 49172 21242 49196 21244
rect 49252 21242 49276 21244
rect 49332 21242 49356 21244
rect 49412 21242 49418 21244
rect 49172 21190 49174 21242
rect 49354 21190 49356 21242
rect 49110 21188 49116 21190
rect 49172 21188 49196 21190
rect 49252 21188 49276 21190
rect 49332 21188 49356 21190
rect 49412 21188 49418 21190
rect 49110 21168 49418 21188
rect 49110 20156 49418 20176
rect 49110 20154 49116 20156
rect 49172 20154 49196 20156
rect 49252 20154 49276 20156
rect 49332 20154 49356 20156
rect 49412 20154 49418 20156
rect 49172 20102 49174 20154
rect 49354 20102 49356 20154
rect 49110 20100 49116 20102
rect 49172 20100 49196 20102
rect 49252 20100 49276 20102
rect 49332 20100 49356 20102
rect 49412 20100 49418 20102
rect 49110 20080 49418 20100
rect 48872 19440 48924 19446
rect 48872 19382 48924 19388
rect 48884 5681 48912 19382
rect 49712 19242 49740 23666
rect 57900 21418 57928 25706
rect 58176 25673 58204 25842
rect 58162 25664 58218 25673
rect 58162 25599 58218 25608
rect 58176 25498 58204 25599
rect 58164 25492 58216 25498
rect 58164 25434 58216 25440
rect 58164 24200 58216 24206
rect 58164 24142 58216 24148
rect 58176 23905 58204 24142
rect 58162 23896 58218 23905
rect 58162 23831 58164 23840
rect 58216 23831 58218 23840
rect 58164 23802 58216 23808
rect 58162 22128 58218 22137
rect 58162 22063 58218 22072
rect 58176 22030 58204 22063
rect 58164 22024 58216 22030
rect 58164 21966 58216 21972
rect 58176 21690 58204 21966
rect 58164 21684 58216 21690
rect 58164 21626 58216 21632
rect 57888 21412 57940 21418
rect 57888 21354 57940 21360
rect 58162 20360 58218 20369
rect 58162 20295 58218 20304
rect 58176 19854 58204 20295
rect 58164 19848 58216 19854
rect 58164 19790 58216 19796
rect 51724 19712 51776 19718
rect 51724 19654 51776 19660
rect 49700 19236 49752 19242
rect 49700 19178 49752 19184
rect 49110 19068 49418 19088
rect 49110 19066 49116 19068
rect 49172 19066 49196 19068
rect 49252 19066 49276 19068
rect 49332 19066 49356 19068
rect 49412 19066 49418 19068
rect 49172 19014 49174 19066
rect 49354 19014 49356 19066
rect 49110 19012 49116 19014
rect 49172 19012 49196 19014
rect 49252 19012 49276 19014
rect 49332 19012 49356 19014
rect 49412 19012 49418 19014
rect 49110 18992 49418 19012
rect 49608 18080 49660 18086
rect 49608 18022 49660 18028
rect 49110 17980 49418 18000
rect 49110 17978 49116 17980
rect 49172 17978 49196 17980
rect 49252 17978 49276 17980
rect 49332 17978 49356 17980
rect 49412 17978 49418 17980
rect 49172 17926 49174 17978
rect 49354 17926 49356 17978
rect 49110 17924 49116 17926
rect 49172 17924 49196 17926
rect 49252 17924 49276 17926
rect 49332 17924 49356 17926
rect 49412 17924 49418 17926
rect 49110 17904 49418 17924
rect 49620 17270 49648 18022
rect 50160 17536 50212 17542
rect 50160 17478 50212 17484
rect 49608 17264 49660 17270
rect 50172 17241 50200 17478
rect 49608 17206 49660 17212
rect 50158 17232 50214 17241
rect 48964 16992 49016 16998
rect 48964 16934 49016 16940
rect 48976 16522 49004 16934
rect 49110 16892 49418 16912
rect 49110 16890 49116 16892
rect 49172 16890 49196 16892
rect 49252 16890 49276 16892
rect 49332 16890 49356 16892
rect 49412 16890 49418 16892
rect 49172 16838 49174 16890
rect 49354 16838 49356 16890
rect 49110 16836 49116 16838
rect 49172 16836 49196 16838
rect 49252 16836 49276 16838
rect 49332 16836 49356 16838
rect 49412 16836 49418 16838
rect 49110 16816 49418 16836
rect 49620 16794 49648 17206
rect 50158 17167 50214 17176
rect 49608 16788 49660 16794
rect 49608 16730 49660 16736
rect 48964 16516 49016 16522
rect 48964 16458 49016 16464
rect 49790 16144 49846 16153
rect 49790 16079 49792 16088
rect 49844 16079 49846 16088
rect 49792 16050 49844 16056
rect 49110 15804 49418 15824
rect 49110 15802 49116 15804
rect 49172 15802 49196 15804
rect 49252 15802 49276 15804
rect 49332 15802 49356 15804
rect 49412 15802 49418 15804
rect 49172 15750 49174 15802
rect 49354 15750 49356 15802
rect 49110 15748 49116 15750
rect 49172 15748 49196 15750
rect 49252 15748 49276 15750
rect 49332 15748 49356 15750
rect 49412 15748 49418 15750
rect 49110 15728 49418 15748
rect 49110 14716 49418 14736
rect 49110 14714 49116 14716
rect 49172 14714 49196 14716
rect 49252 14714 49276 14716
rect 49332 14714 49356 14716
rect 49412 14714 49418 14716
rect 49172 14662 49174 14714
rect 49354 14662 49356 14714
rect 49110 14660 49116 14662
rect 49172 14660 49196 14662
rect 49252 14660 49276 14662
rect 49332 14660 49356 14662
rect 49412 14660 49418 14662
rect 49110 14640 49418 14660
rect 49110 13628 49418 13648
rect 49110 13626 49116 13628
rect 49172 13626 49196 13628
rect 49252 13626 49276 13628
rect 49332 13626 49356 13628
rect 49412 13626 49418 13628
rect 49172 13574 49174 13626
rect 49354 13574 49356 13626
rect 49110 13572 49116 13574
rect 49172 13572 49196 13574
rect 49252 13572 49276 13574
rect 49332 13572 49356 13574
rect 49412 13572 49418 13574
rect 49110 13552 49418 13572
rect 49110 12540 49418 12560
rect 49110 12538 49116 12540
rect 49172 12538 49196 12540
rect 49252 12538 49276 12540
rect 49332 12538 49356 12540
rect 49412 12538 49418 12540
rect 49172 12486 49174 12538
rect 49354 12486 49356 12538
rect 49110 12484 49116 12486
rect 49172 12484 49196 12486
rect 49252 12484 49276 12486
rect 49332 12484 49356 12486
rect 49412 12484 49418 12486
rect 49110 12464 49418 12484
rect 49110 11452 49418 11472
rect 49110 11450 49116 11452
rect 49172 11450 49196 11452
rect 49252 11450 49276 11452
rect 49332 11450 49356 11452
rect 49412 11450 49418 11452
rect 49172 11398 49174 11450
rect 49354 11398 49356 11450
rect 49110 11396 49116 11398
rect 49172 11396 49196 11398
rect 49252 11396 49276 11398
rect 49332 11396 49356 11398
rect 49412 11396 49418 11398
rect 49110 11376 49418 11396
rect 49110 10364 49418 10384
rect 49110 10362 49116 10364
rect 49172 10362 49196 10364
rect 49252 10362 49276 10364
rect 49332 10362 49356 10364
rect 49412 10362 49418 10364
rect 49172 10310 49174 10362
rect 49354 10310 49356 10362
rect 49110 10308 49116 10310
rect 49172 10308 49196 10310
rect 49252 10308 49276 10310
rect 49332 10308 49356 10310
rect 49412 10308 49418 10310
rect 49110 10288 49418 10308
rect 49110 9276 49418 9296
rect 49110 9274 49116 9276
rect 49172 9274 49196 9276
rect 49252 9274 49276 9276
rect 49332 9274 49356 9276
rect 49412 9274 49418 9276
rect 49172 9222 49174 9274
rect 49354 9222 49356 9274
rect 49110 9220 49116 9222
rect 49172 9220 49196 9222
rect 49252 9220 49276 9222
rect 49332 9220 49356 9222
rect 49412 9220 49418 9222
rect 49110 9200 49418 9220
rect 49110 8188 49418 8208
rect 49110 8186 49116 8188
rect 49172 8186 49196 8188
rect 49252 8186 49276 8188
rect 49332 8186 49356 8188
rect 49412 8186 49418 8188
rect 49172 8134 49174 8186
rect 49354 8134 49356 8186
rect 49110 8132 49116 8134
rect 49172 8132 49196 8134
rect 49252 8132 49276 8134
rect 49332 8132 49356 8134
rect 49412 8132 49418 8134
rect 49110 8112 49418 8132
rect 51736 7954 51764 19654
rect 58176 19514 58204 19790
rect 58164 19508 58216 19514
rect 58164 19450 58216 19456
rect 58164 18760 58216 18766
rect 58164 18702 58216 18708
rect 57888 18692 57940 18698
rect 57888 18634 57940 18640
rect 57900 18222 57928 18634
rect 58176 18601 58204 18702
rect 58162 18592 58218 18601
rect 58162 18527 58218 18536
rect 58176 18426 58204 18527
rect 58164 18420 58216 18426
rect 58164 18362 58216 18368
rect 57888 18216 57940 18222
rect 57888 18158 57940 18164
rect 58162 16824 58218 16833
rect 58162 16759 58218 16768
rect 58176 16590 58204 16759
rect 58164 16584 58216 16590
rect 58164 16526 58216 16532
rect 58176 16250 58204 16526
rect 58164 16244 58216 16250
rect 58164 16186 58216 16192
rect 58164 15496 58216 15502
rect 58164 15438 58216 15444
rect 57888 15428 57940 15434
rect 57888 15370 57940 15376
rect 57900 14521 57928 15370
rect 58176 15094 58204 15438
rect 58164 15088 58216 15094
rect 58162 15056 58164 15065
rect 58216 15056 58218 15065
rect 58162 14991 58218 15000
rect 57886 14512 57942 14521
rect 57886 14447 57942 14456
rect 58164 13320 58216 13326
rect 58162 13288 58164 13297
rect 58216 13288 58218 13297
rect 57888 13252 57940 13258
rect 58162 13223 58218 13232
rect 57888 13194 57940 13200
rect 57900 12714 57928 13194
rect 58176 12986 58204 13223
rect 58164 12980 58216 12986
rect 58164 12922 58216 12928
rect 57888 12708 57940 12714
rect 57888 12650 57940 12656
rect 58162 11520 58218 11529
rect 58162 11455 58218 11464
rect 58176 11150 58204 11455
rect 58164 11144 58216 11150
rect 58164 11086 58216 11092
rect 58176 10810 58204 11086
rect 58164 10804 58216 10810
rect 58164 10746 58216 10752
rect 58164 10056 58216 10062
rect 58164 9998 58216 10004
rect 58176 9761 58204 9998
rect 58162 9752 58218 9761
rect 58162 9687 58164 9696
rect 58216 9687 58218 9696
rect 58164 9658 58216 9664
rect 58162 7984 58218 7993
rect 51724 7948 51776 7954
rect 58162 7919 58218 7928
rect 51724 7890 51776 7896
rect 58176 7886 58204 7919
rect 58164 7880 58216 7886
rect 58164 7822 58216 7828
rect 58176 7546 58204 7822
rect 58164 7540 58216 7546
rect 58164 7482 58216 7488
rect 49110 7100 49418 7120
rect 49110 7098 49116 7100
rect 49172 7098 49196 7100
rect 49252 7098 49276 7100
rect 49332 7098 49356 7100
rect 49412 7098 49418 7100
rect 49172 7046 49174 7098
rect 49354 7046 49356 7098
rect 49110 7044 49116 7046
rect 49172 7044 49196 7046
rect 49252 7044 49276 7046
rect 49332 7044 49356 7046
rect 49412 7044 49418 7046
rect 49110 7024 49418 7044
rect 58162 6216 58218 6225
rect 58162 6151 58218 6160
rect 49110 6012 49418 6032
rect 49110 6010 49116 6012
rect 49172 6010 49196 6012
rect 49252 6010 49276 6012
rect 49332 6010 49356 6012
rect 49412 6010 49418 6012
rect 49172 5958 49174 6010
rect 49354 5958 49356 6010
rect 49110 5956 49116 5958
rect 49172 5956 49196 5958
rect 49252 5956 49276 5958
rect 49332 5956 49356 5958
rect 49412 5956 49418 5958
rect 49110 5936 49418 5956
rect 58176 5710 58204 6151
rect 58164 5704 58216 5710
rect 48870 5672 48926 5681
rect 58164 5646 58216 5652
rect 48870 5607 48926 5616
rect 58176 5370 58204 5646
rect 58164 5364 58216 5370
rect 58164 5306 58216 5312
rect 49110 4924 49418 4944
rect 49110 4922 49116 4924
rect 49172 4922 49196 4924
rect 49252 4922 49276 4924
rect 49332 4922 49356 4924
rect 49412 4922 49418 4924
rect 49172 4870 49174 4922
rect 49354 4870 49356 4922
rect 49110 4868 49116 4870
rect 49172 4868 49196 4870
rect 49252 4868 49276 4870
rect 49332 4868 49356 4870
rect 49412 4868 49418 4870
rect 49110 4848 49418 4868
rect 58164 4616 58216 4622
rect 58164 4558 58216 4564
rect 58176 4457 58204 4558
rect 58162 4448 58218 4457
rect 58162 4383 58218 4392
rect 58176 4282 58204 4383
rect 58164 4276 58216 4282
rect 58164 4218 58216 4224
rect 49110 3836 49418 3856
rect 49110 3834 49116 3836
rect 49172 3834 49196 3836
rect 49252 3834 49276 3836
rect 49332 3834 49356 3836
rect 49412 3834 49418 3836
rect 49172 3782 49174 3834
rect 49354 3782 49356 3834
rect 49110 3780 49116 3782
rect 49172 3780 49196 3782
rect 49252 3780 49276 3782
rect 49332 3780 49356 3782
rect 49412 3780 49418 3782
rect 49110 3760 49418 3780
rect 49110 2748 49418 2768
rect 49110 2746 49116 2748
rect 49172 2746 49196 2748
rect 49252 2746 49276 2748
rect 49332 2746 49356 2748
rect 49412 2746 49418 2748
rect 49172 2694 49174 2746
rect 49354 2694 49356 2746
rect 49110 2692 49116 2694
rect 49172 2692 49196 2694
rect 49252 2692 49276 2694
rect 49332 2692 49356 2694
rect 49412 2692 49418 2694
rect 49110 2672 49418 2692
rect 56506 2680 56562 2689
rect 56506 2615 56508 2624
rect 56560 2615 56562 2624
rect 56508 2586 56560 2592
rect 48780 2508 48832 2514
rect 48780 2450 48832 2456
rect 53932 2304 53984 2310
rect 53932 2246 53984 2252
rect 57888 2304 57940 2310
rect 57888 2246 57940 2252
rect 48412 1964 48464 1970
rect 48412 1906 48464 1912
rect 53944 800 53972 2246
rect 57900 921 57928 2246
rect 57886 912 57942 921
rect 57886 847 57942 856
rect 1490 776 1546 785
rect 1490 711 1546 720
rect 5998 0 6054 800
rect 17958 0 18014 800
rect 29918 0 29974 800
rect 41970 0 42026 800
rect 53930 0 53986 800
<< via2 >>
rect 18326 29552 18382 29608
rect 1398 29144 1454 29200
rect 1490 27548 1492 27568
rect 1492 27548 1544 27568
rect 1544 27548 1546 27568
rect 1490 27512 1546 27548
rect 10588 27770 10644 27772
rect 10668 27770 10724 27772
rect 10748 27770 10804 27772
rect 10828 27770 10884 27772
rect 10588 27718 10634 27770
rect 10634 27718 10644 27770
rect 10668 27718 10698 27770
rect 10698 27718 10710 27770
rect 10710 27718 10724 27770
rect 10748 27718 10762 27770
rect 10762 27718 10774 27770
rect 10774 27718 10804 27770
rect 10828 27718 10838 27770
rect 10838 27718 10884 27770
rect 10588 27716 10644 27718
rect 10668 27716 10724 27718
rect 10748 27716 10804 27718
rect 10828 27716 10884 27718
rect 14830 28736 14886 28792
rect 14738 28600 14794 28656
rect 14554 28328 14610 28384
rect 10588 26682 10644 26684
rect 10668 26682 10724 26684
rect 10748 26682 10804 26684
rect 10828 26682 10884 26684
rect 10588 26630 10634 26682
rect 10634 26630 10644 26682
rect 10668 26630 10698 26682
rect 10698 26630 10710 26682
rect 10710 26630 10724 26682
rect 10748 26630 10762 26682
rect 10762 26630 10774 26682
rect 10774 26630 10804 26682
rect 10828 26630 10838 26682
rect 10838 26630 10884 26682
rect 10588 26628 10644 26630
rect 10668 26628 10724 26630
rect 10748 26628 10804 26630
rect 10828 26628 10884 26630
rect 1490 26016 1546 26072
rect 1490 24384 1546 24440
rect 10588 25594 10644 25596
rect 10668 25594 10724 25596
rect 10748 25594 10804 25596
rect 10828 25594 10884 25596
rect 10588 25542 10634 25594
rect 10634 25542 10644 25594
rect 10668 25542 10698 25594
rect 10698 25542 10710 25594
rect 10710 25542 10724 25594
rect 10748 25542 10762 25594
rect 10762 25542 10774 25594
rect 10774 25542 10804 25594
rect 10828 25542 10838 25594
rect 10838 25542 10884 25594
rect 10588 25540 10644 25542
rect 10668 25540 10724 25542
rect 10748 25540 10804 25542
rect 10828 25540 10884 25542
rect 10588 24506 10644 24508
rect 10668 24506 10724 24508
rect 10748 24506 10804 24508
rect 10828 24506 10884 24508
rect 10588 24454 10634 24506
rect 10634 24454 10644 24506
rect 10668 24454 10698 24506
rect 10698 24454 10710 24506
rect 10710 24454 10724 24506
rect 10748 24454 10762 24506
rect 10762 24454 10774 24506
rect 10774 24454 10804 24506
rect 10828 24454 10838 24506
rect 10838 24454 10884 24506
rect 10588 24452 10644 24454
rect 10668 24452 10724 24454
rect 10748 24452 10804 24454
rect 10828 24452 10884 24454
rect 10588 23418 10644 23420
rect 10668 23418 10724 23420
rect 10748 23418 10804 23420
rect 10828 23418 10884 23420
rect 10588 23366 10634 23418
rect 10634 23366 10644 23418
rect 10668 23366 10698 23418
rect 10698 23366 10710 23418
rect 10710 23366 10724 23418
rect 10748 23366 10762 23418
rect 10762 23366 10774 23418
rect 10774 23366 10804 23418
rect 10828 23366 10838 23418
rect 10838 23366 10884 23418
rect 10588 23364 10644 23366
rect 10668 23364 10724 23366
rect 10748 23364 10804 23366
rect 10828 23364 10884 23366
rect 1490 22752 1546 22808
rect 10588 22330 10644 22332
rect 10668 22330 10724 22332
rect 10748 22330 10804 22332
rect 10828 22330 10884 22332
rect 10588 22278 10634 22330
rect 10634 22278 10644 22330
rect 10668 22278 10698 22330
rect 10698 22278 10710 22330
rect 10710 22278 10724 22330
rect 10748 22278 10762 22330
rect 10762 22278 10774 22330
rect 10774 22278 10804 22330
rect 10828 22278 10838 22330
rect 10838 22278 10884 22330
rect 10588 22276 10644 22278
rect 10668 22276 10724 22278
rect 10748 22276 10804 22278
rect 10828 22276 10884 22278
rect 1490 21292 1492 21312
rect 1492 21292 1544 21312
rect 1544 21292 1546 21312
rect 1490 21256 1546 21292
rect 10588 21242 10644 21244
rect 10668 21242 10724 21244
rect 10748 21242 10804 21244
rect 10828 21242 10884 21244
rect 10588 21190 10634 21242
rect 10634 21190 10644 21242
rect 10668 21190 10698 21242
rect 10698 21190 10710 21242
rect 10710 21190 10724 21242
rect 10748 21190 10762 21242
rect 10762 21190 10774 21242
rect 10774 21190 10804 21242
rect 10828 21190 10838 21242
rect 10838 21190 10884 21242
rect 10588 21188 10644 21190
rect 10668 21188 10724 21190
rect 10748 21188 10804 21190
rect 10828 21188 10884 21190
rect 10588 20154 10644 20156
rect 10668 20154 10724 20156
rect 10748 20154 10804 20156
rect 10828 20154 10884 20156
rect 10588 20102 10634 20154
rect 10634 20102 10644 20154
rect 10668 20102 10698 20154
rect 10698 20102 10710 20154
rect 10710 20102 10724 20154
rect 10748 20102 10762 20154
rect 10762 20102 10774 20154
rect 10774 20102 10804 20154
rect 10828 20102 10838 20154
rect 10838 20102 10884 20154
rect 10588 20100 10644 20102
rect 10668 20100 10724 20102
rect 10748 20100 10804 20102
rect 10828 20100 10884 20102
rect 1490 19660 1492 19680
rect 1492 19660 1544 19680
rect 1544 19660 1546 19680
rect 1490 19624 1546 19660
rect 13910 21936 13966 21992
rect 10588 19066 10644 19068
rect 10668 19066 10724 19068
rect 10748 19066 10804 19068
rect 10828 19066 10884 19068
rect 10588 19014 10634 19066
rect 10634 19014 10644 19066
rect 10668 19014 10698 19066
rect 10698 19014 10710 19066
rect 10710 19014 10724 19066
rect 10748 19014 10762 19066
rect 10762 19014 10774 19066
rect 10774 19014 10804 19066
rect 10828 19014 10838 19066
rect 10838 19014 10884 19066
rect 10588 19012 10644 19014
rect 10668 19012 10724 19014
rect 10748 19012 10804 19014
rect 10828 19012 10884 19014
rect 1490 18028 1492 18048
rect 1492 18028 1544 18048
rect 1544 18028 1546 18048
rect 1490 17992 1546 18028
rect 10588 17978 10644 17980
rect 10668 17978 10724 17980
rect 10748 17978 10804 17980
rect 10828 17978 10884 17980
rect 10588 17926 10634 17978
rect 10634 17926 10644 17978
rect 10668 17926 10698 17978
rect 10698 17926 10710 17978
rect 10710 17926 10724 17978
rect 10748 17926 10762 17978
rect 10762 17926 10774 17978
rect 10774 17926 10804 17978
rect 10828 17926 10838 17978
rect 10838 17926 10884 17978
rect 10588 17924 10644 17926
rect 10668 17924 10724 17926
rect 10748 17924 10804 17926
rect 10828 17924 10884 17926
rect 10588 16890 10644 16892
rect 10668 16890 10724 16892
rect 10748 16890 10804 16892
rect 10828 16890 10884 16892
rect 10588 16838 10634 16890
rect 10634 16838 10644 16890
rect 10668 16838 10698 16890
rect 10698 16838 10710 16890
rect 10710 16838 10724 16890
rect 10748 16838 10762 16890
rect 10762 16838 10774 16890
rect 10774 16838 10804 16890
rect 10828 16838 10838 16890
rect 10838 16838 10884 16890
rect 10588 16836 10644 16838
rect 10668 16836 10724 16838
rect 10748 16836 10804 16838
rect 10828 16836 10884 16838
rect 1490 16496 1546 16552
rect 10588 15802 10644 15804
rect 10668 15802 10724 15804
rect 10748 15802 10804 15804
rect 10828 15802 10884 15804
rect 10588 15750 10634 15802
rect 10634 15750 10644 15802
rect 10668 15750 10698 15802
rect 10698 15750 10710 15802
rect 10710 15750 10724 15802
rect 10748 15750 10762 15802
rect 10762 15750 10774 15802
rect 10774 15750 10804 15802
rect 10828 15750 10838 15802
rect 10838 15750 10884 15802
rect 10588 15748 10644 15750
rect 10668 15748 10724 15750
rect 10748 15748 10804 15750
rect 10828 15748 10884 15750
rect 1490 14884 1546 14920
rect 1490 14864 1492 14884
rect 1492 14864 1544 14884
rect 1544 14864 1546 14884
rect 10588 14714 10644 14716
rect 10668 14714 10724 14716
rect 10748 14714 10804 14716
rect 10828 14714 10884 14716
rect 10588 14662 10634 14714
rect 10634 14662 10644 14714
rect 10668 14662 10698 14714
rect 10698 14662 10710 14714
rect 10710 14662 10724 14714
rect 10748 14662 10762 14714
rect 10762 14662 10774 14714
rect 10774 14662 10804 14714
rect 10828 14662 10838 14714
rect 10838 14662 10884 14714
rect 10588 14660 10644 14662
rect 10668 14660 10724 14662
rect 10748 14660 10804 14662
rect 10828 14660 10884 14662
rect 10588 13626 10644 13628
rect 10668 13626 10724 13628
rect 10748 13626 10804 13628
rect 10828 13626 10884 13628
rect 10588 13574 10634 13626
rect 10634 13574 10644 13626
rect 10668 13574 10698 13626
rect 10698 13574 10710 13626
rect 10710 13574 10724 13626
rect 10748 13574 10762 13626
rect 10762 13574 10774 13626
rect 10774 13574 10804 13626
rect 10828 13574 10838 13626
rect 10838 13574 10884 13626
rect 10588 13572 10644 13574
rect 10668 13572 10724 13574
rect 10748 13572 10804 13574
rect 10828 13572 10884 13574
rect 14462 21528 14518 21584
rect 14278 19624 14334 19680
rect 14186 18828 14242 18864
rect 14186 18808 14188 18828
rect 14188 18808 14240 18828
rect 14240 18808 14242 18828
rect 14094 17720 14150 17776
rect 1490 13368 1546 13424
rect 10588 12538 10644 12540
rect 10668 12538 10724 12540
rect 10748 12538 10804 12540
rect 10828 12538 10884 12540
rect 10588 12486 10634 12538
rect 10634 12486 10644 12538
rect 10668 12486 10698 12538
rect 10698 12486 10710 12538
rect 10710 12486 10724 12538
rect 10748 12486 10762 12538
rect 10762 12486 10774 12538
rect 10774 12486 10804 12538
rect 10828 12486 10838 12538
rect 10838 12486 10884 12538
rect 10588 12484 10644 12486
rect 10668 12484 10724 12486
rect 10748 12484 10804 12486
rect 10828 12484 10884 12486
rect 14002 17312 14058 17368
rect 1490 11736 1546 11792
rect 10588 11450 10644 11452
rect 10668 11450 10724 11452
rect 10748 11450 10804 11452
rect 10828 11450 10884 11452
rect 10588 11398 10634 11450
rect 10634 11398 10644 11450
rect 10668 11398 10698 11450
rect 10698 11398 10710 11450
rect 10710 11398 10724 11450
rect 10748 11398 10762 11450
rect 10762 11398 10774 11450
rect 10774 11398 10804 11450
rect 10828 11398 10838 11450
rect 10838 11398 10884 11450
rect 10588 11396 10644 11398
rect 10668 11396 10724 11398
rect 10748 11396 10804 11398
rect 10828 11396 10884 11398
rect 10588 10362 10644 10364
rect 10668 10362 10724 10364
rect 10748 10362 10804 10364
rect 10828 10362 10884 10364
rect 10588 10310 10634 10362
rect 10634 10310 10644 10362
rect 10668 10310 10698 10362
rect 10698 10310 10710 10362
rect 10710 10310 10724 10362
rect 10748 10310 10762 10362
rect 10762 10310 10774 10362
rect 10774 10310 10804 10362
rect 10828 10310 10838 10362
rect 10838 10310 10884 10362
rect 10588 10308 10644 10310
rect 10668 10308 10724 10310
rect 10748 10308 10804 10310
rect 10828 10308 10884 10310
rect 1490 10104 1546 10160
rect 1490 8608 1546 8664
rect 10588 9274 10644 9276
rect 10668 9274 10724 9276
rect 10748 9274 10804 9276
rect 10828 9274 10884 9276
rect 10588 9222 10634 9274
rect 10634 9222 10644 9274
rect 10668 9222 10698 9274
rect 10698 9222 10710 9274
rect 10710 9222 10724 9274
rect 10748 9222 10762 9274
rect 10762 9222 10774 9274
rect 10774 9222 10804 9274
rect 10828 9222 10838 9274
rect 10838 9222 10884 9274
rect 10588 9220 10644 9222
rect 10668 9220 10724 9222
rect 10748 9220 10804 9222
rect 10828 9220 10884 9222
rect 10588 8186 10644 8188
rect 10668 8186 10724 8188
rect 10748 8186 10804 8188
rect 10828 8186 10884 8188
rect 10588 8134 10634 8186
rect 10634 8134 10644 8186
rect 10668 8134 10698 8186
rect 10698 8134 10710 8186
rect 10710 8134 10724 8186
rect 10748 8134 10762 8186
rect 10762 8134 10774 8186
rect 10774 8134 10804 8186
rect 10828 8134 10838 8186
rect 10838 8134 10884 8186
rect 10588 8132 10644 8134
rect 10668 8132 10724 8134
rect 10748 8132 10804 8134
rect 10828 8132 10884 8134
rect 10588 7098 10644 7100
rect 10668 7098 10724 7100
rect 10748 7098 10804 7100
rect 10828 7098 10884 7100
rect 10588 7046 10634 7098
rect 10634 7046 10644 7098
rect 10668 7046 10698 7098
rect 10698 7046 10710 7098
rect 10710 7046 10724 7098
rect 10748 7046 10762 7098
rect 10762 7046 10774 7098
rect 10774 7046 10804 7098
rect 10828 7046 10838 7098
rect 10838 7046 10884 7098
rect 10588 7044 10644 7046
rect 10668 7044 10724 7046
rect 10748 7044 10804 7046
rect 10828 7044 10884 7046
rect 1490 6976 1546 7032
rect 10588 6010 10644 6012
rect 10668 6010 10724 6012
rect 10748 6010 10804 6012
rect 10828 6010 10884 6012
rect 10588 5958 10634 6010
rect 10634 5958 10644 6010
rect 10668 5958 10698 6010
rect 10698 5958 10710 6010
rect 10710 5958 10724 6010
rect 10748 5958 10762 6010
rect 10762 5958 10774 6010
rect 10774 5958 10804 6010
rect 10828 5958 10838 6010
rect 10838 5958 10884 6010
rect 10588 5956 10644 5958
rect 10668 5956 10724 5958
rect 10748 5956 10804 5958
rect 10828 5956 10884 5958
rect 1490 5344 1546 5400
rect 1490 3884 1492 3904
rect 1492 3884 1544 3904
rect 1544 3884 1546 3904
rect 1490 3848 1546 3884
rect 10588 4922 10644 4924
rect 10668 4922 10724 4924
rect 10748 4922 10804 4924
rect 10828 4922 10884 4924
rect 10588 4870 10634 4922
rect 10634 4870 10644 4922
rect 10668 4870 10698 4922
rect 10698 4870 10710 4922
rect 10710 4870 10724 4922
rect 10748 4870 10762 4922
rect 10762 4870 10774 4922
rect 10774 4870 10804 4922
rect 10828 4870 10838 4922
rect 10838 4870 10884 4922
rect 10588 4868 10644 4870
rect 10668 4868 10724 4870
rect 10748 4868 10804 4870
rect 10828 4868 10884 4870
rect 10588 3834 10644 3836
rect 10668 3834 10724 3836
rect 10748 3834 10804 3836
rect 10828 3834 10884 3836
rect 10588 3782 10634 3834
rect 10634 3782 10644 3834
rect 10668 3782 10698 3834
rect 10698 3782 10710 3834
rect 10710 3782 10724 3834
rect 10748 3782 10762 3834
rect 10762 3782 10774 3834
rect 10774 3782 10804 3834
rect 10828 3782 10838 3834
rect 10838 3782 10884 3834
rect 10588 3780 10644 3782
rect 10668 3780 10724 3782
rect 10748 3780 10804 3782
rect 10828 3780 10884 3782
rect 10588 2746 10644 2748
rect 10668 2746 10724 2748
rect 10748 2746 10804 2748
rect 10828 2746 10884 2748
rect 10588 2694 10634 2746
rect 10634 2694 10644 2746
rect 10668 2694 10698 2746
rect 10698 2694 10710 2746
rect 10710 2694 10724 2746
rect 10748 2694 10762 2746
rect 10762 2694 10774 2746
rect 10774 2694 10804 2746
rect 10828 2694 10838 2746
rect 10838 2694 10884 2746
rect 10588 2692 10644 2694
rect 10668 2692 10724 2694
rect 10748 2692 10804 2694
rect 10828 2692 10884 2694
rect 14370 4664 14426 4720
rect 1398 2216 1454 2272
rect 15198 25472 15254 25528
rect 14830 19352 14886 19408
rect 14738 17312 14794 17368
rect 17130 25336 17186 25392
rect 16578 24792 16634 24848
rect 16486 23432 16542 23488
rect 15566 20324 15622 20360
rect 15566 20304 15568 20324
rect 15568 20304 15620 20324
rect 15620 20304 15622 20324
rect 15014 18672 15070 18728
rect 15014 18400 15070 18456
rect 16210 19080 16266 19136
rect 14922 16360 14978 16416
rect 15382 16788 15438 16824
rect 15382 16768 15384 16788
rect 15384 16768 15436 16788
rect 15436 16768 15438 16788
rect 15290 16632 15346 16688
rect 15106 15852 15108 15872
rect 15108 15852 15160 15872
rect 15160 15852 15162 15872
rect 15106 15816 15162 15852
rect 15198 15408 15254 15464
rect 15382 15136 15438 15192
rect 15934 17992 15990 18048
rect 15658 17448 15714 17504
rect 15842 16532 15844 16552
rect 15844 16532 15896 16552
rect 15896 16532 15898 16552
rect 15842 16496 15898 16532
rect 15566 16124 15568 16144
rect 15568 16124 15620 16144
rect 15620 16124 15622 16144
rect 15566 16088 15622 16124
rect 15106 14320 15162 14376
rect 14830 5072 14886 5128
rect 15106 4528 15162 4584
rect 15658 15952 15714 16008
rect 16118 17040 16174 17096
rect 16946 23296 17002 23352
rect 16670 21256 16726 21312
rect 16486 18944 16542 19000
rect 16578 18264 16634 18320
rect 16762 19236 16818 19272
rect 16762 19216 16764 19236
rect 16764 19216 16816 19236
rect 16816 19216 16818 19236
rect 17038 20984 17094 21040
rect 19890 29280 19946 29336
rect 17314 18944 17370 19000
rect 17958 20440 18014 20496
rect 17682 19216 17738 19272
rect 17590 18964 17646 19000
rect 17590 18944 17592 18964
rect 17592 18944 17644 18964
rect 17644 18944 17646 18964
rect 17314 18672 17370 18728
rect 16762 18148 16818 18184
rect 16762 18128 16764 18148
rect 16764 18128 16816 18148
rect 16816 18128 16818 18148
rect 16302 17584 16358 17640
rect 16394 17176 16450 17232
rect 16210 15408 16266 15464
rect 15934 12008 15990 12064
rect 16486 12280 16542 12336
rect 15474 5208 15530 5264
rect 16578 11056 16634 11112
rect 18234 20032 18290 20088
rect 18050 19896 18106 19952
rect 18234 19080 18290 19136
rect 18142 18944 18198 19000
rect 17314 17856 17370 17912
rect 17314 15680 17370 15736
rect 17314 15308 17316 15328
rect 17316 15308 17368 15328
rect 17368 15308 17370 15328
rect 17314 15272 17370 15308
rect 17314 15020 17370 15056
rect 17314 15000 17316 15020
rect 17316 15000 17368 15020
rect 17368 15000 17370 15020
rect 17314 14592 17370 14648
rect 17498 16632 17554 16688
rect 18234 18672 18290 18728
rect 17958 15816 18014 15872
rect 17682 13640 17738 13696
rect 18142 15272 18198 15328
rect 17958 14728 18014 14784
rect 17866 12824 17922 12880
rect 17406 11736 17462 11792
rect 16946 9424 17002 9480
rect 15382 3440 15438 3496
rect 18418 17448 18474 17504
rect 18694 18944 18750 19000
rect 18970 20168 19026 20224
rect 18878 19624 18934 19680
rect 19154 22616 19210 22672
rect 19062 19488 19118 19544
rect 19430 19780 19486 19816
rect 19430 19760 19432 19780
rect 19432 19760 19484 19780
rect 19484 19760 19486 19780
rect 18970 19216 19026 19272
rect 18878 19080 18934 19136
rect 19154 18536 19210 18592
rect 19430 18536 19486 18592
rect 19338 18400 19394 18456
rect 19154 17720 19210 17776
rect 18602 17584 18658 17640
rect 18234 12552 18290 12608
rect 18510 13232 18566 13288
rect 18694 16940 18696 16960
rect 18696 16940 18748 16960
rect 18748 16940 18750 16960
rect 18694 16904 18750 16940
rect 18786 16768 18842 16824
rect 18694 16668 18696 16688
rect 18696 16668 18748 16688
rect 18748 16668 18750 16688
rect 18694 16632 18750 16668
rect 18694 16496 18750 16552
rect 18602 9968 18658 10024
rect 18142 7928 18198 7984
rect 19154 16768 19210 16824
rect 19062 14864 19118 14920
rect 19062 14492 19064 14512
rect 19064 14492 19116 14512
rect 19116 14492 19118 14512
rect 19062 14456 19118 14492
rect 19062 13776 19118 13832
rect 19062 13640 19118 13696
rect 19062 13368 19118 13424
rect 19338 13912 19394 13968
rect 19706 20848 19762 20904
rect 34978 29688 35034 29744
rect 34610 29552 34666 29608
rect 24214 28464 24270 28520
rect 20220 27226 20276 27228
rect 20300 27226 20356 27228
rect 20380 27226 20436 27228
rect 20460 27226 20516 27228
rect 20220 27174 20266 27226
rect 20266 27174 20276 27226
rect 20300 27174 20330 27226
rect 20330 27174 20342 27226
rect 20342 27174 20356 27226
rect 20380 27174 20394 27226
rect 20394 27174 20406 27226
rect 20406 27174 20436 27226
rect 20460 27174 20470 27226
rect 20470 27174 20516 27226
rect 20220 27172 20276 27174
rect 20300 27172 20356 27174
rect 20380 27172 20436 27174
rect 20460 27172 20516 27174
rect 20074 26424 20130 26480
rect 20220 26138 20276 26140
rect 20300 26138 20356 26140
rect 20380 26138 20436 26140
rect 20460 26138 20516 26140
rect 20220 26086 20266 26138
rect 20266 26086 20276 26138
rect 20300 26086 20330 26138
rect 20330 26086 20342 26138
rect 20342 26086 20356 26138
rect 20380 26086 20394 26138
rect 20394 26086 20406 26138
rect 20406 26086 20436 26138
rect 20460 26086 20470 26138
rect 20470 26086 20516 26138
rect 20220 26084 20276 26086
rect 20300 26084 20356 26086
rect 20380 26084 20436 26086
rect 20460 26084 20516 26086
rect 20220 25050 20276 25052
rect 20300 25050 20356 25052
rect 20380 25050 20436 25052
rect 20460 25050 20516 25052
rect 20220 24998 20266 25050
rect 20266 24998 20276 25050
rect 20300 24998 20330 25050
rect 20330 24998 20342 25050
rect 20342 24998 20356 25050
rect 20380 24998 20394 25050
rect 20394 24998 20406 25050
rect 20406 24998 20436 25050
rect 20460 24998 20470 25050
rect 20470 24998 20516 25050
rect 20220 24996 20276 24998
rect 20300 24996 20356 24998
rect 20380 24996 20436 24998
rect 20460 24996 20516 24998
rect 20220 23962 20276 23964
rect 20300 23962 20356 23964
rect 20380 23962 20436 23964
rect 20460 23962 20516 23964
rect 20220 23910 20266 23962
rect 20266 23910 20276 23962
rect 20300 23910 20330 23962
rect 20330 23910 20342 23962
rect 20342 23910 20356 23962
rect 20380 23910 20394 23962
rect 20394 23910 20406 23962
rect 20406 23910 20436 23962
rect 20460 23910 20470 23962
rect 20470 23910 20516 23962
rect 20220 23908 20276 23910
rect 20300 23908 20356 23910
rect 20380 23908 20436 23910
rect 20460 23908 20516 23910
rect 20534 23160 20590 23216
rect 20220 22874 20276 22876
rect 20300 22874 20356 22876
rect 20380 22874 20436 22876
rect 20460 22874 20516 22876
rect 20220 22822 20266 22874
rect 20266 22822 20276 22874
rect 20300 22822 20330 22874
rect 20330 22822 20342 22874
rect 20342 22822 20356 22874
rect 20380 22822 20394 22874
rect 20394 22822 20406 22874
rect 20406 22822 20436 22874
rect 20460 22822 20470 22874
rect 20470 22822 20516 22874
rect 20220 22820 20276 22822
rect 20300 22820 20356 22822
rect 20380 22820 20436 22822
rect 20460 22820 20516 22822
rect 19890 22072 19946 22128
rect 19798 20476 19800 20496
rect 19800 20476 19852 20496
rect 19852 20476 19854 20496
rect 19798 20440 19854 20476
rect 20220 21786 20276 21788
rect 20300 21786 20356 21788
rect 20380 21786 20436 21788
rect 20460 21786 20516 21788
rect 20220 21734 20266 21786
rect 20266 21734 20276 21786
rect 20300 21734 20330 21786
rect 20330 21734 20342 21786
rect 20342 21734 20356 21786
rect 20380 21734 20394 21786
rect 20394 21734 20406 21786
rect 20406 21734 20436 21786
rect 20460 21734 20470 21786
rect 20470 21734 20516 21786
rect 20220 21732 20276 21734
rect 20300 21732 20356 21734
rect 20380 21732 20436 21734
rect 20460 21732 20516 21734
rect 21822 25744 21878 25800
rect 21362 23840 21418 23896
rect 21086 23568 21142 23624
rect 21270 23468 21272 23488
rect 21272 23468 21324 23488
rect 21324 23468 21326 23488
rect 21270 23432 21326 23468
rect 20626 21664 20682 21720
rect 20166 21392 20222 21448
rect 20220 20698 20276 20700
rect 20300 20698 20356 20700
rect 20380 20698 20436 20700
rect 20460 20698 20516 20700
rect 20220 20646 20266 20698
rect 20266 20646 20276 20698
rect 20300 20646 20330 20698
rect 20330 20646 20342 20698
rect 20342 20646 20356 20698
rect 20380 20646 20394 20698
rect 20394 20646 20406 20698
rect 20406 20646 20436 20698
rect 20460 20646 20470 20698
rect 20470 20646 20516 20698
rect 20220 20644 20276 20646
rect 20300 20644 20356 20646
rect 20380 20644 20436 20646
rect 20460 20644 20516 20646
rect 20902 21528 20958 21584
rect 20810 20712 20866 20768
rect 20220 19610 20276 19612
rect 20300 19610 20356 19612
rect 20380 19610 20436 19612
rect 20460 19610 20516 19612
rect 20220 19558 20266 19610
rect 20266 19558 20276 19610
rect 20300 19558 20330 19610
rect 20330 19558 20342 19610
rect 20342 19558 20356 19610
rect 20380 19558 20394 19610
rect 20394 19558 20406 19610
rect 20406 19558 20436 19610
rect 20460 19558 20470 19610
rect 20470 19558 20516 19610
rect 20220 19556 20276 19558
rect 20300 19556 20356 19558
rect 20380 19556 20436 19558
rect 20460 19556 20516 19558
rect 20350 19252 20352 19272
rect 20352 19252 20404 19272
rect 20404 19252 20406 19272
rect 20350 19216 20406 19252
rect 19890 17720 19946 17776
rect 19798 17448 19854 17504
rect 19614 16632 19670 16688
rect 19706 16396 19708 16416
rect 19708 16396 19760 16416
rect 19760 16396 19762 16416
rect 19706 16360 19762 16396
rect 19706 16088 19762 16144
rect 19522 15000 19578 15056
rect 20220 18522 20276 18524
rect 20300 18522 20356 18524
rect 20380 18522 20436 18524
rect 20460 18522 20516 18524
rect 20220 18470 20266 18522
rect 20266 18470 20276 18522
rect 20300 18470 20330 18522
rect 20330 18470 20342 18522
rect 20342 18470 20356 18522
rect 20380 18470 20394 18522
rect 20394 18470 20406 18522
rect 20406 18470 20436 18522
rect 20460 18470 20470 18522
rect 20470 18470 20516 18522
rect 20220 18468 20276 18470
rect 20300 18468 20356 18470
rect 20380 18468 20436 18470
rect 20460 18468 20516 18470
rect 20074 17448 20130 17504
rect 20220 17434 20276 17436
rect 20300 17434 20356 17436
rect 20380 17434 20436 17436
rect 20460 17434 20516 17436
rect 20220 17382 20266 17434
rect 20266 17382 20276 17434
rect 20300 17382 20330 17434
rect 20330 17382 20342 17434
rect 20342 17382 20356 17434
rect 20380 17382 20394 17434
rect 20394 17382 20406 17434
rect 20406 17382 20436 17434
rect 20460 17382 20470 17434
rect 20470 17382 20516 17434
rect 20220 17380 20276 17382
rect 20300 17380 20356 17382
rect 20380 17380 20436 17382
rect 20460 17380 20516 17382
rect 20074 17312 20130 17368
rect 20718 17876 20774 17912
rect 20718 17856 20720 17876
rect 20720 17856 20772 17876
rect 20772 17856 20774 17876
rect 20718 17448 20774 17504
rect 19798 15136 19854 15192
rect 19338 11092 19340 11112
rect 19340 11092 19392 11112
rect 19392 11092 19394 11112
rect 19338 11056 19394 11092
rect 20074 16632 20130 16688
rect 20074 16496 20130 16552
rect 20534 16496 20590 16552
rect 20220 16346 20276 16348
rect 20300 16346 20356 16348
rect 20380 16346 20436 16348
rect 20460 16346 20516 16348
rect 20220 16294 20266 16346
rect 20266 16294 20276 16346
rect 20300 16294 20330 16346
rect 20330 16294 20342 16346
rect 20342 16294 20356 16346
rect 20380 16294 20394 16346
rect 20394 16294 20406 16346
rect 20406 16294 20436 16346
rect 20460 16294 20470 16346
rect 20470 16294 20516 16346
rect 20220 16292 20276 16294
rect 20300 16292 20356 16294
rect 20380 16292 20436 16294
rect 20460 16292 20516 16294
rect 20534 16124 20536 16144
rect 20536 16124 20588 16144
rect 20588 16124 20590 16144
rect 20534 16088 20590 16124
rect 20166 15816 20222 15872
rect 20166 15544 20222 15600
rect 20074 15408 20130 15464
rect 20220 15258 20276 15260
rect 20300 15258 20356 15260
rect 20380 15258 20436 15260
rect 20460 15258 20516 15260
rect 20220 15206 20266 15258
rect 20266 15206 20276 15258
rect 20300 15206 20330 15258
rect 20330 15206 20342 15258
rect 20342 15206 20356 15258
rect 20380 15206 20394 15258
rect 20394 15206 20406 15258
rect 20406 15206 20436 15258
rect 20460 15206 20470 15258
rect 20470 15206 20516 15258
rect 20220 15204 20276 15206
rect 20300 15204 20356 15206
rect 20380 15204 20436 15206
rect 20460 15204 20516 15206
rect 20074 14864 20130 14920
rect 20718 15816 20774 15872
rect 20220 14170 20276 14172
rect 20300 14170 20356 14172
rect 20380 14170 20436 14172
rect 20460 14170 20516 14172
rect 20220 14118 20266 14170
rect 20266 14118 20276 14170
rect 20300 14118 20330 14170
rect 20330 14118 20342 14170
rect 20342 14118 20356 14170
rect 20380 14118 20394 14170
rect 20394 14118 20406 14170
rect 20406 14118 20436 14170
rect 20460 14118 20470 14170
rect 20470 14118 20516 14170
rect 20220 14116 20276 14118
rect 20300 14116 20356 14118
rect 20380 14116 20436 14118
rect 20460 14116 20516 14118
rect 20166 13912 20222 13968
rect 20534 13932 20590 13968
rect 20534 13912 20536 13932
rect 20536 13912 20588 13932
rect 20588 13912 20590 13932
rect 20442 13812 20444 13832
rect 20444 13812 20496 13832
rect 20496 13812 20498 13832
rect 20442 13776 20498 13812
rect 20220 13082 20276 13084
rect 20300 13082 20356 13084
rect 20380 13082 20436 13084
rect 20460 13082 20516 13084
rect 20220 13030 20266 13082
rect 20266 13030 20276 13082
rect 20300 13030 20330 13082
rect 20330 13030 20342 13082
rect 20342 13030 20356 13082
rect 20380 13030 20394 13082
rect 20394 13030 20406 13082
rect 20406 13030 20436 13082
rect 20460 13030 20470 13082
rect 20470 13030 20516 13082
rect 20220 13028 20276 13030
rect 20300 13028 20356 13030
rect 20380 13028 20436 13030
rect 20460 13028 20516 13030
rect 20220 11994 20276 11996
rect 20300 11994 20356 11996
rect 20380 11994 20436 11996
rect 20460 11994 20516 11996
rect 20220 11942 20266 11994
rect 20266 11942 20276 11994
rect 20300 11942 20330 11994
rect 20330 11942 20342 11994
rect 20342 11942 20356 11994
rect 20380 11942 20394 11994
rect 20394 11942 20406 11994
rect 20406 11942 20436 11994
rect 20460 11942 20470 11994
rect 20470 11942 20516 11994
rect 20220 11940 20276 11942
rect 20300 11940 20356 11942
rect 20380 11940 20436 11942
rect 20460 11940 20516 11942
rect 20442 11328 20498 11384
rect 21178 20032 21234 20088
rect 21086 19488 21142 19544
rect 21638 21800 21694 21856
rect 21362 19624 21418 19680
rect 21454 19352 21510 19408
rect 21178 18536 21234 18592
rect 21362 18672 21418 18728
rect 21822 21140 21878 21176
rect 21822 21120 21824 21140
rect 21824 21120 21876 21140
rect 21876 21120 21878 21140
rect 21362 17720 21418 17776
rect 21362 17312 21418 17368
rect 21178 16360 21234 16416
rect 21086 16088 21142 16144
rect 20902 15564 20958 15600
rect 20902 15544 20904 15564
rect 20904 15544 20956 15564
rect 20956 15544 20958 15564
rect 20902 15308 20904 15328
rect 20904 15308 20956 15328
rect 20956 15308 20958 15328
rect 20902 15272 20958 15308
rect 20902 15156 20958 15192
rect 20902 15136 20904 15156
rect 20904 15136 20956 15156
rect 20956 15136 20958 15156
rect 20902 14864 20958 14920
rect 20902 14592 20958 14648
rect 20902 14048 20958 14104
rect 21178 15136 21234 15192
rect 21086 14592 21142 14648
rect 21086 14320 21142 14376
rect 20994 13932 21050 13968
rect 20994 13912 20996 13932
rect 20996 13912 21048 13932
rect 21048 13912 21050 13932
rect 20718 13504 20774 13560
rect 20810 13096 20866 13152
rect 21178 13640 21234 13696
rect 21086 13504 21142 13560
rect 20902 12008 20958 12064
rect 21362 13640 21418 13696
rect 20220 10906 20276 10908
rect 20300 10906 20356 10908
rect 20380 10906 20436 10908
rect 20460 10906 20516 10908
rect 20220 10854 20266 10906
rect 20266 10854 20276 10906
rect 20300 10854 20330 10906
rect 20330 10854 20342 10906
rect 20342 10854 20356 10906
rect 20380 10854 20394 10906
rect 20394 10854 20406 10906
rect 20406 10854 20436 10906
rect 20460 10854 20470 10906
rect 20470 10854 20516 10906
rect 20220 10852 20276 10854
rect 20300 10852 20356 10854
rect 20380 10852 20436 10854
rect 20460 10852 20516 10854
rect 20220 9818 20276 9820
rect 20300 9818 20356 9820
rect 20380 9818 20436 9820
rect 20460 9818 20516 9820
rect 20220 9766 20266 9818
rect 20266 9766 20276 9818
rect 20300 9766 20330 9818
rect 20330 9766 20342 9818
rect 20342 9766 20356 9818
rect 20380 9766 20394 9818
rect 20394 9766 20406 9818
rect 20406 9766 20436 9818
rect 20460 9766 20470 9818
rect 20470 9766 20516 9818
rect 20220 9764 20276 9766
rect 20300 9764 20356 9766
rect 20380 9764 20436 9766
rect 20460 9764 20516 9766
rect 20220 8730 20276 8732
rect 20300 8730 20356 8732
rect 20380 8730 20436 8732
rect 20460 8730 20516 8732
rect 20220 8678 20266 8730
rect 20266 8678 20276 8730
rect 20300 8678 20330 8730
rect 20330 8678 20342 8730
rect 20342 8678 20356 8730
rect 20380 8678 20394 8730
rect 20394 8678 20406 8730
rect 20406 8678 20436 8730
rect 20460 8678 20470 8730
rect 20470 8678 20516 8730
rect 20220 8676 20276 8678
rect 20300 8676 20356 8678
rect 20380 8676 20436 8678
rect 20460 8676 20516 8678
rect 19890 7792 19946 7848
rect 20220 7642 20276 7644
rect 20300 7642 20356 7644
rect 20380 7642 20436 7644
rect 20460 7642 20516 7644
rect 20220 7590 20266 7642
rect 20266 7590 20276 7642
rect 20300 7590 20330 7642
rect 20330 7590 20342 7642
rect 20342 7590 20356 7642
rect 20380 7590 20394 7642
rect 20394 7590 20406 7642
rect 20406 7590 20436 7642
rect 20460 7590 20470 7642
rect 20470 7590 20516 7642
rect 20220 7588 20276 7590
rect 20300 7588 20356 7590
rect 20380 7588 20436 7590
rect 20460 7588 20516 7590
rect 20220 6554 20276 6556
rect 20300 6554 20356 6556
rect 20380 6554 20436 6556
rect 20460 6554 20516 6556
rect 20220 6502 20266 6554
rect 20266 6502 20276 6554
rect 20300 6502 20330 6554
rect 20330 6502 20342 6554
rect 20342 6502 20356 6554
rect 20380 6502 20394 6554
rect 20394 6502 20406 6554
rect 20406 6502 20436 6554
rect 20460 6502 20470 6554
rect 20470 6502 20516 6554
rect 20220 6500 20276 6502
rect 20300 6500 20356 6502
rect 20380 6500 20436 6502
rect 20460 6500 20516 6502
rect 20220 5466 20276 5468
rect 20300 5466 20356 5468
rect 20380 5466 20436 5468
rect 20460 5466 20516 5468
rect 20220 5414 20266 5466
rect 20266 5414 20276 5466
rect 20300 5414 20330 5466
rect 20330 5414 20342 5466
rect 20342 5414 20356 5466
rect 20380 5414 20394 5466
rect 20394 5414 20406 5466
rect 20406 5414 20436 5466
rect 20460 5414 20470 5466
rect 20470 5414 20516 5466
rect 20220 5412 20276 5414
rect 20300 5412 20356 5414
rect 20380 5412 20436 5414
rect 20460 5412 20516 5414
rect 20220 4378 20276 4380
rect 20300 4378 20356 4380
rect 20380 4378 20436 4380
rect 20460 4378 20516 4380
rect 20220 4326 20266 4378
rect 20266 4326 20276 4378
rect 20300 4326 20330 4378
rect 20330 4326 20342 4378
rect 20342 4326 20356 4378
rect 20380 4326 20394 4378
rect 20394 4326 20406 4378
rect 20406 4326 20436 4378
rect 20460 4326 20470 4378
rect 20470 4326 20516 4378
rect 20220 4324 20276 4326
rect 20300 4324 20356 4326
rect 20380 4324 20436 4326
rect 20460 4324 20516 4326
rect 21178 11348 21234 11384
rect 21178 11328 21180 11348
rect 21180 11328 21232 11348
rect 21232 11328 21234 11348
rect 20220 3290 20276 3292
rect 20300 3290 20356 3292
rect 20380 3290 20436 3292
rect 20460 3290 20516 3292
rect 20220 3238 20266 3290
rect 20266 3238 20276 3290
rect 20300 3238 20330 3290
rect 20330 3238 20342 3290
rect 20342 3238 20356 3290
rect 20380 3238 20394 3290
rect 20394 3238 20406 3290
rect 20406 3238 20436 3290
rect 20460 3238 20470 3290
rect 20470 3238 20516 3290
rect 20220 3236 20276 3238
rect 20300 3236 20356 3238
rect 20380 3236 20436 3238
rect 20460 3236 20516 3238
rect 22006 26696 22062 26752
rect 22098 25064 22154 25120
rect 22006 22380 22008 22400
rect 22008 22380 22060 22400
rect 22060 22380 22062 22400
rect 22006 22344 22062 22380
rect 22742 24384 22798 24440
rect 22098 21800 22154 21856
rect 22190 21528 22246 21584
rect 22098 20440 22154 20496
rect 21914 20032 21970 20088
rect 22190 19372 22246 19408
rect 22190 19352 22192 19372
rect 22192 19352 22244 19372
rect 22244 19352 22246 19372
rect 22006 17720 22062 17776
rect 21730 16652 21786 16688
rect 21730 16632 21732 16652
rect 21732 16632 21784 16652
rect 21784 16632 21786 16652
rect 21638 16224 21694 16280
rect 21546 16088 21602 16144
rect 21914 17060 21970 17096
rect 21914 17040 21916 17060
rect 21916 17040 21968 17060
rect 21968 17040 21970 17060
rect 22742 22752 22798 22808
rect 22834 22380 22836 22400
rect 22836 22380 22888 22400
rect 22888 22380 22890 22400
rect 22834 22344 22890 22380
rect 22834 21664 22890 21720
rect 22558 20576 22614 20632
rect 22374 19896 22430 19952
rect 22466 19080 22522 19136
rect 22374 18400 22430 18456
rect 22466 17448 22522 17504
rect 22282 17312 22338 17368
rect 21546 15272 21602 15328
rect 21546 13912 21602 13968
rect 21546 13504 21602 13560
rect 21730 15272 21786 15328
rect 21546 11464 21602 11520
rect 21454 10648 21510 10704
rect 22466 16496 22522 16552
rect 22190 16088 22246 16144
rect 22098 15680 22154 15736
rect 22190 14456 22246 14512
rect 22006 14048 22062 14104
rect 22006 13524 22062 13560
rect 22006 13504 22008 13524
rect 22008 13504 22060 13524
rect 22060 13504 22062 13524
rect 21822 12416 21878 12472
rect 22466 15544 22522 15600
rect 21914 11464 21970 11520
rect 21914 11328 21970 11384
rect 21178 2896 21234 2952
rect 22466 12416 22522 12472
rect 22926 21392 22982 21448
rect 23386 22208 23442 22264
rect 23110 21392 23166 21448
rect 23110 20984 23166 21040
rect 22834 20748 22836 20768
rect 22836 20748 22888 20768
rect 22888 20748 22890 20768
rect 22834 20712 22890 20748
rect 23478 20576 23534 20632
rect 23754 21004 23810 21040
rect 23754 20984 23756 21004
rect 23756 20984 23808 21004
rect 23808 20984 23810 21004
rect 23570 20032 23626 20088
rect 23110 18672 23166 18728
rect 23018 18536 23074 18592
rect 22650 15700 22706 15736
rect 22650 15680 22652 15700
rect 22652 15680 22704 15700
rect 22704 15680 22706 15700
rect 22742 15272 22798 15328
rect 22650 10804 22706 10840
rect 22650 10784 22652 10804
rect 22652 10784 22704 10804
rect 22704 10784 22706 10804
rect 22558 10240 22614 10296
rect 23386 17992 23442 18048
rect 23386 15952 23442 16008
rect 23846 19352 23902 19408
rect 29852 27770 29908 27772
rect 29932 27770 29988 27772
rect 30012 27770 30068 27772
rect 30092 27770 30148 27772
rect 29852 27718 29898 27770
rect 29898 27718 29908 27770
rect 29932 27718 29962 27770
rect 29962 27718 29974 27770
rect 29974 27718 29988 27770
rect 30012 27718 30026 27770
rect 30026 27718 30038 27770
rect 30038 27718 30068 27770
rect 30092 27718 30102 27770
rect 30102 27718 30148 27770
rect 29852 27716 29908 27718
rect 29932 27716 29988 27718
rect 30012 27716 30068 27718
rect 30092 27716 30148 27718
rect 30470 27920 30526 27976
rect 24582 26016 24638 26072
rect 24398 25472 24454 25528
rect 24306 24928 24362 24984
rect 24122 22480 24178 22536
rect 24398 22616 24454 22672
rect 24582 23024 24638 23080
rect 24674 22344 24730 22400
rect 24306 21120 24362 21176
rect 23846 18672 23902 18728
rect 23662 18264 23718 18320
rect 23570 15544 23626 15600
rect 23202 15136 23258 15192
rect 23110 14728 23166 14784
rect 23386 14900 23388 14920
rect 23388 14900 23440 14920
rect 23440 14900 23442 14920
rect 23386 14864 23442 14900
rect 23386 14728 23442 14784
rect 23202 14184 23258 14240
rect 23110 10104 23166 10160
rect 23018 7520 23074 7576
rect 23754 16532 23756 16552
rect 23756 16532 23808 16552
rect 23808 16532 23810 16552
rect 23754 16496 23810 16532
rect 24030 16496 24086 16552
rect 23754 15020 23810 15056
rect 23754 15000 23756 15020
rect 23756 15000 23808 15020
rect 23808 15000 23810 15020
rect 23846 13932 23902 13968
rect 23846 13912 23848 13932
rect 23848 13912 23900 13932
rect 23900 13912 23902 13932
rect 23754 12144 23810 12200
rect 23662 11772 23664 11792
rect 23664 11772 23716 11792
rect 23716 11772 23718 11792
rect 23662 11736 23718 11772
rect 24582 21664 24638 21720
rect 24582 20576 24638 20632
rect 27526 26868 27528 26888
rect 27528 26868 27580 26888
rect 27580 26868 27582 26888
rect 26422 26424 26478 26480
rect 25226 25200 25282 25256
rect 24950 22480 25006 22536
rect 25410 24132 25466 24168
rect 25410 24112 25412 24132
rect 25412 24112 25464 24132
rect 25464 24112 25466 24132
rect 25410 23976 25466 24032
rect 25134 21936 25190 21992
rect 25594 23976 25650 24032
rect 25594 23568 25650 23624
rect 25778 23568 25834 23624
rect 25778 22652 25780 22672
rect 25780 22652 25832 22672
rect 25832 22652 25834 22672
rect 25778 22616 25834 22652
rect 25042 21392 25098 21448
rect 24858 20032 24914 20088
rect 24858 19624 24914 19680
rect 24950 19216 25006 19272
rect 24858 18944 24914 19000
rect 24490 17856 24546 17912
rect 24674 17856 24730 17912
rect 24490 17448 24546 17504
rect 24214 15972 24270 16008
rect 24214 15952 24216 15972
rect 24216 15952 24268 15972
rect 24268 15952 24270 15972
rect 24214 15544 24270 15600
rect 24214 15000 24270 15056
rect 24214 14456 24270 14512
rect 24214 13096 24270 13152
rect 23570 9444 23626 9480
rect 23570 9424 23572 9444
rect 23572 9424 23624 9444
rect 23624 9424 23626 9444
rect 23202 6568 23258 6624
rect 24306 11056 24362 11112
rect 24950 18300 24952 18320
rect 24952 18300 25004 18320
rect 25004 18300 25006 18320
rect 24950 18264 25006 18300
rect 25042 18128 25098 18184
rect 24950 17176 25006 17232
rect 24858 16088 24914 16144
rect 24766 15272 24822 15328
rect 24674 13776 24730 13832
rect 24674 13404 24676 13424
rect 24676 13404 24728 13424
rect 24728 13404 24730 13424
rect 24674 13368 24730 13404
rect 24858 14728 24914 14784
rect 24766 12688 24822 12744
rect 25502 21392 25558 21448
rect 25410 19216 25466 19272
rect 26054 24112 26110 24168
rect 25778 20032 25834 20088
rect 25410 17720 25466 17776
rect 25318 15544 25374 15600
rect 24950 13776 25006 13832
rect 24950 13252 25006 13288
rect 24950 13232 24952 13252
rect 24952 13232 25004 13252
rect 25004 13232 25006 13252
rect 24674 12416 24730 12472
rect 24766 12316 24768 12336
rect 24768 12316 24820 12336
rect 24820 12316 24822 12336
rect 24766 12280 24822 12316
rect 24674 12144 24730 12200
rect 25410 12960 25466 13016
rect 25134 12688 25190 12744
rect 24766 10648 24822 10704
rect 24674 10376 24730 10432
rect 25042 11328 25098 11384
rect 24950 10668 25006 10704
rect 24950 10648 24952 10668
rect 24952 10648 25004 10668
rect 25004 10648 25006 10668
rect 23846 5480 23902 5536
rect 21914 2352 21970 2408
rect 14554 1944 14610 2000
rect 20220 2202 20276 2204
rect 20300 2202 20356 2204
rect 20380 2202 20436 2204
rect 20460 2202 20516 2204
rect 20220 2150 20266 2202
rect 20266 2150 20276 2202
rect 20300 2150 20330 2202
rect 20330 2150 20342 2202
rect 20342 2150 20356 2202
rect 20380 2150 20394 2202
rect 20394 2150 20406 2202
rect 20406 2150 20436 2202
rect 20460 2150 20470 2202
rect 20470 2150 20516 2202
rect 20220 2148 20276 2150
rect 20300 2148 20356 2150
rect 20380 2148 20436 2150
rect 20460 2148 20516 2150
rect 25594 11348 25650 11384
rect 25594 11328 25596 11348
rect 25596 11328 25648 11348
rect 25648 11328 25650 11348
rect 26054 20340 26056 20360
rect 26056 20340 26108 20360
rect 26108 20340 26110 20360
rect 26054 20304 26110 20340
rect 26054 18808 26110 18864
rect 25778 14864 25834 14920
rect 26054 17196 26110 17232
rect 26054 17176 26056 17196
rect 26056 17176 26108 17196
rect 26108 17176 26110 17196
rect 26330 23180 26386 23216
rect 26330 23160 26332 23180
rect 26332 23160 26384 23180
rect 26384 23160 26386 23180
rect 26330 23024 26386 23080
rect 26238 22888 26294 22944
rect 26238 22616 26294 22672
rect 26698 23432 26754 23488
rect 26698 22480 26754 22536
rect 27250 25200 27306 25256
rect 26882 24656 26938 24712
rect 26882 24012 26884 24032
rect 26884 24012 26936 24032
rect 26936 24012 26938 24032
rect 26882 23976 26938 24012
rect 26882 23044 26938 23080
rect 26882 23024 26884 23044
rect 26884 23024 26936 23044
rect 26936 23024 26938 23044
rect 26882 22888 26938 22944
rect 27526 26832 27582 26868
rect 28446 26560 28502 26616
rect 27618 26288 27674 26344
rect 27434 24520 27490 24576
rect 27342 24248 27398 24304
rect 27342 23976 27398 24032
rect 27342 23840 27398 23896
rect 27158 23588 27214 23624
rect 27158 23568 27160 23588
rect 27160 23568 27212 23588
rect 27212 23568 27214 23588
rect 27066 23296 27122 23352
rect 26330 15136 26386 15192
rect 26238 14048 26294 14104
rect 26238 13776 26294 13832
rect 26054 12416 26110 12472
rect 25686 8880 25742 8936
rect 24582 8064 24638 8120
rect 24766 8084 24822 8120
rect 24766 8064 24768 8084
rect 24768 8064 24820 8084
rect 24820 8064 24822 8084
rect 24858 3304 24914 3360
rect 24582 2488 24638 2544
rect 25962 8084 26018 8120
rect 26422 14048 26478 14104
rect 26422 12980 26478 13016
rect 26422 12960 26424 12980
rect 26424 12960 26476 12980
rect 26476 12960 26478 12980
rect 26238 12008 26294 12064
rect 26238 11872 26294 11928
rect 26146 11328 26202 11384
rect 26422 11056 26478 11112
rect 26238 10260 26294 10296
rect 26238 10240 26240 10260
rect 26240 10240 26292 10260
rect 26292 10240 26294 10260
rect 25962 8064 25964 8084
rect 25964 8064 26016 8084
rect 26016 8064 26018 8084
rect 25778 4120 25834 4176
rect 27342 22344 27398 22400
rect 27342 22208 27398 22264
rect 27066 21936 27122 21992
rect 26698 19916 26754 19952
rect 26698 19896 26700 19916
rect 26700 19896 26752 19916
rect 26752 19896 26754 19916
rect 27250 21256 27306 21312
rect 27250 20440 27306 20496
rect 27158 20168 27214 20224
rect 27618 21548 27674 21584
rect 27618 21528 27620 21548
rect 27620 21528 27672 21548
rect 27672 21528 27674 21548
rect 27158 19624 27214 19680
rect 27434 19624 27490 19680
rect 27066 18672 27122 18728
rect 26698 16496 26754 16552
rect 26606 15680 26662 15736
rect 26790 13504 26846 13560
rect 27250 18708 27252 18728
rect 27252 18708 27304 18728
rect 27304 18708 27306 18728
rect 27250 18672 27306 18708
rect 26974 13368 27030 13424
rect 26882 12144 26938 12200
rect 26790 11600 26846 11656
rect 26238 8336 26294 8392
rect 27342 16768 27398 16824
rect 27158 15816 27214 15872
rect 27066 11056 27122 11112
rect 26974 10512 27030 10568
rect 27342 14184 27398 14240
rect 27342 12280 27398 12336
rect 27342 11348 27398 11384
rect 27342 11328 27344 11348
rect 27344 11328 27396 11348
rect 27396 11328 27398 11348
rect 27986 24112 28042 24168
rect 27986 23432 28042 23488
rect 28814 27376 28870 27432
rect 28262 23976 28318 24032
rect 28170 23296 28226 23352
rect 27986 23060 27988 23080
rect 27988 23060 28040 23080
rect 28040 23060 28042 23080
rect 27986 23024 28042 23060
rect 28446 25100 28448 25120
rect 28448 25100 28500 25120
rect 28500 25100 28502 25120
rect 28446 25064 28502 25100
rect 28354 23024 28410 23080
rect 28078 22752 28134 22808
rect 28078 22480 28134 22536
rect 27986 22208 28042 22264
rect 27894 21684 27950 21720
rect 27894 21664 27896 21684
rect 27896 21664 27948 21684
rect 27948 21664 27950 21684
rect 28078 22072 28134 22128
rect 27526 16244 27582 16280
rect 27526 16224 27528 16244
rect 27528 16224 27580 16244
rect 27580 16224 27582 16244
rect 27618 14592 27674 14648
rect 27526 13640 27582 13696
rect 27526 13232 27582 13288
rect 27986 14456 28042 14512
rect 27894 14184 27950 14240
rect 27894 12144 27950 12200
rect 27894 11756 27950 11792
rect 27894 11736 27896 11756
rect 27896 11736 27948 11756
rect 27948 11736 27950 11756
rect 28170 21956 28226 21992
rect 28170 21936 28172 21956
rect 28172 21936 28224 21956
rect 28224 21936 28226 21956
rect 28170 21392 28226 21448
rect 28998 26152 29054 26208
rect 28998 25744 29054 25800
rect 28906 25644 28908 25664
rect 28908 25644 28960 25664
rect 28960 25644 28962 25664
rect 28906 25608 28962 25644
rect 28906 25336 28962 25392
rect 28722 24112 28778 24168
rect 28630 22480 28686 22536
rect 28538 21256 28594 21312
rect 28170 19352 28226 19408
rect 28078 13640 28134 13696
rect 27710 10920 27766 10976
rect 27802 10376 27858 10432
rect 27986 10784 28042 10840
rect 27986 10240 28042 10296
rect 27710 9560 27766 9616
rect 28906 23432 28962 23488
rect 28814 23296 28870 23352
rect 28630 19896 28686 19952
rect 28538 19216 28594 19272
rect 28262 18128 28318 18184
rect 28262 14184 28318 14240
rect 28262 13776 28318 13832
rect 28630 17992 28686 18048
rect 28722 17720 28778 17776
rect 28538 16496 28594 16552
rect 28906 22480 28962 22536
rect 28906 22344 28962 22400
rect 29274 25880 29330 25936
rect 29182 25744 29238 25800
rect 28906 21256 28962 21312
rect 29274 22344 29330 22400
rect 29182 20884 29184 20904
rect 29184 20884 29236 20904
rect 29236 20884 29238 20904
rect 29182 20848 29238 20884
rect 29550 26696 29606 26752
rect 29734 26968 29790 27024
rect 29852 26682 29908 26684
rect 29932 26682 29988 26684
rect 30012 26682 30068 26684
rect 30092 26682 30148 26684
rect 29852 26630 29898 26682
rect 29898 26630 29908 26682
rect 29932 26630 29962 26682
rect 29962 26630 29974 26682
rect 29974 26630 29988 26682
rect 30012 26630 30026 26682
rect 30026 26630 30038 26682
rect 30038 26630 30068 26682
rect 30092 26630 30102 26682
rect 30102 26630 30148 26682
rect 29852 26628 29908 26630
rect 29932 26628 29988 26630
rect 30012 26628 30068 26630
rect 30092 26628 30148 26630
rect 29734 26424 29790 26480
rect 29734 25880 29790 25936
rect 29852 25594 29908 25596
rect 29932 25594 29988 25596
rect 30012 25594 30068 25596
rect 30092 25594 30148 25596
rect 29852 25542 29898 25594
rect 29898 25542 29908 25594
rect 29932 25542 29962 25594
rect 29962 25542 29974 25594
rect 29974 25542 29988 25594
rect 30012 25542 30026 25594
rect 30026 25542 30038 25594
rect 30038 25542 30068 25594
rect 30092 25542 30102 25594
rect 30102 25542 30148 25594
rect 29852 25540 29908 25542
rect 29932 25540 29988 25542
rect 30012 25540 30068 25542
rect 30092 25540 30148 25542
rect 29734 24928 29790 24984
rect 29642 23704 29698 23760
rect 29852 24506 29908 24508
rect 29932 24506 29988 24508
rect 30012 24506 30068 24508
rect 30092 24506 30148 24508
rect 29852 24454 29898 24506
rect 29898 24454 29908 24506
rect 29932 24454 29962 24506
rect 29962 24454 29974 24506
rect 29974 24454 29988 24506
rect 30012 24454 30026 24506
rect 30026 24454 30038 24506
rect 30038 24454 30068 24506
rect 30092 24454 30102 24506
rect 30102 24454 30148 24506
rect 29852 24452 29908 24454
rect 29932 24452 29988 24454
rect 30012 24452 30068 24454
rect 30092 24452 30148 24454
rect 30102 23704 30158 23760
rect 30010 23604 30012 23624
rect 30012 23604 30064 23624
rect 30064 23604 30066 23624
rect 30010 23568 30066 23604
rect 31942 27784 31998 27840
rect 30470 26036 30526 26072
rect 30470 26016 30472 26036
rect 30472 26016 30524 26036
rect 30524 26016 30526 26036
rect 30378 25608 30434 25664
rect 30378 25336 30434 25392
rect 30378 24148 30380 24168
rect 30380 24148 30432 24168
rect 30432 24148 30434 24168
rect 30378 24112 30434 24148
rect 30838 26732 30840 26752
rect 30840 26732 30892 26752
rect 30892 26732 30894 26752
rect 30838 26696 30894 26732
rect 31206 26580 31262 26616
rect 31206 26560 31208 26580
rect 31208 26560 31260 26580
rect 31260 26560 31262 26580
rect 31022 26152 31078 26208
rect 30562 25236 30564 25256
rect 30564 25236 30616 25256
rect 30616 25236 30618 25256
rect 30562 25200 30618 25236
rect 29852 23418 29908 23420
rect 29932 23418 29988 23420
rect 30012 23418 30068 23420
rect 30092 23418 30148 23420
rect 29852 23366 29898 23418
rect 29898 23366 29908 23418
rect 29932 23366 29962 23418
rect 29962 23366 29974 23418
rect 29974 23366 29988 23418
rect 30012 23366 30026 23418
rect 30026 23366 30038 23418
rect 30038 23366 30068 23418
rect 30092 23366 30102 23418
rect 30102 23366 30148 23418
rect 29852 23364 29908 23366
rect 29932 23364 29988 23366
rect 30012 23364 30068 23366
rect 30092 23364 30148 23366
rect 30102 22616 30158 22672
rect 29852 22330 29908 22332
rect 29932 22330 29988 22332
rect 30012 22330 30068 22332
rect 30092 22330 30148 22332
rect 29852 22278 29898 22330
rect 29898 22278 29908 22330
rect 29932 22278 29962 22330
rect 29962 22278 29974 22330
rect 29974 22278 29988 22330
rect 30012 22278 30026 22330
rect 30026 22278 30038 22330
rect 30038 22278 30068 22330
rect 30092 22278 30102 22330
rect 30102 22278 30148 22330
rect 29852 22276 29908 22278
rect 29932 22276 29988 22278
rect 30012 22276 30068 22278
rect 30092 22276 30148 22278
rect 29550 20712 29606 20768
rect 29274 19488 29330 19544
rect 29182 19352 29238 19408
rect 28998 16668 29000 16688
rect 29000 16668 29052 16688
rect 29052 16668 29054 16688
rect 28998 16632 29054 16668
rect 29366 18944 29422 19000
rect 29274 17992 29330 18048
rect 29182 16360 29238 16416
rect 28814 15680 28870 15736
rect 28354 13096 28410 13152
rect 28262 12552 28318 12608
rect 27710 9172 27766 9208
rect 27710 9152 27712 9172
rect 27712 9152 27764 9172
rect 27764 9152 27766 9172
rect 27894 7248 27950 7304
rect 28722 15272 28778 15328
rect 28538 14864 28594 14920
rect 28538 14592 28594 14648
rect 28722 12960 28778 13016
rect 28722 11736 28778 11792
rect 28998 15136 29054 15192
rect 28906 13640 28962 13696
rect 28906 12008 28962 12064
rect 28814 11464 28870 11520
rect 28722 10376 28778 10432
rect 28538 9968 28594 10024
rect 28446 9560 28502 9616
rect 28722 9424 28778 9480
rect 28538 9016 28594 9072
rect 28722 8628 28778 8664
rect 28722 8608 28724 8628
rect 28724 8608 28776 8628
rect 28776 8608 28778 8628
rect 28630 8508 28632 8528
rect 28632 8508 28684 8528
rect 28684 8508 28686 8528
rect 28630 8472 28686 8508
rect 28906 10240 28962 10296
rect 28446 6432 28502 6488
rect 29274 13504 29330 13560
rect 29182 13368 29238 13424
rect 29090 12708 29146 12744
rect 29090 12688 29092 12708
rect 29092 12688 29144 12708
rect 29144 12688 29146 12708
rect 30838 23840 30894 23896
rect 29852 21242 29908 21244
rect 29932 21242 29988 21244
rect 30012 21242 30068 21244
rect 30092 21242 30148 21244
rect 29852 21190 29898 21242
rect 29898 21190 29908 21242
rect 29932 21190 29962 21242
rect 29962 21190 29974 21242
rect 29974 21190 29988 21242
rect 30012 21190 30026 21242
rect 30026 21190 30038 21242
rect 30038 21190 30068 21242
rect 30092 21190 30102 21242
rect 30102 21190 30148 21242
rect 29852 21188 29908 21190
rect 29932 21188 29988 21190
rect 30012 21188 30068 21190
rect 30092 21188 30148 21190
rect 30286 21120 30342 21176
rect 29918 20848 29974 20904
rect 30562 21256 30618 21312
rect 29826 20304 29882 20360
rect 29852 20154 29908 20156
rect 29932 20154 29988 20156
rect 30012 20154 30068 20156
rect 30092 20154 30148 20156
rect 29852 20102 29898 20154
rect 29898 20102 29908 20154
rect 29932 20102 29962 20154
rect 29962 20102 29974 20154
rect 29974 20102 29988 20154
rect 30012 20102 30026 20154
rect 30026 20102 30038 20154
rect 30038 20102 30068 20154
rect 30092 20102 30102 20154
rect 30102 20102 30148 20154
rect 29852 20100 29908 20102
rect 29932 20100 29988 20102
rect 30012 20100 30068 20102
rect 30092 20100 30148 20102
rect 29852 19066 29908 19068
rect 29932 19066 29988 19068
rect 30012 19066 30068 19068
rect 30092 19066 30148 19068
rect 29852 19014 29898 19066
rect 29898 19014 29908 19066
rect 29932 19014 29962 19066
rect 29962 19014 29974 19066
rect 29974 19014 29988 19066
rect 30012 19014 30026 19066
rect 30026 19014 30038 19066
rect 30038 19014 30068 19066
rect 30092 19014 30102 19066
rect 30102 19014 30148 19066
rect 29852 19012 29908 19014
rect 29932 19012 29988 19014
rect 30012 19012 30068 19014
rect 30092 19012 30148 19014
rect 30378 20748 30380 20768
rect 30380 20748 30432 20768
rect 30432 20748 30434 20768
rect 30378 20712 30434 20748
rect 30470 20168 30526 20224
rect 29826 18808 29882 18864
rect 30378 18808 30434 18864
rect 29090 7656 29146 7712
rect 29274 11500 29276 11520
rect 29276 11500 29328 11520
rect 29328 11500 29330 11520
rect 29274 11464 29330 11500
rect 29274 11328 29330 11384
rect 29366 10104 29422 10160
rect 29550 15816 29606 15872
rect 29550 14728 29606 14784
rect 29642 14320 29698 14376
rect 29550 12552 29606 12608
rect 29550 9832 29606 9888
rect 29458 6432 29514 6488
rect 29458 5364 29514 5400
rect 29458 5344 29460 5364
rect 29460 5344 29512 5364
rect 29512 5344 29514 5364
rect 29642 8472 29698 8528
rect 29852 17978 29908 17980
rect 29932 17978 29988 17980
rect 30012 17978 30068 17980
rect 30092 17978 30148 17980
rect 29852 17926 29898 17978
rect 29898 17926 29908 17978
rect 29932 17926 29962 17978
rect 29962 17926 29974 17978
rect 29974 17926 29988 17978
rect 30012 17926 30026 17978
rect 30026 17926 30038 17978
rect 30038 17926 30068 17978
rect 30092 17926 30102 17978
rect 30102 17926 30148 17978
rect 29852 17924 29908 17926
rect 29932 17924 29988 17926
rect 30012 17924 30068 17926
rect 30092 17924 30148 17926
rect 29852 16890 29908 16892
rect 29932 16890 29988 16892
rect 30012 16890 30068 16892
rect 30092 16890 30148 16892
rect 29852 16838 29898 16890
rect 29898 16838 29908 16890
rect 29932 16838 29962 16890
rect 29962 16838 29974 16890
rect 29974 16838 29988 16890
rect 30012 16838 30026 16890
rect 30026 16838 30038 16890
rect 30038 16838 30068 16890
rect 30092 16838 30102 16890
rect 30102 16838 30148 16890
rect 29852 16836 29908 16838
rect 29932 16836 29988 16838
rect 30012 16836 30068 16838
rect 30092 16836 30148 16838
rect 29852 15802 29908 15804
rect 29932 15802 29988 15804
rect 30012 15802 30068 15804
rect 30092 15802 30148 15804
rect 29852 15750 29898 15802
rect 29898 15750 29908 15802
rect 29932 15750 29962 15802
rect 29962 15750 29974 15802
rect 29974 15750 29988 15802
rect 30012 15750 30026 15802
rect 30026 15750 30038 15802
rect 30038 15750 30068 15802
rect 30092 15750 30102 15802
rect 30102 15750 30148 15802
rect 29852 15748 29908 15750
rect 29932 15748 29988 15750
rect 30012 15748 30068 15750
rect 30092 15748 30148 15750
rect 29852 14714 29908 14716
rect 29932 14714 29988 14716
rect 30012 14714 30068 14716
rect 30092 14714 30148 14716
rect 29852 14662 29898 14714
rect 29898 14662 29908 14714
rect 29932 14662 29962 14714
rect 29962 14662 29974 14714
rect 29974 14662 29988 14714
rect 30012 14662 30026 14714
rect 30026 14662 30038 14714
rect 30038 14662 30068 14714
rect 30092 14662 30102 14714
rect 30102 14662 30148 14714
rect 29852 14660 29908 14662
rect 29932 14660 29988 14662
rect 30012 14660 30068 14662
rect 30092 14660 30148 14662
rect 29852 13626 29908 13628
rect 29932 13626 29988 13628
rect 30012 13626 30068 13628
rect 30092 13626 30148 13628
rect 29852 13574 29898 13626
rect 29898 13574 29908 13626
rect 29932 13574 29962 13626
rect 29962 13574 29974 13626
rect 29974 13574 29988 13626
rect 30012 13574 30026 13626
rect 30026 13574 30038 13626
rect 30038 13574 30068 13626
rect 30092 13574 30102 13626
rect 30102 13574 30148 13626
rect 29852 13572 29908 13574
rect 29932 13572 29988 13574
rect 30012 13572 30068 13574
rect 30092 13572 30148 13574
rect 29826 13368 29882 13424
rect 29826 13096 29882 13152
rect 29852 12538 29908 12540
rect 29932 12538 29988 12540
rect 30012 12538 30068 12540
rect 30092 12538 30148 12540
rect 29852 12486 29898 12538
rect 29898 12486 29908 12538
rect 29932 12486 29962 12538
rect 29962 12486 29974 12538
rect 29974 12486 29988 12538
rect 30012 12486 30026 12538
rect 30026 12486 30038 12538
rect 30038 12486 30068 12538
rect 30092 12486 30102 12538
rect 30102 12486 30148 12538
rect 29852 12484 29908 12486
rect 29932 12484 29988 12486
rect 30012 12484 30068 12486
rect 30092 12484 30148 12486
rect 30470 17448 30526 17504
rect 30470 16632 30526 16688
rect 30470 16360 30526 16416
rect 30470 15544 30526 15600
rect 30378 12552 30434 12608
rect 30286 11736 30342 11792
rect 29852 11450 29908 11452
rect 29932 11450 29988 11452
rect 30012 11450 30068 11452
rect 30092 11450 30148 11452
rect 29852 11398 29898 11450
rect 29898 11398 29908 11450
rect 29932 11398 29962 11450
rect 29962 11398 29974 11450
rect 29974 11398 29988 11450
rect 30012 11398 30026 11450
rect 30026 11398 30038 11450
rect 30038 11398 30068 11450
rect 30092 11398 30102 11450
rect 30102 11398 30148 11450
rect 29852 11396 29908 11398
rect 29932 11396 29988 11398
rect 30012 11396 30068 11398
rect 30092 11396 30148 11398
rect 29852 10362 29908 10364
rect 29932 10362 29988 10364
rect 30012 10362 30068 10364
rect 30092 10362 30148 10364
rect 29852 10310 29898 10362
rect 29898 10310 29908 10362
rect 29932 10310 29962 10362
rect 29962 10310 29974 10362
rect 29974 10310 29988 10362
rect 30012 10310 30026 10362
rect 30026 10310 30038 10362
rect 30038 10310 30068 10362
rect 30092 10310 30102 10362
rect 30102 10310 30148 10362
rect 29852 10308 29908 10310
rect 29932 10308 29988 10310
rect 30012 10308 30068 10310
rect 30092 10308 30148 10310
rect 29918 10104 29974 10160
rect 30194 10104 30250 10160
rect 30010 9832 30066 9888
rect 30102 9580 30158 9616
rect 30102 9560 30104 9580
rect 30104 9560 30156 9580
rect 30156 9560 30158 9580
rect 29852 9274 29908 9276
rect 29932 9274 29988 9276
rect 30012 9274 30068 9276
rect 30092 9274 30148 9276
rect 29852 9222 29898 9274
rect 29898 9222 29908 9274
rect 29932 9222 29962 9274
rect 29962 9222 29974 9274
rect 29974 9222 29988 9274
rect 30012 9222 30026 9274
rect 30026 9222 30038 9274
rect 30038 9222 30068 9274
rect 30092 9222 30102 9274
rect 30102 9222 30148 9274
rect 29852 9220 29908 9222
rect 29932 9220 29988 9222
rect 30012 9220 30068 9222
rect 30092 9220 30148 9222
rect 29642 8336 29698 8392
rect 29918 9016 29974 9072
rect 29918 8608 29974 8664
rect 30194 8492 30250 8528
rect 30194 8472 30196 8492
rect 30196 8472 30248 8492
rect 30248 8472 30250 8492
rect 29852 8186 29908 8188
rect 29932 8186 29988 8188
rect 30012 8186 30068 8188
rect 30092 8186 30148 8188
rect 29852 8134 29898 8186
rect 29898 8134 29908 8186
rect 29932 8134 29962 8186
rect 29962 8134 29974 8186
rect 29974 8134 29988 8186
rect 30012 8134 30026 8186
rect 30026 8134 30038 8186
rect 30038 8134 30068 8186
rect 30092 8134 30102 8186
rect 30102 8134 30148 8186
rect 29852 8132 29908 8134
rect 29932 8132 29988 8134
rect 30012 8132 30068 8134
rect 30092 8132 30148 8134
rect 29852 7098 29908 7100
rect 29932 7098 29988 7100
rect 30012 7098 30068 7100
rect 30092 7098 30148 7100
rect 29852 7046 29898 7098
rect 29898 7046 29908 7098
rect 29932 7046 29962 7098
rect 29962 7046 29974 7098
rect 29974 7046 29988 7098
rect 30012 7046 30026 7098
rect 30026 7046 30038 7098
rect 30038 7046 30068 7098
rect 30092 7046 30102 7098
rect 30102 7046 30148 7098
rect 29852 7044 29908 7046
rect 29932 7044 29988 7046
rect 30012 7044 30068 7046
rect 30092 7044 30148 7046
rect 30286 7520 30342 7576
rect 29852 6010 29908 6012
rect 29932 6010 29988 6012
rect 30012 6010 30068 6012
rect 30092 6010 30148 6012
rect 29852 5958 29898 6010
rect 29898 5958 29908 6010
rect 29932 5958 29962 6010
rect 29962 5958 29974 6010
rect 29974 5958 29988 6010
rect 30012 5958 30026 6010
rect 30026 5958 30038 6010
rect 30038 5958 30068 6010
rect 30092 5958 30102 6010
rect 30102 5958 30148 6010
rect 29852 5956 29908 5958
rect 29932 5956 29988 5958
rect 30012 5956 30068 5958
rect 30092 5956 30148 5958
rect 30746 20576 30802 20632
rect 30746 20304 30802 20360
rect 31022 22208 31078 22264
rect 31482 26288 31538 26344
rect 31574 26152 31630 26208
rect 31482 25220 31538 25256
rect 31482 25200 31484 25220
rect 31484 25200 31536 25220
rect 31536 25200 31538 25220
rect 32218 27376 32274 27432
rect 31298 24112 31354 24168
rect 31206 23432 31262 23488
rect 31206 19488 31262 19544
rect 30838 17992 30894 18048
rect 30654 17448 30710 17504
rect 30654 16768 30710 16824
rect 30654 15680 30710 15736
rect 30654 14728 30710 14784
rect 30930 16768 30986 16824
rect 30746 14476 30802 14512
rect 30746 14456 30748 14476
rect 30748 14456 30800 14476
rect 30800 14456 30802 14476
rect 30562 11736 30618 11792
rect 30562 10648 30618 10704
rect 30562 9560 30618 9616
rect 31022 15000 31078 15056
rect 30746 12416 30802 12472
rect 30746 11328 30802 11384
rect 30746 9832 30802 9888
rect 30562 8916 30564 8936
rect 30564 8916 30616 8936
rect 30616 8916 30618 8936
rect 30562 8880 30618 8916
rect 30562 8608 30618 8664
rect 30470 7792 30526 7848
rect 30654 7928 30710 7984
rect 31206 16768 31262 16824
rect 31114 13776 31170 13832
rect 31022 13368 31078 13424
rect 31482 22752 31538 22808
rect 31942 25064 31998 25120
rect 34058 27648 34114 27704
rect 32494 26324 32496 26344
rect 32496 26324 32548 26344
rect 32548 26324 32550 26344
rect 32494 26288 32550 26324
rect 32310 25064 32366 25120
rect 32310 24656 32366 24712
rect 32126 24112 32182 24168
rect 32034 23704 32090 23760
rect 31758 23024 31814 23080
rect 31942 21664 31998 21720
rect 32126 22752 32182 22808
rect 32402 22752 32458 22808
rect 32218 21256 32274 21312
rect 31850 17448 31906 17504
rect 31390 17060 31446 17096
rect 31390 17040 31392 17060
rect 31392 17040 31444 17060
rect 31444 17040 31446 17060
rect 31298 12688 31354 12744
rect 31574 16360 31630 16416
rect 31574 15272 31630 15328
rect 31482 12316 31484 12336
rect 31484 12316 31536 12336
rect 31536 12316 31538 12336
rect 31022 12008 31078 12064
rect 30930 11872 30986 11928
rect 30930 11600 30986 11656
rect 30930 7828 30932 7848
rect 30932 7828 30984 7848
rect 30984 7828 30986 7848
rect 30930 7792 30986 7828
rect 31022 7540 31078 7576
rect 31022 7520 31024 7540
rect 31024 7520 31076 7540
rect 31076 7520 31078 7540
rect 31114 7384 31170 7440
rect 31114 5616 31170 5672
rect 29852 4922 29908 4924
rect 29932 4922 29988 4924
rect 30012 4922 30068 4924
rect 30092 4922 30148 4924
rect 29852 4870 29898 4922
rect 29898 4870 29908 4922
rect 29932 4870 29962 4922
rect 29962 4870 29974 4922
rect 29974 4870 29988 4922
rect 30012 4870 30026 4922
rect 30026 4870 30038 4922
rect 30038 4870 30068 4922
rect 30092 4870 30102 4922
rect 30102 4870 30148 4922
rect 29852 4868 29908 4870
rect 29932 4868 29988 4870
rect 30012 4868 30068 4870
rect 30092 4868 30148 4870
rect 29852 3834 29908 3836
rect 29932 3834 29988 3836
rect 30012 3834 30068 3836
rect 30092 3834 30148 3836
rect 29852 3782 29898 3834
rect 29898 3782 29908 3834
rect 29932 3782 29962 3834
rect 29962 3782 29974 3834
rect 29974 3782 29988 3834
rect 30012 3782 30026 3834
rect 30026 3782 30038 3834
rect 30038 3782 30068 3834
rect 30092 3782 30102 3834
rect 30102 3782 30148 3834
rect 29852 3780 29908 3782
rect 29932 3780 29988 3782
rect 30012 3780 30068 3782
rect 30092 3780 30148 3782
rect 29852 2746 29908 2748
rect 29932 2746 29988 2748
rect 30012 2746 30068 2748
rect 30092 2746 30148 2748
rect 29852 2694 29898 2746
rect 29898 2694 29908 2746
rect 29932 2694 29962 2746
rect 29962 2694 29974 2746
rect 29974 2694 29988 2746
rect 30012 2694 30026 2746
rect 30026 2694 30038 2746
rect 30038 2694 30068 2746
rect 30092 2694 30102 2746
rect 30102 2694 30148 2746
rect 29852 2692 29908 2694
rect 29932 2692 29988 2694
rect 30012 2692 30068 2694
rect 30092 2692 30148 2694
rect 28446 1536 28502 1592
rect 31482 12280 31538 12316
rect 31850 17040 31906 17096
rect 32586 21936 32642 21992
rect 32954 23840 33010 23896
rect 33138 23432 33194 23488
rect 32494 21256 32550 21312
rect 32310 20712 32366 20768
rect 32218 19352 32274 19408
rect 31850 15272 31906 15328
rect 31666 14048 31722 14104
rect 31390 11464 31446 11520
rect 31942 13504 31998 13560
rect 31758 11600 31814 11656
rect 31574 11056 31630 11112
rect 31482 9288 31538 9344
rect 32494 17584 32550 17640
rect 32494 15408 32550 15464
rect 32678 20032 32734 20088
rect 33138 22344 33194 22400
rect 33138 22072 33194 22128
rect 33046 21664 33102 21720
rect 32954 20168 33010 20224
rect 32862 17720 32918 17776
rect 32770 17584 32826 17640
rect 32402 12860 32404 12880
rect 32404 12860 32456 12880
rect 32456 12860 32458 12880
rect 32402 12824 32458 12860
rect 31942 11192 31998 11248
rect 31942 9968 31998 10024
rect 31850 9832 31906 9888
rect 31850 9152 31906 9208
rect 31390 8780 31392 8800
rect 31392 8780 31444 8800
rect 31444 8780 31446 8800
rect 31390 8744 31446 8780
rect 32126 9832 32182 9888
rect 32126 9696 32182 9752
rect 31850 8608 31906 8664
rect 31666 8200 31722 8256
rect 32310 12416 32366 12472
rect 32310 11056 32366 11112
rect 32586 12416 32642 12472
rect 32494 9832 32550 9888
rect 31574 8064 31630 8120
rect 31390 7656 31446 7712
rect 32034 8064 32090 8120
rect 32218 8084 32274 8120
rect 32218 8064 32220 8084
rect 32220 8064 32272 8084
rect 32272 8064 32274 8084
rect 33046 19760 33102 19816
rect 34150 27396 34206 27432
rect 34150 27376 34152 27396
rect 34152 27376 34204 27396
rect 34204 27376 34206 27396
rect 33690 25744 33746 25800
rect 33506 24520 33562 24576
rect 33322 23568 33378 23624
rect 33230 20848 33286 20904
rect 34150 26288 34206 26344
rect 33966 26016 34022 26072
rect 33874 24148 33876 24168
rect 33876 24148 33928 24168
rect 33928 24148 33930 24168
rect 33874 24112 33930 24148
rect 33506 22752 33562 22808
rect 33690 21972 33692 21992
rect 33692 21972 33744 21992
rect 33744 21972 33746 21992
rect 33690 21936 33746 21972
rect 33414 20168 33470 20224
rect 33322 19624 33378 19680
rect 32862 12824 32918 12880
rect 32862 11464 32918 11520
rect 32678 10376 32734 10432
rect 34334 24928 34390 24984
rect 34058 24132 34114 24168
rect 34058 24112 34060 24132
rect 34060 24112 34112 24132
rect 34112 24112 34114 24132
rect 33874 23296 33930 23352
rect 33782 19896 33838 19952
rect 33598 19352 33654 19408
rect 33874 18128 33930 18184
rect 33874 16396 33876 16416
rect 33876 16396 33928 16416
rect 33928 16396 33930 16416
rect 33874 16360 33930 16396
rect 33046 10648 33102 10704
rect 33506 11872 33562 11928
rect 33046 9596 33048 9616
rect 33048 9596 33100 9616
rect 33100 9596 33102 9616
rect 33046 9560 33102 9596
rect 32862 8492 32918 8528
rect 32862 8472 32864 8492
rect 32864 8472 32916 8492
rect 32916 8472 32918 8492
rect 32586 8200 32642 8256
rect 33046 8200 33102 8256
rect 32862 5888 32918 5944
rect 33782 11192 33838 11248
rect 33782 10648 33838 10704
rect 33690 10376 33746 10432
rect 34426 23840 34482 23896
rect 34242 22888 34298 22944
rect 39118 29824 39174 29880
rect 37830 28056 37886 28112
rect 35070 25880 35126 25936
rect 35070 24656 35126 24712
rect 34242 20712 34298 20768
rect 34150 16940 34152 16960
rect 34152 16940 34204 16960
rect 34204 16940 34206 16960
rect 34150 16904 34206 16940
rect 34150 16768 34206 16824
rect 34150 13640 34206 13696
rect 34978 23976 35034 24032
rect 35070 23840 35126 23896
rect 35070 23024 35126 23080
rect 35806 26460 35808 26480
rect 35808 26460 35860 26480
rect 35860 26460 35862 26480
rect 35806 26424 35862 26460
rect 35530 25764 35586 25800
rect 35530 25744 35532 25764
rect 35532 25744 35584 25764
rect 35584 25744 35586 25764
rect 35714 25064 35770 25120
rect 35622 24928 35678 24984
rect 35530 24012 35532 24032
rect 35532 24012 35584 24032
rect 35584 24012 35586 24032
rect 35530 23976 35586 24012
rect 35346 22616 35402 22672
rect 35346 22072 35402 22128
rect 35070 21800 35126 21856
rect 34426 18672 34482 18728
rect 34702 18400 34758 18456
rect 34334 18264 34390 18320
rect 34334 18128 34390 18184
rect 34794 17992 34850 18048
rect 35162 19896 35218 19952
rect 35070 18400 35126 18456
rect 34702 17040 34758 17096
rect 34334 16768 34390 16824
rect 34426 15408 34482 15464
rect 34518 14356 34520 14376
rect 34520 14356 34572 14376
rect 34572 14356 34574 14376
rect 34518 14320 34574 14356
rect 33598 7928 33654 7984
rect 33874 9696 33930 9752
rect 34242 10376 34298 10432
rect 34150 9968 34206 10024
rect 33966 7828 33968 7848
rect 33968 7828 34020 7848
rect 34020 7828 34022 7848
rect 33966 7792 34022 7828
rect 34702 15136 34758 15192
rect 34702 13776 34758 13832
rect 34702 13504 34758 13560
rect 34794 11348 34850 11384
rect 34794 11328 34796 11348
rect 34796 11328 34848 11348
rect 34848 11328 34850 11348
rect 34610 10784 34666 10840
rect 34518 9696 34574 9752
rect 34426 9580 34482 9616
rect 34426 9560 34428 9580
rect 34428 9560 34480 9580
rect 34480 9560 34482 9580
rect 34150 8628 34206 8664
rect 34150 8608 34152 8628
rect 34152 8608 34204 8628
rect 34204 8608 34206 8628
rect 34978 14456 35034 14512
rect 34886 9968 34942 10024
rect 34702 9832 34758 9888
rect 35438 14456 35494 14512
rect 35254 13504 35310 13560
rect 35254 12844 35310 12880
rect 35254 12824 35256 12844
rect 35256 12824 35308 12844
rect 35308 12824 35310 12844
rect 35254 12552 35310 12608
rect 35162 11212 35218 11248
rect 35162 11192 35164 11212
rect 35164 11192 35216 11212
rect 35216 11192 35218 11212
rect 35254 10376 35310 10432
rect 34886 9560 34942 9616
rect 34886 9288 34942 9344
rect 35162 9424 35218 9480
rect 35070 9152 35126 9208
rect 35714 23568 35770 23624
rect 36174 24812 36230 24848
rect 36174 24792 36176 24812
rect 36176 24792 36228 24812
rect 36228 24792 36230 24812
rect 35990 24692 35992 24712
rect 35992 24692 36044 24712
rect 36044 24692 36046 24712
rect 35990 24656 36046 24692
rect 35898 23432 35954 23488
rect 35898 22752 35954 22808
rect 36174 23704 36230 23760
rect 36174 22228 36230 22264
rect 36174 22208 36176 22228
rect 36176 22208 36228 22228
rect 36228 22208 36230 22228
rect 35990 21936 36046 21992
rect 35806 21528 35862 21584
rect 35622 20168 35678 20224
rect 35714 19488 35770 19544
rect 35898 19488 35954 19544
rect 36542 23468 36544 23488
rect 36544 23468 36596 23488
rect 36596 23468 36598 23488
rect 36542 23432 36598 23468
rect 36910 24384 36966 24440
rect 37002 23976 37058 24032
rect 36818 23568 36874 23624
rect 37278 23840 37334 23896
rect 37646 25608 37702 25664
rect 36910 23296 36966 23352
rect 36726 22636 36782 22672
rect 36726 22616 36728 22636
rect 36728 22616 36780 22636
rect 36780 22616 36782 22636
rect 36726 22208 36782 22264
rect 37094 23296 37150 23352
rect 36174 18536 36230 18592
rect 35714 17040 35770 17096
rect 35806 16632 35862 16688
rect 35806 15544 35862 15600
rect 35714 15000 35770 15056
rect 35622 12688 35678 12744
rect 36634 20712 36690 20768
rect 36910 21256 36966 21312
rect 36726 18128 36782 18184
rect 36266 17584 36322 17640
rect 36266 15680 36322 15736
rect 36174 15000 36230 15056
rect 36174 14764 36176 14784
rect 36176 14764 36228 14784
rect 36228 14764 36230 14784
rect 36174 14728 36230 14764
rect 36818 17584 36874 17640
rect 36450 15444 36452 15464
rect 36452 15444 36504 15464
rect 36504 15444 36506 15464
rect 36450 15408 36506 15444
rect 35990 14184 36046 14240
rect 35990 13796 36046 13832
rect 35990 13776 35992 13796
rect 35992 13776 36044 13796
rect 36044 13776 36046 13796
rect 35990 12960 36046 13016
rect 35622 12552 35678 12608
rect 36450 14592 36506 14648
rect 35806 12280 35862 12336
rect 35714 11736 35770 11792
rect 35622 11600 35678 11656
rect 35806 11464 35862 11520
rect 35622 10920 35678 10976
rect 35530 10532 35586 10568
rect 35530 10512 35532 10532
rect 35532 10512 35584 10532
rect 35584 10512 35586 10532
rect 34978 8472 35034 8528
rect 34794 8064 34850 8120
rect 34518 7248 34574 7304
rect 36266 12688 36322 12744
rect 35990 10648 36046 10704
rect 36082 9968 36138 10024
rect 36634 14184 36690 14240
rect 36266 10804 36322 10840
rect 36266 10784 36268 10804
rect 36268 10784 36320 10804
rect 36320 10784 36322 10804
rect 36818 15816 36874 15872
rect 37186 20848 37242 20904
rect 37646 20460 37702 20496
rect 37646 20440 37648 20460
rect 37648 20440 37700 20460
rect 37700 20440 37702 20460
rect 37002 19216 37058 19272
rect 37462 19624 37518 19680
rect 37278 19216 37334 19272
rect 37462 18536 37518 18592
rect 37462 17992 37518 18048
rect 37370 16632 37426 16688
rect 37278 16496 37334 16552
rect 36726 13368 36782 13424
rect 36726 12724 36728 12744
rect 36728 12724 36780 12744
rect 36780 12724 36782 12744
rect 36726 12688 36782 12724
rect 36726 12416 36782 12472
rect 36910 12416 36966 12472
rect 36818 12280 36874 12336
rect 36174 8744 36230 8800
rect 35898 7520 35954 7576
rect 35438 6568 35494 6624
rect 38106 24928 38162 24984
rect 38106 21528 38162 21584
rect 37922 20304 37978 20360
rect 38566 24248 38622 24304
rect 38474 22888 38530 22944
rect 39484 27226 39540 27228
rect 39564 27226 39620 27228
rect 39644 27226 39700 27228
rect 39724 27226 39780 27228
rect 39484 27174 39530 27226
rect 39530 27174 39540 27226
rect 39564 27174 39594 27226
rect 39594 27174 39606 27226
rect 39606 27174 39620 27226
rect 39644 27174 39658 27226
rect 39658 27174 39670 27226
rect 39670 27174 39700 27226
rect 39724 27174 39734 27226
rect 39734 27174 39780 27226
rect 39484 27172 39540 27174
rect 39564 27172 39620 27174
rect 39644 27172 39700 27174
rect 39724 27172 39780 27174
rect 39484 26138 39540 26140
rect 39564 26138 39620 26140
rect 39644 26138 39700 26140
rect 39724 26138 39780 26140
rect 39484 26086 39530 26138
rect 39530 26086 39540 26138
rect 39564 26086 39594 26138
rect 39594 26086 39606 26138
rect 39606 26086 39620 26138
rect 39644 26086 39658 26138
rect 39658 26086 39670 26138
rect 39670 26086 39700 26138
rect 39724 26086 39734 26138
rect 39734 26086 39780 26138
rect 39484 26084 39540 26086
rect 39564 26084 39620 26086
rect 39644 26084 39700 26086
rect 39724 26084 39780 26086
rect 38842 23704 38898 23760
rect 38750 23180 38806 23216
rect 38750 23160 38752 23180
rect 38752 23160 38804 23180
rect 38804 23160 38806 23180
rect 38658 22888 38714 22944
rect 38566 20984 38622 21040
rect 38842 22072 38898 22128
rect 39026 22752 39082 22808
rect 38750 19352 38806 19408
rect 38658 19216 38714 19272
rect 38106 18536 38162 18592
rect 38474 18400 38530 18456
rect 38198 17312 38254 17368
rect 37462 16360 37518 16416
rect 37462 16124 37464 16144
rect 37464 16124 37516 16144
rect 37516 16124 37518 16144
rect 37462 16088 37518 16124
rect 37278 13232 37334 13288
rect 37370 12824 37426 12880
rect 37278 12144 37334 12200
rect 36818 11192 36874 11248
rect 37002 8744 37058 8800
rect 37646 15544 37702 15600
rect 38106 17176 38162 17232
rect 38290 16940 38292 16960
rect 38292 16940 38344 16960
rect 38344 16940 38346 16960
rect 38290 16904 38346 16940
rect 38014 16768 38070 16824
rect 39118 20748 39120 20768
rect 39120 20748 39172 20768
rect 39172 20748 39174 20768
rect 39118 20712 39174 20748
rect 39484 25050 39540 25052
rect 39564 25050 39620 25052
rect 39644 25050 39700 25052
rect 39724 25050 39780 25052
rect 39484 24998 39530 25050
rect 39530 24998 39540 25050
rect 39564 24998 39594 25050
rect 39594 24998 39606 25050
rect 39606 24998 39620 25050
rect 39644 24998 39658 25050
rect 39658 24998 39670 25050
rect 39670 24998 39700 25050
rect 39724 24998 39734 25050
rect 39734 24998 39780 25050
rect 39484 24996 39540 24998
rect 39564 24996 39620 24998
rect 39644 24996 39700 24998
rect 39724 24996 39780 24998
rect 39486 24556 39488 24576
rect 39488 24556 39540 24576
rect 39540 24556 39542 24576
rect 39486 24520 39542 24556
rect 39484 23962 39540 23964
rect 39564 23962 39620 23964
rect 39644 23962 39700 23964
rect 39724 23962 39780 23964
rect 39484 23910 39530 23962
rect 39530 23910 39540 23962
rect 39564 23910 39594 23962
rect 39594 23910 39606 23962
rect 39606 23910 39620 23962
rect 39644 23910 39658 23962
rect 39658 23910 39670 23962
rect 39670 23910 39700 23962
rect 39724 23910 39734 23962
rect 39734 23910 39780 23962
rect 39484 23908 39540 23910
rect 39564 23908 39620 23910
rect 39644 23908 39700 23910
rect 39724 23908 39780 23910
rect 39394 23160 39450 23216
rect 39484 22874 39540 22876
rect 39564 22874 39620 22876
rect 39644 22874 39700 22876
rect 39724 22874 39780 22876
rect 39484 22822 39530 22874
rect 39530 22822 39540 22874
rect 39564 22822 39594 22874
rect 39594 22822 39606 22874
rect 39606 22822 39620 22874
rect 39644 22822 39658 22874
rect 39658 22822 39670 22874
rect 39670 22822 39700 22874
rect 39724 22822 39734 22874
rect 39734 22822 39780 22874
rect 39484 22820 39540 22822
rect 39564 22820 39620 22822
rect 39644 22820 39700 22822
rect 39724 22820 39780 22822
rect 41510 29144 41566 29200
rect 40866 25200 40922 25256
rect 39578 22500 39634 22536
rect 39578 22480 39580 22500
rect 39580 22480 39632 22500
rect 39632 22480 39634 22500
rect 40498 23296 40554 23352
rect 40406 22616 40462 22672
rect 40038 22108 40040 22128
rect 40040 22108 40092 22128
rect 40092 22108 40094 22128
rect 40038 22072 40094 22108
rect 39302 20984 39358 21040
rect 39210 19932 39212 19952
rect 39212 19932 39264 19952
rect 39264 19932 39266 19952
rect 39210 19896 39266 19932
rect 39854 21936 39910 21992
rect 39484 21786 39540 21788
rect 39564 21786 39620 21788
rect 39644 21786 39700 21788
rect 39724 21786 39780 21788
rect 39484 21734 39530 21786
rect 39530 21734 39540 21786
rect 39564 21734 39594 21786
rect 39594 21734 39606 21786
rect 39606 21734 39620 21786
rect 39644 21734 39658 21786
rect 39658 21734 39670 21786
rect 39670 21734 39700 21786
rect 39724 21734 39734 21786
rect 39734 21734 39780 21786
rect 39484 21732 39540 21734
rect 39564 21732 39620 21734
rect 39644 21732 39700 21734
rect 39724 21732 39780 21734
rect 39484 20698 39540 20700
rect 39564 20698 39620 20700
rect 39644 20698 39700 20700
rect 39724 20698 39780 20700
rect 39484 20646 39530 20698
rect 39530 20646 39540 20698
rect 39564 20646 39594 20698
rect 39594 20646 39606 20698
rect 39606 20646 39620 20698
rect 39644 20646 39658 20698
rect 39658 20646 39670 20698
rect 39670 20646 39700 20698
rect 39724 20646 39734 20698
rect 39734 20646 39780 20698
rect 39484 20644 39540 20646
rect 39564 20644 39620 20646
rect 39644 20644 39700 20646
rect 39724 20644 39780 20646
rect 39762 20032 39818 20088
rect 39484 19610 39540 19612
rect 39564 19610 39620 19612
rect 39644 19610 39700 19612
rect 39724 19610 39780 19612
rect 39484 19558 39530 19610
rect 39530 19558 39540 19610
rect 39564 19558 39594 19610
rect 39594 19558 39606 19610
rect 39606 19558 39620 19610
rect 39644 19558 39658 19610
rect 39658 19558 39670 19610
rect 39670 19558 39700 19610
rect 39724 19558 39734 19610
rect 39734 19558 39780 19610
rect 39484 19556 39540 19558
rect 39564 19556 39620 19558
rect 39644 19556 39700 19558
rect 39724 19556 39780 19558
rect 39302 18264 39358 18320
rect 39302 18128 39358 18184
rect 39486 18808 39542 18864
rect 39484 18522 39540 18524
rect 39564 18522 39620 18524
rect 39644 18522 39700 18524
rect 39724 18522 39780 18524
rect 39484 18470 39530 18522
rect 39530 18470 39540 18522
rect 39564 18470 39594 18522
rect 39594 18470 39606 18522
rect 39606 18470 39620 18522
rect 39644 18470 39658 18522
rect 39658 18470 39670 18522
rect 39670 18470 39700 18522
rect 39724 18470 39734 18522
rect 39734 18470 39780 18522
rect 39484 18468 39540 18470
rect 39564 18468 39620 18470
rect 39644 18468 39700 18470
rect 39724 18468 39780 18470
rect 40590 21392 40646 21448
rect 40498 21120 40554 21176
rect 40406 20440 40462 20496
rect 40130 19760 40186 19816
rect 40038 19624 40094 19680
rect 39118 17040 39174 17096
rect 38750 16224 38806 16280
rect 38290 13504 38346 13560
rect 37830 12688 37886 12744
rect 37370 8628 37426 8664
rect 37370 8608 37372 8628
rect 37372 8608 37424 8628
rect 37424 8608 37426 8628
rect 37094 8200 37150 8256
rect 37646 11500 37648 11520
rect 37648 11500 37700 11520
rect 37700 11500 37702 11520
rect 37646 11464 37702 11500
rect 37830 10920 37886 10976
rect 38014 12688 38070 12744
rect 37830 10004 37832 10024
rect 37832 10004 37884 10024
rect 37884 10004 37886 10024
rect 37830 9968 37886 10004
rect 38106 11464 38162 11520
rect 37278 5092 37334 5128
rect 37278 5072 37280 5092
rect 37280 5072 37332 5092
rect 37332 5072 37334 5092
rect 37738 3304 37794 3360
rect 39026 16224 39082 16280
rect 38750 15408 38806 15464
rect 38474 14048 38530 14104
rect 38658 14184 38714 14240
rect 38842 14184 38898 14240
rect 38658 13776 38714 13832
rect 38750 12824 38806 12880
rect 38658 12280 38714 12336
rect 38658 11056 38714 11112
rect 38934 12708 38990 12744
rect 38934 12688 38936 12708
rect 38936 12688 38988 12708
rect 38988 12688 38990 12708
rect 38842 11348 38898 11384
rect 38842 11328 38844 11348
rect 38844 11328 38896 11348
rect 38896 11328 38898 11348
rect 38934 10124 38990 10160
rect 38934 10104 38936 10124
rect 38936 10104 38988 10124
rect 38988 10104 38990 10124
rect 40130 18536 40186 18592
rect 39484 17434 39540 17436
rect 39564 17434 39620 17436
rect 39644 17434 39700 17436
rect 39724 17434 39780 17436
rect 39484 17382 39530 17434
rect 39530 17382 39540 17434
rect 39564 17382 39594 17434
rect 39594 17382 39606 17434
rect 39606 17382 39620 17434
rect 39644 17382 39658 17434
rect 39658 17382 39670 17434
rect 39670 17382 39700 17434
rect 39724 17382 39734 17434
rect 39734 17382 39780 17434
rect 39484 17380 39540 17382
rect 39564 17380 39620 17382
rect 39644 17380 39700 17382
rect 39724 17380 39780 17382
rect 39946 17448 40002 17504
rect 39484 16346 39540 16348
rect 39564 16346 39620 16348
rect 39644 16346 39700 16348
rect 39724 16346 39780 16348
rect 39484 16294 39530 16346
rect 39530 16294 39540 16346
rect 39564 16294 39594 16346
rect 39594 16294 39606 16346
rect 39606 16294 39620 16346
rect 39644 16294 39658 16346
rect 39658 16294 39670 16346
rect 39670 16294 39700 16346
rect 39724 16294 39734 16346
rect 39734 16294 39780 16346
rect 39484 16292 39540 16294
rect 39564 16292 39620 16294
rect 39644 16292 39700 16294
rect 39724 16292 39780 16294
rect 39210 13912 39266 13968
rect 39484 15258 39540 15260
rect 39564 15258 39620 15260
rect 39644 15258 39700 15260
rect 39724 15258 39780 15260
rect 39484 15206 39530 15258
rect 39530 15206 39540 15258
rect 39564 15206 39594 15258
rect 39594 15206 39606 15258
rect 39606 15206 39620 15258
rect 39644 15206 39658 15258
rect 39658 15206 39670 15258
rect 39670 15206 39700 15258
rect 39724 15206 39734 15258
rect 39734 15206 39780 15258
rect 39484 15204 39540 15206
rect 39564 15204 39620 15206
rect 39644 15204 39700 15206
rect 39724 15204 39780 15206
rect 39854 14864 39910 14920
rect 40130 15952 40186 16008
rect 40222 15816 40278 15872
rect 39762 14728 39818 14784
rect 39762 14456 39818 14512
rect 39762 14356 39764 14376
rect 39764 14356 39816 14376
rect 39816 14356 39818 14376
rect 39762 14320 39818 14356
rect 39484 14170 39540 14172
rect 39564 14170 39620 14172
rect 39644 14170 39700 14172
rect 39724 14170 39780 14172
rect 39484 14118 39530 14170
rect 39530 14118 39540 14170
rect 39564 14118 39594 14170
rect 39594 14118 39606 14170
rect 39606 14118 39620 14170
rect 39644 14118 39658 14170
rect 39658 14118 39670 14170
rect 39670 14118 39700 14170
rect 39724 14118 39734 14170
rect 39734 14118 39780 14170
rect 39484 14116 39540 14118
rect 39564 14116 39620 14118
rect 39644 14116 39700 14118
rect 39724 14116 39780 14118
rect 39302 12688 39358 12744
rect 39302 12416 39358 12472
rect 39484 13082 39540 13084
rect 39564 13082 39620 13084
rect 39644 13082 39700 13084
rect 39724 13082 39780 13084
rect 39484 13030 39530 13082
rect 39530 13030 39540 13082
rect 39564 13030 39594 13082
rect 39594 13030 39606 13082
rect 39606 13030 39620 13082
rect 39644 13030 39658 13082
rect 39658 13030 39670 13082
rect 39670 13030 39700 13082
rect 39724 13030 39734 13082
rect 39734 13030 39780 13082
rect 39484 13028 39540 13030
rect 39564 13028 39620 13030
rect 39644 13028 39700 13030
rect 39724 13028 39780 13030
rect 39486 12416 39542 12472
rect 40130 14184 40186 14240
rect 40130 14068 40186 14104
rect 40130 14048 40132 14068
rect 40132 14048 40184 14068
rect 40184 14048 40186 14068
rect 40130 13932 40186 13968
rect 40130 13912 40132 13932
rect 40132 13912 40184 13932
rect 40184 13912 40186 13932
rect 40038 13640 40094 13696
rect 40038 12860 40040 12880
rect 40040 12860 40092 12880
rect 40092 12860 40094 12880
rect 40038 12824 40094 12860
rect 39484 11994 39540 11996
rect 39564 11994 39620 11996
rect 39644 11994 39700 11996
rect 39724 11994 39780 11996
rect 39484 11942 39530 11994
rect 39530 11942 39540 11994
rect 39564 11942 39594 11994
rect 39594 11942 39606 11994
rect 39606 11942 39620 11994
rect 39644 11942 39658 11994
rect 39658 11942 39670 11994
rect 39670 11942 39700 11994
rect 39724 11942 39734 11994
rect 39734 11942 39780 11994
rect 39484 11940 39540 11942
rect 39564 11940 39620 11942
rect 39644 11940 39700 11942
rect 39724 11940 39780 11942
rect 39484 10906 39540 10908
rect 39564 10906 39620 10908
rect 39644 10906 39700 10908
rect 39724 10906 39780 10908
rect 39484 10854 39530 10906
rect 39530 10854 39540 10906
rect 39564 10854 39594 10906
rect 39594 10854 39606 10906
rect 39606 10854 39620 10906
rect 39644 10854 39658 10906
rect 39658 10854 39670 10906
rect 39670 10854 39700 10906
rect 39724 10854 39734 10906
rect 39734 10854 39780 10906
rect 39484 10852 39540 10854
rect 39564 10852 39620 10854
rect 39644 10852 39700 10854
rect 39724 10852 39780 10854
rect 39484 9818 39540 9820
rect 39564 9818 39620 9820
rect 39644 9818 39700 9820
rect 39724 9818 39780 9820
rect 39484 9766 39530 9818
rect 39530 9766 39540 9818
rect 39564 9766 39594 9818
rect 39594 9766 39606 9818
rect 39606 9766 39620 9818
rect 39644 9766 39658 9818
rect 39658 9766 39670 9818
rect 39670 9766 39700 9818
rect 39724 9766 39734 9818
rect 39734 9766 39780 9818
rect 39484 9764 39540 9766
rect 39564 9764 39620 9766
rect 39644 9764 39700 9766
rect 39724 9764 39780 9766
rect 39484 8730 39540 8732
rect 39564 8730 39620 8732
rect 39644 8730 39700 8732
rect 39724 8730 39780 8732
rect 39484 8678 39530 8730
rect 39530 8678 39540 8730
rect 39564 8678 39594 8730
rect 39594 8678 39606 8730
rect 39606 8678 39620 8730
rect 39644 8678 39658 8730
rect 39658 8678 39670 8730
rect 39670 8678 39700 8730
rect 39724 8678 39734 8730
rect 39734 8678 39780 8730
rect 39484 8676 39540 8678
rect 39564 8676 39620 8678
rect 39644 8676 39700 8678
rect 39724 8676 39780 8678
rect 39484 7642 39540 7644
rect 39564 7642 39620 7644
rect 39644 7642 39700 7644
rect 39724 7642 39780 7644
rect 39484 7590 39530 7642
rect 39530 7590 39540 7642
rect 39564 7590 39594 7642
rect 39594 7590 39606 7642
rect 39606 7590 39620 7642
rect 39644 7590 39658 7642
rect 39658 7590 39670 7642
rect 39670 7590 39700 7642
rect 39724 7590 39734 7642
rect 39734 7590 39780 7642
rect 39484 7588 39540 7590
rect 39564 7588 39620 7590
rect 39644 7588 39700 7590
rect 39724 7588 39780 7590
rect 40406 18400 40462 18456
rect 40774 23568 40830 23624
rect 44362 29008 44418 29064
rect 43350 27648 43406 27704
rect 43166 25880 43222 25936
rect 41510 21936 41566 21992
rect 41050 19796 41052 19816
rect 41052 19796 41104 19816
rect 41104 19796 41106 19816
rect 41050 19760 41106 19796
rect 40958 19352 41014 19408
rect 40958 18128 41014 18184
rect 41326 18400 41382 18456
rect 41602 19352 41658 19408
rect 41602 18536 41658 18592
rect 41510 18264 41566 18320
rect 41418 18028 41420 18048
rect 41420 18028 41472 18048
rect 41472 18028 41474 18048
rect 41418 17992 41474 18028
rect 41142 17312 41198 17368
rect 40958 15680 41014 15736
rect 40866 15408 40922 15464
rect 41326 17176 41382 17232
rect 41970 23024 42026 23080
rect 41878 22208 41934 22264
rect 41694 17992 41750 18048
rect 42154 21528 42210 21584
rect 42062 21140 42118 21176
rect 42062 21120 42064 21140
rect 42064 21120 42116 21140
rect 42116 21120 42118 21140
rect 42246 20984 42302 21040
rect 42062 18264 42118 18320
rect 41510 17584 41566 17640
rect 41786 17620 41788 17640
rect 41788 17620 41840 17640
rect 41840 17620 41842 17640
rect 41786 17584 41842 17620
rect 41694 17040 41750 17096
rect 40866 14900 40868 14920
rect 40868 14900 40920 14920
rect 40920 14900 40922 14920
rect 40866 14864 40922 14900
rect 40498 12688 40554 12744
rect 40406 12552 40462 12608
rect 40958 14728 41014 14784
rect 40682 13912 40738 13968
rect 40406 12316 40408 12336
rect 40408 12316 40460 12336
rect 40460 12316 40462 12336
rect 40406 12280 40462 12316
rect 40314 11736 40370 11792
rect 40498 11736 40554 11792
rect 40498 11464 40554 11520
rect 41234 14456 41290 14512
rect 41326 13776 41382 13832
rect 41418 12008 41474 12064
rect 42246 17312 42302 17368
rect 42062 16632 42118 16688
rect 41970 16224 42026 16280
rect 41418 10240 41474 10296
rect 41510 9560 41566 9616
rect 41602 7384 41658 7440
rect 40130 6704 40186 6760
rect 39484 6554 39540 6556
rect 39564 6554 39620 6556
rect 39644 6554 39700 6556
rect 39724 6554 39780 6556
rect 39484 6502 39530 6554
rect 39530 6502 39540 6554
rect 39564 6502 39594 6554
rect 39594 6502 39606 6554
rect 39606 6502 39620 6554
rect 39644 6502 39658 6554
rect 39658 6502 39670 6554
rect 39670 6502 39700 6554
rect 39724 6502 39734 6554
rect 39734 6502 39780 6554
rect 39484 6500 39540 6502
rect 39564 6500 39620 6502
rect 39644 6500 39700 6502
rect 39724 6500 39780 6502
rect 39484 5466 39540 5468
rect 39564 5466 39620 5468
rect 39644 5466 39700 5468
rect 39724 5466 39780 5468
rect 39484 5414 39530 5466
rect 39530 5414 39540 5466
rect 39564 5414 39594 5466
rect 39594 5414 39606 5466
rect 39606 5414 39620 5466
rect 39644 5414 39658 5466
rect 39658 5414 39670 5466
rect 39670 5414 39700 5466
rect 39724 5414 39734 5466
rect 39734 5414 39780 5466
rect 39484 5412 39540 5414
rect 39564 5412 39620 5414
rect 39644 5412 39700 5414
rect 39724 5412 39780 5414
rect 42062 11736 42118 11792
rect 42614 20168 42670 20224
rect 42522 19760 42578 19816
rect 42706 19372 42762 19408
rect 42706 19352 42708 19372
rect 42708 19352 42760 19372
rect 42760 19352 42762 19372
rect 42430 17992 42486 18048
rect 42798 18672 42854 18728
rect 43166 20304 43222 20360
rect 43258 19896 43314 19952
rect 43258 19080 43314 19136
rect 42706 17856 42762 17912
rect 43258 18536 43314 18592
rect 43074 17720 43130 17776
rect 42798 17040 42854 17096
rect 42982 17040 43038 17096
rect 42890 16904 42946 16960
rect 42430 15272 42486 15328
rect 42338 13776 42394 13832
rect 43258 18128 43314 18184
rect 42890 15136 42946 15192
rect 43166 11328 43222 11384
rect 43442 26424 43498 26480
rect 43534 20848 43590 20904
rect 43902 18944 43958 19000
rect 43994 18400 44050 18456
rect 44178 16768 44234 16824
rect 43350 13268 43352 13288
rect 43352 13268 43404 13288
rect 43404 13268 43406 13288
rect 43350 13232 43406 13268
rect 43718 11600 43774 11656
rect 44178 15544 44234 15600
rect 43994 15408 44050 15464
rect 43994 15308 43996 15328
rect 43996 15308 44048 15328
rect 44048 15308 44050 15328
rect 43994 15272 44050 15308
rect 44178 15156 44234 15192
rect 44178 15136 44180 15156
rect 44180 15136 44232 15156
rect 44232 15136 44234 15156
rect 44638 28872 44694 28928
rect 44454 25744 44510 25800
rect 49116 27770 49172 27772
rect 49196 27770 49252 27772
rect 49276 27770 49332 27772
rect 49356 27770 49412 27772
rect 49116 27718 49162 27770
rect 49162 27718 49172 27770
rect 49196 27718 49226 27770
rect 49226 27718 49238 27770
rect 49238 27718 49252 27770
rect 49276 27718 49290 27770
rect 49290 27718 49302 27770
rect 49302 27718 49332 27770
rect 49356 27718 49366 27770
rect 49366 27718 49412 27770
rect 49116 27716 49172 27718
rect 49196 27716 49252 27718
rect 49276 27716 49332 27718
rect 49356 27716 49412 27718
rect 52458 27412 52460 27432
rect 52460 27412 52512 27432
rect 52512 27412 52514 27432
rect 44546 19352 44602 19408
rect 44270 14864 44326 14920
rect 44914 21256 44970 21312
rect 45190 23160 45246 23216
rect 44362 12416 44418 12472
rect 44730 16360 44786 16416
rect 45098 17876 45154 17912
rect 45098 17856 45100 17876
rect 45100 17856 45152 17876
rect 45152 17856 45154 17876
rect 45006 16652 45062 16688
rect 45006 16632 45008 16652
rect 45008 16632 45060 16652
rect 45060 16632 45062 16652
rect 44914 15272 44970 15328
rect 44822 14592 44878 14648
rect 44546 10648 44602 10704
rect 39484 4378 39540 4380
rect 39564 4378 39620 4380
rect 39644 4378 39700 4380
rect 39724 4378 39780 4380
rect 39484 4326 39530 4378
rect 39530 4326 39540 4378
rect 39564 4326 39594 4378
rect 39594 4326 39606 4378
rect 39606 4326 39620 4378
rect 39644 4326 39658 4378
rect 39658 4326 39670 4378
rect 39670 4326 39700 4378
rect 39724 4326 39734 4378
rect 39734 4326 39780 4378
rect 39484 4324 39540 4326
rect 39564 4324 39620 4326
rect 39644 4324 39700 4326
rect 39724 4324 39780 4326
rect 45190 16768 45246 16824
rect 45374 17040 45430 17096
rect 45282 14884 45338 14920
rect 45282 14864 45284 14884
rect 45284 14864 45336 14884
rect 45336 14864 45338 14884
rect 45190 12144 45246 12200
rect 39484 3290 39540 3292
rect 39564 3290 39620 3292
rect 39644 3290 39700 3292
rect 39724 3290 39780 3292
rect 39484 3238 39530 3290
rect 39530 3238 39540 3290
rect 39564 3238 39594 3290
rect 39594 3238 39606 3290
rect 39606 3238 39620 3290
rect 39644 3238 39658 3290
rect 39658 3238 39670 3290
rect 39670 3238 39700 3290
rect 39724 3238 39734 3290
rect 39734 3238 39780 3290
rect 39484 3236 39540 3238
rect 39564 3236 39620 3238
rect 39644 3236 39700 3238
rect 39724 3236 39780 3238
rect 39484 2202 39540 2204
rect 39564 2202 39620 2204
rect 39644 2202 39700 2204
rect 39724 2202 39780 2204
rect 39484 2150 39530 2202
rect 39530 2150 39540 2202
rect 39564 2150 39594 2202
rect 39594 2150 39606 2202
rect 39606 2150 39620 2202
rect 39644 2150 39658 2202
rect 39658 2150 39670 2202
rect 39670 2150 39700 2202
rect 39724 2150 39734 2202
rect 39734 2150 39780 2202
rect 39484 2148 39540 2150
rect 39564 2148 39620 2150
rect 39644 2148 39700 2150
rect 39724 2148 39780 2150
rect 38014 1672 38070 1728
rect 52458 27376 52514 27412
rect 57242 29144 57298 29200
rect 58070 27396 58126 27432
rect 58070 27376 58072 27396
rect 58072 27376 58124 27396
rect 58124 27376 58126 27396
rect 57886 26968 57942 27024
rect 49116 26682 49172 26684
rect 49196 26682 49252 26684
rect 49276 26682 49332 26684
rect 49356 26682 49412 26684
rect 49116 26630 49162 26682
rect 49162 26630 49172 26682
rect 49196 26630 49226 26682
rect 49226 26630 49238 26682
rect 49238 26630 49252 26682
rect 49276 26630 49290 26682
rect 49290 26630 49302 26682
rect 49302 26630 49332 26682
rect 49356 26630 49366 26682
rect 49366 26630 49412 26682
rect 49116 26628 49172 26630
rect 49196 26628 49252 26630
rect 49276 26628 49332 26630
rect 49356 26628 49412 26630
rect 46294 24520 46350 24576
rect 45650 18572 45652 18592
rect 45652 18572 45704 18592
rect 45704 18572 45706 18592
rect 45650 18536 45706 18572
rect 46110 18420 46166 18456
rect 46110 18400 46112 18420
rect 46112 18400 46164 18420
rect 46164 18400 46166 18420
rect 46018 17584 46074 17640
rect 45558 15816 45614 15872
rect 46018 15852 46020 15872
rect 46020 15852 46072 15872
rect 46072 15852 46074 15872
rect 46018 15816 46074 15852
rect 49116 25594 49172 25596
rect 49196 25594 49252 25596
rect 49276 25594 49332 25596
rect 49356 25594 49412 25596
rect 49116 25542 49162 25594
rect 49162 25542 49172 25594
rect 49196 25542 49226 25594
rect 49226 25542 49238 25594
rect 49238 25542 49252 25594
rect 49276 25542 49290 25594
rect 49290 25542 49302 25594
rect 49302 25542 49332 25594
rect 49356 25542 49366 25594
rect 49366 25542 49412 25594
rect 49116 25540 49172 25542
rect 49196 25540 49252 25542
rect 49276 25540 49332 25542
rect 49356 25540 49412 25542
rect 49116 24506 49172 24508
rect 49196 24506 49252 24508
rect 49276 24506 49332 24508
rect 49356 24506 49412 24508
rect 49116 24454 49162 24506
rect 49162 24454 49172 24506
rect 49196 24454 49226 24506
rect 49226 24454 49238 24506
rect 49238 24454 49252 24506
rect 49276 24454 49290 24506
rect 49290 24454 49302 24506
rect 49302 24454 49332 24506
rect 49356 24454 49366 24506
rect 49366 24454 49412 24506
rect 49116 24452 49172 24454
rect 49196 24452 49252 24454
rect 49276 24452 49332 24454
rect 49356 24452 49412 24454
rect 49116 23418 49172 23420
rect 49196 23418 49252 23420
rect 49276 23418 49332 23420
rect 49356 23418 49412 23420
rect 49116 23366 49162 23418
rect 49162 23366 49172 23418
rect 49196 23366 49226 23418
rect 49226 23366 49238 23418
rect 49238 23366 49252 23418
rect 49276 23366 49290 23418
rect 49290 23366 49302 23418
rect 49302 23366 49332 23418
rect 49356 23366 49366 23418
rect 49366 23366 49412 23418
rect 49116 23364 49172 23366
rect 49196 23364 49252 23366
rect 49276 23364 49332 23366
rect 49356 23364 49412 23366
rect 48778 22480 48834 22536
rect 47766 19660 47768 19680
rect 47768 19660 47820 19680
rect 47820 19660 47822 19680
rect 47766 19624 47822 19660
rect 48502 19760 48558 19816
rect 48410 18536 48466 18592
rect 48318 18284 48374 18320
rect 48318 18264 48320 18284
rect 48320 18264 48372 18284
rect 48372 18264 48374 18284
rect 46478 16632 46534 16688
rect 47122 17448 47178 17504
rect 48134 17448 48190 17504
rect 47030 16768 47086 16824
rect 46938 15036 46940 15056
rect 46940 15036 46992 15056
rect 46992 15036 46994 15056
rect 46938 15000 46994 15036
rect 45834 10512 45890 10568
rect 47306 16224 47362 16280
rect 47214 15544 47270 15600
rect 48134 16224 48190 16280
rect 48318 16360 48374 16416
rect 47030 3984 47086 4040
rect 48134 6160 48190 6216
rect 47214 3576 47270 3632
rect 49116 22330 49172 22332
rect 49196 22330 49252 22332
rect 49276 22330 49332 22332
rect 49356 22330 49412 22332
rect 49116 22278 49162 22330
rect 49162 22278 49172 22330
rect 49196 22278 49226 22330
rect 49226 22278 49238 22330
rect 49238 22278 49252 22330
rect 49276 22278 49290 22330
rect 49290 22278 49302 22330
rect 49302 22278 49332 22330
rect 49356 22278 49366 22330
rect 49366 22278 49412 22330
rect 49116 22276 49172 22278
rect 49196 22276 49252 22278
rect 49276 22276 49332 22278
rect 49356 22276 49412 22278
rect 49116 21242 49172 21244
rect 49196 21242 49252 21244
rect 49276 21242 49332 21244
rect 49356 21242 49412 21244
rect 49116 21190 49162 21242
rect 49162 21190 49172 21242
rect 49196 21190 49226 21242
rect 49226 21190 49238 21242
rect 49238 21190 49252 21242
rect 49276 21190 49290 21242
rect 49290 21190 49302 21242
rect 49302 21190 49332 21242
rect 49356 21190 49366 21242
rect 49366 21190 49412 21242
rect 49116 21188 49172 21190
rect 49196 21188 49252 21190
rect 49276 21188 49332 21190
rect 49356 21188 49412 21190
rect 49116 20154 49172 20156
rect 49196 20154 49252 20156
rect 49276 20154 49332 20156
rect 49356 20154 49412 20156
rect 49116 20102 49162 20154
rect 49162 20102 49172 20154
rect 49196 20102 49226 20154
rect 49226 20102 49238 20154
rect 49238 20102 49252 20154
rect 49276 20102 49290 20154
rect 49290 20102 49302 20154
rect 49302 20102 49332 20154
rect 49356 20102 49366 20154
rect 49366 20102 49412 20154
rect 49116 20100 49172 20102
rect 49196 20100 49252 20102
rect 49276 20100 49332 20102
rect 49356 20100 49412 20102
rect 58162 25608 58218 25664
rect 58162 23860 58218 23896
rect 58162 23840 58164 23860
rect 58164 23840 58216 23860
rect 58216 23840 58218 23860
rect 58162 22072 58218 22128
rect 58162 20304 58218 20360
rect 49116 19066 49172 19068
rect 49196 19066 49252 19068
rect 49276 19066 49332 19068
rect 49356 19066 49412 19068
rect 49116 19014 49162 19066
rect 49162 19014 49172 19066
rect 49196 19014 49226 19066
rect 49226 19014 49238 19066
rect 49238 19014 49252 19066
rect 49276 19014 49290 19066
rect 49290 19014 49302 19066
rect 49302 19014 49332 19066
rect 49356 19014 49366 19066
rect 49366 19014 49412 19066
rect 49116 19012 49172 19014
rect 49196 19012 49252 19014
rect 49276 19012 49332 19014
rect 49356 19012 49412 19014
rect 49116 17978 49172 17980
rect 49196 17978 49252 17980
rect 49276 17978 49332 17980
rect 49356 17978 49412 17980
rect 49116 17926 49162 17978
rect 49162 17926 49172 17978
rect 49196 17926 49226 17978
rect 49226 17926 49238 17978
rect 49238 17926 49252 17978
rect 49276 17926 49290 17978
rect 49290 17926 49302 17978
rect 49302 17926 49332 17978
rect 49356 17926 49366 17978
rect 49366 17926 49412 17978
rect 49116 17924 49172 17926
rect 49196 17924 49252 17926
rect 49276 17924 49332 17926
rect 49356 17924 49412 17926
rect 49116 16890 49172 16892
rect 49196 16890 49252 16892
rect 49276 16890 49332 16892
rect 49356 16890 49412 16892
rect 49116 16838 49162 16890
rect 49162 16838 49172 16890
rect 49196 16838 49226 16890
rect 49226 16838 49238 16890
rect 49238 16838 49252 16890
rect 49276 16838 49290 16890
rect 49290 16838 49302 16890
rect 49302 16838 49332 16890
rect 49356 16838 49366 16890
rect 49366 16838 49412 16890
rect 49116 16836 49172 16838
rect 49196 16836 49252 16838
rect 49276 16836 49332 16838
rect 49356 16836 49412 16838
rect 50158 17176 50214 17232
rect 49790 16108 49846 16144
rect 49790 16088 49792 16108
rect 49792 16088 49844 16108
rect 49844 16088 49846 16108
rect 49116 15802 49172 15804
rect 49196 15802 49252 15804
rect 49276 15802 49332 15804
rect 49356 15802 49412 15804
rect 49116 15750 49162 15802
rect 49162 15750 49172 15802
rect 49196 15750 49226 15802
rect 49226 15750 49238 15802
rect 49238 15750 49252 15802
rect 49276 15750 49290 15802
rect 49290 15750 49302 15802
rect 49302 15750 49332 15802
rect 49356 15750 49366 15802
rect 49366 15750 49412 15802
rect 49116 15748 49172 15750
rect 49196 15748 49252 15750
rect 49276 15748 49332 15750
rect 49356 15748 49412 15750
rect 49116 14714 49172 14716
rect 49196 14714 49252 14716
rect 49276 14714 49332 14716
rect 49356 14714 49412 14716
rect 49116 14662 49162 14714
rect 49162 14662 49172 14714
rect 49196 14662 49226 14714
rect 49226 14662 49238 14714
rect 49238 14662 49252 14714
rect 49276 14662 49290 14714
rect 49290 14662 49302 14714
rect 49302 14662 49332 14714
rect 49356 14662 49366 14714
rect 49366 14662 49412 14714
rect 49116 14660 49172 14662
rect 49196 14660 49252 14662
rect 49276 14660 49332 14662
rect 49356 14660 49412 14662
rect 49116 13626 49172 13628
rect 49196 13626 49252 13628
rect 49276 13626 49332 13628
rect 49356 13626 49412 13628
rect 49116 13574 49162 13626
rect 49162 13574 49172 13626
rect 49196 13574 49226 13626
rect 49226 13574 49238 13626
rect 49238 13574 49252 13626
rect 49276 13574 49290 13626
rect 49290 13574 49302 13626
rect 49302 13574 49332 13626
rect 49356 13574 49366 13626
rect 49366 13574 49412 13626
rect 49116 13572 49172 13574
rect 49196 13572 49252 13574
rect 49276 13572 49332 13574
rect 49356 13572 49412 13574
rect 49116 12538 49172 12540
rect 49196 12538 49252 12540
rect 49276 12538 49332 12540
rect 49356 12538 49412 12540
rect 49116 12486 49162 12538
rect 49162 12486 49172 12538
rect 49196 12486 49226 12538
rect 49226 12486 49238 12538
rect 49238 12486 49252 12538
rect 49276 12486 49290 12538
rect 49290 12486 49302 12538
rect 49302 12486 49332 12538
rect 49356 12486 49366 12538
rect 49366 12486 49412 12538
rect 49116 12484 49172 12486
rect 49196 12484 49252 12486
rect 49276 12484 49332 12486
rect 49356 12484 49412 12486
rect 49116 11450 49172 11452
rect 49196 11450 49252 11452
rect 49276 11450 49332 11452
rect 49356 11450 49412 11452
rect 49116 11398 49162 11450
rect 49162 11398 49172 11450
rect 49196 11398 49226 11450
rect 49226 11398 49238 11450
rect 49238 11398 49252 11450
rect 49276 11398 49290 11450
rect 49290 11398 49302 11450
rect 49302 11398 49332 11450
rect 49356 11398 49366 11450
rect 49366 11398 49412 11450
rect 49116 11396 49172 11398
rect 49196 11396 49252 11398
rect 49276 11396 49332 11398
rect 49356 11396 49412 11398
rect 49116 10362 49172 10364
rect 49196 10362 49252 10364
rect 49276 10362 49332 10364
rect 49356 10362 49412 10364
rect 49116 10310 49162 10362
rect 49162 10310 49172 10362
rect 49196 10310 49226 10362
rect 49226 10310 49238 10362
rect 49238 10310 49252 10362
rect 49276 10310 49290 10362
rect 49290 10310 49302 10362
rect 49302 10310 49332 10362
rect 49356 10310 49366 10362
rect 49366 10310 49412 10362
rect 49116 10308 49172 10310
rect 49196 10308 49252 10310
rect 49276 10308 49332 10310
rect 49356 10308 49412 10310
rect 49116 9274 49172 9276
rect 49196 9274 49252 9276
rect 49276 9274 49332 9276
rect 49356 9274 49412 9276
rect 49116 9222 49162 9274
rect 49162 9222 49172 9274
rect 49196 9222 49226 9274
rect 49226 9222 49238 9274
rect 49238 9222 49252 9274
rect 49276 9222 49290 9274
rect 49290 9222 49302 9274
rect 49302 9222 49332 9274
rect 49356 9222 49366 9274
rect 49366 9222 49412 9274
rect 49116 9220 49172 9222
rect 49196 9220 49252 9222
rect 49276 9220 49332 9222
rect 49356 9220 49412 9222
rect 49116 8186 49172 8188
rect 49196 8186 49252 8188
rect 49276 8186 49332 8188
rect 49356 8186 49412 8188
rect 49116 8134 49162 8186
rect 49162 8134 49172 8186
rect 49196 8134 49226 8186
rect 49226 8134 49238 8186
rect 49238 8134 49252 8186
rect 49276 8134 49290 8186
rect 49290 8134 49302 8186
rect 49302 8134 49332 8186
rect 49356 8134 49366 8186
rect 49366 8134 49412 8186
rect 49116 8132 49172 8134
rect 49196 8132 49252 8134
rect 49276 8132 49332 8134
rect 49356 8132 49412 8134
rect 58162 18536 58218 18592
rect 58162 16768 58218 16824
rect 58162 15036 58164 15056
rect 58164 15036 58216 15056
rect 58216 15036 58218 15056
rect 58162 15000 58218 15036
rect 57886 14456 57942 14512
rect 58162 13268 58164 13288
rect 58164 13268 58216 13288
rect 58216 13268 58218 13288
rect 58162 13232 58218 13268
rect 58162 11464 58218 11520
rect 58162 9716 58218 9752
rect 58162 9696 58164 9716
rect 58164 9696 58216 9716
rect 58216 9696 58218 9716
rect 58162 7928 58218 7984
rect 49116 7098 49172 7100
rect 49196 7098 49252 7100
rect 49276 7098 49332 7100
rect 49356 7098 49412 7100
rect 49116 7046 49162 7098
rect 49162 7046 49172 7098
rect 49196 7046 49226 7098
rect 49226 7046 49238 7098
rect 49238 7046 49252 7098
rect 49276 7046 49290 7098
rect 49290 7046 49302 7098
rect 49302 7046 49332 7098
rect 49356 7046 49366 7098
rect 49366 7046 49412 7098
rect 49116 7044 49172 7046
rect 49196 7044 49252 7046
rect 49276 7044 49332 7046
rect 49356 7044 49412 7046
rect 58162 6160 58218 6216
rect 49116 6010 49172 6012
rect 49196 6010 49252 6012
rect 49276 6010 49332 6012
rect 49356 6010 49412 6012
rect 49116 5958 49162 6010
rect 49162 5958 49172 6010
rect 49196 5958 49226 6010
rect 49226 5958 49238 6010
rect 49238 5958 49252 6010
rect 49276 5958 49290 6010
rect 49290 5958 49302 6010
rect 49302 5958 49332 6010
rect 49356 5958 49366 6010
rect 49366 5958 49412 6010
rect 49116 5956 49172 5958
rect 49196 5956 49252 5958
rect 49276 5956 49332 5958
rect 49356 5956 49412 5958
rect 48870 5616 48926 5672
rect 49116 4922 49172 4924
rect 49196 4922 49252 4924
rect 49276 4922 49332 4924
rect 49356 4922 49412 4924
rect 49116 4870 49162 4922
rect 49162 4870 49172 4922
rect 49196 4870 49226 4922
rect 49226 4870 49238 4922
rect 49238 4870 49252 4922
rect 49276 4870 49290 4922
rect 49290 4870 49302 4922
rect 49302 4870 49332 4922
rect 49356 4870 49366 4922
rect 49366 4870 49412 4922
rect 49116 4868 49172 4870
rect 49196 4868 49252 4870
rect 49276 4868 49332 4870
rect 49356 4868 49412 4870
rect 58162 4392 58218 4448
rect 49116 3834 49172 3836
rect 49196 3834 49252 3836
rect 49276 3834 49332 3836
rect 49356 3834 49412 3836
rect 49116 3782 49162 3834
rect 49162 3782 49172 3834
rect 49196 3782 49226 3834
rect 49226 3782 49238 3834
rect 49238 3782 49252 3834
rect 49276 3782 49290 3834
rect 49290 3782 49302 3834
rect 49302 3782 49332 3834
rect 49356 3782 49366 3834
rect 49366 3782 49412 3834
rect 49116 3780 49172 3782
rect 49196 3780 49252 3782
rect 49276 3780 49332 3782
rect 49356 3780 49412 3782
rect 49116 2746 49172 2748
rect 49196 2746 49252 2748
rect 49276 2746 49332 2748
rect 49356 2746 49412 2748
rect 49116 2694 49162 2746
rect 49162 2694 49172 2746
rect 49196 2694 49226 2746
rect 49226 2694 49238 2746
rect 49238 2694 49252 2746
rect 49276 2694 49290 2746
rect 49290 2694 49302 2746
rect 49302 2694 49332 2746
rect 49356 2694 49366 2746
rect 49366 2694 49412 2746
rect 49116 2692 49172 2694
rect 49196 2692 49252 2694
rect 49276 2692 49332 2694
rect 49356 2692 49412 2694
rect 56506 2644 56562 2680
rect 56506 2624 56508 2644
rect 56508 2624 56560 2644
rect 56560 2624 56562 2644
rect 57886 856 57942 912
rect 1490 720 1546 776
<< metal3 >>
rect 24342 29820 24348 29884
rect 24412 29882 24418 29884
rect 39113 29882 39179 29885
rect 24412 29880 39179 29882
rect 24412 29824 39118 29880
rect 39174 29824 39179 29880
rect 24412 29822 39179 29824
rect 24412 29820 24418 29822
rect 39113 29819 39179 29822
rect 19190 29684 19196 29748
rect 19260 29746 19266 29748
rect 34973 29746 35039 29749
rect 19260 29744 35039 29746
rect 19260 29688 34978 29744
rect 35034 29688 35039 29744
rect 19260 29686 35039 29688
rect 19260 29684 19266 29686
rect 34973 29683 35039 29686
rect 18321 29610 18387 29613
rect 34605 29610 34671 29613
rect 18321 29608 34671 29610
rect 18321 29552 18326 29608
rect 18382 29552 34610 29608
rect 34666 29552 34671 29608
rect 18321 29550 34671 29552
rect 18321 29547 18387 29550
rect 34605 29547 34671 29550
rect 19885 29338 19951 29341
rect 40166 29338 40172 29340
rect 19885 29336 40172 29338
rect 19885 29280 19890 29336
rect 19946 29280 40172 29336
rect 19885 29278 40172 29280
rect 19885 29275 19951 29278
rect 40166 29276 40172 29278
rect 40236 29276 40242 29340
rect 0 29202 800 29232
rect 1393 29202 1459 29205
rect 0 29200 1459 29202
rect 0 29144 1398 29200
rect 1454 29144 1459 29200
rect 0 29142 1459 29144
rect 0 29112 800 29142
rect 1393 29139 1459 29142
rect 16798 29140 16804 29204
rect 16868 29202 16874 29204
rect 41505 29202 41571 29205
rect 16868 29200 41571 29202
rect 16868 29144 41510 29200
rect 41566 29144 41571 29200
rect 16868 29142 41571 29144
rect 16868 29140 16874 29142
rect 41505 29139 41571 29142
rect 57237 29202 57303 29205
rect 59200 29202 60000 29232
rect 57237 29200 60000 29202
rect 57237 29144 57242 29200
rect 57298 29144 60000 29200
rect 57237 29142 60000 29144
rect 57237 29139 57303 29142
rect 59200 29112 60000 29142
rect 17534 29004 17540 29068
rect 17604 29066 17610 29068
rect 44357 29066 44423 29069
rect 17604 29064 44423 29066
rect 17604 29008 44362 29064
rect 44418 29008 44423 29064
rect 17604 29006 44423 29008
rect 17604 29004 17610 29006
rect 44357 29003 44423 29006
rect 21214 28868 21220 28932
rect 21284 28930 21290 28932
rect 44633 28930 44699 28933
rect 21284 28928 44699 28930
rect 21284 28872 44638 28928
rect 44694 28872 44699 28928
rect 21284 28870 44699 28872
rect 21284 28868 21290 28870
rect 44633 28867 44699 28870
rect 14825 28794 14891 28797
rect 42742 28794 42748 28796
rect 14825 28792 42748 28794
rect 14825 28736 14830 28792
rect 14886 28736 42748 28792
rect 14825 28734 42748 28736
rect 14825 28731 14891 28734
rect 42742 28732 42748 28734
rect 42812 28732 42818 28796
rect 14733 28658 14799 28661
rect 45134 28658 45140 28660
rect 14733 28656 45140 28658
rect 14733 28600 14738 28656
rect 14794 28600 45140 28656
rect 14733 28598 45140 28600
rect 14733 28595 14799 28598
rect 45134 28596 45140 28598
rect 45204 28596 45210 28660
rect 24209 28522 24275 28525
rect 40350 28522 40356 28524
rect 24209 28520 40356 28522
rect 24209 28464 24214 28520
rect 24270 28464 40356 28520
rect 24209 28462 40356 28464
rect 24209 28459 24275 28462
rect 40350 28460 40356 28462
rect 40420 28460 40426 28524
rect 14549 28386 14615 28389
rect 37590 28386 37596 28388
rect 14549 28384 37596 28386
rect 14549 28328 14554 28384
rect 14610 28328 37596 28384
rect 14549 28326 37596 28328
rect 14549 28323 14615 28326
rect 37590 28324 37596 28326
rect 37660 28324 37666 28388
rect 19006 28188 19012 28252
rect 19076 28250 19082 28252
rect 42006 28250 42012 28252
rect 19076 28190 42012 28250
rect 19076 28188 19082 28190
rect 42006 28188 42012 28190
rect 42076 28188 42082 28252
rect 21766 28052 21772 28116
rect 21836 28114 21842 28116
rect 37825 28114 37891 28117
rect 21836 28112 37891 28114
rect 21836 28056 37830 28112
rect 37886 28056 37891 28112
rect 21836 28054 37891 28056
rect 21836 28052 21842 28054
rect 37825 28051 37891 28054
rect 30465 27978 30531 27981
rect 38326 27978 38332 27980
rect 30465 27976 38332 27978
rect 30465 27920 30470 27976
rect 30526 27920 38332 27976
rect 30465 27918 38332 27920
rect 30465 27915 30531 27918
rect 38326 27916 38332 27918
rect 38396 27916 38402 27980
rect 31937 27842 32003 27845
rect 40902 27842 40908 27844
rect 31937 27840 40908 27842
rect 31937 27784 31942 27840
rect 31998 27784 40908 27840
rect 31937 27782 40908 27784
rect 31937 27779 32003 27782
rect 40902 27780 40908 27782
rect 40972 27780 40978 27844
rect 10576 27776 10896 27777
rect 10576 27712 10584 27776
rect 10648 27712 10664 27776
rect 10728 27712 10744 27776
rect 10808 27712 10824 27776
rect 10888 27712 10896 27776
rect 10576 27711 10896 27712
rect 29840 27776 30160 27777
rect 29840 27712 29848 27776
rect 29912 27712 29928 27776
rect 29992 27712 30008 27776
rect 30072 27712 30088 27776
rect 30152 27712 30160 27776
rect 29840 27711 30160 27712
rect 49104 27776 49424 27777
rect 49104 27712 49112 27776
rect 49176 27712 49192 27776
rect 49256 27712 49272 27776
rect 49336 27712 49352 27776
rect 49416 27712 49424 27776
rect 49104 27711 49424 27712
rect 34053 27706 34119 27709
rect 43345 27706 43411 27709
rect 34053 27704 43411 27706
rect 34053 27648 34058 27704
rect 34114 27648 43350 27704
rect 43406 27648 43411 27704
rect 34053 27646 43411 27648
rect 34053 27643 34119 27646
rect 43345 27643 43411 27646
rect 0 27570 800 27600
rect 1485 27570 1551 27573
rect 0 27568 1551 27570
rect 0 27512 1490 27568
rect 1546 27512 1551 27568
rect 0 27510 1551 27512
rect 0 27480 800 27510
rect 1485 27507 1551 27510
rect 19742 27508 19748 27572
rect 19812 27570 19818 27572
rect 39246 27570 39252 27572
rect 19812 27510 39252 27570
rect 19812 27508 19818 27510
rect 39246 27508 39252 27510
rect 39316 27508 39322 27572
rect 28809 27434 28875 27437
rect 32213 27434 32279 27437
rect 34145 27434 34211 27437
rect 52453 27434 52519 27437
rect 28809 27432 52519 27434
rect 28809 27376 28814 27432
rect 28870 27376 32218 27432
rect 32274 27376 34150 27432
rect 34206 27376 52458 27432
rect 52514 27376 52519 27432
rect 28809 27374 52519 27376
rect 28809 27371 28875 27374
rect 32213 27371 32279 27374
rect 34145 27371 34211 27374
rect 52453 27371 52519 27374
rect 58065 27434 58131 27437
rect 59200 27434 60000 27464
rect 58065 27432 60000 27434
rect 58065 27376 58070 27432
rect 58126 27376 60000 27432
rect 58065 27374 60000 27376
rect 58065 27371 58131 27374
rect 59200 27344 60000 27374
rect 20208 27232 20528 27233
rect 20208 27168 20216 27232
rect 20280 27168 20296 27232
rect 20360 27168 20376 27232
rect 20440 27168 20456 27232
rect 20520 27168 20528 27232
rect 20208 27167 20528 27168
rect 39472 27232 39792 27233
rect 39472 27168 39480 27232
rect 39544 27168 39560 27232
rect 39624 27168 39640 27232
rect 39704 27168 39720 27232
rect 39784 27168 39792 27232
rect 39472 27167 39792 27168
rect 29729 27026 29795 27029
rect 57881 27026 57947 27029
rect 29729 27024 57947 27026
rect 29729 26968 29734 27024
rect 29790 26968 57886 27024
rect 57942 26968 57947 27024
rect 29729 26966 57947 26968
rect 29729 26963 29795 26966
rect 57881 26963 57947 26966
rect 27521 26890 27587 26893
rect 27521 26888 30298 26890
rect 27521 26832 27526 26888
rect 27582 26832 30298 26888
rect 27521 26830 30298 26832
rect 27521 26827 27587 26830
rect 22001 26754 22067 26757
rect 29545 26754 29611 26757
rect 22001 26752 29611 26754
rect 22001 26696 22006 26752
rect 22062 26696 29550 26752
rect 29606 26696 29611 26752
rect 22001 26694 29611 26696
rect 22001 26691 22067 26694
rect 29545 26691 29611 26694
rect 10576 26688 10896 26689
rect 10576 26624 10584 26688
rect 10648 26624 10664 26688
rect 10728 26624 10744 26688
rect 10808 26624 10824 26688
rect 10888 26624 10896 26688
rect 10576 26623 10896 26624
rect 29840 26688 30160 26689
rect 29840 26624 29848 26688
rect 29912 26624 29928 26688
rect 29992 26624 30008 26688
rect 30072 26624 30088 26688
rect 30152 26624 30160 26688
rect 29840 26623 30160 26624
rect 28441 26618 28507 26621
rect 22050 26616 28507 26618
rect 22050 26560 28446 26616
rect 28502 26560 28507 26616
rect 22050 26558 28507 26560
rect 20069 26482 20135 26485
rect 22050 26482 22110 26558
rect 28441 26555 28507 26558
rect 20069 26480 22110 26482
rect 20069 26424 20074 26480
rect 20130 26424 22110 26480
rect 20069 26422 22110 26424
rect 26417 26482 26483 26485
rect 29729 26482 29795 26485
rect 26417 26480 29795 26482
rect 26417 26424 26422 26480
rect 26478 26424 29734 26480
rect 29790 26424 29795 26480
rect 26417 26422 29795 26424
rect 30238 26482 30298 26830
rect 30833 26754 30899 26757
rect 38694 26754 38700 26756
rect 30833 26752 38700 26754
rect 30833 26696 30838 26752
rect 30894 26696 38700 26752
rect 30833 26694 38700 26696
rect 30833 26691 30899 26694
rect 38694 26692 38700 26694
rect 38764 26692 38770 26756
rect 49104 26688 49424 26689
rect 49104 26624 49112 26688
rect 49176 26624 49192 26688
rect 49256 26624 49272 26688
rect 49336 26624 49352 26688
rect 49416 26624 49424 26688
rect 49104 26623 49424 26624
rect 31201 26618 31267 26621
rect 37406 26618 37412 26620
rect 31201 26616 37412 26618
rect 31201 26560 31206 26616
rect 31262 26560 37412 26616
rect 31201 26558 37412 26560
rect 31201 26555 31267 26558
rect 37406 26556 37412 26558
rect 37476 26556 37482 26620
rect 35801 26482 35867 26485
rect 43437 26482 43503 26485
rect 30238 26480 35867 26482
rect 30238 26424 35806 26480
rect 35862 26424 35867 26480
rect 30238 26422 35867 26424
rect 20069 26419 20135 26422
rect 26417 26419 26483 26422
rect 29729 26419 29795 26422
rect 35801 26419 35867 26422
rect 41370 26480 43503 26482
rect 41370 26424 43442 26480
rect 43498 26424 43503 26480
rect 41370 26422 43503 26424
rect 21950 26284 21956 26348
rect 22020 26346 22026 26348
rect 27613 26346 27679 26349
rect 22020 26344 27679 26346
rect 22020 26288 27618 26344
rect 27674 26288 27679 26344
rect 22020 26286 27679 26288
rect 22020 26284 22026 26286
rect 27613 26283 27679 26286
rect 30782 26284 30788 26348
rect 30852 26346 30858 26348
rect 31477 26346 31543 26349
rect 30852 26344 31543 26346
rect 30852 26288 31482 26344
rect 31538 26288 31543 26344
rect 30852 26286 31543 26288
rect 30852 26284 30858 26286
rect 31477 26283 31543 26286
rect 32489 26346 32555 26349
rect 32622 26346 32628 26348
rect 32489 26344 32628 26346
rect 32489 26288 32494 26344
rect 32550 26288 32628 26344
rect 32489 26286 32628 26288
rect 32489 26283 32555 26286
rect 32622 26284 32628 26286
rect 32692 26284 32698 26348
rect 34145 26346 34211 26349
rect 41370 26346 41430 26422
rect 43437 26419 43503 26422
rect 34145 26344 41430 26346
rect 34145 26288 34150 26344
rect 34206 26288 41430 26344
rect 34145 26286 41430 26288
rect 34145 26283 34211 26286
rect 28993 26210 29059 26213
rect 31017 26210 31083 26213
rect 31569 26210 31635 26213
rect 28993 26208 31635 26210
rect 28993 26152 28998 26208
rect 29054 26152 31022 26208
rect 31078 26152 31574 26208
rect 31630 26152 31635 26208
rect 28993 26150 31635 26152
rect 28993 26147 29059 26150
rect 31017 26147 31083 26150
rect 31569 26147 31635 26150
rect 20208 26144 20528 26145
rect 0 26074 800 26104
rect 20208 26080 20216 26144
rect 20280 26080 20296 26144
rect 20360 26080 20376 26144
rect 20440 26080 20456 26144
rect 20520 26080 20528 26144
rect 20208 26079 20528 26080
rect 39472 26144 39792 26145
rect 39472 26080 39480 26144
rect 39544 26080 39560 26144
rect 39624 26080 39640 26144
rect 39704 26080 39720 26144
rect 39784 26080 39792 26144
rect 39472 26079 39792 26080
rect 1485 26074 1551 26077
rect 0 26072 1551 26074
rect 0 26016 1490 26072
rect 1546 26016 1551 26072
rect 0 26014 1551 26016
rect 0 25984 800 26014
rect 1485 26011 1551 26014
rect 24577 26074 24643 26077
rect 30465 26074 30531 26077
rect 33961 26074 34027 26077
rect 24577 26072 30531 26074
rect 24577 26016 24582 26072
rect 24638 26016 30470 26072
rect 30526 26016 30531 26072
rect 24577 26014 30531 26016
rect 24577 26011 24643 26014
rect 30465 26011 30531 26014
rect 31710 26072 34027 26074
rect 31710 26016 33966 26072
rect 34022 26016 34027 26072
rect 31710 26014 34027 26016
rect 17902 25876 17908 25940
rect 17972 25938 17978 25940
rect 29269 25938 29335 25941
rect 17972 25936 29335 25938
rect 17972 25880 29274 25936
rect 29330 25880 29335 25936
rect 17972 25878 29335 25880
rect 17972 25876 17978 25878
rect 29269 25875 29335 25878
rect 29729 25938 29795 25941
rect 31710 25938 31770 26014
rect 33961 26011 34027 26014
rect 29729 25936 31770 25938
rect 29729 25880 29734 25936
rect 29790 25880 31770 25936
rect 29729 25878 31770 25880
rect 35065 25938 35131 25941
rect 43161 25938 43227 25941
rect 35065 25936 43227 25938
rect 35065 25880 35070 25936
rect 35126 25880 43166 25936
rect 43222 25880 43227 25936
rect 35065 25878 43227 25880
rect 29729 25875 29795 25878
rect 35065 25875 35131 25878
rect 43161 25875 43227 25878
rect 21817 25802 21883 25805
rect 28993 25802 29059 25805
rect 21817 25800 29059 25802
rect 21817 25744 21822 25800
rect 21878 25744 28998 25800
rect 29054 25744 29059 25800
rect 21817 25742 29059 25744
rect 21817 25739 21883 25742
rect 28993 25739 29059 25742
rect 29177 25802 29243 25805
rect 33685 25802 33751 25805
rect 29177 25800 33751 25802
rect 29177 25744 29182 25800
rect 29238 25744 33690 25800
rect 33746 25744 33751 25800
rect 29177 25742 33751 25744
rect 29177 25739 29243 25742
rect 33685 25739 33751 25742
rect 35525 25802 35591 25805
rect 44449 25802 44515 25805
rect 35525 25800 44515 25802
rect 35525 25744 35530 25800
rect 35586 25744 44454 25800
rect 44510 25744 44515 25800
rect 35525 25742 44515 25744
rect 35525 25739 35591 25742
rect 44449 25739 44515 25742
rect 19006 25604 19012 25668
rect 19076 25666 19082 25668
rect 28901 25666 28967 25669
rect 19076 25664 28967 25666
rect 19076 25608 28906 25664
rect 28962 25608 28967 25664
rect 19076 25606 28967 25608
rect 19076 25604 19082 25606
rect 28901 25603 28967 25606
rect 30373 25666 30439 25669
rect 37641 25666 37707 25669
rect 30373 25664 37707 25666
rect 30373 25608 30378 25664
rect 30434 25608 37646 25664
rect 37702 25608 37707 25664
rect 30373 25606 37707 25608
rect 30373 25603 30439 25606
rect 37641 25603 37707 25606
rect 58157 25666 58223 25669
rect 59200 25666 60000 25696
rect 58157 25664 60000 25666
rect 58157 25608 58162 25664
rect 58218 25608 60000 25664
rect 58157 25606 60000 25608
rect 58157 25603 58223 25606
rect 10576 25600 10896 25601
rect 10576 25536 10584 25600
rect 10648 25536 10664 25600
rect 10728 25536 10744 25600
rect 10808 25536 10824 25600
rect 10888 25536 10896 25600
rect 10576 25535 10896 25536
rect 29840 25600 30160 25601
rect 29840 25536 29848 25600
rect 29912 25536 29928 25600
rect 29992 25536 30008 25600
rect 30072 25536 30088 25600
rect 30152 25536 30160 25600
rect 29840 25535 30160 25536
rect 49104 25600 49424 25601
rect 49104 25536 49112 25600
rect 49176 25536 49192 25600
rect 49256 25536 49272 25600
rect 49336 25536 49352 25600
rect 49416 25536 49424 25600
rect 59200 25576 60000 25606
rect 49104 25535 49424 25536
rect 15193 25530 15259 25533
rect 24393 25530 24459 25533
rect 27470 25530 27476 25532
rect 15193 25528 27476 25530
rect 15193 25472 15198 25528
rect 15254 25472 24398 25528
rect 24454 25472 27476 25528
rect 15193 25470 27476 25472
rect 15193 25467 15259 25470
rect 24393 25467 24459 25470
rect 27470 25468 27476 25470
rect 27540 25468 27546 25532
rect 17125 25394 17191 25397
rect 28206 25394 28212 25396
rect 17125 25392 28212 25394
rect 17125 25336 17130 25392
rect 17186 25336 28212 25392
rect 17125 25334 28212 25336
rect 17125 25331 17191 25334
rect 28206 25332 28212 25334
rect 28276 25332 28282 25396
rect 28901 25394 28967 25397
rect 30373 25394 30439 25397
rect 28901 25392 30439 25394
rect 28901 25336 28906 25392
rect 28962 25336 30378 25392
rect 30434 25336 30439 25392
rect 28901 25334 30439 25336
rect 28901 25331 28967 25334
rect 30373 25331 30439 25334
rect 25221 25260 25287 25261
rect 25221 25256 25268 25260
rect 25332 25258 25338 25260
rect 27245 25258 27311 25261
rect 28390 25258 28396 25260
rect 25221 25200 25226 25256
rect 25221 25196 25268 25200
rect 25332 25198 25378 25258
rect 27245 25256 28396 25258
rect 27245 25200 27250 25256
rect 27306 25200 28396 25256
rect 27245 25198 28396 25200
rect 25332 25196 25338 25198
rect 25221 25195 25287 25196
rect 27245 25195 27311 25198
rect 28390 25196 28396 25198
rect 28460 25196 28466 25260
rect 29678 25196 29684 25260
rect 29748 25258 29754 25260
rect 30557 25258 30623 25261
rect 29748 25256 30623 25258
rect 29748 25200 30562 25256
rect 30618 25200 30623 25256
rect 29748 25198 30623 25200
rect 29748 25196 29754 25198
rect 30557 25195 30623 25198
rect 31477 25258 31543 25261
rect 40861 25258 40927 25261
rect 31477 25256 40927 25258
rect 31477 25200 31482 25256
rect 31538 25200 40866 25256
rect 40922 25200 40927 25256
rect 31477 25198 40927 25200
rect 31477 25195 31543 25198
rect 40861 25195 40927 25198
rect 22093 25122 22159 25125
rect 28441 25122 28507 25125
rect 22093 25120 28507 25122
rect 22093 25064 22098 25120
rect 22154 25064 28446 25120
rect 28502 25064 28507 25120
rect 22093 25062 28507 25064
rect 22093 25059 22159 25062
rect 28441 25059 28507 25062
rect 29310 25060 29316 25124
rect 29380 25122 29386 25124
rect 31937 25122 32003 25125
rect 29380 25120 32003 25122
rect 29380 25064 31942 25120
rect 31998 25064 32003 25120
rect 29380 25062 32003 25064
rect 29380 25060 29386 25062
rect 31937 25059 32003 25062
rect 32305 25122 32371 25125
rect 35709 25122 35775 25125
rect 32305 25120 35775 25122
rect 32305 25064 32310 25120
rect 32366 25064 35714 25120
rect 35770 25064 35775 25120
rect 32305 25062 35775 25064
rect 32305 25059 32371 25062
rect 35709 25059 35775 25062
rect 20208 25056 20528 25057
rect 20208 24992 20216 25056
rect 20280 24992 20296 25056
rect 20360 24992 20376 25056
rect 20440 24992 20456 25056
rect 20520 24992 20528 25056
rect 20208 24991 20528 24992
rect 39472 25056 39792 25057
rect 39472 24992 39480 25056
rect 39544 24992 39560 25056
rect 39624 24992 39640 25056
rect 39704 24992 39720 25056
rect 39784 24992 39792 25056
rect 39472 24991 39792 24992
rect 24301 24986 24367 24989
rect 29729 24986 29795 24989
rect 34329 24988 34395 24989
rect 24301 24984 29795 24986
rect 24301 24928 24306 24984
rect 24362 24928 29734 24984
rect 29790 24928 29795 24984
rect 24301 24926 29795 24928
rect 24301 24923 24367 24926
rect 29729 24923 29795 24926
rect 34278 24924 34284 24988
rect 34348 24986 34395 24988
rect 35617 24986 35683 24989
rect 38101 24986 38167 24989
rect 34348 24984 34440 24986
rect 34390 24928 34440 24984
rect 34348 24926 34440 24928
rect 35617 24984 38167 24986
rect 35617 24928 35622 24984
rect 35678 24928 38106 24984
rect 38162 24928 38167 24984
rect 35617 24926 38167 24928
rect 34348 24924 34395 24926
rect 34329 24923 34395 24924
rect 35617 24923 35683 24926
rect 38101 24923 38167 24926
rect 16573 24850 16639 24853
rect 36169 24850 36235 24853
rect 16573 24848 36235 24850
rect 16573 24792 16578 24848
rect 16634 24792 36174 24848
rect 36230 24792 36235 24848
rect 16573 24790 36235 24792
rect 16573 24787 16639 24790
rect 36169 24787 36235 24790
rect 26877 24714 26943 24717
rect 32305 24714 32371 24717
rect 35065 24714 35131 24717
rect 26877 24712 32184 24714
rect 26877 24656 26882 24712
rect 26938 24656 32184 24712
rect 26877 24654 32184 24656
rect 26877 24651 26943 24654
rect 27429 24578 27495 24581
rect 28758 24578 28764 24580
rect 27429 24576 28764 24578
rect 27429 24520 27434 24576
rect 27490 24520 28764 24576
rect 27429 24518 28764 24520
rect 27429 24515 27495 24518
rect 28758 24516 28764 24518
rect 28828 24516 28834 24580
rect 10576 24512 10896 24513
rect 0 24442 800 24472
rect 10576 24448 10584 24512
rect 10648 24448 10664 24512
rect 10728 24448 10744 24512
rect 10808 24448 10824 24512
rect 10888 24448 10896 24512
rect 10576 24447 10896 24448
rect 29840 24512 30160 24513
rect 29840 24448 29848 24512
rect 29912 24448 29928 24512
rect 29992 24448 30008 24512
rect 30072 24448 30088 24512
rect 30152 24448 30160 24512
rect 29840 24447 30160 24448
rect 1485 24442 1551 24445
rect 0 24440 1551 24442
rect 0 24384 1490 24440
rect 1546 24384 1551 24440
rect 0 24382 1551 24384
rect 0 24352 800 24382
rect 1485 24379 1551 24382
rect 22737 24442 22803 24445
rect 29310 24442 29316 24444
rect 22737 24440 29316 24442
rect 22737 24384 22742 24440
rect 22798 24384 29316 24440
rect 22737 24382 29316 24384
rect 22737 24379 22803 24382
rect 29310 24380 29316 24382
rect 29380 24380 29386 24444
rect 32124 24442 32184 24654
rect 32305 24712 35131 24714
rect 32305 24656 32310 24712
rect 32366 24656 35070 24712
rect 35126 24656 35131 24712
rect 32305 24654 35131 24656
rect 32305 24651 32371 24654
rect 35065 24651 35131 24654
rect 35985 24714 36051 24717
rect 37958 24714 37964 24716
rect 35985 24712 37964 24714
rect 35985 24656 35990 24712
rect 36046 24656 37964 24712
rect 35985 24654 37964 24656
rect 35985 24651 36051 24654
rect 37958 24652 37964 24654
rect 38028 24652 38034 24716
rect 33358 24516 33364 24580
rect 33428 24578 33434 24580
rect 33501 24578 33567 24581
rect 33428 24576 33567 24578
rect 33428 24520 33506 24576
rect 33562 24520 33567 24576
rect 33428 24518 33567 24520
rect 33428 24516 33434 24518
rect 33501 24515 33567 24518
rect 36670 24516 36676 24580
rect 36740 24578 36746 24580
rect 39481 24578 39547 24581
rect 46289 24578 46355 24581
rect 36740 24576 46355 24578
rect 36740 24520 39486 24576
rect 39542 24520 46294 24576
rect 46350 24520 46355 24576
rect 36740 24518 46355 24520
rect 36740 24516 36746 24518
rect 39481 24515 39547 24518
rect 46289 24515 46355 24518
rect 49104 24512 49424 24513
rect 49104 24448 49112 24512
rect 49176 24448 49192 24512
rect 49256 24448 49272 24512
rect 49336 24448 49352 24512
rect 49416 24448 49424 24512
rect 49104 24447 49424 24448
rect 36905 24442 36971 24445
rect 32124 24440 36971 24442
rect 32124 24384 36910 24440
rect 36966 24384 36971 24440
rect 32124 24382 36971 24384
rect 36905 24379 36971 24382
rect 27337 24306 27403 24309
rect 38561 24306 38627 24309
rect 27337 24304 38627 24306
rect 27337 24248 27342 24304
rect 27398 24248 38566 24304
rect 38622 24248 38627 24304
rect 27337 24246 38627 24248
rect 27337 24243 27403 24246
rect 38561 24243 38627 24246
rect 25405 24170 25471 24173
rect 26049 24170 26115 24173
rect 27981 24170 28047 24173
rect 25405 24168 28047 24170
rect 25405 24112 25410 24168
rect 25466 24112 26054 24168
rect 26110 24112 27986 24168
rect 28042 24112 28047 24168
rect 25405 24110 28047 24112
rect 25405 24107 25471 24110
rect 26049 24107 26115 24110
rect 27981 24107 28047 24110
rect 28574 24108 28580 24172
rect 28644 24170 28650 24172
rect 28717 24170 28783 24173
rect 28644 24168 28783 24170
rect 28644 24112 28722 24168
rect 28778 24112 28783 24168
rect 28644 24110 28783 24112
rect 28644 24108 28650 24110
rect 28717 24107 28783 24110
rect 30373 24170 30439 24173
rect 31293 24170 31359 24173
rect 30373 24168 31359 24170
rect 30373 24112 30378 24168
rect 30434 24112 31298 24168
rect 31354 24112 31359 24168
rect 30373 24110 31359 24112
rect 30373 24107 30439 24110
rect 31293 24107 31359 24110
rect 32121 24170 32187 24173
rect 33869 24170 33935 24173
rect 32121 24168 33935 24170
rect 32121 24112 32126 24168
rect 32182 24112 33874 24168
rect 33930 24112 33935 24168
rect 32121 24110 33935 24112
rect 32121 24107 32187 24110
rect 33869 24107 33935 24110
rect 34053 24170 34119 24173
rect 41086 24170 41092 24172
rect 34053 24168 41092 24170
rect 34053 24112 34058 24168
rect 34114 24112 41092 24168
rect 34053 24110 41092 24112
rect 34053 24107 34119 24110
rect 41086 24108 41092 24110
rect 41156 24108 41162 24172
rect 25405 24034 25471 24037
rect 25589 24034 25655 24037
rect 25405 24032 25655 24034
rect 25405 23976 25410 24032
rect 25466 23976 25594 24032
rect 25650 23976 25655 24032
rect 25405 23974 25655 23976
rect 25405 23971 25471 23974
rect 25589 23971 25655 23974
rect 25814 23972 25820 24036
rect 25884 24034 25890 24036
rect 26877 24034 26943 24037
rect 27337 24036 27403 24037
rect 27286 24034 27292 24036
rect 25884 24032 26943 24034
rect 25884 23976 26882 24032
rect 26938 23976 26943 24032
rect 25884 23974 26943 23976
rect 27246 23974 27292 24034
rect 27356 24032 27403 24036
rect 27398 23976 27403 24032
rect 25884 23972 25890 23974
rect 26877 23971 26943 23974
rect 27286 23972 27292 23974
rect 27356 23972 27403 23976
rect 27337 23971 27403 23972
rect 28257 24034 28323 24037
rect 34973 24034 35039 24037
rect 28257 24032 35039 24034
rect 28257 23976 28262 24032
rect 28318 23976 34978 24032
rect 35034 23976 35039 24032
rect 28257 23974 35039 23976
rect 28257 23971 28323 23974
rect 34973 23971 35039 23974
rect 35525 24034 35591 24037
rect 36997 24034 37063 24037
rect 35525 24032 37063 24034
rect 35525 23976 35530 24032
rect 35586 23976 37002 24032
rect 37058 23976 37063 24032
rect 35525 23974 37063 23976
rect 35525 23971 35591 23974
rect 36997 23971 37063 23974
rect 20208 23968 20528 23969
rect 20208 23904 20216 23968
rect 20280 23904 20296 23968
rect 20360 23904 20376 23968
rect 20440 23904 20456 23968
rect 20520 23904 20528 23968
rect 20208 23903 20528 23904
rect 39472 23968 39792 23969
rect 39472 23904 39480 23968
rect 39544 23904 39560 23968
rect 39624 23904 39640 23968
rect 39704 23904 39720 23968
rect 39784 23904 39792 23968
rect 39472 23903 39792 23904
rect 21357 23898 21423 23901
rect 27337 23898 27403 23901
rect 21357 23896 27403 23898
rect 21357 23840 21362 23896
rect 21418 23840 27342 23896
rect 27398 23840 27403 23896
rect 21357 23838 27403 23840
rect 21357 23835 21423 23838
rect 27337 23835 27403 23838
rect 28022 23836 28028 23900
rect 28092 23898 28098 23900
rect 30833 23898 30899 23901
rect 32949 23900 33015 23901
rect 32949 23898 32996 23900
rect 28092 23896 30899 23898
rect 28092 23840 30838 23896
rect 30894 23840 30899 23896
rect 28092 23838 30899 23840
rect 32904 23896 32996 23898
rect 32904 23840 32954 23896
rect 32904 23838 32996 23840
rect 28092 23836 28098 23838
rect 30833 23835 30899 23838
rect 32949 23836 32996 23838
rect 33060 23836 33066 23900
rect 34421 23898 34487 23901
rect 34830 23898 34836 23900
rect 34421 23896 34836 23898
rect 34421 23840 34426 23896
rect 34482 23840 34836 23896
rect 34421 23838 34836 23840
rect 32949 23835 33015 23836
rect 34421 23835 34487 23838
rect 34830 23836 34836 23838
rect 34900 23836 34906 23900
rect 35065 23898 35131 23901
rect 37273 23898 37339 23901
rect 35065 23896 37339 23898
rect 35065 23840 35070 23896
rect 35126 23840 37278 23896
rect 37334 23840 37339 23896
rect 35065 23838 37339 23840
rect 35065 23835 35131 23838
rect 37273 23835 37339 23838
rect 58157 23898 58223 23901
rect 59200 23898 60000 23928
rect 58157 23896 60000 23898
rect 58157 23840 58162 23896
rect 58218 23840 60000 23896
rect 58157 23838 60000 23840
rect 58157 23835 58223 23838
rect 59200 23808 60000 23838
rect 24894 23762 24900 23764
rect 16622 23702 24900 23762
rect 16481 23490 16547 23493
rect 16622 23490 16682 23702
rect 24894 23700 24900 23702
rect 24964 23700 24970 23764
rect 27102 23700 27108 23764
rect 27172 23762 27178 23764
rect 29637 23762 29703 23765
rect 27172 23760 29703 23762
rect 27172 23704 29642 23760
rect 29698 23704 29703 23760
rect 27172 23702 29703 23704
rect 27172 23700 27178 23702
rect 29637 23699 29703 23702
rect 30097 23762 30163 23765
rect 32029 23762 32095 23765
rect 36169 23762 36235 23765
rect 38837 23762 38903 23765
rect 30097 23760 32095 23762
rect 30097 23704 30102 23760
rect 30158 23704 32034 23760
rect 32090 23704 32095 23760
rect 30097 23702 32095 23704
rect 30097 23699 30163 23702
rect 32029 23699 32095 23702
rect 32262 23760 36235 23762
rect 32262 23704 36174 23760
rect 36230 23704 36235 23760
rect 32262 23702 36235 23704
rect 21081 23626 21147 23629
rect 25589 23626 25655 23629
rect 21081 23624 25655 23626
rect 21081 23568 21086 23624
rect 21142 23568 25594 23624
rect 25650 23568 25655 23624
rect 21081 23566 25655 23568
rect 21081 23563 21147 23566
rect 25589 23563 25655 23566
rect 25773 23626 25839 23629
rect 27153 23626 27219 23629
rect 25773 23624 27219 23626
rect 25773 23568 25778 23624
rect 25834 23568 27158 23624
rect 27214 23568 27219 23624
rect 25773 23566 27219 23568
rect 25773 23563 25839 23566
rect 27153 23563 27219 23566
rect 30005 23626 30071 23629
rect 30414 23626 30420 23628
rect 30005 23624 30420 23626
rect 30005 23568 30010 23624
rect 30066 23568 30420 23624
rect 30005 23566 30420 23568
rect 30005 23563 30071 23566
rect 30414 23564 30420 23566
rect 30484 23564 30490 23628
rect 30966 23564 30972 23628
rect 31036 23626 31042 23628
rect 32262 23626 32322 23702
rect 36169 23699 36235 23702
rect 36310 23760 38903 23762
rect 36310 23704 38842 23760
rect 38898 23704 38903 23760
rect 36310 23702 38903 23704
rect 33317 23626 33383 23629
rect 35709 23628 35775 23629
rect 35709 23626 35756 23628
rect 31036 23566 32322 23626
rect 32446 23624 33383 23626
rect 32446 23568 33322 23624
rect 33378 23568 33383 23624
rect 32446 23566 33383 23568
rect 35664 23624 35756 23626
rect 35664 23568 35714 23624
rect 35664 23566 35756 23568
rect 31036 23564 31042 23566
rect 16481 23488 16682 23490
rect 16481 23432 16486 23488
rect 16542 23432 16682 23488
rect 16481 23430 16682 23432
rect 21265 23490 21331 23493
rect 22318 23490 22324 23492
rect 21265 23488 22324 23490
rect 21265 23432 21270 23488
rect 21326 23432 22324 23488
rect 21265 23430 22324 23432
rect 16481 23427 16547 23430
rect 21265 23427 21331 23430
rect 22318 23428 22324 23430
rect 22388 23428 22394 23492
rect 24710 23428 24716 23492
rect 24780 23490 24786 23492
rect 26693 23490 26759 23493
rect 24780 23488 26759 23490
rect 24780 23432 26698 23488
rect 26754 23432 26759 23488
rect 24780 23430 26759 23432
rect 24780 23428 24786 23430
rect 26693 23427 26759 23430
rect 27981 23490 28047 23493
rect 28901 23490 28967 23493
rect 27981 23488 28967 23490
rect 27981 23432 27986 23488
rect 28042 23432 28906 23488
rect 28962 23432 28967 23488
rect 27981 23430 28967 23432
rect 27981 23427 28047 23430
rect 28901 23427 28967 23430
rect 31201 23490 31267 23493
rect 32446 23490 32506 23566
rect 33317 23563 33383 23566
rect 35709 23564 35756 23566
rect 35820 23564 35826 23628
rect 36310 23626 36370 23702
rect 38837 23699 38903 23702
rect 35896 23566 36370 23626
rect 36813 23626 36879 23629
rect 40769 23626 40835 23629
rect 36813 23624 40835 23626
rect 36813 23568 36818 23624
rect 36874 23568 40774 23624
rect 40830 23568 40835 23624
rect 36813 23566 40835 23568
rect 35709 23563 35775 23564
rect 35896 23493 35956 23566
rect 36813 23563 36879 23566
rect 40769 23563 40835 23566
rect 31201 23488 32506 23490
rect 31201 23432 31206 23488
rect 31262 23432 32506 23488
rect 31201 23430 32506 23432
rect 33133 23492 33199 23493
rect 33133 23488 33180 23492
rect 33244 23490 33250 23492
rect 33133 23432 33138 23488
rect 31201 23427 31267 23430
rect 33133 23428 33180 23432
rect 33244 23430 33290 23490
rect 35893 23488 35959 23493
rect 35893 23432 35898 23488
rect 35954 23432 35959 23488
rect 33244 23428 33250 23430
rect 33133 23427 33199 23428
rect 35893 23427 35959 23432
rect 36537 23490 36603 23493
rect 37222 23490 37228 23492
rect 36537 23488 37228 23490
rect 36537 23432 36542 23488
rect 36598 23432 37228 23488
rect 36537 23430 37228 23432
rect 36537 23427 36603 23430
rect 37222 23428 37228 23430
rect 37292 23428 37298 23492
rect 10576 23424 10896 23425
rect 10576 23360 10584 23424
rect 10648 23360 10664 23424
rect 10728 23360 10744 23424
rect 10808 23360 10824 23424
rect 10888 23360 10896 23424
rect 10576 23359 10896 23360
rect 29840 23424 30160 23425
rect 29840 23360 29848 23424
rect 29912 23360 29928 23424
rect 29992 23360 30008 23424
rect 30072 23360 30088 23424
rect 30152 23360 30160 23424
rect 29840 23359 30160 23360
rect 49104 23424 49424 23425
rect 49104 23360 49112 23424
rect 49176 23360 49192 23424
rect 49256 23360 49272 23424
rect 49336 23360 49352 23424
rect 49416 23360 49424 23424
rect 49104 23359 49424 23360
rect 16941 23354 17007 23357
rect 27061 23354 27127 23357
rect 16941 23352 27127 23354
rect 16941 23296 16946 23352
rect 17002 23296 27066 23352
rect 27122 23296 27127 23352
rect 16941 23294 27127 23296
rect 16941 23291 17007 23294
rect 27061 23291 27127 23294
rect 28165 23354 28231 23357
rect 28809 23354 28875 23357
rect 28165 23352 28875 23354
rect 28165 23296 28170 23352
rect 28226 23296 28814 23352
rect 28870 23296 28875 23352
rect 28165 23294 28875 23296
rect 28165 23291 28231 23294
rect 28809 23291 28875 23294
rect 33869 23354 33935 23357
rect 36905 23354 36971 23357
rect 33869 23352 36971 23354
rect 33869 23296 33874 23352
rect 33930 23296 36910 23352
rect 36966 23296 36971 23352
rect 33869 23294 36971 23296
rect 33869 23291 33935 23294
rect 36905 23291 36971 23294
rect 37089 23354 37155 23357
rect 40493 23354 40559 23357
rect 37089 23352 40559 23354
rect 37089 23296 37094 23352
rect 37150 23296 40498 23352
rect 40554 23296 40559 23352
rect 37089 23294 40559 23296
rect 37089 23291 37155 23294
rect 40493 23291 40559 23294
rect 19558 23156 19564 23220
rect 19628 23218 19634 23220
rect 20529 23218 20595 23221
rect 19628 23216 20595 23218
rect 19628 23160 20534 23216
rect 20590 23160 20595 23216
rect 19628 23158 20595 23160
rect 19628 23156 19634 23158
rect 20529 23155 20595 23158
rect 26325 23218 26391 23221
rect 38745 23218 38811 23221
rect 26325 23216 38811 23218
rect 26325 23160 26330 23216
rect 26386 23160 38750 23216
rect 38806 23160 38811 23216
rect 26325 23158 38811 23160
rect 26325 23155 26391 23158
rect 38745 23155 38811 23158
rect 39389 23218 39455 23221
rect 45185 23218 45251 23221
rect 39389 23216 45251 23218
rect 39389 23160 39394 23216
rect 39450 23160 45190 23216
rect 45246 23160 45251 23216
rect 39389 23158 45251 23160
rect 39389 23155 39455 23158
rect 45185 23155 45251 23158
rect 21398 23020 21404 23084
rect 21468 23082 21474 23084
rect 24577 23082 24643 23085
rect 26325 23082 26391 23085
rect 21468 23080 26391 23082
rect 21468 23024 24582 23080
rect 24638 23024 26330 23080
rect 26386 23024 26391 23080
rect 21468 23022 26391 23024
rect 21468 23020 21474 23022
rect 24577 23019 24643 23022
rect 26325 23019 26391 23022
rect 26877 23082 26943 23085
rect 26877 23080 27354 23082
rect 26877 23024 26882 23080
rect 26938 23024 27354 23080
rect 26877 23022 27354 23024
rect 26877 23019 26943 23022
rect 26233 22946 26299 22949
rect 26877 22946 26943 22949
rect 26233 22944 26943 22946
rect 26233 22888 26238 22944
rect 26294 22888 26882 22944
rect 26938 22888 26943 22944
rect 26233 22886 26943 22888
rect 27294 22946 27354 23022
rect 27838 23020 27844 23084
rect 27908 23082 27914 23084
rect 27981 23082 28047 23085
rect 27908 23080 28047 23082
rect 27908 23024 27986 23080
rect 28042 23024 28047 23080
rect 27908 23022 28047 23024
rect 27908 23020 27914 23022
rect 27981 23019 28047 23022
rect 28349 23082 28415 23085
rect 30598 23082 30604 23084
rect 28349 23080 30604 23082
rect 28349 23024 28354 23080
rect 28410 23024 30604 23080
rect 28349 23022 30604 23024
rect 28349 23019 28415 23022
rect 30598 23020 30604 23022
rect 30668 23020 30674 23084
rect 31753 23082 31819 23085
rect 35065 23082 35131 23085
rect 41965 23082 42031 23085
rect 31753 23080 34898 23082
rect 31753 23024 31758 23080
rect 31814 23024 34898 23080
rect 31753 23022 34898 23024
rect 31753 23019 31819 23022
rect 34237 22946 34303 22949
rect 27294 22944 34303 22946
rect 27294 22888 34242 22944
rect 34298 22888 34303 22944
rect 27294 22886 34303 22888
rect 34838 22946 34898 23022
rect 35065 23080 42031 23082
rect 35065 23024 35070 23080
rect 35126 23024 41970 23080
rect 42026 23024 42031 23080
rect 35065 23022 42031 23024
rect 35065 23019 35131 23022
rect 41965 23019 42031 23022
rect 38469 22946 38535 22949
rect 34838 22944 38535 22946
rect 34838 22888 38474 22944
rect 38530 22888 38535 22944
rect 34838 22886 38535 22888
rect 26233 22883 26299 22886
rect 26877 22883 26943 22886
rect 34237 22883 34303 22886
rect 38469 22883 38535 22886
rect 38653 22946 38719 22949
rect 38878 22946 38884 22948
rect 38653 22944 38884 22946
rect 38653 22888 38658 22944
rect 38714 22888 38884 22944
rect 38653 22886 38884 22888
rect 38653 22883 38719 22886
rect 38878 22884 38884 22886
rect 38948 22884 38954 22948
rect 20208 22880 20528 22881
rect 0 22810 800 22840
rect 20208 22816 20216 22880
rect 20280 22816 20296 22880
rect 20360 22816 20376 22880
rect 20440 22816 20456 22880
rect 20520 22816 20528 22880
rect 20208 22815 20528 22816
rect 1485 22810 1551 22813
rect 0 22808 1551 22810
rect 0 22752 1490 22808
rect 1546 22752 1551 22808
rect 0 22750 1551 22752
rect 0 22720 800 22750
rect 1485 22747 1551 22750
rect 22737 22810 22803 22813
rect 26236 22810 26296 22883
rect 39472 22880 39792 22881
rect 39472 22816 39480 22880
rect 39544 22816 39560 22880
rect 39624 22816 39640 22880
rect 39704 22816 39720 22880
rect 39784 22816 39792 22880
rect 39472 22815 39792 22816
rect 22737 22808 26296 22810
rect 22737 22752 22742 22808
rect 22798 22752 26296 22808
rect 22737 22750 26296 22752
rect 28073 22810 28139 22813
rect 28390 22810 28396 22812
rect 28073 22808 28396 22810
rect 28073 22752 28078 22808
rect 28134 22752 28396 22808
rect 28073 22750 28396 22752
rect 22737 22747 22803 22750
rect 28073 22747 28139 22750
rect 28390 22748 28396 22750
rect 28460 22810 28466 22812
rect 31477 22810 31543 22813
rect 28460 22808 31543 22810
rect 28460 22752 31482 22808
rect 31538 22752 31543 22808
rect 28460 22750 31543 22752
rect 28460 22748 28466 22750
rect 31477 22747 31543 22750
rect 32121 22810 32187 22813
rect 32397 22810 32463 22813
rect 32121 22808 32463 22810
rect 32121 22752 32126 22808
rect 32182 22752 32402 22808
rect 32458 22752 32463 22808
rect 32121 22750 32463 22752
rect 32121 22747 32187 22750
rect 32397 22747 32463 22750
rect 33501 22810 33567 22813
rect 35893 22810 35959 22813
rect 39021 22810 39087 22813
rect 33501 22808 35634 22810
rect 33501 22752 33506 22808
rect 33562 22752 35634 22808
rect 33501 22750 35634 22752
rect 33501 22747 33567 22750
rect 19149 22674 19215 22677
rect 24393 22674 24459 22677
rect 25773 22676 25839 22677
rect 25773 22674 25820 22676
rect 19149 22672 24459 22674
rect 19149 22616 19154 22672
rect 19210 22616 24398 22672
rect 24454 22616 24459 22672
rect 19149 22614 24459 22616
rect 25728 22672 25820 22674
rect 25728 22616 25778 22672
rect 25728 22614 25820 22616
rect 19149 22611 19215 22614
rect 24393 22611 24459 22614
rect 25773 22612 25820 22614
rect 25884 22612 25890 22676
rect 26233 22674 26299 22677
rect 28574 22674 28580 22676
rect 26233 22672 28580 22674
rect 26233 22616 26238 22672
rect 26294 22616 28580 22672
rect 26233 22614 28580 22616
rect 25773 22611 25839 22612
rect 26233 22611 26299 22614
rect 28574 22612 28580 22614
rect 28644 22674 28650 22676
rect 29126 22674 29132 22676
rect 28644 22614 29132 22674
rect 28644 22612 28650 22614
rect 29126 22612 29132 22614
rect 29196 22612 29202 22676
rect 30097 22674 30163 22677
rect 35341 22674 35407 22677
rect 30097 22672 35407 22674
rect 30097 22616 30102 22672
rect 30158 22616 35346 22672
rect 35402 22616 35407 22672
rect 30097 22614 35407 22616
rect 30097 22611 30163 22614
rect 35341 22611 35407 22614
rect 24117 22540 24183 22541
rect 24117 22538 24164 22540
rect 24072 22536 24164 22538
rect 24072 22480 24122 22536
rect 24072 22478 24164 22480
rect 24117 22476 24164 22478
rect 24228 22476 24234 22540
rect 24945 22538 25011 22541
rect 25078 22538 25084 22540
rect 24945 22536 25084 22538
rect 24945 22480 24950 22536
rect 25006 22480 25084 22536
rect 24945 22478 25084 22480
rect 24117 22475 24183 22476
rect 24945 22475 25011 22478
rect 25078 22476 25084 22478
rect 25148 22476 25154 22540
rect 26693 22538 26759 22541
rect 28073 22538 28139 22541
rect 26693 22536 28139 22538
rect 26693 22480 26698 22536
rect 26754 22480 28078 22536
rect 28134 22480 28139 22536
rect 26693 22478 28139 22480
rect 26693 22475 26759 22478
rect 28073 22475 28139 22478
rect 28625 22538 28691 22541
rect 28901 22538 28967 22541
rect 34646 22538 34652 22540
rect 28625 22536 28826 22538
rect 28625 22480 28630 22536
rect 28686 22480 28826 22536
rect 28625 22478 28826 22480
rect 28625 22475 28691 22478
rect 21582 22340 21588 22404
rect 21652 22402 21658 22404
rect 22001 22402 22067 22405
rect 21652 22400 22067 22402
rect 21652 22344 22006 22400
rect 22062 22344 22067 22400
rect 21652 22342 22067 22344
rect 21652 22340 21658 22342
rect 22001 22339 22067 22342
rect 22829 22402 22895 22405
rect 24342 22402 24348 22404
rect 22829 22400 24348 22402
rect 22829 22344 22834 22400
rect 22890 22344 24348 22400
rect 22829 22342 24348 22344
rect 22829 22339 22895 22342
rect 24342 22340 24348 22342
rect 24412 22340 24418 22404
rect 24669 22402 24735 22405
rect 27337 22402 27403 22405
rect 28766 22402 28826 22478
rect 28901 22536 34652 22538
rect 28901 22480 28906 22536
rect 28962 22480 34652 22536
rect 28901 22478 34652 22480
rect 28901 22475 28967 22478
rect 34646 22476 34652 22478
rect 34716 22476 34722 22540
rect 28901 22402 28967 22405
rect 29269 22404 29335 22405
rect 29269 22402 29316 22404
rect 24669 22400 27538 22402
rect 24669 22344 24674 22400
rect 24730 22344 27342 22400
rect 27398 22344 27538 22400
rect 24669 22342 27538 22344
rect 28766 22400 28967 22402
rect 28766 22344 28906 22400
rect 28962 22344 28967 22400
rect 28766 22342 28967 22344
rect 29224 22400 29316 22402
rect 29224 22344 29274 22400
rect 29224 22342 29316 22344
rect 24669 22339 24735 22342
rect 27337 22339 27403 22342
rect 10576 22336 10896 22337
rect 10576 22272 10584 22336
rect 10648 22272 10664 22336
rect 10728 22272 10744 22336
rect 10808 22272 10824 22336
rect 10888 22272 10896 22336
rect 10576 22271 10896 22272
rect 20662 22204 20668 22268
rect 20732 22266 20738 22268
rect 23381 22266 23447 22269
rect 27337 22266 27403 22269
rect 20732 22206 23306 22266
rect 20732 22204 20738 22206
rect 19885 22132 19951 22133
rect 19885 22128 19932 22132
rect 19996 22130 20002 22132
rect 23246 22130 23306 22206
rect 23381 22264 27403 22266
rect 23381 22208 23386 22264
rect 23442 22208 27342 22264
rect 27398 22208 27403 22264
rect 23381 22206 27403 22208
rect 27478 22266 27538 22342
rect 28901 22339 28967 22342
rect 29269 22340 29316 22342
rect 29380 22340 29386 22404
rect 33133 22402 33199 22405
rect 34462 22402 34468 22404
rect 33133 22400 34468 22402
rect 33133 22344 33138 22400
rect 33194 22344 34468 22400
rect 33133 22342 34468 22344
rect 29269 22339 29335 22340
rect 33133 22339 33199 22342
rect 34462 22340 34468 22342
rect 34532 22340 34538 22404
rect 35574 22402 35634 22750
rect 35893 22808 39087 22810
rect 35893 22752 35898 22808
rect 35954 22752 39026 22808
rect 39082 22752 39087 22808
rect 35893 22750 39087 22752
rect 35893 22747 35959 22750
rect 39021 22747 39087 22750
rect 36721 22674 36787 22677
rect 40401 22674 40467 22677
rect 36721 22672 40467 22674
rect 36721 22616 36726 22672
rect 36782 22616 40406 22672
rect 40462 22616 40467 22672
rect 36721 22614 40467 22616
rect 36721 22611 36787 22614
rect 40401 22611 40467 22614
rect 39573 22538 39639 22541
rect 48773 22538 48839 22541
rect 39573 22536 48839 22538
rect 39573 22480 39578 22536
rect 39634 22480 48778 22536
rect 48834 22480 48839 22536
rect 39573 22478 48839 22480
rect 39573 22475 39639 22478
rect 48773 22475 48839 22478
rect 35574 22342 41430 22402
rect 29840 22336 30160 22337
rect 29840 22272 29848 22336
rect 29912 22272 29928 22336
rect 29992 22272 30008 22336
rect 30072 22272 30088 22336
rect 30152 22272 30160 22336
rect 29840 22271 30160 22272
rect 27981 22266 28047 22269
rect 29494 22266 29500 22268
rect 27478 22264 29500 22266
rect 27478 22208 27986 22264
rect 28042 22208 29500 22264
rect 27478 22206 29500 22208
rect 23381 22203 23447 22206
rect 27337 22203 27403 22206
rect 27981 22203 28047 22206
rect 29494 22204 29500 22206
rect 29564 22204 29570 22268
rect 31017 22266 31083 22269
rect 36169 22266 36235 22269
rect 31017 22264 36235 22266
rect 31017 22208 31022 22264
rect 31078 22208 36174 22264
rect 36230 22208 36235 22264
rect 31017 22206 36235 22208
rect 31017 22203 31083 22206
rect 36169 22203 36235 22206
rect 36721 22266 36787 22269
rect 37038 22266 37044 22268
rect 36721 22264 37044 22266
rect 36721 22208 36726 22264
rect 36782 22208 37044 22264
rect 36721 22206 37044 22208
rect 36721 22203 36787 22206
rect 37038 22204 37044 22206
rect 37108 22204 37114 22268
rect 41370 22266 41430 22342
rect 49104 22336 49424 22337
rect 49104 22272 49112 22336
rect 49176 22272 49192 22336
rect 49256 22272 49272 22336
rect 49336 22272 49352 22336
rect 49416 22272 49424 22336
rect 49104 22271 49424 22272
rect 41873 22266 41939 22269
rect 41370 22264 41939 22266
rect 41370 22208 41878 22264
rect 41934 22208 41939 22264
rect 41370 22206 41939 22208
rect 41873 22203 41939 22206
rect 28073 22130 28139 22133
rect 19885 22072 19890 22128
rect 19885 22068 19932 22072
rect 19996 22070 20042 22130
rect 21406 22070 21834 22130
rect 23246 22128 28139 22130
rect 23246 22072 28078 22128
rect 28134 22072 28139 22128
rect 23246 22070 28139 22072
rect 19996 22068 20002 22070
rect 19885 22067 19951 22068
rect 13905 21994 13971 21997
rect 21406 21994 21466 22070
rect 13905 21992 21466 21994
rect 13905 21936 13910 21992
rect 13966 21936 21466 21992
rect 13905 21934 21466 21936
rect 21774 21994 21834 22070
rect 28073 22067 28139 22070
rect 33133 22130 33199 22133
rect 35341 22130 35407 22133
rect 37774 22130 37780 22132
rect 33133 22128 35266 22130
rect 33133 22072 33138 22128
rect 33194 22072 35266 22128
rect 33133 22070 35266 22072
rect 33133 22067 33199 22070
rect 25129 21994 25195 21997
rect 21774 21992 25195 21994
rect 21774 21936 25134 21992
rect 25190 21936 25195 21992
rect 21774 21934 25195 21936
rect 13905 21931 13971 21934
rect 25129 21931 25195 21934
rect 27061 21994 27127 21997
rect 28165 21994 28231 21997
rect 27061 21992 28231 21994
rect 27061 21936 27066 21992
rect 27122 21936 28170 21992
rect 28226 21936 28231 21992
rect 27061 21934 28231 21936
rect 27061 21931 27127 21934
rect 28165 21931 28231 21934
rect 29126 21932 29132 21996
rect 29196 21994 29202 21996
rect 32581 21994 32647 21997
rect 29196 21992 32647 21994
rect 29196 21936 32586 21992
rect 32642 21936 32647 21992
rect 29196 21934 32647 21936
rect 29196 21932 29202 21934
rect 32581 21931 32647 21934
rect 33685 21996 33751 21997
rect 33685 21992 33732 21996
rect 33796 21994 33802 21996
rect 35206 21994 35266 22070
rect 35341 22128 36738 22130
rect 35341 22072 35346 22128
rect 35402 22072 36738 22128
rect 35341 22070 36738 22072
rect 35341 22067 35407 22070
rect 35985 21994 36051 21997
rect 33685 21936 33690 21992
rect 33685 21932 33732 21936
rect 33796 21934 33842 21994
rect 35206 21992 36051 21994
rect 35206 21936 35990 21992
rect 36046 21936 36051 21992
rect 35206 21934 36051 21936
rect 36678 21994 36738 22070
rect 37046 22070 37780 22130
rect 37046 21994 37106 22070
rect 37774 22068 37780 22070
rect 37844 22130 37850 22132
rect 38837 22130 38903 22133
rect 40033 22130 40099 22133
rect 37844 22128 38903 22130
rect 37844 22072 38842 22128
rect 38898 22072 38903 22128
rect 37844 22070 38903 22072
rect 37844 22068 37850 22070
rect 38837 22067 38903 22070
rect 39254 22128 40099 22130
rect 39254 22072 40038 22128
rect 40094 22072 40099 22128
rect 39254 22070 40099 22072
rect 36678 21934 37106 21994
rect 33796 21932 33802 21934
rect 33685 21931 33751 21932
rect 35985 21931 36051 21934
rect 37590 21932 37596 21996
rect 37660 21994 37666 21996
rect 39254 21994 39314 22070
rect 40033 22067 40099 22070
rect 58157 22130 58223 22133
rect 59200 22130 60000 22160
rect 58157 22128 60000 22130
rect 58157 22072 58162 22128
rect 58218 22072 60000 22128
rect 58157 22070 60000 22072
rect 58157 22067 58223 22070
rect 59200 22040 60000 22070
rect 37660 21934 39314 21994
rect 39849 21994 39915 21997
rect 41505 21994 41571 21997
rect 39849 21992 41571 21994
rect 39849 21936 39854 21992
rect 39910 21936 41510 21992
rect 41566 21936 41571 21992
rect 39849 21934 41571 21936
rect 37660 21932 37666 21934
rect 39849 21931 39915 21934
rect 41505 21931 41571 21934
rect 21633 21858 21699 21861
rect 21766 21858 21772 21860
rect 21633 21856 21772 21858
rect 21633 21800 21638 21856
rect 21694 21800 21772 21856
rect 21633 21798 21772 21800
rect 21633 21795 21699 21798
rect 21766 21796 21772 21798
rect 21836 21796 21842 21860
rect 22093 21858 22159 21861
rect 22093 21856 24824 21858
rect 22093 21800 22098 21856
rect 22154 21800 24824 21856
rect 22093 21798 24824 21800
rect 22093 21795 22159 21798
rect 20208 21792 20528 21793
rect 20208 21728 20216 21792
rect 20280 21728 20296 21792
rect 20360 21728 20376 21792
rect 20440 21728 20456 21792
rect 20520 21728 20528 21792
rect 20208 21727 20528 21728
rect 20621 21722 20687 21725
rect 22829 21722 22895 21725
rect 20621 21720 22895 21722
rect 20621 21664 20626 21720
rect 20682 21664 22834 21720
rect 22890 21664 22895 21720
rect 20621 21662 22895 21664
rect 20621 21659 20687 21662
rect 22829 21659 22895 21662
rect 24342 21660 24348 21724
rect 24412 21722 24418 21724
rect 24577 21722 24643 21725
rect 24412 21720 24643 21722
rect 24412 21664 24582 21720
rect 24638 21664 24643 21720
rect 24412 21662 24643 21664
rect 24764 21722 24824 21798
rect 24894 21796 24900 21860
rect 24964 21858 24970 21860
rect 35065 21858 35131 21861
rect 24964 21856 35131 21858
rect 24964 21800 35070 21856
rect 35126 21800 35131 21856
rect 24964 21798 35131 21800
rect 24964 21796 24970 21798
rect 35065 21795 35131 21798
rect 39472 21792 39792 21793
rect 39472 21728 39480 21792
rect 39544 21728 39560 21792
rect 39624 21728 39640 21792
rect 39704 21728 39720 21792
rect 39784 21728 39792 21792
rect 39472 21727 39792 21728
rect 27889 21724 27955 21725
rect 27838 21722 27844 21724
rect 24764 21662 27844 21722
rect 27908 21720 27955 21724
rect 27950 21664 27955 21720
rect 24412 21660 24418 21662
rect 24577 21659 24643 21662
rect 27838 21660 27844 21662
rect 27908 21660 27955 21664
rect 30966 21660 30972 21724
rect 31036 21722 31042 21724
rect 31937 21722 32003 21725
rect 31036 21720 32003 21722
rect 31036 21664 31942 21720
rect 31998 21664 32003 21720
rect 31036 21662 32003 21664
rect 31036 21660 31042 21662
rect 27889 21659 27955 21660
rect 31937 21659 32003 21662
rect 33041 21722 33107 21725
rect 33358 21722 33364 21724
rect 33041 21720 33364 21722
rect 33041 21664 33046 21720
rect 33102 21664 33364 21720
rect 33041 21662 33364 21664
rect 33041 21659 33107 21662
rect 33358 21660 33364 21662
rect 33428 21660 33434 21724
rect 14457 21586 14523 21589
rect 20897 21586 20963 21589
rect 22185 21586 22251 21589
rect 14457 21584 22251 21586
rect 14457 21528 14462 21584
rect 14518 21528 20902 21584
rect 20958 21528 22190 21584
rect 22246 21528 22251 21584
rect 14457 21526 22251 21528
rect 14457 21523 14523 21526
rect 20897 21523 20963 21526
rect 22185 21523 22251 21526
rect 22686 21524 22692 21588
rect 22756 21586 22762 21588
rect 26550 21586 26556 21588
rect 22756 21526 26556 21586
rect 22756 21524 22762 21526
rect 26550 21524 26556 21526
rect 26620 21524 26626 21588
rect 27470 21524 27476 21588
rect 27540 21586 27546 21588
rect 27613 21586 27679 21589
rect 35801 21586 35867 21589
rect 38101 21586 38167 21589
rect 42149 21586 42215 21589
rect 27540 21584 42215 21586
rect 27540 21528 27618 21584
rect 27674 21528 35806 21584
rect 35862 21528 38106 21584
rect 38162 21528 42154 21584
rect 42210 21528 42215 21584
rect 27540 21526 42215 21528
rect 27540 21524 27546 21526
rect 27613 21523 27679 21526
rect 35801 21523 35867 21526
rect 38101 21523 38167 21526
rect 42149 21523 42215 21526
rect 18270 21388 18276 21452
rect 18340 21450 18346 21452
rect 20161 21450 20227 21453
rect 22921 21450 22987 21453
rect 18340 21448 22987 21450
rect 18340 21392 20166 21448
rect 20222 21392 22926 21448
rect 22982 21392 22987 21448
rect 18340 21390 22987 21392
rect 18340 21388 18346 21390
rect 20161 21387 20227 21390
rect 22921 21387 22987 21390
rect 23105 21450 23171 21453
rect 25037 21450 25103 21453
rect 23105 21448 25103 21450
rect 23105 21392 23110 21448
rect 23166 21392 25042 21448
rect 25098 21392 25103 21448
rect 23105 21390 25103 21392
rect 23105 21387 23171 21390
rect 25037 21387 25103 21390
rect 25497 21450 25563 21453
rect 28165 21450 28231 21453
rect 25497 21448 28231 21450
rect 25497 21392 25502 21448
rect 25558 21392 28170 21448
rect 28226 21392 28231 21448
rect 25497 21390 28231 21392
rect 25497 21387 25563 21390
rect 28165 21387 28231 21390
rect 29494 21388 29500 21452
rect 29564 21450 29570 21452
rect 29564 21390 35450 21450
rect 29564 21388 29570 21390
rect 0 21314 800 21344
rect 1485 21314 1551 21317
rect 0 21312 1551 21314
rect 0 21256 1490 21312
rect 1546 21256 1551 21312
rect 0 21254 1551 21256
rect 0 21224 800 21254
rect 1485 21251 1551 21254
rect 16665 21314 16731 21317
rect 27245 21314 27311 21317
rect 16665 21312 27311 21314
rect 16665 21256 16670 21312
rect 16726 21256 27250 21312
rect 27306 21256 27311 21312
rect 16665 21254 27311 21256
rect 16665 21251 16731 21254
rect 27245 21251 27311 21254
rect 28533 21314 28599 21317
rect 28901 21314 28967 21317
rect 28533 21312 28967 21314
rect 28533 21256 28538 21312
rect 28594 21256 28906 21312
rect 28962 21256 28967 21312
rect 28533 21254 28967 21256
rect 28533 21251 28599 21254
rect 28901 21251 28967 21254
rect 30557 21314 30623 21317
rect 30782 21314 30788 21316
rect 30557 21312 30788 21314
rect 30557 21256 30562 21312
rect 30618 21256 30788 21312
rect 30557 21254 30788 21256
rect 30557 21251 30623 21254
rect 30782 21252 30788 21254
rect 30852 21252 30858 21316
rect 32213 21314 32279 21317
rect 32489 21314 32555 21317
rect 32213 21312 32555 21314
rect 32213 21256 32218 21312
rect 32274 21256 32494 21312
rect 32550 21256 32555 21312
rect 32213 21254 32555 21256
rect 35390 21314 35450 21390
rect 35566 21388 35572 21452
rect 35636 21450 35642 21452
rect 40585 21450 40651 21453
rect 35636 21448 40651 21450
rect 35636 21392 40590 21448
rect 40646 21392 40651 21448
rect 35636 21390 40651 21392
rect 35636 21388 35642 21390
rect 40585 21387 40651 21390
rect 36905 21314 36971 21317
rect 35390 21312 36971 21314
rect 35390 21256 36910 21312
rect 36966 21256 36971 21312
rect 35390 21254 36971 21256
rect 32213 21251 32279 21254
rect 32489 21251 32555 21254
rect 36905 21251 36971 21254
rect 37958 21252 37964 21316
rect 38028 21314 38034 21316
rect 44909 21314 44975 21317
rect 38028 21312 44975 21314
rect 38028 21256 44914 21312
rect 44970 21256 44975 21312
rect 38028 21254 44975 21256
rect 38028 21252 38034 21254
rect 44909 21251 44975 21254
rect 10576 21248 10896 21249
rect 10576 21184 10584 21248
rect 10648 21184 10664 21248
rect 10728 21184 10744 21248
rect 10808 21184 10824 21248
rect 10888 21184 10896 21248
rect 10576 21183 10896 21184
rect 29840 21248 30160 21249
rect 29840 21184 29848 21248
rect 29912 21184 29928 21248
rect 29992 21184 30008 21248
rect 30072 21184 30088 21248
rect 30152 21184 30160 21248
rect 29840 21183 30160 21184
rect 49104 21248 49424 21249
rect 49104 21184 49112 21248
rect 49176 21184 49192 21248
rect 49256 21184 49272 21248
rect 49336 21184 49352 21248
rect 49416 21184 49424 21248
rect 49104 21183 49424 21184
rect 21817 21178 21883 21181
rect 24301 21178 24367 21181
rect 21817 21176 24367 21178
rect 21817 21120 21822 21176
rect 21878 21120 24306 21176
rect 24362 21120 24367 21176
rect 21817 21118 24367 21120
rect 21817 21115 21883 21118
rect 24301 21115 24367 21118
rect 30281 21178 30347 21181
rect 40493 21178 40559 21181
rect 42057 21180 42123 21181
rect 30281 21176 40559 21178
rect 30281 21120 30286 21176
rect 30342 21120 40498 21176
rect 40554 21120 40559 21176
rect 30281 21118 40559 21120
rect 30281 21115 30347 21118
rect 40493 21115 40559 21118
rect 42006 21116 42012 21180
rect 42076 21178 42123 21180
rect 42076 21176 42168 21178
rect 42118 21120 42168 21176
rect 42076 21118 42168 21120
rect 42076 21116 42123 21118
rect 42057 21115 42123 21116
rect 17033 21042 17099 21045
rect 23105 21042 23171 21045
rect 17033 21040 23171 21042
rect 17033 20984 17038 21040
rect 17094 20984 23110 21040
rect 23166 20984 23171 21040
rect 17033 20982 23171 20984
rect 17033 20979 17099 20982
rect 23105 20979 23171 20982
rect 23749 21042 23815 21045
rect 38561 21042 38627 21045
rect 23749 21040 38627 21042
rect 23749 20984 23754 21040
rect 23810 20984 38566 21040
rect 38622 20984 38627 21040
rect 23749 20982 38627 20984
rect 23749 20979 23815 20982
rect 38561 20979 38627 20982
rect 39297 21042 39363 21045
rect 42241 21042 42307 21045
rect 39297 21040 42307 21042
rect 39297 20984 39302 21040
rect 39358 20984 42246 21040
rect 42302 20984 42307 21040
rect 39297 20982 42307 20984
rect 39297 20979 39363 20982
rect 42241 20979 42307 20982
rect 19701 20906 19767 20909
rect 29177 20906 29243 20909
rect 19701 20904 29243 20906
rect 19701 20848 19706 20904
rect 19762 20848 29182 20904
rect 29238 20848 29243 20904
rect 19701 20846 29243 20848
rect 19701 20843 19767 20846
rect 29177 20843 29243 20846
rect 29913 20906 29979 20909
rect 33225 20906 33291 20909
rect 29913 20904 33291 20906
rect 29913 20848 29918 20904
rect 29974 20848 33230 20904
rect 33286 20848 33291 20904
rect 29913 20846 33291 20848
rect 29913 20843 29979 20846
rect 33225 20843 33291 20846
rect 37181 20906 37247 20909
rect 43529 20906 43595 20909
rect 37181 20904 43595 20906
rect 37181 20848 37186 20904
rect 37242 20848 43534 20904
rect 43590 20848 43595 20904
rect 37181 20846 43595 20848
rect 37181 20843 37247 20846
rect 43529 20843 43595 20846
rect 20805 20770 20871 20773
rect 22686 20770 22692 20772
rect 20805 20768 22692 20770
rect 20805 20712 20810 20768
rect 20866 20712 22692 20768
rect 20805 20710 22692 20712
rect 20805 20707 20871 20710
rect 22686 20708 22692 20710
rect 22756 20708 22762 20772
rect 22829 20770 22895 20773
rect 29545 20770 29611 20773
rect 22829 20768 29611 20770
rect 22829 20712 22834 20768
rect 22890 20712 29550 20768
rect 29606 20712 29611 20768
rect 22829 20710 29611 20712
rect 22829 20707 22895 20710
rect 29545 20707 29611 20710
rect 30373 20770 30439 20773
rect 32305 20772 32371 20773
rect 30782 20770 30788 20772
rect 30373 20768 30788 20770
rect 30373 20712 30378 20768
rect 30434 20712 30788 20768
rect 30373 20710 30788 20712
rect 30373 20707 30439 20710
rect 30782 20708 30788 20710
rect 30852 20708 30858 20772
rect 32254 20770 32260 20772
rect 32214 20710 32260 20770
rect 32324 20768 32371 20772
rect 32366 20712 32371 20768
rect 32254 20708 32260 20710
rect 32324 20708 32371 20712
rect 32305 20707 32371 20708
rect 34237 20770 34303 20773
rect 36629 20770 36695 20773
rect 34237 20768 36695 20770
rect 34237 20712 34242 20768
rect 34298 20712 36634 20768
rect 36690 20712 36695 20768
rect 34237 20710 36695 20712
rect 34237 20707 34303 20710
rect 36629 20707 36695 20710
rect 36854 20708 36860 20772
rect 36924 20770 36930 20772
rect 39113 20770 39179 20773
rect 36924 20768 39179 20770
rect 36924 20712 39118 20768
rect 39174 20712 39179 20768
rect 36924 20710 39179 20712
rect 36924 20708 36930 20710
rect 39113 20707 39179 20710
rect 20208 20704 20528 20705
rect 20208 20640 20216 20704
rect 20280 20640 20296 20704
rect 20360 20640 20376 20704
rect 20440 20640 20456 20704
rect 20520 20640 20528 20704
rect 20208 20639 20528 20640
rect 39472 20704 39792 20705
rect 39472 20640 39480 20704
rect 39544 20640 39560 20704
rect 39624 20640 39640 20704
rect 39704 20640 39720 20704
rect 39784 20640 39792 20704
rect 39472 20639 39792 20640
rect 22553 20634 22619 20637
rect 23473 20634 23539 20637
rect 22553 20632 23539 20634
rect 22553 20576 22558 20632
rect 22614 20576 23478 20632
rect 23534 20576 23539 20632
rect 22553 20574 23539 20576
rect 22553 20571 22619 20574
rect 23473 20571 23539 20574
rect 24577 20634 24643 20637
rect 30741 20634 30807 20637
rect 24577 20632 30807 20634
rect 24577 20576 24582 20632
rect 24638 20576 30746 20632
rect 30802 20576 30807 20632
rect 24577 20574 30807 20576
rect 24577 20571 24643 20574
rect 30741 20571 30807 20574
rect 17953 20498 18019 20501
rect 19190 20498 19196 20500
rect 17953 20496 19196 20498
rect 17953 20440 17958 20496
rect 18014 20440 19196 20496
rect 17953 20438 19196 20440
rect 17953 20435 18019 20438
rect 19190 20436 19196 20438
rect 19260 20436 19266 20500
rect 19793 20498 19859 20501
rect 20662 20498 20668 20500
rect 19793 20496 20668 20498
rect 19793 20440 19798 20496
rect 19854 20440 20668 20496
rect 19793 20438 20668 20440
rect 19793 20435 19859 20438
rect 20662 20436 20668 20438
rect 20732 20436 20738 20500
rect 22093 20498 22159 20501
rect 27102 20498 27108 20500
rect 22093 20496 27108 20498
rect 22093 20440 22098 20496
rect 22154 20440 27108 20496
rect 22093 20438 27108 20440
rect 22093 20435 22159 20438
rect 27102 20436 27108 20438
rect 27172 20436 27178 20500
rect 27245 20498 27311 20501
rect 37641 20498 37707 20501
rect 40401 20498 40467 20501
rect 27245 20496 40467 20498
rect 27245 20440 27250 20496
rect 27306 20440 37646 20496
rect 37702 20440 40406 20496
rect 40462 20440 40467 20496
rect 27245 20438 40467 20440
rect 27245 20435 27311 20438
rect 37641 20435 37707 20438
rect 40401 20435 40467 20438
rect 15561 20362 15627 20365
rect 26049 20362 26115 20365
rect 15561 20360 26115 20362
rect 15561 20304 15566 20360
rect 15622 20304 26054 20360
rect 26110 20304 26115 20360
rect 15561 20302 26115 20304
rect 15561 20299 15627 20302
rect 26049 20299 26115 20302
rect 28390 20300 28396 20364
rect 28460 20362 28466 20364
rect 29821 20362 29887 20365
rect 30741 20362 30807 20365
rect 37917 20362 37983 20365
rect 43161 20362 43227 20365
rect 28460 20360 30298 20362
rect 28460 20304 29826 20360
rect 29882 20304 30298 20360
rect 28460 20302 30298 20304
rect 28460 20300 28466 20302
rect 29821 20299 29887 20302
rect 18965 20226 19031 20229
rect 27153 20226 27219 20229
rect 18965 20224 27219 20226
rect 18965 20168 18970 20224
rect 19026 20168 27158 20224
rect 27214 20168 27219 20224
rect 18965 20166 27219 20168
rect 18965 20163 19031 20166
rect 27153 20163 27219 20166
rect 10576 20160 10896 20161
rect 10576 20096 10584 20160
rect 10648 20096 10664 20160
rect 10728 20096 10744 20160
rect 10808 20096 10824 20160
rect 10888 20096 10896 20160
rect 10576 20095 10896 20096
rect 29840 20160 30160 20161
rect 29840 20096 29848 20160
rect 29912 20096 29928 20160
rect 29992 20096 30008 20160
rect 30072 20096 30088 20160
rect 30152 20096 30160 20160
rect 29840 20095 30160 20096
rect 18229 20090 18295 20093
rect 21173 20092 21239 20093
rect 20846 20090 20852 20092
rect 18229 20088 20852 20090
rect 18229 20032 18234 20088
rect 18290 20032 20852 20088
rect 18229 20030 20852 20032
rect 18229 20027 18295 20030
rect 20846 20028 20852 20030
rect 20916 20028 20922 20092
rect 21173 20090 21220 20092
rect 21128 20088 21220 20090
rect 21128 20032 21178 20088
rect 21128 20030 21220 20032
rect 21173 20028 21220 20030
rect 21284 20028 21290 20092
rect 21909 20090 21975 20093
rect 23565 20090 23631 20093
rect 21909 20088 23631 20090
rect 21909 20032 21914 20088
rect 21970 20032 23570 20088
rect 23626 20032 23631 20088
rect 21909 20030 23631 20032
rect 21173 20027 21239 20028
rect 21909 20027 21975 20030
rect 23565 20027 23631 20030
rect 24853 20090 24919 20093
rect 25773 20090 25839 20093
rect 24853 20088 25839 20090
rect 24853 20032 24858 20088
rect 24914 20032 25778 20088
rect 25834 20032 25839 20088
rect 24853 20030 25839 20032
rect 30238 20090 30298 20302
rect 30741 20360 43227 20362
rect 30741 20304 30746 20360
rect 30802 20304 37922 20360
rect 37978 20304 43166 20360
rect 43222 20304 43227 20360
rect 30741 20302 43227 20304
rect 30741 20299 30807 20302
rect 37917 20299 37983 20302
rect 43161 20299 43227 20302
rect 58157 20362 58223 20365
rect 59200 20362 60000 20392
rect 58157 20360 60000 20362
rect 58157 20304 58162 20360
rect 58218 20304 60000 20360
rect 58157 20302 60000 20304
rect 58157 20299 58223 20302
rect 59200 20272 60000 20302
rect 30465 20226 30531 20229
rect 32949 20226 33015 20229
rect 30465 20224 33015 20226
rect 30465 20168 30470 20224
rect 30526 20168 32954 20224
rect 33010 20168 33015 20224
rect 30465 20166 33015 20168
rect 30465 20163 30531 20166
rect 32949 20163 33015 20166
rect 33409 20226 33475 20229
rect 35617 20226 35683 20229
rect 33409 20224 35683 20226
rect 33409 20168 33414 20224
rect 33470 20168 35622 20224
rect 35678 20168 35683 20224
rect 33409 20166 35683 20168
rect 33409 20163 33475 20166
rect 35617 20163 35683 20166
rect 35934 20164 35940 20228
rect 36004 20226 36010 20228
rect 42609 20226 42675 20229
rect 36004 20224 42675 20226
rect 36004 20168 42614 20224
rect 42670 20168 42675 20224
rect 36004 20166 42675 20168
rect 36004 20164 36010 20166
rect 42609 20163 42675 20166
rect 49104 20160 49424 20161
rect 49104 20096 49112 20160
rect 49176 20096 49192 20160
rect 49256 20096 49272 20160
rect 49336 20096 49352 20160
rect 49416 20096 49424 20160
rect 49104 20095 49424 20096
rect 32673 20090 32739 20093
rect 34278 20090 34284 20092
rect 30238 20088 34284 20090
rect 30238 20032 32678 20088
rect 32734 20032 34284 20088
rect 30238 20030 34284 20032
rect 24853 20027 24919 20030
rect 25773 20027 25839 20030
rect 32673 20027 32739 20030
rect 34278 20028 34284 20030
rect 34348 20090 34354 20092
rect 39757 20090 39823 20093
rect 34348 20088 39823 20090
rect 34348 20032 39762 20088
rect 39818 20032 39823 20088
rect 34348 20030 39823 20032
rect 34348 20028 34354 20030
rect 39757 20027 39823 20030
rect 18045 19954 18111 19957
rect 21030 19954 21036 19956
rect 18045 19952 21036 19954
rect 18045 19896 18050 19952
rect 18106 19896 21036 19952
rect 18045 19894 21036 19896
rect 18045 19891 18111 19894
rect 21030 19892 21036 19894
rect 21100 19954 21106 19956
rect 22369 19954 22435 19957
rect 21100 19952 22435 19954
rect 21100 19896 22374 19952
rect 22430 19896 22435 19952
rect 21100 19894 22435 19896
rect 21100 19892 21106 19894
rect 22369 19891 22435 19894
rect 22502 19892 22508 19956
rect 22572 19954 22578 19956
rect 26693 19954 26759 19957
rect 22572 19952 26759 19954
rect 22572 19896 26698 19952
rect 26754 19896 26759 19952
rect 22572 19894 26759 19896
rect 22572 19892 22578 19894
rect 26693 19891 26759 19894
rect 28625 19954 28691 19957
rect 28758 19954 28764 19956
rect 28625 19952 28764 19954
rect 28625 19896 28630 19952
rect 28686 19896 28764 19952
rect 28625 19894 28764 19896
rect 28625 19891 28691 19894
rect 28758 19892 28764 19894
rect 28828 19892 28834 19956
rect 33777 19954 33843 19957
rect 35157 19954 35223 19957
rect 33777 19952 35223 19954
rect 33777 19896 33782 19952
rect 33838 19896 35162 19952
rect 35218 19896 35223 19952
rect 33777 19894 35223 19896
rect 33777 19891 33843 19894
rect 35157 19891 35223 19894
rect 39205 19954 39271 19957
rect 43253 19954 43319 19957
rect 39205 19952 43319 19954
rect 39205 19896 39210 19952
rect 39266 19896 43258 19952
rect 43314 19896 43319 19952
rect 39205 19894 43319 19896
rect 39205 19891 39271 19894
rect 43253 19891 43319 19894
rect 18638 19756 18644 19820
rect 18708 19818 18714 19820
rect 19425 19818 19491 19821
rect 27838 19818 27844 19820
rect 18708 19758 19258 19818
rect 18708 19756 18714 19758
rect 0 19682 800 19712
rect 1485 19682 1551 19685
rect 0 19680 1551 19682
rect 0 19624 1490 19680
rect 1546 19624 1551 19680
rect 0 19622 1551 19624
rect 0 19592 800 19622
rect 1485 19619 1551 19622
rect 14273 19682 14339 19685
rect 18873 19682 18939 19685
rect 14273 19680 18939 19682
rect 14273 19624 14278 19680
rect 14334 19624 18878 19680
rect 18934 19624 18939 19680
rect 14273 19622 18939 19624
rect 14273 19619 14339 19622
rect 18873 19619 18939 19622
rect 18822 19484 18828 19548
rect 18892 19546 18898 19548
rect 19057 19546 19123 19549
rect 18892 19544 19123 19546
rect 18892 19488 19062 19544
rect 19118 19488 19123 19544
rect 18892 19486 19123 19488
rect 18892 19484 18898 19486
rect 19057 19483 19123 19486
rect 14825 19410 14891 19413
rect 18638 19410 18644 19412
rect 14825 19408 18644 19410
rect 14825 19352 14830 19408
rect 14886 19352 18644 19408
rect 14825 19350 18644 19352
rect 14825 19347 14891 19350
rect 18638 19348 18644 19350
rect 18708 19348 18714 19412
rect 19198 19410 19258 19758
rect 19425 19816 27844 19818
rect 19425 19760 19430 19816
rect 19486 19760 27844 19816
rect 19425 19758 27844 19760
rect 19425 19755 19491 19758
rect 27838 19756 27844 19758
rect 27908 19756 27914 19820
rect 33041 19818 33107 19821
rect 40125 19818 40191 19821
rect 41045 19818 41111 19821
rect 33041 19816 41111 19818
rect 33041 19760 33046 19816
rect 33102 19760 40130 19816
rect 40186 19760 41050 19816
rect 41106 19760 41111 19816
rect 33041 19758 41111 19760
rect 33041 19755 33107 19758
rect 40125 19755 40191 19758
rect 41045 19755 41111 19758
rect 42517 19818 42583 19821
rect 48497 19818 48563 19821
rect 42517 19816 48563 19818
rect 42517 19760 42522 19816
rect 42578 19760 48502 19816
rect 48558 19760 48563 19816
rect 42517 19758 48563 19760
rect 42517 19755 42583 19758
rect 48497 19755 48563 19758
rect 21357 19682 21423 19685
rect 24853 19682 24919 19685
rect 27153 19684 27219 19685
rect 21357 19680 24919 19682
rect 21357 19624 21362 19680
rect 21418 19624 24858 19680
rect 24914 19624 24919 19680
rect 21357 19622 24919 19624
rect 21357 19619 21423 19622
rect 24853 19619 24919 19622
rect 27102 19620 27108 19684
rect 27172 19682 27219 19684
rect 27429 19682 27495 19685
rect 33317 19682 33383 19685
rect 27172 19680 27264 19682
rect 27214 19624 27264 19680
rect 27172 19622 27264 19624
rect 27429 19680 33383 19682
rect 27429 19624 27434 19680
rect 27490 19624 33322 19680
rect 33378 19624 33383 19680
rect 27429 19622 33383 19624
rect 27172 19620 27219 19622
rect 27153 19619 27219 19620
rect 27429 19619 27495 19622
rect 33317 19619 33383 19622
rect 34646 19620 34652 19684
rect 34716 19682 34722 19684
rect 37457 19682 37523 19685
rect 34716 19680 37523 19682
rect 34716 19624 37462 19680
rect 37518 19624 37523 19680
rect 34716 19622 37523 19624
rect 34716 19620 34722 19622
rect 37457 19619 37523 19622
rect 40033 19682 40099 19685
rect 47761 19682 47827 19685
rect 40033 19680 47827 19682
rect 40033 19624 40038 19680
rect 40094 19624 47766 19680
rect 47822 19624 47827 19680
rect 40033 19622 47827 19624
rect 40033 19619 40099 19622
rect 47761 19619 47827 19622
rect 20208 19616 20528 19617
rect 20208 19552 20216 19616
rect 20280 19552 20296 19616
rect 20360 19552 20376 19616
rect 20440 19552 20456 19616
rect 20520 19552 20528 19616
rect 20208 19551 20528 19552
rect 39472 19616 39792 19617
rect 39472 19552 39480 19616
rect 39544 19552 39560 19616
rect 39624 19552 39640 19616
rect 39704 19552 39720 19616
rect 39784 19552 39792 19616
rect 39472 19551 39792 19552
rect 20662 19484 20668 19548
rect 20732 19546 20738 19548
rect 21081 19546 21147 19549
rect 27102 19546 27108 19548
rect 20732 19544 21147 19546
rect 20732 19488 21086 19544
rect 21142 19488 21147 19544
rect 20732 19486 21147 19488
rect 20732 19484 20738 19486
rect 21081 19483 21147 19486
rect 23384 19486 27108 19546
rect 21449 19410 21515 19413
rect 22185 19412 22251 19413
rect 19198 19408 21515 19410
rect 19198 19352 21454 19408
rect 21510 19352 21515 19408
rect 19198 19350 21515 19352
rect 21449 19347 21515 19350
rect 22134 19348 22140 19412
rect 22204 19410 22251 19412
rect 23384 19410 23444 19486
rect 27102 19484 27108 19486
rect 27172 19546 27178 19548
rect 29269 19546 29335 19549
rect 27172 19544 29335 19546
rect 27172 19488 29274 19544
rect 29330 19488 29335 19544
rect 27172 19486 29335 19488
rect 27172 19484 27178 19486
rect 29269 19483 29335 19486
rect 29494 19484 29500 19548
rect 29564 19546 29570 19548
rect 31201 19546 31267 19549
rect 35709 19546 35775 19549
rect 29564 19544 31267 19546
rect 29564 19488 31206 19544
rect 31262 19488 31267 19544
rect 29564 19486 31267 19488
rect 29564 19484 29570 19486
rect 31201 19483 31267 19486
rect 32078 19544 35775 19546
rect 32078 19488 35714 19544
rect 35770 19488 35775 19544
rect 32078 19486 35775 19488
rect 22204 19408 23444 19410
rect 22246 19352 23444 19408
rect 22204 19350 23444 19352
rect 23841 19410 23907 19413
rect 27286 19410 27292 19412
rect 23841 19408 27292 19410
rect 23841 19352 23846 19408
rect 23902 19352 27292 19408
rect 23841 19350 27292 19352
rect 22204 19348 22251 19350
rect 22185 19347 22251 19348
rect 23841 19347 23907 19350
rect 27286 19348 27292 19350
rect 27356 19348 27362 19412
rect 28022 19348 28028 19412
rect 28092 19410 28098 19412
rect 28165 19410 28231 19413
rect 28092 19408 28231 19410
rect 28092 19352 28170 19408
rect 28226 19352 28231 19408
rect 28092 19350 28231 19352
rect 28092 19348 28098 19350
rect 28165 19347 28231 19350
rect 29177 19410 29243 19413
rect 32078 19410 32138 19486
rect 35709 19483 35775 19486
rect 35893 19546 35959 19549
rect 36670 19546 36676 19548
rect 35893 19544 36676 19546
rect 35893 19488 35898 19544
rect 35954 19488 36676 19544
rect 35893 19486 36676 19488
rect 35893 19483 35959 19486
rect 36670 19484 36676 19486
rect 36740 19484 36746 19548
rect 39944 19486 42626 19546
rect 29177 19408 32138 19410
rect 29177 19352 29182 19408
rect 29238 19352 32138 19408
rect 29177 19350 32138 19352
rect 32213 19410 32279 19413
rect 33593 19410 33659 19413
rect 32213 19408 33659 19410
rect 32213 19352 32218 19408
rect 32274 19352 33598 19408
rect 33654 19352 33659 19408
rect 32213 19350 33659 19352
rect 29177 19347 29243 19350
rect 32213 19347 32279 19350
rect 33593 19347 33659 19350
rect 38745 19410 38811 19413
rect 39944 19410 40004 19486
rect 40953 19412 41019 19413
rect 38745 19408 40004 19410
rect 38745 19352 38750 19408
rect 38806 19352 40004 19408
rect 38745 19350 40004 19352
rect 38745 19347 38811 19350
rect 40902 19348 40908 19412
rect 40972 19410 41019 19412
rect 41597 19412 41663 19413
rect 40972 19408 41064 19410
rect 41014 19352 41064 19408
rect 40972 19350 41064 19352
rect 41597 19408 41644 19412
rect 41708 19410 41714 19412
rect 42566 19410 42626 19486
rect 42701 19412 42767 19413
rect 42701 19410 42748 19412
rect 41597 19352 41602 19408
rect 40972 19348 41019 19350
rect 40953 19347 41019 19348
rect 41597 19348 41644 19352
rect 41708 19350 41754 19410
rect 42566 19408 42748 19410
rect 42812 19410 42818 19412
rect 44541 19410 44607 19413
rect 42812 19408 44607 19410
rect 42566 19352 42706 19408
rect 42812 19352 44546 19408
rect 44602 19352 44607 19408
rect 42566 19350 42748 19352
rect 41708 19348 41714 19350
rect 42701 19348 42748 19350
rect 42812 19350 44607 19352
rect 42812 19348 42818 19350
rect 41597 19347 41663 19348
rect 42701 19347 42767 19348
rect 44541 19347 44607 19350
rect 16757 19276 16823 19277
rect 16757 19274 16804 19276
rect 16712 19272 16804 19274
rect 16712 19216 16762 19272
rect 16712 19214 16804 19216
rect 16757 19212 16804 19214
rect 16868 19212 16874 19276
rect 17166 19212 17172 19276
rect 17236 19274 17242 19276
rect 17677 19274 17743 19277
rect 17236 19272 17743 19274
rect 17236 19216 17682 19272
rect 17738 19216 17743 19272
rect 17236 19214 17743 19216
rect 17236 19212 17242 19214
rect 16757 19211 16823 19212
rect 17677 19211 17743 19214
rect 18086 19212 18092 19276
rect 18156 19274 18162 19276
rect 18965 19274 19031 19277
rect 18156 19272 19031 19274
rect 18156 19216 18970 19272
rect 19026 19216 19031 19272
rect 18156 19214 19031 19216
rect 18156 19212 18162 19214
rect 18965 19211 19031 19214
rect 19926 19212 19932 19276
rect 19996 19274 20002 19276
rect 20345 19274 20411 19277
rect 19996 19272 20411 19274
rect 19996 19216 20350 19272
rect 20406 19216 20411 19272
rect 19996 19214 20411 19216
rect 19996 19212 20002 19214
rect 20345 19211 20411 19214
rect 20846 19212 20852 19276
rect 20916 19274 20922 19276
rect 24945 19274 25011 19277
rect 20916 19272 25011 19274
rect 20916 19216 24950 19272
rect 25006 19216 25011 19272
rect 20916 19214 25011 19216
rect 20916 19212 20922 19214
rect 24945 19211 25011 19214
rect 25262 19212 25268 19276
rect 25332 19274 25338 19276
rect 25405 19274 25471 19277
rect 25332 19272 25471 19274
rect 25332 19216 25410 19272
rect 25466 19216 25471 19272
rect 25332 19214 25471 19216
rect 25332 19212 25338 19214
rect 25405 19211 25471 19214
rect 28533 19274 28599 19277
rect 28533 19272 31770 19274
rect 28533 19216 28538 19272
rect 28594 19216 31770 19272
rect 28533 19214 31770 19216
rect 28533 19211 28599 19214
rect 16205 19138 16271 19141
rect 18229 19138 18295 19141
rect 16205 19136 18295 19138
rect 16205 19080 16210 19136
rect 16266 19080 18234 19136
rect 18290 19080 18295 19136
rect 16205 19078 18295 19080
rect 16205 19075 16271 19078
rect 18229 19075 18295 19078
rect 18873 19138 18939 19141
rect 19006 19138 19012 19140
rect 18873 19136 19012 19138
rect 18873 19080 18878 19136
rect 18934 19080 19012 19136
rect 18873 19078 19012 19080
rect 18873 19075 18939 19078
rect 19006 19076 19012 19078
rect 19076 19076 19082 19140
rect 19190 19076 19196 19140
rect 19260 19138 19266 19140
rect 22461 19138 22527 19141
rect 25078 19138 25084 19140
rect 19260 19136 22527 19138
rect 19260 19080 22466 19136
rect 22522 19080 22527 19136
rect 19260 19078 22527 19080
rect 19260 19076 19266 19078
rect 22461 19075 22527 19078
rect 22648 19078 25084 19138
rect 10576 19072 10896 19073
rect 10576 19008 10584 19072
rect 10648 19008 10664 19072
rect 10728 19008 10744 19072
rect 10808 19008 10824 19072
rect 10888 19008 10896 19072
rect 10576 19007 10896 19008
rect 16481 19002 16547 19005
rect 17309 19002 17375 19005
rect 16481 19000 17375 19002
rect 16481 18944 16486 19000
rect 16542 18944 17314 19000
rect 17370 18944 17375 19000
rect 16481 18942 17375 18944
rect 16481 18939 16547 18942
rect 17309 18939 17375 18942
rect 17585 19002 17651 19005
rect 17902 19002 17908 19004
rect 17585 19000 17908 19002
rect 17585 18944 17590 19000
rect 17646 18944 17908 19000
rect 17585 18942 17908 18944
rect 17585 18939 17651 18942
rect 17902 18940 17908 18942
rect 17972 18940 17978 19004
rect 18137 19002 18203 19005
rect 18270 19002 18276 19004
rect 18137 19000 18276 19002
rect 18137 18944 18142 19000
rect 18198 18944 18276 19000
rect 18137 18942 18276 18944
rect 18137 18939 18203 18942
rect 18270 18940 18276 18942
rect 18340 18940 18346 19004
rect 18689 19002 18755 19005
rect 22648 19002 22708 19078
rect 25078 19076 25084 19078
rect 25148 19138 25154 19140
rect 29494 19138 29500 19140
rect 25148 19078 29500 19138
rect 25148 19076 25154 19078
rect 29494 19076 29500 19078
rect 29564 19076 29570 19140
rect 31710 19138 31770 19214
rect 33726 19212 33732 19276
rect 33796 19274 33802 19276
rect 36997 19274 37063 19277
rect 33796 19272 37063 19274
rect 33796 19216 37002 19272
rect 37058 19216 37063 19272
rect 33796 19214 37063 19216
rect 33796 19212 33802 19214
rect 36997 19211 37063 19214
rect 37273 19274 37339 19277
rect 38653 19276 38719 19277
rect 37406 19274 37412 19276
rect 37273 19272 37412 19274
rect 37273 19216 37278 19272
rect 37334 19216 37412 19272
rect 37273 19214 37412 19216
rect 37273 19211 37339 19214
rect 37406 19212 37412 19214
rect 37476 19212 37482 19276
rect 38653 19272 38700 19276
rect 38764 19274 38770 19276
rect 38653 19216 38658 19272
rect 38653 19212 38700 19216
rect 38764 19214 38810 19274
rect 38764 19212 38770 19214
rect 38653 19211 38719 19212
rect 43253 19138 43319 19141
rect 31710 19136 43319 19138
rect 31710 19080 43258 19136
rect 43314 19080 43319 19136
rect 31710 19078 43319 19080
rect 43253 19075 43319 19078
rect 29840 19072 30160 19073
rect 29840 19008 29848 19072
rect 29912 19008 29928 19072
rect 29992 19008 30008 19072
rect 30072 19008 30088 19072
rect 30152 19008 30160 19072
rect 29840 19007 30160 19008
rect 49104 19072 49424 19073
rect 49104 19008 49112 19072
rect 49176 19008 49192 19072
rect 49256 19008 49272 19072
rect 49336 19008 49352 19072
rect 49416 19008 49424 19072
rect 49104 19007 49424 19008
rect 18689 19000 22708 19002
rect 18689 18944 18694 19000
rect 18750 18944 22708 19000
rect 18689 18942 22708 18944
rect 24853 19002 24919 19005
rect 29361 19002 29427 19005
rect 24853 19000 29427 19002
rect 24853 18944 24858 19000
rect 24914 18944 29366 19000
rect 29422 18944 29427 19000
rect 24853 18942 29427 18944
rect 18689 18939 18755 18942
rect 24853 18939 24919 18942
rect 29361 18939 29427 18942
rect 30598 18940 30604 19004
rect 30668 19002 30674 19004
rect 43897 19002 43963 19005
rect 30668 19000 43963 19002
rect 30668 18944 43902 19000
rect 43958 18944 43963 19000
rect 30668 18942 43963 18944
rect 30668 18940 30674 18942
rect 43897 18939 43963 18942
rect 14181 18866 14247 18869
rect 26049 18866 26115 18869
rect 14181 18864 26115 18866
rect 14181 18808 14186 18864
rect 14242 18808 26054 18864
rect 26110 18808 26115 18864
rect 14181 18806 26115 18808
rect 14181 18803 14247 18806
rect 26049 18803 26115 18806
rect 29678 18804 29684 18868
rect 29748 18866 29754 18868
rect 29821 18866 29887 18869
rect 29748 18864 29887 18866
rect 29748 18808 29826 18864
rect 29882 18808 29887 18864
rect 29748 18806 29887 18808
rect 29748 18804 29754 18806
rect 29821 18803 29887 18806
rect 30373 18866 30439 18869
rect 39481 18866 39547 18869
rect 30373 18864 39547 18866
rect 30373 18808 30378 18864
rect 30434 18808 39486 18864
rect 39542 18808 39547 18864
rect 30373 18806 39547 18808
rect 30373 18803 30439 18806
rect 39481 18803 39547 18806
rect 15009 18730 15075 18733
rect 17309 18730 17375 18733
rect 15009 18728 17375 18730
rect 15009 18672 15014 18728
rect 15070 18672 17314 18728
rect 17370 18672 17375 18728
rect 15009 18670 17375 18672
rect 15009 18667 15075 18670
rect 17309 18667 17375 18670
rect 18229 18730 18295 18733
rect 21357 18730 21423 18733
rect 23105 18730 23171 18733
rect 18229 18728 21423 18730
rect 18229 18672 18234 18728
rect 18290 18672 21362 18728
rect 21418 18672 21423 18728
rect 18229 18670 21423 18672
rect 18229 18667 18295 18670
rect 21357 18667 21423 18670
rect 21544 18728 23171 18730
rect 21544 18672 23110 18728
rect 23166 18672 23171 18728
rect 21544 18670 23171 18672
rect 16430 18532 16436 18596
rect 16500 18594 16506 18596
rect 19149 18594 19215 18597
rect 19425 18596 19491 18597
rect 16500 18592 19215 18594
rect 16500 18536 19154 18592
rect 19210 18536 19215 18592
rect 16500 18534 19215 18536
rect 16500 18532 16506 18534
rect 19149 18531 19215 18534
rect 19374 18532 19380 18596
rect 19444 18594 19491 18596
rect 19444 18592 19536 18594
rect 19486 18536 19536 18592
rect 19444 18534 19536 18536
rect 19444 18532 19491 18534
rect 20846 18532 20852 18596
rect 20916 18594 20922 18596
rect 21173 18594 21239 18597
rect 21544 18594 21604 18670
rect 23105 18667 23171 18670
rect 23841 18730 23907 18733
rect 27061 18730 27127 18733
rect 23841 18728 27127 18730
rect 23841 18672 23846 18728
rect 23902 18672 27066 18728
rect 27122 18672 27127 18728
rect 23841 18670 27127 18672
rect 23841 18667 23907 18670
rect 27061 18667 27127 18670
rect 27245 18730 27311 18733
rect 34094 18730 34100 18732
rect 27245 18728 34100 18730
rect 27245 18672 27250 18728
rect 27306 18672 34100 18728
rect 27245 18670 34100 18672
rect 27245 18667 27311 18670
rect 34094 18668 34100 18670
rect 34164 18668 34170 18732
rect 34421 18730 34487 18733
rect 42793 18730 42859 18733
rect 34421 18728 42859 18730
rect 34421 18672 34426 18728
rect 34482 18672 42798 18728
rect 42854 18672 42859 18728
rect 34421 18670 42859 18672
rect 34421 18667 34487 18670
rect 42793 18667 42859 18670
rect 20916 18592 21604 18594
rect 20916 18536 21178 18592
rect 21234 18536 21604 18592
rect 20916 18534 21604 18536
rect 23013 18594 23079 18597
rect 36169 18594 36235 18597
rect 23013 18592 36235 18594
rect 23013 18536 23018 18592
rect 23074 18536 36174 18592
rect 36230 18536 36235 18592
rect 23013 18534 36235 18536
rect 20916 18532 20922 18534
rect 19425 18531 19491 18532
rect 21173 18531 21239 18534
rect 23013 18531 23079 18534
rect 36169 18531 36235 18534
rect 37457 18594 37523 18597
rect 38101 18594 38167 18597
rect 37457 18592 38167 18594
rect 37457 18536 37462 18592
rect 37518 18536 38106 18592
rect 38162 18536 38167 18592
rect 37457 18534 38167 18536
rect 37457 18531 37523 18534
rect 38101 18531 38167 18534
rect 40125 18594 40191 18597
rect 41597 18594 41663 18597
rect 40125 18592 41663 18594
rect 40125 18536 40130 18592
rect 40186 18536 41602 18592
rect 41658 18536 41663 18592
rect 40125 18534 41663 18536
rect 40125 18531 40191 18534
rect 41597 18531 41663 18534
rect 43253 18594 43319 18597
rect 45645 18594 45711 18597
rect 48405 18594 48471 18597
rect 43253 18592 48471 18594
rect 43253 18536 43258 18592
rect 43314 18536 45650 18592
rect 45706 18536 48410 18592
rect 48466 18536 48471 18592
rect 43253 18534 48471 18536
rect 43253 18531 43319 18534
rect 45645 18531 45711 18534
rect 48405 18531 48471 18534
rect 58157 18594 58223 18597
rect 59200 18594 60000 18624
rect 58157 18592 60000 18594
rect 58157 18536 58162 18592
rect 58218 18536 60000 18592
rect 58157 18534 60000 18536
rect 58157 18531 58223 18534
rect 20208 18528 20528 18529
rect 20208 18464 20216 18528
rect 20280 18464 20296 18528
rect 20360 18464 20376 18528
rect 20440 18464 20456 18528
rect 20520 18464 20528 18528
rect 20208 18463 20528 18464
rect 39472 18528 39792 18529
rect 39472 18464 39480 18528
rect 39544 18464 39560 18528
rect 39624 18464 39640 18528
rect 39704 18464 39720 18528
rect 39784 18464 39792 18528
rect 59200 18504 60000 18534
rect 39472 18463 39792 18464
rect 15009 18458 15075 18461
rect 19333 18458 19399 18461
rect 15009 18456 19399 18458
rect 15009 18400 15014 18456
rect 15070 18400 19338 18456
rect 19394 18400 19399 18456
rect 15009 18398 19399 18400
rect 15009 18395 15075 18398
rect 19333 18395 19399 18398
rect 22369 18458 22435 18461
rect 34697 18460 34763 18461
rect 32622 18458 32628 18460
rect 22369 18456 32628 18458
rect 22369 18400 22374 18456
rect 22430 18400 32628 18456
rect 22369 18398 32628 18400
rect 22369 18395 22435 18398
rect 32622 18396 32628 18398
rect 32692 18396 32698 18460
rect 34646 18396 34652 18460
rect 34716 18458 34763 18460
rect 35065 18458 35131 18461
rect 38469 18458 38535 18461
rect 34716 18456 34808 18458
rect 34758 18400 34808 18456
rect 34716 18398 34808 18400
rect 35065 18456 38535 18458
rect 35065 18400 35070 18456
rect 35126 18400 38474 18456
rect 38530 18400 38535 18456
rect 35065 18398 38535 18400
rect 34716 18396 34763 18398
rect 34697 18395 34763 18396
rect 35065 18395 35131 18398
rect 38469 18395 38535 18398
rect 40401 18458 40467 18461
rect 41321 18458 41387 18461
rect 43989 18458 44055 18461
rect 46105 18458 46171 18461
rect 40401 18456 46171 18458
rect 40401 18400 40406 18456
rect 40462 18400 41326 18456
rect 41382 18400 43994 18456
rect 44050 18400 46110 18456
rect 46166 18400 46171 18456
rect 40401 18398 46171 18400
rect 40401 18395 40467 18398
rect 41321 18395 41387 18398
rect 43989 18395 44055 18398
rect 46105 18395 46171 18398
rect 16573 18322 16639 18325
rect 23657 18322 23723 18325
rect 16573 18320 23723 18322
rect 16573 18264 16578 18320
rect 16634 18264 23662 18320
rect 23718 18264 23723 18320
rect 16573 18262 23723 18264
rect 16573 18259 16639 18262
rect 23657 18259 23723 18262
rect 24945 18322 25011 18325
rect 33174 18322 33180 18324
rect 24945 18320 33180 18322
rect 24945 18264 24950 18320
rect 25006 18264 33180 18320
rect 24945 18262 33180 18264
rect 24945 18259 25011 18262
rect 33174 18260 33180 18262
rect 33244 18260 33250 18324
rect 34329 18322 34395 18325
rect 39297 18322 39363 18325
rect 34329 18320 39363 18322
rect 34329 18264 34334 18320
rect 34390 18264 39302 18320
rect 39358 18264 39363 18320
rect 34329 18262 39363 18264
rect 34329 18259 34395 18262
rect 39297 18259 39363 18262
rect 41505 18322 41571 18325
rect 42057 18322 42123 18325
rect 48313 18322 48379 18325
rect 41505 18320 48379 18322
rect 41505 18264 41510 18320
rect 41566 18264 42062 18320
rect 42118 18264 48318 18320
rect 48374 18264 48379 18320
rect 41505 18262 48379 18264
rect 41505 18259 41571 18262
rect 42057 18259 42123 18262
rect 48313 18259 48379 18262
rect 16757 18186 16823 18189
rect 25037 18186 25103 18189
rect 16757 18184 25103 18186
rect 16757 18128 16762 18184
rect 16818 18128 25042 18184
rect 25098 18128 25103 18184
rect 16757 18126 25103 18128
rect 16757 18123 16823 18126
rect 25037 18123 25103 18126
rect 28257 18186 28323 18189
rect 33869 18186 33935 18189
rect 28257 18184 33935 18186
rect 28257 18128 28262 18184
rect 28318 18128 33874 18184
rect 33930 18128 33935 18184
rect 28257 18126 33935 18128
rect 28257 18123 28323 18126
rect 33869 18123 33935 18126
rect 34329 18186 34395 18189
rect 35566 18186 35572 18188
rect 34329 18184 35572 18186
rect 34329 18128 34334 18184
rect 34390 18128 35572 18184
rect 34329 18126 35572 18128
rect 34329 18123 34395 18126
rect 35566 18124 35572 18126
rect 35636 18124 35642 18188
rect 36721 18186 36787 18189
rect 39297 18186 39363 18189
rect 36721 18184 39363 18186
rect 36721 18128 36726 18184
rect 36782 18128 39302 18184
rect 39358 18128 39363 18184
rect 36721 18126 39363 18128
rect 36721 18123 36787 18126
rect 39297 18123 39363 18126
rect 40953 18186 41019 18189
rect 43253 18186 43319 18189
rect 40953 18184 43319 18186
rect 40953 18128 40958 18184
rect 41014 18128 43258 18184
rect 43314 18128 43319 18184
rect 40953 18126 43319 18128
rect 40953 18123 41019 18126
rect 43253 18123 43319 18126
rect 0 18050 800 18080
rect 1485 18050 1551 18053
rect 0 18048 1551 18050
rect 0 17992 1490 18048
rect 1546 17992 1551 18048
rect 0 17990 1551 17992
rect 0 17960 800 17990
rect 1485 17987 1551 17990
rect 15929 18050 15995 18053
rect 23381 18050 23447 18053
rect 28625 18050 28691 18053
rect 15929 18048 22202 18050
rect 15929 17992 15934 18048
rect 15990 17992 22202 18048
rect 15929 17990 22202 17992
rect 15929 17987 15995 17990
rect 10576 17984 10896 17985
rect 10576 17920 10584 17984
rect 10648 17920 10664 17984
rect 10728 17920 10744 17984
rect 10808 17920 10824 17984
rect 10888 17920 10896 17984
rect 10576 17919 10896 17920
rect 17309 17914 17375 17917
rect 17534 17914 17540 17916
rect 17309 17912 17540 17914
rect 17309 17856 17314 17912
rect 17370 17856 17540 17912
rect 17309 17854 17540 17856
rect 17309 17851 17375 17854
rect 17534 17852 17540 17854
rect 17604 17852 17610 17916
rect 20713 17914 20779 17917
rect 21950 17914 21956 17916
rect 20713 17912 21956 17914
rect 20713 17856 20718 17912
rect 20774 17856 21956 17912
rect 20713 17854 21956 17856
rect 20713 17851 20779 17854
rect 21950 17852 21956 17854
rect 22020 17852 22026 17916
rect 22142 17914 22202 17990
rect 23381 18048 28691 18050
rect 23381 17992 23386 18048
rect 23442 17992 28630 18048
rect 28686 17992 28691 18048
rect 23381 17990 28691 17992
rect 23381 17987 23447 17990
rect 28625 17987 28691 17990
rect 29269 18050 29335 18053
rect 29678 18050 29684 18052
rect 29269 18048 29684 18050
rect 29269 17992 29274 18048
rect 29330 17992 29684 18048
rect 29269 17990 29684 17992
rect 29269 17987 29335 17990
rect 29678 17988 29684 17990
rect 29748 17988 29754 18052
rect 30833 18050 30899 18053
rect 34789 18050 34855 18053
rect 30833 18048 34855 18050
rect 30833 17992 30838 18048
rect 30894 17992 34794 18048
rect 34850 17992 34855 18048
rect 30833 17990 34855 17992
rect 30833 17987 30899 17990
rect 34789 17987 34855 17990
rect 37457 18050 37523 18053
rect 41413 18050 41479 18053
rect 37457 18048 41479 18050
rect 37457 17992 37462 18048
rect 37518 17992 41418 18048
rect 41474 17992 41479 18048
rect 37457 17990 41479 17992
rect 37457 17987 37523 17990
rect 41413 17987 41479 17990
rect 41689 18050 41755 18053
rect 42425 18050 42491 18053
rect 41689 18048 42491 18050
rect 41689 17992 41694 18048
rect 41750 17992 42430 18048
rect 42486 17992 42491 18048
rect 41689 17990 42491 17992
rect 41689 17987 41755 17990
rect 42425 17987 42491 17990
rect 29840 17984 30160 17985
rect 29840 17920 29848 17984
rect 29912 17920 29928 17984
rect 29992 17920 30008 17984
rect 30072 17920 30088 17984
rect 30152 17920 30160 17984
rect 29840 17919 30160 17920
rect 49104 17984 49424 17985
rect 49104 17920 49112 17984
rect 49176 17920 49192 17984
rect 49256 17920 49272 17984
rect 49336 17920 49352 17984
rect 49416 17920 49424 17984
rect 49104 17919 49424 17920
rect 24485 17914 24551 17917
rect 22142 17912 24551 17914
rect 22142 17856 24490 17912
rect 24546 17856 24551 17912
rect 22142 17854 24551 17856
rect 24485 17851 24551 17854
rect 24669 17916 24735 17917
rect 24669 17912 24716 17916
rect 24780 17914 24786 17916
rect 42701 17914 42767 17917
rect 24669 17856 24674 17912
rect 24669 17852 24716 17856
rect 24780 17854 24826 17914
rect 31710 17912 42767 17914
rect 31710 17856 42706 17912
rect 42762 17856 42767 17912
rect 31710 17854 42767 17856
rect 24780 17852 24786 17854
rect 24669 17851 24735 17852
rect 14089 17778 14155 17781
rect 19149 17778 19215 17781
rect 14089 17776 19215 17778
rect 14089 17720 14094 17776
rect 14150 17720 19154 17776
rect 19210 17720 19215 17776
rect 14089 17718 19215 17720
rect 14089 17715 14155 17718
rect 19149 17715 19215 17718
rect 19885 17778 19951 17781
rect 21214 17778 21220 17780
rect 19885 17776 21220 17778
rect 19885 17720 19890 17776
rect 19946 17720 21220 17776
rect 19885 17718 21220 17720
rect 19885 17715 19951 17718
rect 21214 17716 21220 17718
rect 21284 17778 21290 17780
rect 21357 17778 21423 17781
rect 21284 17776 21423 17778
rect 21284 17720 21362 17776
rect 21418 17720 21423 17776
rect 21284 17718 21423 17720
rect 21284 17716 21290 17718
rect 21357 17715 21423 17718
rect 22001 17778 22067 17781
rect 25405 17778 25471 17781
rect 22001 17776 25471 17778
rect 22001 17720 22006 17776
rect 22062 17720 25410 17776
rect 25466 17720 25471 17776
rect 22001 17718 25471 17720
rect 22001 17715 22067 17718
rect 25405 17715 25471 17718
rect 28717 17778 28783 17781
rect 31710 17778 31770 17854
rect 42701 17851 42767 17854
rect 45093 17916 45159 17917
rect 45093 17912 45140 17916
rect 45204 17914 45210 17916
rect 45093 17856 45098 17912
rect 45093 17852 45140 17856
rect 45204 17854 45250 17914
rect 45204 17852 45210 17854
rect 45093 17851 45159 17852
rect 28717 17776 31770 17778
rect 28717 17720 28722 17776
rect 28778 17720 31770 17776
rect 28717 17718 31770 17720
rect 32857 17778 32923 17781
rect 43069 17778 43135 17781
rect 32857 17776 43135 17778
rect 32857 17720 32862 17776
rect 32918 17720 43074 17776
rect 43130 17720 43135 17776
rect 32857 17718 43135 17720
rect 28717 17715 28783 17718
rect 32857 17715 32923 17718
rect 43069 17715 43135 17718
rect 16297 17642 16363 17645
rect 18086 17642 18092 17644
rect 16297 17640 18092 17642
rect 16297 17584 16302 17640
rect 16358 17584 18092 17640
rect 16297 17582 18092 17584
rect 16297 17579 16363 17582
rect 18086 17580 18092 17582
rect 18156 17580 18162 17644
rect 18597 17642 18663 17645
rect 32489 17642 32555 17645
rect 18597 17640 32555 17642
rect 18597 17584 18602 17640
rect 18658 17584 32494 17640
rect 32550 17584 32555 17640
rect 18597 17582 32555 17584
rect 18597 17579 18663 17582
rect 32489 17579 32555 17582
rect 32765 17642 32831 17645
rect 36261 17642 36327 17645
rect 32765 17640 36327 17642
rect 32765 17584 32770 17640
rect 32826 17584 36266 17640
rect 36322 17584 36327 17640
rect 32765 17582 36327 17584
rect 32765 17579 32831 17582
rect 36261 17579 36327 17582
rect 36813 17642 36879 17645
rect 41505 17642 41571 17645
rect 36813 17640 41571 17642
rect 36813 17584 36818 17640
rect 36874 17584 41510 17640
rect 41566 17584 41571 17640
rect 36813 17582 41571 17584
rect 36813 17579 36879 17582
rect 41505 17579 41571 17582
rect 41781 17642 41847 17645
rect 46013 17642 46079 17645
rect 41781 17640 46079 17642
rect 41781 17584 41786 17640
rect 41842 17584 46018 17640
rect 46074 17584 46079 17640
rect 41781 17582 46079 17584
rect 41781 17579 41847 17582
rect 46013 17579 46079 17582
rect 15653 17506 15719 17509
rect 18413 17506 18479 17509
rect 15653 17504 18479 17506
rect 15653 17448 15658 17504
rect 15714 17448 18418 17504
rect 18474 17448 18479 17504
rect 15653 17446 18479 17448
rect 15653 17443 15719 17446
rect 18413 17443 18479 17446
rect 19793 17506 19859 17509
rect 20069 17506 20135 17509
rect 19793 17504 20135 17506
rect 19793 17448 19798 17504
rect 19854 17448 20074 17504
rect 20130 17448 20135 17504
rect 19793 17446 20135 17448
rect 19793 17443 19859 17446
rect 20069 17443 20135 17446
rect 20713 17506 20779 17509
rect 22461 17506 22527 17509
rect 20713 17504 22527 17506
rect 20713 17448 20718 17504
rect 20774 17448 22466 17504
rect 22522 17448 22527 17504
rect 20713 17446 22527 17448
rect 20713 17443 20779 17446
rect 22461 17443 22527 17446
rect 24485 17506 24551 17509
rect 30465 17506 30531 17509
rect 24485 17504 30531 17506
rect 24485 17448 24490 17504
rect 24546 17448 30470 17504
rect 30526 17448 30531 17504
rect 24485 17446 30531 17448
rect 24485 17443 24551 17446
rect 30465 17443 30531 17446
rect 30649 17506 30715 17509
rect 31845 17506 31911 17509
rect 30649 17504 31911 17506
rect 30649 17448 30654 17504
rect 30710 17448 31850 17504
rect 31906 17448 31911 17504
rect 30649 17446 31911 17448
rect 30649 17443 30715 17446
rect 31845 17443 31911 17446
rect 39941 17506 40007 17509
rect 47117 17506 47183 17509
rect 48129 17506 48195 17509
rect 39941 17504 48195 17506
rect 39941 17448 39946 17504
rect 40002 17448 47122 17504
rect 47178 17448 48134 17504
rect 48190 17448 48195 17504
rect 39941 17446 48195 17448
rect 39941 17443 40007 17446
rect 47117 17443 47183 17446
rect 48129 17443 48195 17446
rect 20208 17440 20528 17441
rect 20208 17376 20216 17440
rect 20280 17376 20296 17440
rect 20360 17376 20376 17440
rect 20440 17376 20456 17440
rect 20520 17376 20528 17440
rect 20208 17375 20528 17376
rect 39472 17440 39792 17441
rect 39472 17376 39480 17440
rect 39544 17376 39560 17440
rect 39624 17376 39640 17440
rect 39704 17376 39720 17440
rect 39784 17376 39792 17440
rect 39472 17375 39792 17376
rect 13997 17370 14063 17373
rect 14733 17370 14799 17373
rect 20069 17370 20135 17373
rect 13997 17368 20135 17370
rect 13997 17312 14002 17368
rect 14058 17312 14738 17368
rect 14794 17312 20074 17368
rect 20130 17312 20135 17368
rect 13997 17310 20135 17312
rect 13997 17307 14063 17310
rect 14733 17307 14799 17310
rect 20069 17307 20135 17310
rect 21357 17370 21423 17373
rect 22277 17370 22343 17373
rect 38193 17370 38259 17373
rect 41137 17372 41203 17373
rect 41086 17370 41092 17372
rect 21357 17368 22343 17370
rect 21357 17312 21362 17368
rect 21418 17312 22282 17368
rect 22338 17312 22343 17368
rect 21357 17310 22343 17312
rect 21357 17307 21423 17310
rect 22277 17307 22343 17310
rect 25822 17368 38259 17370
rect 25822 17312 38198 17368
rect 38254 17312 38259 17368
rect 25822 17310 38259 17312
rect 41046 17310 41092 17370
rect 41156 17368 41203 17372
rect 41198 17312 41203 17368
rect 16389 17234 16455 17237
rect 20846 17234 20852 17236
rect 16389 17232 20852 17234
rect 16389 17176 16394 17232
rect 16450 17176 20852 17232
rect 16389 17174 20852 17176
rect 16389 17171 16455 17174
rect 20846 17172 20852 17174
rect 20916 17172 20922 17236
rect 24945 17234 25011 17237
rect 21774 17232 25011 17234
rect 21774 17176 24950 17232
rect 25006 17176 25011 17232
rect 21774 17174 25011 17176
rect 16113 17098 16179 17101
rect 21774 17098 21834 17174
rect 24945 17171 25011 17174
rect 16113 17096 21834 17098
rect 16113 17040 16118 17096
rect 16174 17040 21834 17096
rect 16113 17038 21834 17040
rect 21909 17098 21975 17101
rect 25822 17098 25882 17310
rect 38193 17307 38259 17310
rect 41086 17308 41092 17310
rect 41156 17308 41203 17312
rect 41137 17307 41203 17308
rect 42241 17370 42307 17373
rect 46054 17370 46060 17372
rect 42241 17368 46060 17370
rect 42241 17312 42246 17368
rect 42302 17312 46060 17368
rect 42241 17310 46060 17312
rect 42241 17307 42307 17310
rect 46054 17308 46060 17310
rect 46124 17308 46130 17372
rect 26049 17234 26115 17237
rect 36854 17234 36860 17236
rect 26049 17232 36860 17234
rect 26049 17176 26054 17232
rect 26110 17176 36860 17232
rect 26049 17174 36860 17176
rect 26049 17171 26115 17174
rect 36854 17172 36860 17174
rect 36924 17172 36930 17236
rect 37222 17172 37228 17236
rect 37292 17234 37298 17236
rect 37774 17234 37780 17236
rect 37292 17174 37780 17234
rect 37292 17172 37298 17174
rect 37774 17172 37780 17174
rect 37844 17172 37850 17236
rect 38101 17234 38167 17237
rect 41321 17234 41387 17237
rect 50153 17234 50219 17237
rect 38101 17232 50219 17234
rect 38101 17176 38106 17232
rect 38162 17176 41326 17232
rect 41382 17176 50158 17232
rect 50214 17176 50219 17232
rect 38101 17174 50219 17176
rect 38101 17171 38167 17174
rect 41321 17171 41387 17174
rect 50153 17171 50219 17174
rect 31385 17098 31451 17101
rect 21909 17096 25882 17098
rect 21909 17040 21914 17096
rect 21970 17040 25882 17096
rect 21909 17038 25882 17040
rect 26926 17096 31451 17098
rect 26926 17040 31390 17096
rect 31446 17040 31451 17096
rect 26926 17038 31451 17040
rect 16113 17035 16179 17038
rect 21909 17035 21975 17038
rect 18689 16962 18755 16965
rect 26926 16962 26986 17038
rect 31385 17035 31451 17038
rect 31845 17098 31911 17101
rect 34697 17098 34763 17101
rect 31845 17096 34763 17098
rect 31845 17040 31850 17096
rect 31906 17040 34702 17096
rect 34758 17040 34763 17096
rect 31845 17038 34763 17040
rect 31845 17035 31911 17038
rect 34697 17035 34763 17038
rect 35709 17098 35775 17101
rect 39113 17098 39179 17101
rect 35709 17096 39179 17098
rect 35709 17040 35714 17096
rect 35770 17040 39118 17096
rect 39174 17040 39179 17096
rect 35709 17038 39179 17040
rect 35709 17035 35775 17038
rect 39113 17035 39179 17038
rect 41689 17098 41755 17101
rect 42793 17098 42859 17101
rect 41689 17096 42859 17098
rect 41689 17040 41694 17096
rect 41750 17040 42798 17096
rect 42854 17040 42859 17096
rect 41689 17038 42859 17040
rect 41689 17035 41755 17038
rect 42793 17035 42859 17038
rect 42977 17098 43043 17101
rect 45369 17098 45435 17101
rect 42977 17096 45435 17098
rect 42977 17040 42982 17096
rect 43038 17040 45374 17096
rect 45430 17040 45435 17096
rect 42977 17038 45435 17040
rect 42977 17035 43043 17038
rect 45369 17035 45435 17038
rect 18689 16960 26986 16962
rect 18689 16904 18694 16960
rect 18750 16904 26986 16960
rect 18689 16902 26986 16904
rect 18689 16899 18755 16902
rect 32438 16900 32444 16964
rect 32508 16962 32514 16964
rect 34145 16962 34211 16965
rect 32508 16960 34211 16962
rect 32508 16904 34150 16960
rect 34206 16904 34211 16960
rect 32508 16902 34211 16904
rect 32508 16900 32514 16902
rect 34145 16899 34211 16902
rect 37038 16900 37044 16964
rect 37108 16962 37114 16964
rect 38285 16962 38351 16965
rect 42885 16962 42951 16965
rect 37108 16902 38210 16962
rect 37108 16900 37114 16902
rect 10576 16896 10896 16897
rect 10576 16832 10584 16896
rect 10648 16832 10664 16896
rect 10728 16832 10744 16896
rect 10808 16832 10824 16896
rect 10888 16832 10896 16896
rect 10576 16831 10896 16832
rect 29840 16896 30160 16897
rect 29840 16832 29848 16896
rect 29912 16832 29928 16896
rect 29992 16832 30008 16896
rect 30072 16832 30088 16896
rect 30152 16832 30160 16896
rect 29840 16831 30160 16832
rect 15377 16826 15443 16829
rect 18781 16826 18847 16829
rect 15377 16824 18847 16826
rect 15377 16768 15382 16824
rect 15438 16768 18786 16824
rect 18842 16768 18847 16824
rect 15377 16766 18847 16768
rect 15377 16763 15443 16766
rect 18781 16763 18847 16766
rect 19149 16826 19215 16829
rect 27337 16826 27403 16829
rect 30649 16826 30715 16829
rect 19149 16824 27403 16826
rect 19149 16768 19154 16824
rect 19210 16768 27342 16824
rect 27398 16768 27403 16824
rect 19149 16766 27403 16768
rect 19149 16763 19215 16766
rect 27337 16763 27403 16766
rect 30238 16824 30715 16826
rect 30238 16768 30654 16824
rect 30710 16768 30715 16824
rect 30238 16766 30715 16768
rect 15285 16692 15351 16693
rect 17493 16692 17559 16693
rect 15285 16688 15332 16692
rect 15396 16690 15402 16692
rect 15285 16632 15290 16688
rect 15285 16628 15332 16632
rect 15396 16630 15442 16690
rect 17493 16688 17540 16692
rect 17604 16690 17610 16692
rect 18689 16690 18755 16693
rect 18822 16690 18828 16692
rect 17493 16632 17498 16688
rect 15396 16628 15402 16630
rect 17493 16628 17540 16632
rect 17604 16630 17650 16690
rect 18689 16688 18828 16690
rect 18689 16632 18694 16688
rect 18750 16632 18828 16688
rect 18689 16630 18828 16632
rect 17604 16628 17610 16630
rect 15285 16627 15351 16628
rect 17493 16627 17559 16628
rect 18689 16627 18755 16630
rect 18822 16628 18828 16630
rect 18892 16628 18898 16692
rect 19609 16690 19675 16693
rect 19742 16690 19748 16692
rect 19609 16688 19748 16690
rect 19609 16632 19614 16688
rect 19670 16632 19748 16688
rect 19609 16630 19748 16632
rect 19609 16627 19675 16630
rect 19742 16628 19748 16630
rect 19812 16628 19818 16692
rect 20069 16690 20135 16693
rect 21725 16690 21791 16693
rect 26366 16690 26372 16692
rect 20069 16688 21791 16690
rect 20069 16632 20074 16688
rect 20130 16632 21730 16688
rect 21786 16632 21791 16688
rect 20069 16630 21791 16632
rect 20069 16627 20135 16630
rect 21725 16627 21791 16630
rect 22326 16630 26372 16690
rect 0 16554 800 16584
rect 1485 16554 1551 16557
rect 0 16552 1551 16554
rect 0 16496 1490 16552
rect 1546 16496 1551 16552
rect 0 16494 1551 16496
rect 0 16464 800 16494
rect 1485 16491 1551 16494
rect 15837 16554 15903 16557
rect 18454 16554 18460 16556
rect 15837 16552 18460 16554
rect 15837 16496 15842 16552
rect 15898 16496 18460 16552
rect 15837 16494 18460 16496
rect 15837 16491 15903 16494
rect 18454 16492 18460 16494
rect 18524 16492 18530 16556
rect 18689 16554 18755 16557
rect 19006 16554 19012 16556
rect 18689 16552 19012 16554
rect 18689 16496 18694 16552
rect 18750 16496 19012 16552
rect 18689 16494 19012 16496
rect 18689 16491 18755 16494
rect 19006 16492 19012 16494
rect 19076 16492 19082 16556
rect 19926 16492 19932 16556
rect 19996 16554 20002 16556
rect 20069 16554 20135 16557
rect 19996 16552 20135 16554
rect 19996 16496 20074 16552
rect 20130 16496 20135 16552
rect 19996 16494 20135 16496
rect 19996 16492 20002 16494
rect 20069 16491 20135 16494
rect 20529 16554 20595 16557
rect 22326 16554 22386 16630
rect 26366 16628 26372 16630
rect 26436 16628 26442 16692
rect 28993 16690 29059 16693
rect 30238 16690 30298 16766
rect 30649 16763 30715 16766
rect 30925 16826 30991 16829
rect 31201 16826 31267 16829
rect 30925 16824 31267 16826
rect 30925 16768 30930 16824
rect 30986 16768 31206 16824
rect 31262 16768 31267 16824
rect 30925 16766 31267 16768
rect 30925 16763 30991 16766
rect 31201 16763 31267 16766
rect 31886 16764 31892 16828
rect 31956 16826 31962 16828
rect 34145 16826 34211 16829
rect 34329 16826 34395 16829
rect 31956 16824 34395 16826
rect 31956 16768 34150 16824
rect 34206 16768 34334 16824
rect 34390 16768 34395 16824
rect 31956 16766 34395 16768
rect 31956 16764 31962 16766
rect 34145 16763 34211 16766
rect 34329 16763 34395 16766
rect 34462 16764 34468 16828
rect 34532 16826 34538 16828
rect 38009 16826 38075 16829
rect 34532 16824 38075 16826
rect 34532 16768 38014 16824
rect 38070 16768 38075 16824
rect 34532 16766 38075 16768
rect 38150 16826 38210 16902
rect 38285 16960 42951 16962
rect 38285 16904 38290 16960
rect 38346 16904 42890 16960
rect 42946 16904 42951 16960
rect 38285 16902 42951 16904
rect 38285 16899 38351 16902
rect 42885 16899 42951 16902
rect 49104 16896 49424 16897
rect 49104 16832 49112 16896
rect 49176 16832 49192 16896
rect 49256 16832 49272 16896
rect 49336 16832 49352 16896
rect 49416 16832 49424 16896
rect 49104 16831 49424 16832
rect 44173 16826 44239 16829
rect 38150 16824 44239 16826
rect 38150 16768 44178 16824
rect 44234 16768 44239 16824
rect 38150 16766 44239 16768
rect 34532 16764 34538 16766
rect 38009 16763 38075 16766
rect 44173 16763 44239 16766
rect 45185 16826 45251 16829
rect 47025 16826 47091 16829
rect 45185 16824 47091 16826
rect 45185 16768 45190 16824
rect 45246 16768 47030 16824
rect 47086 16768 47091 16824
rect 45185 16766 47091 16768
rect 45185 16763 45251 16766
rect 47025 16763 47091 16766
rect 58157 16826 58223 16829
rect 59200 16826 60000 16856
rect 58157 16824 60000 16826
rect 58157 16768 58162 16824
rect 58218 16768 60000 16824
rect 58157 16766 60000 16768
rect 58157 16763 58223 16766
rect 59200 16736 60000 16766
rect 28993 16688 30298 16690
rect 28993 16632 28998 16688
rect 29054 16632 30298 16688
rect 28993 16630 30298 16632
rect 30465 16690 30531 16693
rect 35801 16690 35867 16693
rect 30465 16688 35867 16690
rect 30465 16632 30470 16688
rect 30526 16632 35806 16688
rect 35862 16632 35867 16688
rect 30465 16630 35867 16632
rect 28993 16627 29059 16630
rect 30465 16627 30531 16630
rect 35801 16627 35867 16630
rect 37365 16690 37431 16693
rect 42057 16690 42123 16693
rect 42190 16690 42196 16692
rect 37365 16688 41936 16690
rect 37365 16632 37370 16688
rect 37426 16632 41936 16688
rect 37365 16630 41936 16632
rect 37365 16627 37431 16630
rect 20529 16552 22386 16554
rect 20529 16496 20534 16552
rect 20590 16496 22386 16552
rect 20529 16494 22386 16496
rect 22461 16554 22527 16557
rect 23749 16554 23815 16557
rect 22461 16552 23815 16554
rect 22461 16496 22466 16552
rect 22522 16496 23754 16552
rect 23810 16496 23815 16552
rect 22461 16494 23815 16496
rect 20529 16491 20595 16494
rect 22461 16491 22527 16494
rect 23749 16491 23815 16494
rect 24025 16554 24091 16557
rect 25446 16554 25452 16556
rect 24025 16552 25452 16554
rect 24025 16496 24030 16552
rect 24086 16496 25452 16552
rect 24025 16494 25452 16496
rect 24025 16491 24091 16494
rect 25446 16492 25452 16494
rect 25516 16492 25522 16556
rect 26550 16492 26556 16556
rect 26620 16554 26626 16556
rect 26693 16554 26759 16557
rect 26620 16552 26759 16554
rect 26620 16496 26698 16552
rect 26754 16496 26759 16552
rect 26620 16494 26759 16496
rect 26620 16492 26626 16494
rect 26693 16491 26759 16494
rect 28533 16554 28599 16557
rect 37273 16554 37339 16557
rect 41876 16554 41936 16630
rect 42057 16688 42196 16690
rect 42057 16632 42062 16688
rect 42118 16632 42196 16688
rect 42057 16630 42196 16632
rect 42057 16627 42123 16630
rect 42190 16628 42196 16630
rect 42260 16628 42266 16692
rect 45001 16690 45067 16693
rect 42382 16688 45067 16690
rect 42382 16632 45006 16688
rect 45062 16632 45067 16688
rect 42382 16630 45067 16632
rect 42382 16554 42442 16630
rect 45001 16627 45067 16630
rect 46473 16690 46539 16693
rect 46606 16690 46612 16692
rect 46473 16688 46612 16690
rect 46473 16632 46478 16688
rect 46534 16632 46612 16688
rect 46473 16630 46612 16632
rect 46473 16627 46539 16630
rect 46606 16628 46612 16630
rect 46676 16628 46682 16692
rect 28533 16552 36554 16554
rect 28533 16496 28538 16552
rect 28594 16496 36554 16552
rect 28533 16494 36554 16496
rect 28533 16491 28599 16494
rect 14917 16418 14983 16421
rect 19701 16418 19767 16421
rect 20846 16418 20852 16420
rect 14917 16416 19767 16418
rect 14917 16360 14922 16416
rect 14978 16360 19706 16416
rect 19762 16360 19767 16416
rect 14917 16358 19767 16360
rect 14917 16355 14983 16358
rect 19701 16355 19767 16358
rect 20670 16358 20852 16418
rect 20208 16352 20528 16353
rect 20208 16288 20216 16352
rect 20280 16288 20296 16352
rect 20360 16288 20376 16352
rect 20440 16288 20456 16352
rect 20520 16288 20528 16352
rect 20208 16287 20528 16288
rect 15561 16146 15627 16149
rect 19701 16146 19767 16149
rect 15561 16144 19767 16146
rect 15561 16088 15566 16144
rect 15622 16088 19706 16144
rect 19762 16088 19767 16144
rect 15561 16086 19767 16088
rect 15561 16083 15627 16086
rect 19701 16083 19767 16086
rect 20529 16146 20595 16149
rect 20670 16146 20730 16358
rect 20846 16356 20852 16358
rect 20916 16356 20922 16420
rect 21173 16418 21239 16421
rect 21173 16416 25100 16418
rect 21173 16360 21178 16416
rect 21234 16360 25100 16416
rect 21173 16358 25100 16360
rect 21173 16355 21239 16358
rect 21176 16282 21236 16355
rect 20529 16144 20730 16146
rect 20529 16088 20534 16144
rect 20590 16088 20730 16144
rect 20529 16086 20730 16088
rect 20900 16222 21236 16282
rect 21633 16282 21699 16285
rect 22134 16282 22140 16284
rect 21633 16280 22140 16282
rect 21633 16224 21638 16280
rect 21694 16224 22140 16280
rect 21633 16222 22140 16224
rect 20529 16083 20595 16086
rect 15653 16010 15719 16013
rect 20900 16010 20960 16222
rect 21633 16219 21699 16222
rect 22134 16220 22140 16222
rect 22204 16220 22210 16284
rect 21081 16148 21147 16149
rect 21030 16084 21036 16148
rect 21100 16146 21147 16148
rect 21541 16148 21607 16149
rect 21541 16146 21588 16148
rect 21100 16144 21192 16146
rect 21142 16088 21192 16144
rect 21100 16086 21192 16088
rect 21496 16144 21588 16146
rect 21496 16088 21546 16144
rect 21496 16086 21588 16088
rect 21100 16084 21147 16086
rect 21081 16083 21147 16084
rect 21541 16084 21588 16086
rect 21652 16084 21658 16148
rect 22185 16146 22251 16149
rect 24526 16146 24532 16148
rect 22185 16144 24532 16146
rect 22185 16088 22190 16144
rect 22246 16088 24532 16144
rect 22185 16086 24532 16088
rect 21541 16083 21607 16084
rect 22185 16083 22251 16086
rect 24526 16084 24532 16086
rect 24596 16146 24602 16148
rect 24853 16146 24919 16149
rect 24596 16144 24919 16146
rect 24596 16088 24858 16144
rect 24914 16088 24919 16144
rect 24596 16086 24919 16088
rect 25040 16146 25100 16358
rect 28206 16356 28212 16420
rect 28276 16418 28282 16420
rect 29177 16418 29243 16421
rect 28276 16416 29243 16418
rect 28276 16360 29182 16416
rect 29238 16360 29243 16416
rect 28276 16358 29243 16360
rect 28276 16356 28282 16358
rect 29177 16355 29243 16358
rect 30465 16418 30531 16421
rect 31569 16418 31635 16421
rect 30465 16416 31635 16418
rect 30465 16360 30470 16416
rect 30526 16360 31574 16416
rect 31630 16360 31635 16416
rect 30465 16358 31635 16360
rect 30465 16355 30531 16358
rect 31569 16355 31635 16358
rect 33869 16418 33935 16421
rect 36118 16418 36124 16420
rect 33869 16416 36124 16418
rect 33869 16360 33874 16416
rect 33930 16360 36124 16416
rect 33869 16358 36124 16360
rect 33869 16355 33935 16358
rect 36118 16356 36124 16358
rect 36188 16356 36194 16420
rect 36494 16418 36554 16494
rect 37273 16552 41430 16554
rect 37273 16496 37278 16552
rect 37334 16496 41430 16552
rect 37273 16494 41430 16496
rect 41876 16494 42442 16554
rect 37273 16491 37339 16494
rect 37457 16418 37523 16421
rect 36494 16416 37523 16418
rect 36494 16360 37462 16416
rect 37518 16360 37523 16416
rect 36494 16358 37523 16360
rect 41370 16418 41430 16494
rect 44725 16418 44791 16421
rect 48313 16418 48379 16421
rect 41370 16416 48379 16418
rect 41370 16360 44730 16416
rect 44786 16360 48318 16416
rect 48374 16360 48379 16416
rect 41370 16358 48379 16360
rect 37457 16355 37523 16358
rect 44725 16355 44791 16358
rect 48313 16355 48379 16358
rect 39472 16352 39792 16353
rect 39472 16288 39480 16352
rect 39544 16288 39560 16352
rect 39624 16288 39640 16352
rect 39704 16288 39720 16352
rect 39784 16288 39792 16352
rect 39472 16287 39792 16288
rect 27521 16282 27587 16285
rect 38745 16282 38811 16285
rect 27521 16280 38811 16282
rect 27521 16224 27526 16280
rect 27582 16224 38750 16280
rect 38806 16224 38811 16280
rect 27521 16222 38811 16224
rect 27521 16219 27587 16222
rect 38745 16219 38811 16222
rect 38878 16220 38884 16284
rect 38948 16282 38954 16284
rect 39021 16282 39087 16285
rect 38948 16280 39087 16282
rect 38948 16224 39026 16280
rect 39082 16224 39087 16280
rect 38948 16222 39087 16224
rect 38948 16220 38954 16222
rect 39021 16219 39087 16222
rect 41965 16282 42031 16285
rect 47301 16282 47367 16285
rect 48129 16282 48195 16285
rect 41965 16280 48195 16282
rect 41965 16224 41970 16280
rect 42026 16224 47306 16280
rect 47362 16224 48134 16280
rect 48190 16224 48195 16280
rect 41965 16222 48195 16224
rect 41965 16219 42031 16222
rect 47301 16219 47367 16222
rect 48129 16219 48195 16222
rect 30966 16146 30972 16148
rect 25040 16086 30972 16146
rect 24596 16084 24602 16086
rect 24853 16083 24919 16086
rect 30966 16084 30972 16086
rect 31036 16084 31042 16148
rect 37457 16146 37523 16149
rect 49785 16146 49851 16149
rect 37457 16144 49851 16146
rect 37457 16088 37462 16144
rect 37518 16088 49790 16144
rect 49846 16088 49851 16144
rect 37457 16086 49851 16088
rect 37457 16083 37523 16086
rect 49785 16083 49851 16086
rect 23381 16010 23447 16013
rect 15653 16008 20960 16010
rect 15653 15952 15658 16008
rect 15714 15952 20960 16008
rect 15653 15950 20960 15952
rect 21038 16008 23447 16010
rect 21038 15952 23386 16008
rect 23442 15952 23447 16008
rect 21038 15950 23447 15952
rect 15653 15947 15719 15950
rect 15101 15874 15167 15877
rect 17953 15874 18019 15877
rect 20161 15874 20227 15877
rect 15101 15872 20227 15874
rect 15101 15816 15106 15872
rect 15162 15816 17958 15872
rect 18014 15816 20166 15872
rect 20222 15816 20227 15872
rect 15101 15814 20227 15816
rect 15101 15811 15167 15814
rect 17953 15811 18019 15814
rect 20161 15811 20227 15814
rect 20713 15874 20779 15877
rect 21038 15874 21098 15950
rect 23381 15947 23447 15950
rect 24209 16010 24275 16013
rect 32070 16010 32076 16012
rect 24209 16008 32076 16010
rect 24209 15952 24214 16008
rect 24270 15952 32076 16008
rect 24209 15950 32076 15952
rect 24209 15947 24275 15950
rect 32070 15948 32076 15950
rect 32140 16010 32146 16012
rect 40125 16010 40191 16013
rect 32140 16008 40418 16010
rect 32140 15952 40130 16008
rect 40186 15952 40418 16008
rect 32140 15950 40418 15952
rect 32140 15948 32146 15950
rect 40125 15947 40191 15950
rect 27153 15874 27219 15877
rect 29545 15876 29611 15877
rect 20713 15872 21098 15874
rect 20713 15816 20718 15872
rect 20774 15816 21098 15872
rect 20713 15814 21098 15816
rect 22326 15872 27219 15874
rect 22326 15816 27158 15872
rect 27214 15816 27219 15872
rect 22326 15814 27219 15816
rect 20713 15811 20779 15814
rect 10576 15808 10896 15809
rect 10576 15744 10584 15808
rect 10648 15744 10664 15808
rect 10728 15744 10744 15808
rect 10808 15744 10824 15808
rect 10888 15744 10896 15808
rect 10576 15743 10896 15744
rect 17309 15738 17375 15741
rect 22093 15738 22159 15741
rect 17309 15736 22159 15738
rect 17309 15680 17314 15736
rect 17370 15680 22098 15736
rect 22154 15680 22159 15736
rect 17309 15678 22159 15680
rect 17309 15675 17375 15678
rect 22093 15675 22159 15678
rect 20161 15602 20227 15605
rect 19290 15600 20227 15602
rect 19290 15544 20166 15600
rect 20222 15544 20227 15600
rect 19290 15542 20227 15544
rect 15193 15466 15259 15469
rect 16205 15466 16271 15469
rect 19290 15466 19350 15542
rect 20161 15539 20227 15542
rect 20897 15602 20963 15605
rect 22326 15602 22386 15814
rect 27153 15811 27219 15814
rect 29494 15812 29500 15876
rect 29564 15874 29611 15876
rect 36813 15874 36879 15877
rect 40217 15874 40283 15877
rect 29564 15872 29656 15874
rect 29606 15816 29656 15872
rect 29564 15814 29656 15816
rect 30238 15872 40283 15874
rect 30238 15816 36818 15872
rect 36874 15816 40222 15872
rect 40278 15816 40283 15872
rect 30238 15814 40283 15816
rect 40358 15874 40418 15950
rect 45553 15874 45619 15877
rect 46013 15876 46079 15877
rect 46013 15874 46060 15876
rect 40358 15872 45619 15874
rect 40358 15816 45558 15872
rect 45614 15816 45619 15872
rect 40358 15814 45619 15816
rect 45968 15872 46060 15874
rect 45968 15816 46018 15872
rect 45968 15814 46060 15816
rect 29564 15812 29611 15814
rect 29545 15811 29611 15812
rect 29840 15808 30160 15809
rect 29840 15744 29848 15808
rect 29912 15744 29928 15808
rect 29992 15744 30008 15808
rect 30072 15744 30088 15808
rect 30152 15744 30160 15808
rect 29840 15743 30160 15744
rect 22645 15738 22711 15741
rect 26601 15738 26667 15741
rect 22645 15736 26667 15738
rect 22645 15680 22650 15736
rect 22706 15680 26606 15736
rect 26662 15680 26667 15736
rect 22645 15678 26667 15680
rect 22645 15675 22711 15678
rect 26601 15675 26667 15678
rect 28809 15738 28875 15741
rect 28809 15736 29746 15738
rect 28809 15680 28814 15736
rect 28870 15680 29746 15736
rect 28809 15678 29746 15680
rect 28809 15675 28875 15678
rect 20897 15600 22386 15602
rect 20897 15544 20902 15600
rect 20958 15544 22386 15600
rect 20897 15542 22386 15544
rect 22461 15602 22527 15605
rect 23422 15602 23428 15604
rect 22461 15600 23428 15602
rect 22461 15544 22466 15600
rect 22522 15544 23428 15600
rect 22461 15542 23428 15544
rect 20897 15539 20963 15542
rect 22461 15539 22527 15542
rect 23422 15540 23428 15542
rect 23492 15540 23498 15604
rect 23565 15602 23631 15605
rect 24209 15602 24275 15605
rect 23565 15600 24275 15602
rect 23565 15544 23570 15600
rect 23626 15544 24214 15600
rect 24270 15544 24275 15600
rect 23565 15542 24275 15544
rect 23565 15539 23631 15542
rect 24209 15539 24275 15542
rect 25313 15602 25379 15605
rect 28942 15602 28948 15604
rect 25313 15600 28948 15602
rect 25313 15544 25318 15600
rect 25374 15544 28948 15600
rect 25313 15542 28948 15544
rect 25313 15539 25379 15542
rect 28942 15540 28948 15542
rect 29012 15540 29018 15604
rect 29686 15602 29746 15678
rect 30238 15602 30298 15814
rect 36813 15811 36879 15814
rect 40217 15811 40283 15814
rect 45553 15811 45619 15814
rect 46013 15812 46060 15814
rect 46124 15812 46130 15876
rect 46013 15811 46079 15812
rect 49104 15808 49424 15809
rect 49104 15744 49112 15808
rect 49176 15744 49192 15808
rect 49256 15744 49272 15808
rect 49336 15744 49352 15808
rect 49416 15744 49424 15808
rect 49104 15743 49424 15744
rect 30649 15738 30715 15741
rect 36261 15738 36327 15741
rect 40953 15738 41019 15741
rect 30649 15736 36002 15738
rect 30649 15680 30654 15736
rect 30710 15680 36002 15736
rect 30649 15678 36002 15680
rect 30649 15675 30715 15678
rect 29686 15542 30298 15602
rect 30465 15602 30531 15605
rect 35801 15602 35867 15605
rect 30465 15600 35867 15602
rect 30465 15544 30470 15600
rect 30526 15544 35806 15600
rect 35862 15544 35867 15600
rect 30465 15542 35867 15544
rect 35942 15602 36002 15678
rect 36261 15736 41019 15738
rect 36261 15680 36266 15736
rect 36322 15680 40958 15736
rect 41014 15680 41019 15736
rect 36261 15678 41019 15680
rect 36261 15675 36327 15678
rect 40953 15675 41019 15678
rect 37641 15602 37707 15605
rect 35942 15600 37707 15602
rect 35942 15544 37646 15600
rect 37702 15544 37707 15600
rect 35942 15542 37707 15544
rect 30465 15539 30531 15542
rect 35801 15539 35867 15542
rect 37641 15539 37707 15542
rect 44173 15602 44239 15605
rect 47209 15602 47275 15605
rect 44173 15600 47275 15602
rect 44173 15544 44178 15600
rect 44234 15544 47214 15600
rect 47270 15544 47275 15600
rect 44173 15542 47275 15544
rect 44173 15539 44239 15542
rect 47209 15539 47275 15542
rect 15193 15464 19350 15466
rect 15193 15408 15198 15464
rect 15254 15408 16210 15464
rect 16266 15408 19350 15464
rect 15193 15406 19350 15408
rect 20069 15466 20135 15469
rect 32489 15466 32555 15469
rect 20069 15464 32555 15466
rect 20069 15408 20074 15464
rect 20130 15408 32494 15464
rect 32550 15408 32555 15464
rect 20069 15406 32555 15408
rect 15193 15403 15259 15406
rect 16205 15403 16271 15406
rect 20069 15403 20135 15406
rect 32489 15403 32555 15406
rect 34421 15466 34487 15469
rect 36445 15466 36511 15469
rect 38745 15468 38811 15469
rect 38694 15466 38700 15468
rect 34421 15464 36511 15466
rect 34421 15408 34426 15464
rect 34482 15408 36450 15464
rect 36506 15408 36511 15464
rect 34421 15406 36511 15408
rect 38654 15406 38700 15466
rect 38764 15464 38811 15468
rect 40861 15466 40927 15469
rect 38806 15408 38811 15464
rect 34421 15403 34487 15406
rect 36445 15403 36511 15406
rect 38694 15404 38700 15406
rect 38764 15404 38811 15408
rect 38745 15403 38811 15404
rect 39300 15464 40927 15466
rect 39300 15408 40866 15464
rect 40922 15408 40927 15464
rect 39300 15406 40927 15408
rect 17309 15332 17375 15333
rect 18137 15332 18203 15333
rect 17309 15330 17356 15332
rect 17264 15328 17356 15330
rect 17264 15272 17314 15328
rect 17264 15270 17356 15272
rect 17309 15268 17356 15270
rect 17420 15268 17426 15332
rect 18086 15330 18092 15332
rect 18046 15270 18092 15330
rect 18156 15328 18203 15332
rect 20897 15330 20963 15333
rect 21541 15330 21607 15333
rect 18198 15272 18203 15328
rect 18086 15268 18092 15270
rect 18156 15268 18203 15272
rect 17309 15267 17375 15268
rect 18137 15267 18203 15268
rect 20716 15328 20963 15330
rect 20716 15272 20902 15328
rect 20958 15272 20963 15328
rect 20716 15270 20963 15272
rect 20208 15264 20528 15265
rect 20208 15200 20216 15264
rect 20280 15200 20296 15264
rect 20360 15200 20376 15264
rect 20440 15200 20456 15264
rect 20520 15200 20528 15264
rect 20208 15199 20528 15200
rect 15377 15194 15443 15197
rect 19793 15194 19859 15197
rect 15377 15192 19859 15194
rect 15377 15136 15382 15192
rect 15438 15136 19798 15192
rect 19854 15136 19859 15192
rect 15377 15134 19859 15136
rect 15377 15131 15443 15134
rect 19793 15131 19859 15134
rect 17166 14996 17172 15060
rect 17236 15058 17242 15060
rect 17309 15058 17375 15061
rect 17236 15056 17375 15058
rect 17236 15000 17314 15056
rect 17370 15000 17375 15056
rect 17236 14998 17375 15000
rect 17236 14996 17242 14998
rect 17309 14995 17375 14998
rect 19517 15058 19583 15061
rect 20716 15058 20776 15270
rect 20897 15267 20963 15270
rect 21038 15328 21607 15330
rect 21038 15272 21546 15328
rect 21602 15272 21607 15328
rect 21038 15270 21607 15272
rect 20897 15194 20963 15197
rect 21038 15194 21098 15270
rect 21541 15267 21607 15270
rect 21725 15332 21791 15333
rect 21725 15328 21772 15332
rect 21836 15330 21842 15332
rect 21725 15272 21730 15328
rect 21725 15268 21772 15272
rect 21836 15270 21882 15330
rect 21836 15268 21842 15270
rect 22134 15268 22140 15332
rect 22204 15330 22210 15332
rect 22737 15330 22803 15333
rect 24761 15330 24827 15333
rect 22204 15328 22803 15330
rect 22204 15272 22742 15328
rect 22798 15272 22803 15328
rect 22204 15270 22803 15272
rect 22204 15268 22210 15270
rect 21725 15267 21791 15268
rect 22737 15267 22803 15270
rect 22878 15328 24827 15330
rect 22878 15272 24766 15328
rect 24822 15272 24827 15328
rect 22878 15270 24827 15272
rect 20897 15192 21098 15194
rect 20897 15136 20902 15192
rect 20958 15136 21098 15192
rect 20897 15134 21098 15136
rect 21173 15194 21239 15197
rect 22878 15194 22938 15270
rect 24761 15267 24827 15270
rect 28717 15332 28783 15333
rect 28717 15328 28764 15332
rect 28828 15330 28834 15332
rect 28717 15272 28722 15328
rect 28717 15268 28764 15272
rect 28828 15270 28874 15330
rect 28828 15268 28834 15270
rect 30598 15268 30604 15332
rect 30668 15330 30674 15332
rect 31569 15330 31635 15333
rect 30668 15328 31635 15330
rect 30668 15272 31574 15328
rect 31630 15272 31635 15328
rect 30668 15270 31635 15272
rect 30668 15268 30674 15270
rect 28717 15267 28783 15268
rect 31569 15267 31635 15270
rect 31845 15330 31911 15333
rect 38878 15330 38884 15332
rect 31845 15328 38884 15330
rect 31845 15272 31850 15328
rect 31906 15272 38884 15328
rect 31845 15270 38884 15272
rect 31845 15267 31911 15270
rect 38878 15268 38884 15270
rect 38948 15268 38954 15332
rect 21173 15192 22938 15194
rect 21173 15136 21178 15192
rect 21234 15136 22938 15192
rect 21173 15134 22938 15136
rect 23197 15194 23263 15197
rect 26325 15194 26391 15197
rect 23197 15192 26391 15194
rect 23197 15136 23202 15192
rect 23258 15136 26330 15192
rect 26386 15136 26391 15192
rect 23197 15134 26391 15136
rect 20897 15131 20963 15134
rect 21173 15131 21239 15134
rect 23197 15131 23263 15134
rect 26325 15131 26391 15134
rect 28993 15194 29059 15197
rect 34697 15194 34763 15197
rect 39300 15194 39360 15406
rect 40861 15403 40927 15406
rect 43989 15466 44055 15469
rect 44398 15466 44404 15468
rect 43989 15464 44404 15466
rect 43989 15408 43994 15464
rect 44050 15408 44404 15464
rect 43989 15406 44404 15408
rect 43989 15403 44055 15406
rect 44398 15404 44404 15406
rect 44468 15404 44474 15468
rect 42425 15330 42491 15333
rect 42558 15330 42564 15332
rect 42425 15328 42564 15330
rect 42425 15272 42430 15328
rect 42486 15272 42564 15328
rect 42425 15270 42564 15272
rect 42425 15267 42491 15270
rect 42558 15268 42564 15270
rect 42628 15268 42634 15332
rect 43989 15330 44055 15333
rect 44909 15332 44975 15333
rect 44214 15330 44220 15332
rect 43989 15328 44220 15330
rect 43989 15272 43994 15328
rect 44050 15272 44220 15328
rect 43989 15270 44220 15272
rect 43989 15267 44055 15270
rect 44214 15268 44220 15270
rect 44284 15268 44290 15332
rect 44909 15328 44956 15332
rect 45020 15330 45026 15332
rect 44909 15272 44914 15328
rect 44909 15268 44956 15272
rect 45020 15270 45066 15330
rect 45020 15268 45026 15270
rect 44909 15267 44975 15268
rect 39472 15264 39792 15265
rect 39472 15200 39480 15264
rect 39544 15200 39560 15264
rect 39624 15200 39640 15264
rect 39704 15200 39720 15264
rect 39784 15200 39792 15264
rect 39472 15199 39792 15200
rect 28993 15192 32874 15194
rect 28993 15136 28998 15192
rect 29054 15136 32874 15192
rect 28993 15134 32874 15136
rect 28993 15131 29059 15134
rect 23749 15058 23815 15061
rect 19517 15056 23815 15058
rect 19517 15000 19522 15056
rect 19578 15000 23754 15056
rect 23810 15000 23815 15056
rect 19517 14998 23815 15000
rect 19517 14995 19583 14998
rect 23749 14995 23815 14998
rect 24209 15058 24275 15061
rect 31017 15058 31083 15061
rect 24209 15056 31083 15058
rect 24209 15000 24214 15056
rect 24270 15000 31022 15056
rect 31078 15000 31083 15056
rect 24209 14998 31083 15000
rect 32814 15058 32874 15134
rect 34697 15192 39360 15194
rect 34697 15136 34702 15192
rect 34758 15136 39360 15192
rect 34697 15134 39360 15136
rect 42885 15194 42951 15197
rect 44173 15194 44239 15197
rect 42885 15192 44239 15194
rect 42885 15136 42890 15192
rect 42946 15136 44178 15192
rect 44234 15136 44239 15192
rect 42885 15134 44239 15136
rect 34697 15131 34763 15134
rect 42885 15131 42951 15134
rect 44173 15131 44239 15134
rect 35709 15058 35775 15061
rect 32814 15056 35775 15058
rect 32814 15000 35714 15056
rect 35770 15000 35775 15056
rect 32814 14998 35775 15000
rect 24209 14995 24275 14998
rect 31017 14995 31083 14998
rect 35709 14995 35775 14998
rect 36169 15058 36235 15061
rect 46933 15058 46999 15061
rect 36169 15056 46999 15058
rect 36169 15000 36174 15056
rect 36230 15000 46938 15056
rect 46994 15000 46999 15056
rect 36169 14998 46999 15000
rect 36169 14995 36235 14998
rect 46933 14995 46999 14998
rect 58157 15058 58223 15061
rect 59200 15058 60000 15088
rect 58157 15056 60000 15058
rect 58157 15000 58162 15056
rect 58218 15000 60000 15056
rect 58157 14998 60000 15000
rect 58157 14995 58223 14998
rect 59200 14968 60000 14998
rect 0 14922 800 14952
rect 1485 14922 1551 14925
rect 0 14920 1551 14922
rect 0 14864 1490 14920
rect 1546 14864 1551 14920
rect 0 14862 1551 14864
rect 0 14832 800 14862
rect 1485 14859 1551 14862
rect 19057 14922 19123 14925
rect 19558 14922 19564 14924
rect 19057 14920 19564 14922
rect 19057 14864 19062 14920
rect 19118 14864 19564 14920
rect 19057 14862 19564 14864
rect 19057 14859 19123 14862
rect 19558 14860 19564 14862
rect 19628 14860 19634 14924
rect 20069 14922 20135 14925
rect 20662 14922 20668 14924
rect 20069 14920 20668 14922
rect 20069 14864 20074 14920
rect 20130 14864 20668 14920
rect 20069 14862 20668 14864
rect 20069 14859 20135 14862
rect 20662 14860 20668 14862
rect 20732 14860 20738 14924
rect 20897 14922 20963 14925
rect 23381 14922 23447 14925
rect 23974 14922 23980 14924
rect 20897 14920 23980 14922
rect 20897 14864 20902 14920
rect 20958 14864 23386 14920
rect 23442 14864 23980 14920
rect 20897 14862 23980 14864
rect 20897 14859 20963 14862
rect 23381 14859 23447 14862
rect 23974 14860 23980 14862
rect 24044 14860 24050 14924
rect 25773 14922 25839 14925
rect 27470 14922 27476 14924
rect 25773 14920 27476 14922
rect 25773 14864 25778 14920
rect 25834 14864 27476 14920
rect 25773 14862 27476 14864
rect 25773 14859 25839 14862
rect 27470 14860 27476 14862
rect 27540 14860 27546 14924
rect 28533 14922 28599 14925
rect 39849 14922 39915 14925
rect 28533 14920 39915 14922
rect 28533 14864 28538 14920
rect 28594 14864 39854 14920
rect 39910 14864 39915 14920
rect 28533 14862 39915 14864
rect 28533 14859 28599 14862
rect 39849 14859 39915 14862
rect 40861 14922 40927 14925
rect 44265 14922 44331 14925
rect 45277 14922 45343 14925
rect 40861 14920 45343 14922
rect 40861 14864 40866 14920
rect 40922 14864 44270 14920
rect 44326 14864 45282 14920
rect 45338 14864 45343 14920
rect 40861 14862 45343 14864
rect 40861 14859 40927 14862
rect 44265 14859 44331 14862
rect 45277 14859 45343 14862
rect 17953 14786 18019 14789
rect 23105 14786 23171 14789
rect 17953 14784 23171 14786
rect 17953 14728 17958 14784
rect 18014 14728 23110 14784
rect 23166 14728 23171 14784
rect 17953 14726 23171 14728
rect 17953 14723 18019 14726
rect 23105 14723 23171 14726
rect 23381 14786 23447 14789
rect 24853 14786 24919 14789
rect 29545 14786 29611 14789
rect 23381 14784 29611 14786
rect 23381 14728 23386 14784
rect 23442 14728 24858 14784
rect 24914 14728 29550 14784
rect 29606 14728 29611 14784
rect 23381 14726 29611 14728
rect 23381 14723 23447 14726
rect 24853 14723 24919 14726
rect 29545 14723 29611 14726
rect 30230 14724 30236 14788
rect 30300 14786 30306 14788
rect 30649 14786 30715 14789
rect 30300 14784 30715 14786
rect 30300 14728 30654 14784
rect 30710 14728 30715 14784
rect 30300 14726 30715 14728
rect 30300 14724 30306 14726
rect 30649 14723 30715 14726
rect 30782 14724 30788 14788
rect 30852 14786 30858 14788
rect 36169 14786 36235 14789
rect 36302 14786 36308 14788
rect 30852 14784 36308 14786
rect 30852 14728 36174 14784
rect 36230 14728 36308 14784
rect 30852 14726 36308 14728
rect 30852 14724 30858 14726
rect 36169 14723 36235 14726
rect 36302 14724 36308 14726
rect 36372 14724 36378 14788
rect 39757 14786 39823 14789
rect 40953 14786 41019 14789
rect 39757 14784 41019 14786
rect 39757 14728 39762 14784
rect 39818 14728 40958 14784
rect 41014 14728 41019 14784
rect 39757 14726 41019 14728
rect 39757 14723 39823 14726
rect 40953 14723 41019 14726
rect 10576 14720 10896 14721
rect 10576 14656 10584 14720
rect 10648 14656 10664 14720
rect 10728 14656 10744 14720
rect 10808 14656 10824 14720
rect 10888 14656 10896 14720
rect 10576 14655 10896 14656
rect 29840 14720 30160 14721
rect 29840 14656 29848 14720
rect 29912 14656 29928 14720
rect 29992 14656 30008 14720
rect 30072 14656 30088 14720
rect 30152 14656 30160 14720
rect 29840 14655 30160 14656
rect 49104 14720 49424 14721
rect 49104 14656 49112 14720
rect 49176 14656 49192 14720
rect 49256 14656 49272 14720
rect 49336 14656 49352 14720
rect 49416 14656 49424 14720
rect 49104 14655 49424 14656
rect 17309 14650 17375 14653
rect 20897 14650 20963 14653
rect 17309 14648 20963 14650
rect 17309 14592 17314 14648
rect 17370 14592 20902 14648
rect 20958 14592 20963 14648
rect 17309 14590 20963 14592
rect 17309 14587 17375 14590
rect 20897 14587 20963 14590
rect 21081 14650 21147 14653
rect 27613 14650 27679 14653
rect 28533 14650 28599 14653
rect 36445 14652 36511 14653
rect 21081 14648 27679 14650
rect 21081 14592 21086 14648
rect 21142 14592 27618 14648
rect 27674 14592 27679 14648
rect 21081 14590 27679 14592
rect 21081 14587 21147 14590
rect 27613 14587 27679 14590
rect 27846 14648 28599 14650
rect 27846 14592 28538 14648
rect 28594 14592 28599 14648
rect 27846 14590 28599 14592
rect 19057 14514 19123 14517
rect 22185 14514 22251 14517
rect 19057 14512 22251 14514
rect 19057 14456 19062 14512
rect 19118 14456 22190 14512
rect 22246 14456 22251 14512
rect 19057 14454 22251 14456
rect 19057 14451 19123 14454
rect 22185 14451 22251 14454
rect 24209 14514 24275 14517
rect 27846 14514 27906 14590
rect 28533 14587 28599 14590
rect 33174 14588 33180 14652
rect 33244 14650 33250 14652
rect 35934 14650 35940 14652
rect 33244 14590 35940 14650
rect 33244 14588 33250 14590
rect 35934 14588 35940 14590
rect 36004 14588 36010 14652
rect 36445 14650 36492 14652
rect 36364 14648 36492 14650
rect 36556 14650 36562 14652
rect 44817 14650 44883 14653
rect 36556 14648 44883 14650
rect 36364 14592 36450 14648
rect 36556 14592 44822 14648
rect 44878 14592 44883 14648
rect 36364 14590 36492 14592
rect 36445 14588 36492 14590
rect 36556 14590 44883 14592
rect 36556 14588 36562 14590
rect 36445 14587 36511 14588
rect 44817 14587 44883 14590
rect 24209 14512 27906 14514
rect 24209 14456 24214 14512
rect 24270 14456 27906 14512
rect 24209 14454 27906 14456
rect 27981 14514 28047 14517
rect 30741 14516 30807 14517
rect 30741 14514 30788 14516
rect 27981 14512 30788 14514
rect 27981 14456 27986 14512
rect 28042 14456 30746 14512
rect 27981 14454 30788 14456
rect 24209 14451 24275 14454
rect 27981 14451 28047 14454
rect 30741 14452 30788 14454
rect 30852 14452 30858 14516
rect 34973 14512 35039 14517
rect 34973 14456 34978 14512
rect 35034 14456 35039 14512
rect 30741 14451 30807 14452
rect 34973 14451 35039 14456
rect 35433 14514 35499 14517
rect 39757 14514 39823 14517
rect 35433 14512 39823 14514
rect 35433 14456 35438 14512
rect 35494 14456 39762 14512
rect 39818 14456 39823 14512
rect 35433 14454 39823 14456
rect 35433 14451 35499 14454
rect 39757 14451 39823 14454
rect 41229 14514 41295 14517
rect 57881 14514 57947 14517
rect 41229 14512 57947 14514
rect 41229 14456 41234 14512
rect 41290 14456 57886 14512
rect 57942 14456 57947 14512
rect 41229 14454 57947 14456
rect 41229 14451 41295 14454
rect 57881 14451 57947 14454
rect 15101 14378 15167 14381
rect 21081 14378 21147 14381
rect 29637 14378 29703 14381
rect 15101 14376 21147 14378
rect 15101 14320 15106 14376
rect 15162 14320 21086 14376
rect 21142 14320 21147 14376
rect 15101 14318 21147 14320
rect 15101 14315 15167 14318
rect 21081 14315 21147 14318
rect 22050 14376 29703 14378
rect 22050 14320 29642 14376
rect 29698 14320 29703 14376
rect 22050 14318 29703 14320
rect 22050 14242 22110 14318
rect 29637 14315 29703 14318
rect 34513 14378 34579 14381
rect 34976 14378 35036 14451
rect 39757 14378 39823 14381
rect 34513 14376 39823 14378
rect 34513 14320 34518 14376
rect 34574 14320 39762 14376
rect 39818 14320 39823 14376
rect 34513 14318 39823 14320
rect 34513 14315 34579 14318
rect 38840 14245 38900 14318
rect 39757 14315 39823 14318
rect 20670 14182 22110 14242
rect 23197 14242 23263 14245
rect 27337 14242 27403 14245
rect 23197 14240 27403 14242
rect 23197 14184 23202 14240
rect 23258 14184 27342 14240
rect 27398 14184 27403 14240
rect 23197 14182 27403 14184
rect 20208 14176 20528 14177
rect 20208 14112 20216 14176
rect 20280 14112 20296 14176
rect 20360 14112 20376 14176
rect 20440 14112 20456 14176
rect 20520 14112 20528 14176
rect 20208 14111 20528 14112
rect 19333 13970 19399 13973
rect 20161 13970 20227 13973
rect 19333 13968 20227 13970
rect 19333 13912 19338 13968
rect 19394 13912 20166 13968
rect 20222 13912 20227 13968
rect 19333 13910 20227 13912
rect 19333 13907 19399 13910
rect 20161 13907 20227 13910
rect 20529 13970 20595 13973
rect 20670 13970 20730 14182
rect 23197 14179 23263 14182
rect 27337 14179 27403 14182
rect 27889 14242 27955 14245
rect 28022 14242 28028 14244
rect 27889 14240 28028 14242
rect 27889 14184 27894 14240
rect 27950 14184 28028 14240
rect 27889 14182 28028 14184
rect 27889 14179 27955 14182
rect 28022 14180 28028 14182
rect 28092 14180 28098 14244
rect 28257 14242 28323 14245
rect 28390 14242 28396 14244
rect 28257 14240 28396 14242
rect 28257 14184 28262 14240
rect 28318 14184 28396 14240
rect 28257 14182 28396 14184
rect 28257 14179 28323 14182
rect 28390 14180 28396 14182
rect 28460 14180 28466 14244
rect 35985 14242 36051 14245
rect 28628 14240 36051 14242
rect 28628 14184 35990 14240
rect 36046 14184 36051 14240
rect 28628 14182 36051 14184
rect 20897 14106 20963 14109
rect 21766 14106 21772 14108
rect 20897 14104 21772 14106
rect 20897 14048 20902 14104
rect 20958 14048 21772 14104
rect 20897 14046 21772 14048
rect 20897 14043 20963 14046
rect 21766 14044 21772 14046
rect 21836 14044 21842 14108
rect 22001 14106 22067 14109
rect 22318 14106 22324 14108
rect 22001 14104 22324 14106
rect 22001 14048 22006 14104
rect 22062 14048 22324 14104
rect 22001 14046 22324 14048
rect 22001 14043 22067 14046
rect 22318 14044 22324 14046
rect 22388 14044 22394 14108
rect 26233 14106 26299 14109
rect 23660 14104 26299 14106
rect 23660 14048 26238 14104
rect 26294 14048 26299 14104
rect 23660 14046 26299 14048
rect 20529 13968 20730 13970
rect 20529 13912 20534 13968
rect 20590 13912 20730 13968
rect 20529 13910 20730 13912
rect 20989 13970 21055 13973
rect 21398 13970 21404 13972
rect 20989 13968 21404 13970
rect 20989 13912 20994 13968
rect 21050 13912 21404 13968
rect 20989 13910 21404 13912
rect 20529 13907 20595 13910
rect 20989 13907 21055 13910
rect 21398 13908 21404 13910
rect 21468 13908 21474 13972
rect 21541 13970 21607 13973
rect 21950 13970 21956 13972
rect 21541 13968 21956 13970
rect 21541 13912 21546 13968
rect 21602 13912 21956 13968
rect 21541 13910 21956 13912
rect 21541 13907 21607 13910
rect 21950 13908 21956 13910
rect 22020 13908 22026 13972
rect 19057 13834 19123 13837
rect 20437 13834 20503 13837
rect 23660 13834 23720 14046
rect 26233 14043 26299 14046
rect 26417 14106 26483 14109
rect 28628 14106 28688 14182
rect 35985 14179 36051 14182
rect 36629 14242 36695 14245
rect 38653 14242 38719 14245
rect 36629 14240 38719 14242
rect 36629 14184 36634 14240
rect 36690 14184 38658 14240
rect 38714 14184 38719 14240
rect 36629 14182 38719 14184
rect 36629 14179 36695 14182
rect 38653 14179 38719 14182
rect 38837 14240 38903 14245
rect 38837 14184 38842 14240
rect 38898 14184 38903 14240
rect 38837 14179 38903 14184
rect 40125 14242 40191 14245
rect 40125 14240 40556 14242
rect 40125 14184 40130 14240
rect 40186 14184 40556 14240
rect 40125 14182 40556 14184
rect 40125 14179 40191 14182
rect 39472 14176 39792 14177
rect 39472 14112 39480 14176
rect 39544 14112 39560 14176
rect 39624 14112 39640 14176
rect 39704 14112 39720 14176
rect 39784 14112 39792 14176
rect 39472 14111 39792 14112
rect 26417 14104 28688 14106
rect 26417 14048 26422 14104
rect 26478 14048 28688 14104
rect 26417 14046 28688 14048
rect 31661 14106 31727 14109
rect 38469 14106 38535 14109
rect 40125 14108 40191 14109
rect 40125 14106 40172 14108
rect 31661 14104 38535 14106
rect 31661 14048 31666 14104
rect 31722 14048 38474 14104
rect 38530 14048 38535 14104
rect 31661 14046 38535 14048
rect 40080 14104 40172 14106
rect 40080 14048 40130 14104
rect 40080 14046 40172 14048
rect 26417 14043 26483 14046
rect 31661 14043 31727 14046
rect 38469 14043 38535 14046
rect 40125 14044 40172 14046
rect 40236 14044 40242 14108
rect 40125 14043 40191 14044
rect 23841 13970 23907 13973
rect 39205 13972 39271 13973
rect 34830 13970 34836 13972
rect 23841 13968 34836 13970
rect 23841 13912 23846 13968
rect 23902 13912 34836 13968
rect 23841 13910 34836 13912
rect 23841 13907 23907 13910
rect 34830 13908 34836 13910
rect 34900 13908 34906 13972
rect 39205 13970 39252 13972
rect 39160 13968 39252 13970
rect 39316 13970 39322 13972
rect 39982 13970 39988 13972
rect 39160 13912 39210 13968
rect 39160 13910 39252 13912
rect 39205 13908 39252 13910
rect 39316 13910 39988 13970
rect 39316 13908 39322 13910
rect 39982 13908 39988 13910
rect 40052 13908 40058 13972
rect 40125 13970 40191 13973
rect 40350 13970 40356 13972
rect 40125 13968 40356 13970
rect 40125 13912 40130 13968
rect 40186 13912 40356 13968
rect 40125 13910 40356 13912
rect 39205 13907 39271 13908
rect 40125 13907 40191 13910
rect 40350 13908 40356 13910
rect 40420 13908 40426 13972
rect 19057 13832 19258 13834
rect 19057 13776 19062 13832
rect 19118 13776 19258 13832
rect 19057 13774 19258 13776
rect 19057 13771 19123 13774
rect 17677 13698 17743 13701
rect 19057 13698 19123 13701
rect 17677 13696 19123 13698
rect 17677 13640 17682 13696
rect 17738 13640 19062 13696
rect 19118 13640 19123 13696
rect 17677 13638 19123 13640
rect 19198 13698 19258 13774
rect 20437 13832 23720 13834
rect 20437 13776 20442 13832
rect 20498 13776 23720 13832
rect 20437 13774 23720 13776
rect 24669 13836 24735 13837
rect 24945 13836 25011 13837
rect 24669 13832 24716 13836
rect 24780 13834 24786 13836
rect 24669 13776 24674 13832
rect 20437 13771 20503 13774
rect 24669 13772 24716 13776
rect 24780 13774 24826 13834
rect 24780 13772 24786 13774
rect 24894 13772 24900 13836
rect 24964 13834 25011 13836
rect 26233 13834 26299 13837
rect 28257 13834 28323 13837
rect 24964 13832 25056 13834
rect 25006 13776 25056 13832
rect 24964 13774 25056 13776
rect 26233 13832 28323 13834
rect 26233 13776 26238 13832
rect 26294 13776 28262 13832
rect 28318 13776 28323 13832
rect 26233 13774 28323 13776
rect 24964 13772 25011 13774
rect 24669 13771 24735 13772
rect 24945 13771 25011 13772
rect 26233 13771 26299 13774
rect 28257 13771 28323 13774
rect 28942 13772 28948 13836
rect 29012 13834 29018 13836
rect 31109 13834 31175 13837
rect 29012 13832 31175 13834
rect 29012 13776 31114 13832
rect 31170 13776 31175 13832
rect 29012 13774 31175 13776
rect 29012 13772 29018 13774
rect 31109 13771 31175 13774
rect 34697 13834 34763 13837
rect 35985 13836 36051 13837
rect 35198 13834 35204 13836
rect 34697 13832 35204 13834
rect 34697 13776 34702 13832
rect 34758 13776 35204 13832
rect 34697 13774 35204 13776
rect 34697 13771 34763 13774
rect 35198 13772 35204 13774
rect 35268 13772 35274 13836
rect 35934 13772 35940 13836
rect 36004 13834 36051 13836
rect 38653 13834 38719 13837
rect 40496 13834 40556 14182
rect 40677 13970 40743 13973
rect 42926 13970 42932 13972
rect 40677 13968 42932 13970
rect 40677 13912 40682 13968
rect 40738 13912 42932 13968
rect 40677 13910 42932 13912
rect 40677 13907 40743 13910
rect 42926 13908 42932 13910
rect 42996 13908 43002 13972
rect 41321 13834 41387 13837
rect 36004 13832 36096 13834
rect 36046 13776 36096 13832
rect 36004 13774 36096 13776
rect 38653 13832 41387 13834
rect 38653 13776 38658 13832
rect 38714 13776 41326 13832
rect 41382 13776 41387 13832
rect 38653 13774 41387 13776
rect 36004 13772 36051 13774
rect 35985 13771 36051 13772
rect 38653 13771 38719 13774
rect 41321 13771 41387 13774
rect 42333 13834 42399 13837
rect 42742 13834 42748 13836
rect 42333 13832 42748 13834
rect 42333 13776 42338 13832
rect 42394 13776 42748 13832
rect 42333 13774 42748 13776
rect 42333 13771 42399 13774
rect 42742 13772 42748 13774
rect 42812 13772 42818 13836
rect 21030 13698 21036 13700
rect 19198 13638 21036 13698
rect 17677 13635 17743 13638
rect 19057 13635 19123 13638
rect 21030 13636 21036 13638
rect 21100 13698 21106 13700
rect 21173 13698 21239 13701
rect 21100 13696 21239 13698
rect 21100 13640 21178 13696
rect 21234 13640 21239 13696
rect 21100 13638 21239 13640
rect 21100 13636 21106 13638
rect 21173 13635 21239 13638
rect 21357 13698 21423 13701
rect 27521 13698 27587 13701
rect 21357 13696 27587 13698
rect 21357 13640 21362 13696
rect 21418 13640 27526 13696
rect 27582 13640 27587 13696
rect 21357 13638 27587 13640
rect 21357 13635 21423 13638
rect 27521 13635 27587 13638
rect 28073 13698 28139 13701
rect 28901 13698 28967 13701
rect 28073 13696 28967 13698
rect 28073 13640 28078 13696
rect 28134 13640 28906 13696
rect 28962 13640 28967 13696
rect 28073 13638 28967 13640
rect 28073 13635 28139 13638
rect 28901 13635 28967 13638
rect 34145 13698 34211 13701
rect 40033 13698 40099 13701
rect 34145 13696 40099 13698
rect 34145 13640 34150 13696
rect 34206 13640 40038 13696
rect 40094 13640 40099 13696
rect 34145 13638 40099 13640
rect 34145 13635 34211 13638
rect 40033 13635 40099 13638
rect 10576 13632 10896 13633
rect 10576 13568 10584 13632
rect 10648 13568 10664 13632
rect 10728 13568 10744 13632
rect 10808 13568 10824 13632
rect 10888 13568 10896 13632
rect 10576 13567 10896 13568
rect 29840 13632 30160 13633
rect 29840 13568 29848 13632
rect 29912 13568 29928 13632
rect 29992 13568 30008 13632
rect 30072 13568 30088 13632
rect 30152 13568 30160 13632
rect 29840 13567 30160 13568
rect 49104 13632 49424 13633
rect 49104 13568 49112 13632
rect 49176 13568 49192 13632
rect 49256 13568 49272 13632
rect 49336 13568 49352 13632
rect 49416 13568 49424 13632
rect 49104 13567 49424 13568
rect 19374 13500 19380 13564
rect 19444 13562 19450 13564
rect 20713 13562 20779 13565
rect 19444 13560 20779 13562
rect 19444 13504 20718 13560
rect 20774 13504 20779 13560
rect 19444 13502 20779 13504
rect 19444 13500 19450 13502
rect 20713 13499 20779 13502
rect 21081 13562 21147 13565
rect 21541 13562 21607 13565
rect 21081 13560 21607 13562
rect 21081 13504 21086 13560
rect 21142 13504 21546 13560
rect 21602 13504 21607 13560
rect 21081 13502 21607 13504
rect 21081 13499 21147 13502
rect 21541 13499 21607 13502
rect 22001 13562 22067 13565
rect 26785 13562 26851 13565
rect 29269 13562 29335 13565
rect 22001 13560 24916 13562
rect 22001 13504 22006 13560
rect 22062 13504 24916 13560
rect 22001 13502 24916 13504
rect 22001 13499 22067 13502
rect 0 13426 800 13456
rect 1485 13426 1551 13429
rect 0 13424 1551 13426
rect 0 13368 1490 13424
rect 1546 13368 1551 13424
rect 0 13366 1551 13368
rect 0 13336 800 13366
rect 1485 13363 1551 13366
rect 19057 13426 19123 13429
rect 24669 13426 24735 13429
rect 19057 13424 24735 13426
rect 19057 13368 19062 13424
rect 19118 13368 24674 13424
rect 24730 13368 24735 13424
rect 19057 13366 24735 13368
rect 24856 13426 24916 13502
rect 26785 13560 29335 13562
rect 26785 13504 26790 13560
rect 26846 13504 29274 13560
rect 29330 13504 29335 13560
rect 26785 13502 29335 13504
rect 26785 13499 26851 13502
rect 29269 13499 29335 13502
rect 31937 13562 32003 13565
rect 34697 13562 34763 13565
rect 35249 13562 35315 13565
rect 38285 13564 38351 13565
rect 38285 13562 38332 13564
rect 31937 13560 34576 13562
rect 31937 13504 31942 13560
rect 31998 13504 34576 13560
rect 31937 13502 34576 13504
rect 31937 13499 32003 13502
rect 26969 13426 27035 13429
rect 29177 13426 29243 13429
rect 29821 13426 29887 13429
rect 24856 13424 27035 13426
rect 24856 13368 26974 13424
rect 27030 13368 27035 13424
rect 24856 13366 27035 13368
rect 19057 13363 19123 13366
rect 24669 13363 24735 13366
rect 26969 13363 27035 13366
rect 27110 13424 29887 13426
rect 27110 13368 29182 13424
rect 29238 13368 29826 13424
rect 29882 13368 29887 13424
rect 27110 13366 29887 13368
rect 18505 13290 18571 13293
rect 24945 13290 25011 13293
rect 25262 13290 25268 13292
rect 18505 13288 25268 13290
rect 18505 13232 18510 13288
rect 18566 13232 24950 13288
rect 25006 13232 25268 13288
rect 18505 13230 25268 13232
rect 18505 13227 18571 13230
rect 24945 13227 25011 13230
rect 25262 13228 25268 13230
rect 25332 13228 25338 13292
rect 20805 13154 20871 13157
rect 24209 13154 24275 13157
rect 27110 13154 27170 13366
rect 29177 13363 29243 13366
rect 29821 13363 29887 13366
rect 31017 13426 31083 13429
rect 33726 13426 33732 13428
rect 31017 13424 33732 13426
rect 31017 13368 31022 13424
rect 31078 13368 33732 13424
rect 31017 13366 33732 13368
rect 31017 13363 31083 13366
rect 33726 13364 33732 13366
rect 33796 13364 33802 13428
rect 34516 13426 34576 13502
rect 34697 13560 37474 13562
rect 34697 13504 34702 13560
rect 34758 13504 35254 13560
rect 35310 13504 37474 13560
rect 34697 13502 37474 13504
rect 38240 13560 38332 13562
rect 38240 13504 38290 13560
rect 38240 13502 38332 13504
rect 34697 13499 34763 13502
rect 35249 13499 35315 13502
rect 36721 13426 36787 13429
rect 34516 13424 36787 13426
rect 34516 13368 36726 13424
rect 36782 13368 36787 13424
rect 34516 13366 36787 13368
rect 36721 13363 36787 13366
rect 27521 13290 27587 13293
rect 37273 13290 37339 13293
rect 27521 13288 37339 13290
rect 27521 13232 27526 13288
rect 27582 13232 37278 13288
rect 37334 13232 37339 13288
rect 27521 13230 37339 13232
rect 37414 13290 37474 13502
rect 38285 13500 38332 13502
rect 38396 13500 38402 13564
rect 38285 13499 38351 13500
rect 43345 13290 43411 13293
rect 37414 13288 43411 13290
rect 37414 13232 43350 13288
rect 43406 13232 43411 13288
rect 37414 13230 43411 13232
rect 27521 13227 27587 13230
rect 37273 13227 37339 13230
rect 43345 13227 43411 13230
rect 58157 13290 58223 13293
rect 59200 13290 60000 13320
rect 58157 13288 60000 13290
rect 58157 13232 58162 13288
rect 58218 13232 60000 13288
rect 58157 13230 60000 13232
rect 58157 13227 58223 13230
rect 59200 13200 60000 13230
rect 20805 13152 27170 13154
rect 20805 13096 20810 13152
rect 20866 13096 24214 13152
rect 24270 13096 27170 13152
rect 20805 13094 27170 13096
rect 28349 13154 28415 13157
rect 29821 13154 29887 13157
rect 28349 13152 29010 13154
rect 28349 13096 28354 13152
rect 28410 13096 29010 13152
rect 28349 13094 29010 13096
rect 20805 13091 20871 13094
rect 24209 13091 24275 13094
rect 28349 13091 28415 13094
rect 20208 13088 20528 13089
rect 20208 13024 20216 13088
rect 20280 13024 20296 13088
rect 20360 13024 20376 13088
rect 20440 13024 20456 13088
rect 20520 13024 20528 13088
rect 20208 13023 20528 13024
rect 21214 12956 21220 13020
rect 21284 13018 21290 13020
rect 25405 13018 25471 13021
rect 26417 13020 26483 13021
rect 21284 13016 25471 13018
rect 21284 12960 25410 13016
rect 25466 12960 25471 13016
rect 21284 12958 25471 12960
rect 21284 12956 21290 12958
rect 25405 12955 25471 12958
rect 26366 12956 26372 13020
rect 26436 13018 26483 13020
rect 26436 13016 26528 13018
rect 26478 12960 26528 13016
rect 26436 12958 26528 12960
rect 26436 12956 26483 12958
rect 27654 12956 27660 13020
rect 27724 13018 27730 13020
rect 28717 13018 28783 13021
rect 27724 13016 28783 13018
rect 27724 12960 28722 13016
rect 28778 12960 28783 13016
rect 27724 12958 28783 12960
rect 28950 13018 29010 13094
rect 29821 13152 39314 13154
rect 29821 13096 29826 13152
rect 29882 13096 39314 13152
rect 29821 13094 39314 13096
rect 29821 13091 29887 13094
rect 35985 13018 36051 13021
rect 28950 13016 36051 13018
rect 28950 12960 35990 13016
rect 36046 12960 36051 13016
rect 28950 12958 36051 12960
rect 27724 12956 27730 12958
rect 26417 12955 26483 12956
rect 28717 12955 28783 12958
rect 35985 12955 36051 12958
rect 17861 12882 17927 12885
rect 32397 12882 32463 12885
rect 17861 12880 32463 12882
rect 17861 12824 17866 12880
rect 17922 12824 32402 12880
rect 32458 12824 32463 12880
rect 17861 12822 32463 12824
rect 17861 12819 17927 12822
rect 32397 12819 32463 12822
rect 32857 12882 32923 12885
rect 35249 12882 35315 12885
rect 37365 12882 37431 12885
rect 38745 12884 38811 12885
rect 32857 12880 37431 12882
rect 32857 12824 32862 12880
rect 32918 12824 35254 12880
rect 35310 12824 37370 12880
rect 37426 12824 37431 12880
rect 32857 12822 37431 12824
rect 32857 12819 32923 12822
rect 35249 12819 35315 12822
rect 37365 12819 37431 12822
rect 38694 12820 38700 12884
rect 38764 12882 38811 12884
rect 39254 12882 39314 13094
rect 39472 13088 39792 13089
rect 39472 13024 39480 13088
rect 39544 13024 39560 13088
rect 39624 13024 39640 13088
rect 39704 13024 39720 13088
rect 39784 13024 39792 13088
rect 39472 13023 39792 13024
rect 40033 12882 40099 12885
rect 38764 12880 38856 12882
rect 38806 12824 38856 12880
rect 38764 12822 38856 12824
rect 39254 12880 40099 12882
rect 39254 12824 40038 12880
rect 40094 12824 40099 12880
rect 39254 12822 40099 12824
rect 38764 12820 38811 12822
rect 38745 12819 38811 12820
rect 40033 12819 40099 12822
rect 20662 12684 20668 12748
rect 20732 12746 20738 12748
rect 24761 12746 24827 12749
rect 20732 12744 24827 12746
rect 20732 12688 24766 12744
rect 24822 12688 24827 12744
rect 20732 12686 24827 12688
rect 20732 12684 20738 12686
rect 24761 12683 24827 12686
rect 25129 12746 25195 12749
rect 25814 12746 25820 12748
rect 25129 12744 25820 12746
rect 25129 12688 25134 12744
rect 25190 12688 25820 12744
rect 25129 12686 25820 12688
rect 25129 12683 25195 12686
rect 25814 12684 25820 12686
rect 25884 12684 25890 12748
rect 27838 12684 27844 12748
rect 27908 12746 27914 12748
rect 29085 12746 29151 12749
rect 27908 12744 29151 12746
rect 27908 12688 29090 12744
rect 29146 12688 29151 12744
rect 27908 12686 29151 12688
rect 27908 12684 27914 12686
rect 29085 12683 29151 12686
rect 29318 12686 30850 12746
rect 18229 12610 18295 12613
rect 18229 12608 24962 12610
rect 18229 12552 18234 12608
rect 18290 12552 24962 12608
rect 18229 12550 24962 12552
rect 18229 12547 18295 12550
rect 10576 12544 10896 12545
rect 10576 12480 10584 12544
rect 10648 12480 10664 12544
rect 10728 12480 10744 12544
rect 10808 12480 10824 12544
rect 10888 12480 10896 12544
rect 10576 12479 10896 12480
rect 21582 12412 21588 12476
rect 21652 12474 21658 12476
rect 21817 12474 21883 12477
rect 21652 12472 21883 12474
rect 21652 12416 21822 12472
rect 21878 12416 21883 12472
rect 21652 12414 21883 12416
rect 21652 12412 21658 12414
rect 21817 12411 21883 12414
rect 22461 12474 22527 12477
rect 24669 12474 24735 12477
rect 22461 12472 24735 12474
rect 22461 12416 22466 12472
rect 22522 12416 24674 12472
rect 24730 12416 24735 12472
rect 22461 12414 24735 12416
rect 22461 12411 22527 12414
rect 24669 12411 24735 12414
rect 16481 12338 16547 12341
rect 16481 12336 24410 12338
rect 16481 12280 16486 12336
rect 16542 12280 24410 12336
rect 16481 12278 24410 12280
rect 16481 12275 16547 12278
rect 23749 12202 23815 12205
rect 19934 12200 23815 12202
rect 19934 12144 23754 12200
rect 23810 12144 23815 12200
rect 19934 12142 23815 12144
rect 24350 12202 24410 12278
rect 24526 12276 24532 12340
rect 24596 12338 24602 12340
rect 24761 12338 24827 12341
rect 24596 12336 24827 12338
rect 24596 12280 24766 12336
rect 24822 12280 24827 12336
rect 24596 12278 24827 12280
rect 24902 12338 24962 12550
rect 28022 12548 28028 12612
rect 28092 12610 28098 12612
rect 28257 12610 28323 12613
rect 28092 12608 28323 12610
rect 28092 12552 28262 12608
rect 28318 12552 28323 12608
rect 28092 12550 28323 12552
rect 28092 12548 28098 12550
rect 28257 12547 28323 12550
rect 26049 12474 26115 12477
rect 29318 12474 29378 12686
rect 29545 12612 29611 12613
rect 29494 12610 29500 12612
rect 29454 12550 29500 12610
rect 29564 12608 29611 12612
rect 29606 12552 29611 12608
rect 29494 12548 29500 12550
rect 29564 12548 29611 12552
rect 29545 12547 29611 12548
rect 30373 12610 30439 12613
rect 30790 12610 30850 12686
rect 30966 12684 30972 12748
rect 31036 12746 31042 12748
rect 31293 12746 31359 12749
rect 31036 12744 31359 12746
rect 31036 12688 31298 12744
rect 31354 12688 31359 12744
rect 31036 12686 31359 12688
rect 31036 12684 31042 12686
rect 31293 12683 31359 12686
rect 35617 12746 35683 12749
rect 36261 12746 36327 12749
rect 35617 12744 36327 12746
rect 35617 12688 35622 12744
rect 35678 12688 36266 12744
rect 36322 12688 36327 12744
rect 35617 12686 36327 12688
rect 35617 12683 35683 12686
rect 36261 12683 36327 12686
rect 36721 12746 36787 12749
rect 37825 12746 37891 12749
rect 36721 12744 37891 12746
rect 36721 12688 36726 12744
rect 36782 12688 37830 12744
rect 37886 12688 37891 12744
rect 36721 12686 37891 12688
rect 36721 12683 36787 12686
rect 37825 12683 37891 12686
rect 38009 12746 38075 12749
rect 38929 12748 38995 12749
rect 38878 12746 38884 12748
rect 38009 12744 38884 12746
rect 38948 12746 38995 12748
rect 39297 12746 39363 12749
rect 40493 12746 40559 12749
rect 38948 12744 39040 12746
rect 38009 12688 38014 12744
rect 38070 12688 38884 12744
rect 38990 12688 39040 12744
rect 38009 12686 38884 12688
rect 38009 12683 38075 12686
rect 38878 12684 38884 12686
rect 38948 12686 39040 12688
rect 39297 12744 40559 12746
rect 39297 12688 39302 12744
rect 39358 12688 40498 12744
rect 40554 12688 40559 12744
rect 39297 12686 40559 12688
rect 38948 12684 38995 12686
rect 38929 12683 38995 12684
rect 39297 12683 39363 12686
rect 40493 12683 40559 12686
rect 30373 12608 30666 12610
rect 30373 12552 30378 12608
rect 30434 12552 30666 12608
rect 30373 12550 30666 12552
rect 30790 12550 33058 12610
rect 30373 12547 30439 12550
rect 29840 12544 30160 12545
rect 29840 12480 29848 12544
rect 29912 12480 29928 12544
rect 29992 12480 30008 12544
rect 30072 12480 30088 12544
rect 30152 12480 30160 12544
rect 29840 12479 30160 12480
rect 26049 12472 29378 12474
rect 26049 12416 26054 12472
rect 26110 12416 29378 12472
rect 26049 12414 29378 12416
rect 30606 12474 30666 12550
rect 30741 12474 30807 12477
rect 32305 12474 32371 12477
rect 32581 12474 32647 12477
rect 30606 12472 30807 12474
rect 30606 12416 30746 12472
rect 30802 12416 30807 12472
rect 30606 12414 30807 12416
rect 26049 12411 26115 12414
rect 30741 12411 30807 12414
rect 31342 12414 32184 12474
rect 27337 12338 27403 12341
rect 31342 12338 31402 12414
rect 24902 12336 27403 12338
rect 24902 12280 27342 12336
rect 27398 12280 27403 12336
rect 24902 12278 27403 12280
rect 24596 12276 24602 12278
rect 24761 12275 24827 12278
rect 27337 12275 27403 12278
rect 27478 12278 31402 12338
rect 31477 12338 31543 12341
rect 31886 12338 31892 12340
rect 31477 12336 31892 12338
rect 31477 12280 31482 12336
rect 31538 12280 31892 12336
rect 31477 12278 31892 12280
rect 24669 12202 24735 12205
rect 24350 12200 24735 12202
rect 24350 12144 24674 12200
rect 24730 12144 24735 12200
rect 24350 12142 24735 12144
rect 15929 12066 15995 12069
rect 19934 12066 19994 12142
rect 23749 12139 23815 12142
rect 24669 12139 24735 12142
rect 26877 12202 26943 12205
rect 27478 12202 27538 12278
rect 31477 12275 31543 12278
rect 31886 12276 31892 12278
rect 31956 12276 31962 12340
rect 32124 12338 32184 12414
rect 32305 12472 32647 12474
rect 32305 12416 32310 12472
rect 32366 12416 32586 12472
rect 32642 12416 32647 12472
rect 32305 12414 32647 12416
rect 32998 12474 33058 12550
rect 33726 12548 33732 12612
rect 33796 12610 33802 12612
rect 35249 12610 35315 12613
rect 33796 12608 35315 12610
rect 33796 12552 35254 12608
rect 35310 12552 35315 12608
rect 33796 12550 35315 12552
rect 33796 12548 33802 12550
rect 35249 12547 35315 12550
rect 35617 12610 35683 12613
rect 40401 12610 40467 12613
rect 35617 12608 40467 12610
rect 35617 12552 35622 12608
rect 35678 12552 40406 12608
rect 40462 12552 40467 12608
rect 35617 12550 40467 12552
rect 35617 12547 35683 12550
rect 40401 12547 40467 12550
rect 49104 12544 49424 12545
rect 49104 12480 49112 12544
rect 49176 12480 49192 12544
rect 49256 12480 49272 12544
rect 49336 12480 49352 12544
rect 49416 12480 49424 12544
rect 49104 12479 49424 12480
rect 36721 12474 36787 12477
rect 32998 12472 36787 12474
rect 32998 12416 36726 12472
rect 36782 12416 36787 12472
rect 32998 12414 36787 12416
rect 32305 12411 32371 12414
rect 32581 12411 32647 12414
rect 36721 12411 36787 12414
rect 36905 12474 36971 12477
rect 39297 12474 39363 12477
rect 36905 12472 39363 12474
rect 36905 12416 36910 12472
rect 36966 12416 39302 12472
rect 39358 12416 39363 12472
rect 36905 12414 39363 12416
rect 36905 12411 36971 12414
rect 39297 12411 39363 12414
rect 39481 12474 39547 12477
rect 44357 12474 44423 12477
rect 39481 12472 44423 12474
rect 39481 12416 39486 12472
rect 39542 12416 44362 12472
rect 44418 12416 44423 12472
rect 39481 12414 44423 12416
rect 39481 12411 39547 12414
rect 44357 12411 44423 12414
rect 35801 12338 35867 12341
rect 32124 12336 35867 12338
rect 32124 12280 35806 12336
rect 35862 12280 35867 12336
rect 32124 12278 35867 12280
rect 35801 12275 35867 12278
rect 36813 12338 36879 12341
rect 38653 12338 38719 12341
rect 40401 12340 40467 12341
rect 40350 12338 40356 12340
rect 36813 12336 38719 12338
rect 36813 12280 36818 12336
rect 36874 12280 38658 12336
rect 38714 12280 38719 12336
rect 36813 12278 38719 12280
rect 40310 12278 40356 12338
rect 40420 12336 40467 12340
rect 40462 12280 40467 12336
rect 36813 12275 36879 12278
rect 38653 12275 38719 12278
rect 40350 12276 40356 12278
rect 40420 12276 40467 12280
rect 40401 12275 40467 12276
rect 26877 12200 27538 12202
rect 26877 12144 26882 12200
rect 26938 12144 27538 12200
rect 26877 12142 27538 12144
rect 27889 12202 27955 12205
rect 37273 12202 37339 12205
rect 45185 12202 45251 12205
rect 27889 12200 37339 12202
rect 27889 12144 27894 12200
rect 27950 12144 37278 12200
rect 37334 12144 37339 12200
rect 27889 12142 37339 12144
rect 26877 12139 26943 12142
rect 27889 12139 27955 12142
rect 37273 12139 37339 12142
rect 37414 12200 45251 12202
rect 37414 12144 45190 12200
rect 45246 12144 45251 12200
rect 37414 12142 45251 12144
rect 20897 12068 20963 12069
rect 20846 12066 20852 12068
rect 15929 12064 19994 12066
rect 15929 12008 15934 12064
rect 15990 12008 19994 12064
rect 15929 12006 19994 12008
rect 20806 12006 20852 12066
rect 20916 12064 20963 12068
rect 20958 12008 20963 12064
rect 15929 12003 15995 12006
rect 20846 12004 20852 12006
rect 20916 12004 20963 12008
rect 20897 12003 20963 12004
rect 26233 12066 26299 12069
rect 28574 12066 28580 12068
rect 26233 12064 28580 12066
rect 26233 12008 26238 12064
rect 26294 12008 28580 12064
rect 26233 12006 28580 12008
rect 26233 12003 26299 12006
rect 28574 12004 28580 12006
rect 28644 12004 28650 12068
rect 28901 12066 28967 12069
rect 30230 12066 30236 12068
rect 28901 12064 30236 12066
rect 28901 12008 28906 12064
rect 28962 12008 30236 12064
rect 28901 12006 30236 12008
rect 28901 12003 28967 12006
rect 30230 12004 30236 12006
rect 30300 12004 30306 12068
rect 31017 12066 31083 12069
rect 34646 12066 34652 12068
rect 31017 12064 34652 12066
rect 31017 12008 31022 12064
rect 31078 12008 34652 12064
rect 31017 12006 34652 12008
rect 31017 12003 31083 12006
rect 34646 12004 34652 12006
rect 34716 12004 34722 12068
rect 20208 12000 20528 12001
rect 20208 11936 20216 12000
rect 20280 11936 20296 12000
rect 20360 11936 20376 12000
rect 20440 11936 20456 12000
rect 20520 11936 20528 12000
rect 20208 11935 20528 11936
rect 26233 11930 26299 11933
rect 30925 11930 30991 11933
rect 26233 11928 30991 11930
rect 26233 11872 26238 11928
rect 26294 11872 30930 11928
rect 30986 11872 30991 11928
rect 26233 11870 30991 11872
rect 26233 11867 26299 11870
rect 30925 11867 30991 11870
rect 33501 11930 33567 11933
rect 37414 11930 37474 12142
rect 45185 12139 45251 12142
rect 39982 12004 39988 12068
rect 40052 12066 40058 12068
rect 41413 12066 41479 12069
rect 40052 12064 41479 12066
rect 40052 12008 41418 12064
rect 41474 12008 41479 12064
rect 40052 12006 41479 12008
rect 40052 12004 40058 12006
rect 41413 12003 41479 12006
rect 39472 12000 39792 12001
rect 39472 11936 39480 12000
rect 39544 11936 39560 12000
rect 39624 11936 39640 12000
rect 39704 11936 39720 12000
rect 39784 11936 39792 12000
rect 39472 11935 39792 11936
rect 33501 11928 37474 11930
rect 33501 11872 33506 11928
rect 33562 11872 37474 11928
rect 33501 11870 37474 11872
rect 33501 11867 33567 11870
rect 0 11794 800 11824
rect 1485 11794 1551 11797
rect 0 11792 1551 11794
rect 0 11736 1490 11792
rect 1546 11736 1551 11792
rect 0 11734 1551 11736
rect 0 11704 800 11734
rect 1485 11731 1551 11734
rect 17401 11794 17467 11797
rect 23657 11794 23723 11797
rect 17401 11792 23723 11794
rect 17401 11736 17406 11792
rect 17462 11736 23662 11792
rect 23718 11736 23723 11792
rect 17401 11734 23723 11736
rect 17401 11731 17467 11734
rect 23657 11731 23723 11734
rect 27889 11794 27955 11797
rect 28717 11794 28783 11797
rect 27889 11792 28783 11794
rect 27889 11736 27894 11792
rect 27950 11736 28722 11792
rect 28778 11736 28783 11792
rect 27889 11734 28783 11736
rect 27889 11731 27955 11734
rect 28717 11731 28783 11734
rect 29310 11732 29316 11796
rect 29380 11794 29386 11796
rect 30281 11794 30347 11797
rect 29380 11792 30347 11794
rect 29380 11736 30286 11792
rect 30342 11736 30347 11792
rect 29380 11734 30347 11736
rect 29380 11732 29386 11734
rect 30281 11731 30347 11734
rect 30557 11794 30623 11797
rect 35709 11794 35775 11797
rect 40309 11794 40375 11797
rect 30557 11792 35775 11794
rect 30557 11736 30562 11792
rect 30618 11736 35714 11792
rect 35770 11736 35775 11792
rect 30557 11734 35775 11736
rect 30557 11731 30623 11734
rect 35709 11731 35775 11734
rect 35942 11792 40375 11794
rect 35942 11736 40314 11792
rect 40370 11736 40375 11792
rect 35942 11734 40375 11736
rect 26785 11658 26851 11661
rect 30414 11658 30420 11660
rect 26785 11656 30420 11658
rect 26785 11600 26790 11656
rect 26846 11600 30420 11656
rect 26785 11598 30420 11600
rect 26785 11595 26851 11598
rect 30414 11596 30420 11598
rect 30484 11596 30490 11660
rect 30925 11658 30991 11661
rect 31753 11658 31819 11661
rect 30925 11656 31819 11658
rect 30925 11600 30930 11656
rect 30986 11600 31758 11656
rect 31814 11600 31819 11656
rect 30925 11598 31819 11600
rect 30925 11595 30991 11598
rect 31753 11595 31819 11598
rect 35617 11658 35683 11661
rect 35942 11658 36002 11734
rect 40309 11731 40375 11734
rect 40493 11794 40559 11797
rect 42057 11794 42123 11797
rect 40493 11792 42123 11794
rect 40493 11736 40498 11792
rect 40554 11736 42062 11792
rect 42118 11736 42123 11792
rect 40493 11734 42123 11736
rect 40493 11731 40559 11734
rect 42057 11731 42123 11734
rect 35617 11656 36002 11658
rect 35617 11600 35622 11656
rect 35678 11600 36002 11656
rect 35617 11598 36002 11600
rect 35617 11595 35683 11598
rect 36302 11596 36308 11660
rect 36372 11658 36378 11660
rect 43713 11658 43779 11661
rect 36372 11656 43779 11658
rect 36372 11600 43718 11656
rect 43774 11600 43779 11656
rect 36372 11598 43779 11600
rect 36372 11596 36378 11598
rect 43713 11595 43779 11598
rect 21214 11460 21220 11524
rect 21284 11522 21290 11524
rect 21541 11522 21607 11525
rect 21284 11520 21607 11522
rect 21284 11464 21546 11520
rect 21602 11464 21607 11520
rect 21284 11462 21607 11464
rect 21284 11460 21290 11462
rect 21541 11459 21607 11462
rect 21909 11522 21975 11525
rect 28809 11522 28875 11525
rect 21909 11520 28875 11522
rect 21909 11464 21914 11520
rect 21970 11464 28814 11520
rect 28870 11464 28875 11520
rect 21909 11462 28875 11464
rect 21909 11459 21975 11462
rect 28809 11459 28875 11462
rect 29269 11524 29335 11525
rect 29269 11520 29316 11524
rect 29380 11522 29386 11524
rect 29269 11464 29274 11520
rect 29269 11460 29316 11464
rect 29380 11462 29426 11522
rect 29380 11460 29386 11462
rect 30230 11460 30236 11524
rect 30300 11522 30306 11524
rect 31385 11522 31451 11525
rect 30300 11520 31451 11522
rect 30300 11464 31390 11520
rect 31446 11464 31451 11520
rect 30300 11462 31451 11464
rect 30300 11460 30306 11462
rect 29269 11459 29335 11460
rect 31385 11459 31451 11462
rect 32857 11522 32923 11525
rect 35801 11524 35867 11525
rect 37641 11524 37707 11525
rect 35750 11522 35756 11524
rect 32857 11520 35756 11522
rect 35820 11520 35867 11524
rect 37590 11522 37596 11524
rect 32857 11464 32862 11520
rect 32918 11464 35756 11520
rect 35862 11464 35867 11520
rect 32857 11462 35756 11464
rect 32857 11459 32923 11462
rect 35750 11460 35756 11462
rect 35820 11460 35867 11464
rect 37550 11462 37596 11522
rect 37660 11520 37707 11524
rect 37702 11464 37707 11520
rect 37590 11460 37596 11462
rect 37660 11460 37707 11464
rect 35801 11459 35867 11460
rect 37641 11459 37707 11460
rect 38101 11522 38167 11525
rect 40493 11522 40559 11525
rect 38101 11520 40559 11522
rect 38101 11464 38106 11520
rect 38162 11464 40498 11520
rect 40554 11464 40559 11520
rect 38101 11462 40559 11464
rect 38101 11459 38167 11462
rect 40493 11459 40559 11462
rect 58157 11522 58223 11525
rect 59200 11522 60000 11552
rect 58157 11520 60000 11522
rect 58157 11464 58162 11520
rect 58218 11464 60000 11520
rect 58157 11462 60000 11464
rect 58157 11459 58223 11462
rect 10576 11456 10896 11457
rect 10576 11392 10584 11456
rect 10648 11392 10664 11456
rect 10728 11392 10744 11456
rect 10808 11392 10824 11456
rect 10888 11392 10896 11456
rect 10576 11391 10896 11392
rect 29840 11456 30160 11457
rect 29840 11392 29848 11456
rect 29912 11392 29928 11456
rect 29992 11392 30008 11456
rect 30072 11392 30088 11456
rect 30152 11392 30160 11456
rect 29840 11391 30160 11392
rect 49104 11456 49424 11457
rect 49104 11392 49112 11456
rect 49176 11392 49192 11456
rect 49256 11392 49272 11456
rect 49336 11392 49352 11456
rect 49416 11392 49424 11456
rect 59200 11432 60000 11462
rect 49104 11391 49424 11392
rect 20437 11386 20503 11389
rect 20662 11386 20668 11388
rect 20437 11384 20668 11386
rect 20437 11328 20442 11384
rect 20498 11328 20668 11384
rect 20437 11326 20668 11328
rect 20437 11323 20503 11326
rect 20662 11324 20668 11326
rect 20732 11324 20738 11388
rect 21173 11386 21239 11389
rect 21909 11386 21975 11389
rect 22134 11386 22140 11388
rect 21173 11384 22140 11386
rect 21173 11328 21178 11384
rect 21234 11328 21914 11384
rect 21970 11328 22140 11384
rect 21173 11326 22140 11328
rect 21173 11323 21239 11326
rect 21909 11323 21975 11326
rect 22134 11324 22140 11326
rect 22204 11324 22210 11388
rect 24158 11324 24164 11388
rect 24228 11386 24234 11388
rect 25037 11386 25103 11389
rect 24228 11384 25103 11386
rect 24228 11328 25042 11384
rect 25098 11328 25103 11384
rect 24228 11326 25103 11328
rect 24228 11324 24234 11326
rect 25037 11323 25103 11326
rect 25446 11324 25452 11388
rect 25516 11386 25522 11388
rect 25589 11386 25655 11389
rect 26141 11386 26207 11389
rect 25516 11384 26207 11386
rect 25516 11328 25594 11384
rect 25650 11328 26146 11384
rect 26202 11328 26207 11384
rect 25516 11326 26207 11328
rect 25516 11324 25522 11326
rect 25589 11323 25655 11326
rect 26141 11323 26207 11326
rect 27102 11324 27108 11388
rect 27172 11386 27178 11388
rect 27337 11386 27403 11389
rect 27172 11384 27403 11386
rect 27172 11328 27342 11384
rect 27398 11328 27403 11384
rect 27172 11326 27403 11328
rect 27172 11324 27178 11326
rect 27337 11323 27403 11326
rect 28574 11324 28580 11388
rect 28644 11386 28650 11388
rect 29269 11386 29335 11389
rect 28644 11384 29335 11386
rect 28644 11328 29274 11384
rect 29330 11328 29335 11384
rect 28644 11326 29335 11328
rect 28644 11324 28650 11326
rect 29269 11323 29335 11326
rect 30741 11386 30807 11389
rect 34789 11386 34855 11389
rect 38837 11386 38903 11389
rect 43161 11386 43227 11389
rect 30741 11384 38903 11386
rect 30741 11328 30746 11384
rect 30802 11328 34794 11384
rect 34850 11328 38842 11384
rect 38898 11328 38903 11384
rect 30741 11326 38903 11328
rect 30741 11323 30807 11326
rect 34789 11323 34855 11326
rect 38837 11323 38903 11326
rect 41370 11384 43227 11386
rect 41370 11328 43166 11384
rect 43222 11328 43227 11384
rect 41370 11326 43227 11328
rect 31937 11250 32003 11253
rect 22050 11248 32003 11250
rect 22050 11192 31942 11248
rect 31998 11192 32003 11248
rect 22050 11190 32003 11192
rect 16573 11114 16639 11117
rect 19333 11114 19399 11117
rect 22050 11114 22110 11190
rect 31937 11187 32003 11190
rect 32078 11190 33426 11250
rect 16573 11112 22110 11114
rect 16573 11056 16578 11112
rect 16634 11056 19338 11112
rect 19394 11056 22110 11112
rect 16573 11054 22110 11056
rect 16573 11051 16639 11054
rect 19333 11051 19399 11054
rect 23974 11052 23980 11116
rect 24044 11114 24050 11116
rect 24301 11114 24367 11117
rect 24044 11112 24367 11114
rect 24044 11056 24306 11112
rect 24362 11056 24367 11112
rect 24044 11054 24367 11056
rect 24044 11052 24050 11054
rect 24301 11051 24367 11054
rect 26417 11114 26483 11117
rect 26918 11114 26924 11116
rect 26417 11112 26924 11114
rect 26417 11056 26422 11112
rect 26478 11056 26924 11112
rect 26417 11054 26924 11056
rect 26417 11051 26483 11054
rect 26918 11052 26924 11054
rect 26988 11052 26994 11116
rect 27061 11114 27127 11117
rect 28942 11114 28948 11116
rect 27061 11112 28948 11114
rect 27061 11056 27066 11112
rect 27122 11056 28948 11112
rect 27061 11054 28948 11056
rect 27061 11051 27127 11054
rect 28942 11052 28948 11054
rect 29012 11052 29018 11116
rect 31569 11114 31635 11117
rect 32078 11114 32138 11190
rect 31569 11112 32138 11114
rect 31569 11056 31574 11112
rect 31630 11056 32138 11112
rect 31569 11054 32138 11056
rect 32305 11114 32371 11117
rect 32806 11114 32812 11116
rect 32305 11112 32812 11114
rect 32305 11056 32310 11112
rect 32366 11056 32812 11112
rect 32305 11054 32812 11056
rect 31569 11051 31635 11054
rect 32305 11051 32371 11054
rect 32806 11052 32812 11054
rect 32876 11052 32882 11116
rect 33366 11114 33426 11190
rect 33542 11188 33548 11252
rect 33612 11250 33618 11252
rect 33777 11250 33843 11253
rect 33612 11248 33843 11250
rect 33612 11192 33782 11248
rect 33838 11192 33843 11248
rect 33612 11190 33843 11192
rect 33612 11188 33618 11190
rect 33777 11187 33843 11190
rect 35157 11250 35223 11253
rect 35934 11250 35940 11252
rect 35157 11248 35940 11250
rect 35157 11192 35162 11248
rect 35218 11192 35940 11248
rect 35157 11190 35940 11192
rect 35157 11187 35223 11190
rect 35934 11188 35940 11190
rect 36004 11188 36010 11252
rect 36813 11250 36879 11253
rect 41370 11250 41430 11326
rect 43161 11323 43227 11326
rect 36813 11248 41430 11250
rect 36813 11192 36818 11248
rect 36874 11192 41430 11248
rect 36813 11190 41430 11192
rect 36813 11187 36879 11190
rect 38653 11114 38719 11117
rect 33366 11112 38719 11114
rect 33366 11056 38658 11112
rect 38714 11056 38719 11112
rect 33366 11054 38719 11056
rect 38653 11051 38719 11054
rect 27705 10978 27771 10981
rect 33174 10978 33180 10980
rect 25086 10976 33180 10978
rect 25086 10920 27710 10976
rect 27766 10920 33180 10976
rect 25086 10918 33180 10920
rect 20208 10912 20528 10913
rect 20208 10848 20216 10912
rect 20280 10848 20296 10912
rect 20360 10848 20376 10912
rect 20440 10848 20456 10912
rect 20520 10848 20528 10912
rect 20208 10847 20528 10848
rect 22645 10842 22711 10845
rect 25086 10842 25146 10918
rect 27705 10915 27771 10918
rect 33174 10916 33180 10918
rect 33244 10916 33250 10980
rect 35617 10978 35683 10981
rect 37825 10978 37891 10981
rect 35617 10976 37891 10978
rect 35617 10920 35622 10976
rect 35678 10920 37830 10976
rect 37886 10920 37891 10976
rect 35617 10918 37891 10920
rect 35617 10915 35683 10918
rect 37825 10915 37891 10918
rect 39472 10912 39792 10913
rect 39472 10848 39480 10912
rect 39544 10848 39560 10912
rect 39624 10848 39640 10912
rect 39704 10848 39720 10912
rect 39784 10848 39792 10912
rect 39472 10847 39792 10848
rect 22645 10840 25146 10842
rect 22645 10784 22650 10840
rect 22706 10784 25146 10840
rect 22645 10782 25146 10784
rect 27981 10842 28047 10845
rect 34605 10842 34671 10845
rect 27981 10840 34671 10842
rect 27981 10784 27986 10840
rect 28042 10784 34610 10840
rect 34666 10784 34671 10840
rect 27981 10782 34671 10784
rect 22645 10779 22711 10782
rect 27981 10779 28047 10782
rect 34605 10779 34671 10782
rect 36118 10780 36124 10844
rect 36188 10842 36194 10844
rect 36261 10842 36327 10845
rect 36188 10840 36327 10842
rect 36188 10784 36266 10840
rect 36322 10784 36327 10840
rect 36188 10782 36327 10784
rect 36188 10780 36194 10782
rect 36261 10779 36327 10782
rect 21449 10706 21515 10709
rect 24761 10706 24827 10709
rect 21449 10704 24827 10706
rect 21449 10648 21454 10704
rect 21510 10648 24766 10704
rect 24822 10648 24827 10704
rect 21449 10646 24827 10648
rect 21449 10643 21515 10646
rect 24761 10643 24827 10646
rect 24945 10706 25011 10709
rect 29126 10706 29132 10708
rect 24945 10704 29132 10706
rect 24945 10648 24950 10704
rect 25006 10648 29132 10704
rect 24945 10646 29132 10648
rect 24945 10643 25011 10646
rect 29126 10644 29132 10646
rect 29196 10644 29202 10708
rect 30557 10706 30623 10709
rect 33041 10706 33107 10709
rect 33777 10708 33843 10709
rect 30557 10704 33107 10706
rect 30557 10648 30562 10704
rect 30618 10648 33046 10704
rect 33102 10648 33107 10704
rect 30557 10646 33107 10648
rect 30557 10643 30623 10646
rect 33041 10643 33107 10646
rect 33726 10644 33732 10708
rect 33796 10706 33843 10708
rect 35985 10706 36051 10709
rect 44541 10706 44607 10709
rect 33796 10704 33888 10706
rect 33838 10648 33888 10704
rect 33796 10646 33888 10648
rect 35985 10704 44607 10706
rect 35985 10648 35990 10704
rect 36046 10648 44546 10704
rect 44602 10648 44607 10704
rect 35985 10646 44607 10648
rect 33796 10644 33843 10646
rect 33777 10643 33843 10644
rect 35985 10643 36051 10646
rect 44541 10643 44607 10646
rect 26969 10570 27035 10573
rect 35525 10570 35591 10573
rect 45829 10570 45895 10573
rect 26969 10568 45895 10570
rect 26969 10512 26974 10568
rect 27030 10512 35530 10568
rect 35586 10512 45834 10568
rect 45890 10512 45895 10568
rect 26969 10510 45895 10512
rect 26969 10507 27035 10510
rect 35525 10507 35591 10510
rect 45829 10507 45895 10510
rect 24669 10434 24735 10437
rect 27797 10434 27863 10437
rect 28717 10434 28783 10437
rect 24669 10432 28783 10434
rect 24669 10376 24674 10432
rect 24730 10376 27802 10432
rect 27858 10376 28722 10432
rect 28778 10376 28783 10432
rect 24669 10374 28783 10376
rect 24669 10371 24735 10374
rect 27797 10371 27863 10374
rect 28717 10371 28783 10374
rect 32673 10434 32739 10437
rect 33685 10434 33751 10437
rect 32673 10432 33751 10434
rect 32673 10376 32678 10432
rect 32734 10376 33690 10432
rect 33746 10376 33751 10432
rect 32673 10374 33751 10376
rect 32673 10371 32739 10374
rect 33685 10371 33751 10374
rect 34237 10434 34303 10437
rect 35249 10434 35315 10437
rect 37222 10434 37228 10436
rect 34237 10432 37228 10434
rect 34237 10376 34242 10432
rect 34298 10376 35254 10432
rect 35310 10376 37228 10432
rect 34237 10374 37228 10376
rect 34237 10371 34303 10374
rect 35249 10371 35315 10374
rect 37222 10372 37228 10374
rect 37292 10372 37298 10436
rect 10576 10368 10896 10369
rect 10576 10304 10584 10368
rect 10648 10304 10664 10368
rect 10728 10304 10744 10368
rect 10808 10304 10824 10368
rect 10888 10304 10896 10368
rect 10576 10303 10896 10304
rect 29840 10368 30160 10369
rect 29840 10304 29848 10368
rect 29912 10304 29928 10368
rect 29992 10304 30008 10368
rect 30072 10304 30088 10368
rect 30152 10304 30160 10368
rect 29840 10303 30160 10304
rect 49104 10368 49424 10369
rect 49104 10304 49112 10368
rect 49176 10304 49192 10368
rect 49256 10304 49272 10368
rect 49336 10304 49352 10368
rect 49416 10304 49424 10368
rect 49104 10303 49424 10304
rect 22553 10298 22619 10301
rect 26233 10298 26299 10301
rect 22553 10296 26299 10298
rect 22553 10240 22558 10296
rect 22614 10240 26238 10296
rect 26294 10240 26299 10296
rect 22553 10238 26299 10240
rect 22553 10235 22619 10238
rect 26233 10235 26299 10238
rect 27981 10298 28047 10301
rect 28901 10298 28967 10301
rect 41413 10298 41479 10301
rect 27981 10296 28967 10298
rect 27981 10240 27986 10296
rect 28042 10240 28906 10296
rect 28962 10240 28967 10296
rect 27981 10238 28967 10240
rect 27981 10235 28047 10238
rect 28901 10235 28967 10238
rect 31710 10296 41479 10298
rect 31710 10240 41418 10296
rect 41474 10240 41479 10296
rect 31710 10238 41479 10240
rect 0 10162 800 10192
rect 1485 10162 1551 10165
rect 0 10160 1551 10162
rect 0 10104 1490 10160
rect 1546 10104 1551 10160
rect 0 10102 1551 10104
rect 0 10072 800 10102
rect 1485 10099 1551 10102
rect 23105 10162 23171 10165
rect 29361 10162 29427 10165
rect 29913 10162 29979 10165
rect 23105 10160 28826 10162
rect 23105 10104 23110 10160
rect 23166 10104 28826 10160
rect 23105 10102 28826 10104
rect 23105 10099 23171 10102
rect 18597 10026 18663 10029
rect 18597 10024 20730 10026
rect 18597 9968 18602 10024
rect 18658 9968 20730 10024
rect 18597 9966 20730 9968
rect 18597 9963 18663 9966
rect 20670 9890 20730 9966
rect 25262 9964 25268 10028
rect 25332 10026 25338 10028
rect 28533 10026 28599 10029
rect 25332 10024 28599 10026
rect 25332 9968 28538 10024
rect 28594 9968 28599 10024
rect 25332 9966 28599 9968
rect 28766 10026 28826 10102
rect 29361 10160 29979 10162
rect 29361 10104 29366 10160
rect 29422 10104 29918 10160
rect 29974 10104 29979 10160
rect 29361 10102 29979 10104
rect 29361 10099 29427 10102
rect 29913 10099 29979 10102
rect 30189 10162 30255 10165
rect 31710 10162 31770 10238
rect 41413 10235 41479 10238
rect 30189 10160 31770 10162
rect 30189 10104 30194 10160
rect 30250 10104 31770 10160
rect 30189 10102 31770 10104
rect 30189 10099 30255 10102
rect 35750 10100 35756 10164
rect 35820 10162 35826 10164
rect 38929 10162 38995 10165
rect 35820 10160 38995 10162
rect 35820 10104 38934 10160
rect 38990 10104 38995 10160
rect 35820 10102 38995 10104
rect 35820 10100 35826 10102
rect 38929 10099 38995 10102
rect 31937 10026 32003 10029
rect 34145 10026 34211 10029
rect 34881 10026 34947 10029
rect 28766 10024 34211 10026
rect 28766 9968 31942 10024
rect 31998 9968 34150 10024
rect 34206 9968 34211 10024
rect 28766 9966 34211 9968
rect 25332 9964 25338 9966
rect 28533 9963 28599 9966
rect 31937 9963 32003 9966
rect 34145 9963 34211 9966
rect 34838 10024 34947 10026
rect 34838 9968 34886 10024
rect 34942 9968 34947 10024
rect 34838 9963 34947 9968
rect 36077 10026 36143 10029
rect 37825 10026 37891 10029
rect 36077 10024 37891 10026
rect 36077 9968 36082 10024
rect 36138 9968 37830 10024
rect 37886 9968 37891 10024
rect 36077 9966 37891 9968
rect 36077 9963 36143 9966
rect 37825 9963 37891 9966
rect 29545 9890 29611 9893
rect 30005 9890 30071 9893
rect 20670 9888 30071 9890
rect 20670 9832 29550 9888
rect 29606 9832 30010 9888
rect 30066 9832 30071 9888
rect 20670 9830 30071 9832
rect 29545 9827 29611 9830
rect 30005 9827 30071 9830
rect 30741 9890 30807 9893
rect 31845 9890 31911 9893
rect 30741 9888 31911 9890
rect 30741 9832 30746 9888
rect 30802 9832 31850 9888
rect 31906 9832 31911 9888
rect 30741 9830 31911 9832
rect 30741 9827 30807 9830
rect 31845 9827 31911 9830
rect 32121 9890 32187 9893
rect 32489 9890 32555 9893
rect 34697 9890 34763 9893
rect 32121 9888 34763 9890
rect 32121 9832 32126 9888
rect 32182 9832 32494 9888
rect 32550 9832 34702 9888
rect 34758 9832 34763 9888
rect 32121 9830 34763 9832
rect 32121 9827 32187 9830
rect 32489 9827 32555 9830
rect 34697 9827 34763 9830
rect 20208 9824 20528 9825
rect 20208 9760 20216 9824
rect 20280 9760 20296 9824
rect 20360 9760 20376 9824
rect 20440 9760 20456 9824
rect 20520 9760 20528 9824
rect 20208 9759 20528 9760
rect 32121 9756 32187 9757
rect 21950 9692 21956 9756
rect 22020 9754 22026 9756
rect 30230 9754 30236 9756
rect 22020 9694 30236 9754
rect 22020 9692 22026 9694
rect 30230 9692 30236 9694
rect 30300 9692 30306 9756
rect 32070 9692 32076 9756
rect 32140 9754 32187 9756
rect 32990 9754 32996 9756
rect 32140 9752 32232 9754
rect 32182 9696 32232 9752
rect 32140 9694 32232 9696
rect 32308 9694 32996 9754
rect 32140 9692 32187 9694
rect 32121 9691 32187 9692
rect 27705 9618 27771 9621
rect 28441 9618 28507 9621
rect 27705 9616 28507 9618
rect 27705 9560 27710 9616
rect 27766 9560 28446 9616
rect 28502 9560 28507 9616
rect 27705 9558 28507 9560
rect 27705 9555 27771 9558
rect 28441 9555 28507 9558
rect 29678 9556 29684 9620
rect 29748 9618 29754 9620
rect 30097 9618 30163 9621
rect 29748 9616 30163 9618
rect 29748 9560 30102 9616
rect 30158 9560 30163 9616
rect 29748 9558 30163 9560
rect 29748 9556 29754 9558
rect 30097 9555 30163 9558
rect 30557 9618 30623 9621
rect 32308 9618 32368 9694
rect 32990 9692 32996 9694
rect 33060 9754 33066 9756
rect 33869 9754 33935 9757
rect 34513 9756 34579 9757
rect 34462 9754 34468 9756
rect 33060 9752 33935 9754
rect 33060 9696 33874 9752
rect 33930 9696 33935 9752
rect 33060 9694 33935 9696
rect 34422 9694 34468 9754
rect 34532 9752 34579 9756
rect 34574 9696 34579 9752
rect 33060 9692 33066 9694
rect 33869 9691 33935 9694
rect 34462 9692 34468 9694
rect 34532 9692 34579 9696
rect 34513 9691 34579 9692
rect 34838 9621 34898 9963
rect 39472 9824 39792 9825
rect 39472 9760 39480 9824
rect 39544 9760 39560 9824
rect 39624 9760 39640 9824
rect 39704 9760 39720 9824
rect 39784 9760 39792 9824
rect 39472 9759 39792 9760
rect 58157 9754 58223 9757
rect 59200 9754 60000 9784
rect 58157 9752 60000 9754
rect 58157 9696 58162 9752
rect 58218 9696 60000 9752
rect 58157 9694 60000 9696
rect 58157 9691 58223 9694
rect 59200 9664 60000 9694
rect 30557 9616 32368 9618
rect 30557 9560 30562 9616
rect 30618 9560 32368 9616
rect 30557 9558 32368 9560
rect 30557 9555 30623 9558
rect 32438 9556 32444 9620
rect 32508 9618 32514 9620
rect 33041 9618 33107 9621
rect 32508 9616 33107 9618
rect 32508 9560 33046 9616
rect 33102 9560 33107 9616
rect 32508 9558 33107 9560
rect 32508 9556 32514 9558
rect 33041 9555 33107 9558
rect 34094 9556 34100 9620
rect 34164 9618 34170 9620
rect 34421 9618 34487 9621
rect 34164 9616 34487 9618
rect 34164 9560 34426 9616
rect 34482 9560 34487 9616
rect 34164 9558 34487 9560
rect 34838 9616 34947 9621
rect 34838 9560 34886 9616
rect 34942 9560 34947 9616
rect 34838 9558 34947 9560
rect 34164 9556 34170 9558
rect 34421 9555 34487 9558
rect 34881 9555 34947 9558
rect 35014 9556 35020 9620
rect 35084 9618 35090 9620
rect 41505 9618 41571 9621
rect 35084 9616 41571 9618
rect 35084 9560 41510 9616
rect 41566 9560 41571 9616
rect 35084 9558 41571 9560
rect 35084 9556 35090 9558
rect 41505 9555 41571 9558
rect 16941 9482 17007 9485
rect 23565 9482 23631 9485
rect 24894 9482 24900 9484
rect 16941 9480 22110 9482
rect 16941 9424 16946 9480
rect 17002 9424 22110 9480
rect 16941 9422 22110 9424
rect 16941 9419 17007 9422
rect 10576 9280 10896 9281
rect 10576 9216 10584 9280
rect 10648 9216 10664 9280
rect 10728 9216 10744 9280
rect 10808 9216 10824 9280
rect 10888 9216 10896 9280
rect 10576 9215 10896 9216
rect 22050 8802 22110 9422
rect 23565 9480 24900 9482
rect 23565 9424 23570 9480
rect 23626 9424 24900 9480
rect 23565 9422 24900 9424
rect 23565 9419 23631 9422
rect 24894 9420 24900 9422
rect 24964 9420 24970 9484
rect 28717 9482 28783 9485
rect 30966 9482 30972 9484
rect 28717 9480 30972 9482
rect 28717 9424 28722 9480
rect 28778 9424 30972 9480
rect 28717 9422 30972 9424
rect 28717 9419 28783 9422
rect 30966 9420 30972 9422
rect 31036 9420 31042 9484
rect 32254 9420 32260 9484
rect 32324 9482 32330 9484
rect 35157 9482 35223 9485
rect 32324 9480 35223 9482
rect 32324 9424 35162 9480
rect 35218 9424 35223 9480
rect 32324 9422 35223 9424
rect 32324 9420 32330 9422
rect 35157 9419 35223 9422
rect 31477 9346 31543 9349
rect 34881 9346 34947 9349
rect 31477 9344 34947 9346
rect 31477 9288 31482 9344
rect 31538 9288 34886 9344
rect 34942 9288 34947 9344
rect 31477 9286 34947 9288
rect 31477 9283 31543 9286
rect 34881 9283 34947 9286
rect 29840 9280 30160 9281
rect 29840 9216 29848 9280
rect 29912 9216 29928 9280
rect 29992 9216 30008 9280
rect 30072 9216 30088 9280
rect 30152 9216 30160 9280
rect 29840 9215 30160 9216
rect 49104 9280 49424 9281
rect 49104 9216 49112 9280
rect 49176 9216 49192 9280
rect 49256 9216 49272 9280
rect 49336 9216 49352 9280
rect 49416 9216 49424 9280
rect 49104 9215 49424 9216
rect 26550 9148 26556 9212
rect 26620 9210 26626 9212
rect 27705 9210 27771 9213
rect 26620 9208 27771 9210
rect 26620 9152 27710 9208
rect 27766 9152 27771 9208
rect 26620 9150 27771 9152
rect 26620 9148 26626 9150
rect 27705 9147 27771 9150
rect 31845 9210 31911 9213
rect 35065 9210 35131 9213
rect 31845 9208 35131 9210
rect 31845 9152 31850 9208
rect 31906 9152 35070 9208
rect 35126 9152 35131 9208
rect 31845 9150 35131 9152
rect 31845 9147 31911 9150
rect 35065 9147 35131 9150
rect 27470 9012 27476 9076
rect 27540 9074 27546 9076
rect 28533 9074 28599 9077
rect 27540 9072 28599 9074
rect 27540 9016 28538 9072
rect 28594 9016 28599 9072
rect 27540 9014 28599 9016
rect 27540 9012 27546 9014
rect 28533 9011 28599 9014
rect 29913 9074 29979 9077
rect 37406 9074 37412 9076
rect 29913 9072 37412 9074
rect 29913 9016 29918 9072
rect 29974 9016 37412 9072
rect 29913 9014 37412 9016
rect 29913 9011 29979 9014
rect 37406 9012 37412 9014
rect 37476 9012 37482 9076
rect 25681 8938 25747 8941
rect 30557 8938 30623 8941
rect 25681 8936 30623 8938
rect 25681 8880 25686 8936
rect 25742 8880 30562 8936
rect 30618 8880 30623 8936
rect 25681 8878 30623 8880
rect 25681 8875 25747 8878
rect 30557 8875 30623 8878
rect 30598 8802 30604 8804
rect 22050 8742 30604 8802
rect 30598 8740 30604 8742
rect 30668 8740 30674 8804
rect 31385 8802 31451 8805
rect 36169 8802 36235 8805
rect 36997 8802 37063 8805
rect 31385 8800 37063 8802
rect 31385 8744 31390 8800
rect 31446 8744 36174 8800
rect 36230 8744 37002 8800
rect 37058 8744 37063 8800
rect 31385 8742 37063 8744
rect 31385 8739 31451 8742
rect 36169 8739 36235 8742
rect 36997 8739 37063 8742
rect 20208 8736 20528 8737
rect 0 8666 800 8696
rect 20208 8672 20216 8736
rect 20280 8672 20296 8736
rect 20360 8672 20376 8736
rect 20440 8672 20456 8736
rect 20520 8672 20528 8736
rect 20208 8671 20528 8672
rect 39472 8736 39792 8737
rect 39472 8672 39480 8736
rect 39544 8672 39560 8736
rect 39624 8672 39640 8736
rect 39704 8672 39720 8736
rect 39784 8672 39792 8736
rect 39472 8671 39792 8672
rect 1485 8666 1551 8669
rect 0 8664 1551 8666
rect 0 8608 1490 8664
rect 1546 8608 1551 8664
rect 0 8606 1551 8608
rect 0 8576 800 8606
rect 1485 8603 1551 8606
rect 23422 8604 23428 8668
rect 23492 8666 23498 8668
rect 28717 8666 28783 8669
rect 29913 8666 29979 8669
rect 23492 8664 28783 8666
rect 23492 8608 28722 8664
rect 28778 8608 28783 8664
rect 23492 8606 28783 8608
rect 23492 8604 23498 8606
rect 28717 8603 28783 8606
rect 28904 8664 29979 8666
rect 28904 8608 29918 8664
rect 29974 8608 29979 8664
rect 28904 8606 29979 8608
rect 28625 8530 28691 8533
rect 28904 8530 28964 8606
rect 29913 8603 29979 8606
rect 30557 8666 30623 8669
rect 31845 8666 31911 8669
rect 30557 8664 31911 8666
rect 30557 8608 30562 8664
rect 30618 8608 31850 8664
rect 31906 8608 31911 8664
rect 30557 8606 31911 8608
rect 30557 8603 30623 8606
rect 31845 8603 31911 8606
rect 34145 8666 34211 8669
rect 37365 8666 37431 8669
rect 34145 8664 37431 8666
rect 34145 8608 34150 8664
rect 34206 8608 37370 8664
rect 37426 8608 37431 8664
rect 34145 8606 37431 8608
rect 34145 8603 34211 8606
rect 37365 8603 37431 8606
rect 28625 8528 28964 8530
rect 28625 8472 28630 8528
rect 28686 8472 28964 8528
rect 28625 8470 28964 8472
rect 29637 8530 29703 8533
rect 30189 8530 30255 8533
rect 29637 8528 30255 8530
rect 29637 8472 29642 8528
rect 29698 8472 30194 8528
rect 30250 8472 30255 8528
rect 29637 8470 30255 8472
rect 28625 8467 28691 8470
rect 29637 8467 29703 8470
rect 30189 8467 30255 8470
rect 32857 8530 32923 8533
rect 34973 8530 35039 8533
rect 32857 8528 35039 8530
rect 32857 8472 32862 8528
rect 32918 8472 34978 8528
rect 35034 8472 35039 8528
rect 32857 8470 35039 8472
rect 32857 8467 32923 8470
rect 34973 8467 35039 8470
rect 26233 8394 26299 8397
rect 27654 8394 27660 8396
rect 26233 8392 27660 8394
rect 26233 8336 26238 8392
rect 26294 8336 27660 8392
rect 26233 8334 27660 8336
rect 26233 8331 26299 8334
rect 27654 8332 27660 8334
rect 27724 8332 27730 8396
rect 28942 8332 28948 8396
rect 29012 8394 29018 8396
rect 29637 8394 29703 8397
rect 29012 8392 29703 8394
rect 29012 8336 29642 8392
rect 29698 8336 29703 8392
rect 29012 8334 29703 8336
rect 29012 8332 29018 8334
rect 29637 8331 29703 8334
rect 15326 8196 15332 8260
rect 15396 8258 15402 8260
rect 29494 8258 29500 8260
rect 15396 8198 29500 8258
rect 15396 8196 15402 8198
rect 29494 8196 29500 8198
rect 29564 8196 29570 8260
rect 31661 8258 31727 8261
rect 32581 8258 32647 8261
rect 31661 8256 32647 8258
rect 31661 8200 31666 8256
rect 31722 8200 32586 8256
rect 32642 8200 32647 8256
rect 31661 8198 32647 8200
rect 31661 8195 31727 8198
rect 32581 8195 32647 8198
rect 33041 8258 33107 8261
rect 37089 8258 37155 8261
rect 33041 8256 37155 8258
rect 33041 8200 33046 8256
rect 33102 8200 37094 8256
rect 37150 8200 37155 8256
rect 33041 8198 37155 8200
rect 33041 8195 33107 8198
rect 37089 8195 37155 8198
rect 10576 8192 10896 8193
rect 10576 8128 10584 8192
rect 10648 8128 10664 8192
rect 10728 8128 10744 8192
rect 10808 8128 10824 8192
rect 10888 8128 10896 8192
rect 10576 8127 10896 8128
rect 29840 8192 30160 8193
rect 29840 8128 29848 8192
rect 29912 8128 29928 8192
rect 29992 8128 30008 8192
rect 30072 8128 30088 8192
rect 30152 8128 30160 8192
rect 29840 8127 30160 8128
rect 49104 8192 49424 8193
rect 49104 8128 49112 8192
rect 49176 8128 49192 8192
rect 49256 8128 49272 8192
rect 49336 8128 49352 8192
rect 49416 8128 49424 8192
rect 49104 8127 49424 8128
rect 19742 8060 19748 8124
rect 19812 8122 19818 8124
rect 24577 8122 24643 8125
rect 24761 8124 24827 8125
rect 19812 8120 24643 8122
rect 19812 8064 24582 8120
rect 24638 8064 24643 8120
rect 19812 8062 24643 8064
rect 19812 8060 19818 8062
rect 24577 8059 24643 8062
rect 24710 8060 24716 8124
rect 24780 8122 24827 8124
rect 24780 8120 24872 8122
rect 24822 8064 24872 8120
rect 24780 8062 24872 8064
rect 24780 8060 24827 8062
rect 25814 8060 25820 8124
rect 25884 8122 25890 8124
rect 25957 8122 26023 8125
rect 25884 8120 26023 8122
rect 25884 8064 25962 8120
rect 26018 8064 26023 8120
rect 25884 8062 26023 8064
rect 25884 8060 25890 8062
rect 24761 8059 24827 8060
rect 25957 8059 26023 8062
rect 31569 8122 31635 8125
rect 32029 8122 32095 8125
rect 31569 8120 32095 8122
rect 31569 8064 31574 8120
rect 31630 8064 32034 8120
rect 32090 8064 32095 8120
rect 31569 8062 32095 8064
rect 31569 8059 31635 8062
rect 32029 8059 32095 8062
rect 32213 8122 32279 8125
rect 34789 8122 34855 8125
rect 32213 8120 34855 8122
rect 32213 8064 32218 8120
rect 32274 8064 34794 8120
rect 34850 8064 34855 8120
rect 32213 8062 34855 8064
rect 32213 8059 32279 8062
rect 34789 8059 34855 8062
rect 18137 7986 18203 7989
rect 30649 7986 30715 7989
rect 33593 7986 33659 7989
rect 18137 7984 33659 7986
rect 18137 7928 18142 7984
rect 18198 7928 30654 7984
rect 30710 7928 33598 7984
rect 33654 7928 33659 7984
rect 18137 7926 33659 7928
rect 18137 7923 18203 7926
rect 30649 7923 30715 7926
rect 33593 7923 33659 7926
rect 58157 7986 58223 7989
rect 59200 7986 60000 8016
rect 58157 7984 60000 7986
rect 58157 7928 58162 7984
rect 58218 7928 60000 7984
rect 58157 7926 60000 7928
rect 58157 7923 58223 7926
rect 59200 7896 60000 7926
rect 19885 7850 19951 7853
rect 19885 7848 21650 7850
rect 19885 7792 19890 7848
rect 19946 7792 21650 7848
rect 19885 7790 21650 7792
rect 19885 7787 19951 7790
rect 21590 7714 21650 7790
rect 21766 7788 21772 7852
rect 21836 7850 21842 7852
rect 30465 7850 30531 7853
rect 21836 7848 30531 7850
rect 21836 7792 30470 7848
rect 30526 7792 30531 7848
rect 21836 7790 30531 7792
rect 21836 7788 21842 7790
rect 30465 7787 30531 7790
rect 30925 7850 30991 7853
rect 33961 7850 34027 7853
rect 30925 7848 34027 7850
rect 30925 7792 30930 7848
rect 30986 7792 33966 7848
rect 34022 7792 34027 7848
rect 30925 7790 34027 7792
rect 30925 7787 30991 7790
rect 33961 7787 34027 7790
rect 29085 7714 29151 7717
rect 31385 7714 31451 7717
rect 21590 7712 29151 7714
rect 21590 7656 29090 7712
rect 29146 7656 29151 7712
rect 21590 7654 29151 7656
rect 29085 7651 29151 7654
rect 29318 7712 31451 7714
rect 29318 7656 31390 7712
rect 31446 7656 31451 7712
rect 29318 7654 31451 7656
rect 20208 7648 20528 7649
rect 20208 7584 20216 7648
rect 20280 7584 20296 7648
rect 20360 7584 20376 7648
rect 20440 7584 20456 7648
rect 20520 7584 20528 7648
rect 20208 7583 20528 7584
rect 23013 7578 23079 7581
rect 29318 7578 29378 7654
rect 31385 7651 31451 7654
rect 39472 7648 39792 7649
rect 39472 7584 39480 7648
rect 39544 7584 39560 7648
rect 39624 7584 39640 7648
rect 39704 7584 39720 7648
rect 39784 7584 39792 7648
rect 39472 7583 39792 7584
rect 30281 7580 30347 7581
rect 30230 7578 30236 7580
rect 23013 7576 29378 7578
rect 23013 7520 23018 7576
rect 23074 7520 29378 7576
rect 23013 7518 29378 7520
rect 30190 7518 30236 7578
rect 30300 7576 30347 7580
rect 30342 7520 30347 7576
rect 23013 7515 23079 7518
rect 30230 7516 30236 7518
rect 30300 7516 30347 7520
rect 30281 7515 30347 7516
rect 31017 7578 31083 7581
rect 35893 7578 35959 7581
rect 31017 7576 35959 7578
rect 31017 7520 31022 7576
rect 31078 7520 35898 7576
rect 35954 7520 35959 7576
rect 31017 7518 35959 7520
rect 31017 7515 31083 7518
rect 35893 7515 35959 7518
rect 28758 7380 28764 7444
rect 28828 7442 28834 7444
rect 31109 7442 31175 7445
rect 28828 7440 31175 7442
rect 28828 7384 31114 7440
rect 31170 7384 31175 7440
rect 28828 7382 31175 7384
rect 28828 7380 28834 7382
rect 31109 7379 31175 7382
rect 33542 7380 33548 7444
rect 33612 7442 33618 7444
rect 41597 7442 41663 7445
rect 33612 7440 41663 7442
rect 33612 7384 41602 7440
rect 41658 7384 41663 7440
rect 33612 7382 41663 7384
rect 33612 7380 33618 7382
rect 41597 7379 41663 7382
rect 27889 7306 27955 7309
rect 34513 7306 34579 7309
rect 27889 7304 34579 7306
rect 27889 7248 27894 7304
rect 27950 7248 34518 7304
rect 34574 7248 34579 7304
rect 27889 7246 34579 7248
rect 27889 7243 27955 7246
rect 34513 7243 34579 7246
rect 10576 7104 10896 7105
rect 0 7034 800 7064
rect 10576 7040 10584 7104
rect 10648 7040 10664 7104
rect 10728 7040 10744 7104
rect 10808 7040 10824 7104
rect 10888 7040 10896 7104
rect 10576 7039 10896 7040
rect 29840 7104 30160 7105
rect 29840 7040 29848 7104
rect 29912 7040 29928 7104
rect 29992 7040 30008 7104
rect 30072 7040 30088 7104
rect 30152 7040 30160 7104
rect 29840 7039 30160 7040
rect 49104 7104 49424 7105
rect 49104 7040 49112 7104
rect 49176 7040 49192 7104
rect 49256 7040 49272 7104
rect 49336 7040 49352 7104
rect 49416 7040 49424 7104
rect 49104 7039 49424 7040
rect 1485 7034 1551 7037
rect 0 7032 1551 7034
rect 0 6976 1490 7032
rect 1546 6976 1551 7032
rect 0 6974 1551 6976
rect 0 6944 800 6974
rect 1485 6971 1551 6974
rect 17534 6836 17540 6900
rect 17604 6898 17610 6900
rect 32806 6898 32812 6900
rect 17604 6838 32812 6898
rect 17604 6836 17610 6838
rect 32806 6836 32812 6838
rect 32876 6836 32882 6900
rect 18454 6700 18460 6764
rect 18524 6762 18530 6764
rect 36486 6762 36492 6764
rect 18524 6702 36492 6762
rect 18524 6700 18530 6702
rect 36486 6700 36492 6702
rect 36556 6700 36562 6764
rect 40125 6762 40191 6765
rect 36678 6760 40191 6762
rect 36678 6704 40130 6760
rect 40186 6704 40191 6760
rect 36678 6702 40191 6704
rect 23197 6626 23263 6629
rect 35433 6626 35499 6629
rect 23197 6624 35499 6626
rect 23197 6568 23202 6624
rect 23258 6568 35438 6624
rect 35494 6568 35499 6624
rect 23197 6566 35499 6568
rect 23197 6563 23263 6566
rect 35433 6563 35499 6566
rect 20208 6560 20528 6561
rect 20208 6496 20216 6560
rect 20280 6496 20296 6560
rect 20360 6496 20376 6560
rect 20440 6496 20456 6560
rect 20520 6496 20528 6560
rect 20208 6495 20528 6496
rect 28441 6492 28507 6493
rect 28390 6428 28396 6492
rect 28460 6490 28507 6492
rect 29453 6490 29519 6493
rect 36678 6490 36738 6702
rect 40125 6699 40191 6702
rect 39472 6560 39792 6561
rect 39472 6496 39480 6560
rect 39544 6496 39560 6560
rect 39624 6496 39640 6560
rect 39704 6496 39720 6560
rect 39784 6496 39792 6560
rect 39472 6495 39792 6496
rect 28460 6488 28552 6490
rect 28502 6432 28552 6488
rect 28460 6430 28552 6432
rect 29453 6488 36738 6490
rect 29453 6432 29458 6488
rect 29514 6432 36738 6488
rect 29453 6430 36738 6432
rect 28460 6428 28507 6430
rect 28441 6427 28507 6428
rect 29453 6427 29519 6430
rect 17350 6292 17356 6356
rect 17420 6354 17426 6356
rect 42558 6354 42564 6356
rect 17420 6294 42564 6354
rect 17420 6292 17426 6294
rect 42558 6292 42564 6294
rect 42628 6292 42634 6356
rect 30230 6156 30236 6220
rect 30300 6218 30306 6220
rect 48129 6218 48195 6221
rect 30300 6216 48195 6218
rect 30300 6160 48134 6216
rect 48190 6160 48195 6216
rect 30300 6158 48195 6160
rect 30300 6156 30306 6158
rect 48129 6155 48195 6158
rect 58157 6218 58223 6221
rect 59200 6218 60000 6248
rect 58157 6216 60000 6218
rect 58157 6160 58162 6216
rect 58218 6160 60000 6216
rect 58157 6158 60000 6160
rect 58157 6155 58223 6158
rect 59200 6128 60000 6158
rect 10576 6016 10896 6017
rect 10576 5952 10584 6016
rect 10648 5952 10664 6016
rect 10728 5952 10744 6016
rect 10808 5952 10824 6016
rect 10888 5952 10896 6016
rect 10576 5951 10896 5952
rect 29840 6016 30160 6017
rect 29840 5952 29848 6016
rect 29912 5952 29928 6016
rect 29992 5952 30008 6016
rect 30072 5952 30088 6016
rect 30152 5952 30160 6016
rect 29840 5951 30160 5952
rect 49104 6016 49424 6017
rect 49104 5952 49112 6016
rect 49176 5952 49192 6016
rect 49256 5952 49272 6016
rect 49336 5952 49352 6016
rect 49416 5952 49424 6016
rect 49104 5951 49424 5952
rect 32857 5948 32923 5949
rect 32806 5884 32812 5948
rect 32876 5946 32923 5948
rect 32876 5944 32968 5946
rect 32918 5888 32968 5944
rect 32876 5886 32968 5888
rect 32876 5884 32923 5886
rect 32857 5883 32923 5884
rect 31109 5674 31175 5677
rect 48865 5674 48931 5677
rect 31109 5672 48931 5674
rect 31109 5616 31114 5672
rect 31170 5616 48870 5672
rect 48926 5616 48931 5672
rect 31109 5614 48931 5616
rect 31109 5611 31175 5614
rect 48865 5611 48931 5614
rect 23841 5538 23907 5541
rect 23841 5536 31770 5538
rect 23841 5480 23846 5536
rect 23902 5480 31770 5536
rect 23841 5478 31770 5480
rect 23841 5475 23907 5478
rect 20208 5472 20528 5473
rect 0 5402 800 5432
rect 20208 5408 20216 5472
rect 20280 5408 20296 5472
rect 20360 5408 20376 5472
rect 20440 5408 20456 5472
rect 20520 5408 20528 5472
rect 20208 5407 20528 5408
rect 1485 5402 1551 5405
rect 29453 5404 29519 5405
rect 29453 5402 29500 5404
rect 0 5400 1551 5402
rect 0 5344 1490 5400
rect 1546 5344 1551 5400
rect 0 5342 1551 5344
rect 29408 5400 29500 5402
rect 29408 5344 29458 5400
rect 29408 5342 29500 5344
rect 0 5312 800 5342
rect 1485 5339 1551 5342
rect 29453 5340 29500 5342
rect 29564 5340 29570 5404
rect 31710 5402 31770 5478
rect 39472 5472 39792 5473
rect 39472 5408 39480 5472
rect 39544 5408 39560 5472
rect 39624 5408 39640 5472
rect 39704 5408 39720 5472
rect 39784 5408 39792 5472
rect 39472 5407 39792 5408
rect 31710 5342 36554 5402
rect 29453 5339 29519 5340
rect 15469 5266 15535 5269
rect 35934 5266 35940 5268
rect 15469 5264 35940 5266
rect 15469 5208 15474 5264
rect 15530 5208 35940 5264
rect 15469 5206 35940 5208
rect 15469 5203 15535 5206
rect 35934 5204 35940 5206
rect 36004 5204 36010 5268
rect 36494 5266 36554 5342
rect 42190 5266 42196 5268
rect 36494 5206 42196 5266
rect 42190 5204 42196 5206
rect 42260 5204 42266 5268
rect 14825 5130 14891 5133
rect 33542 5130 33548 5132
rect 14825 5128 33548 5130
rect 14825 5072 14830 5128
rect 14886 5072 33548 5128
rect 14825 5070 33548 5072
rect 14825 5067 14891 5070
rect 33542 5068 33548 5070
rect 33612 5068 33618 5132
rect 37273 5130 37339 5133
rect 37590 5130 37596 5132
rect 37273 5128 37596 5130
rect 37273 5072 37278 5128
rect 37334 5072 37596 5128
rect 37273 5070 37596 5072
rect 37273 5067 37339 5070
rect 37590 5068 37596 5070
rect 37660 5068 37666 5132
rect 10576 4928 10896 4929
rect 10576 4864 10584 4928
rect 10648 4864 10664 4928
rect 10728 4864 10744 4928
rect 10808 4864 10824 4928
rect 10888 4864 10896 4928
rect 10576 4863 10896 4864
rect 29840 4928 30160 4929
rect 29840 4864 29848 4928
rect 29912 4864 29928 4928
rect 29992 4864 30008 4928
rect 30072 4864 30088 4928
rect 30152 4864 30160 4928
rect 29840 4863 30160 4864
rect 49104 4928 49424 4929
rect 49104 4864 49112 4928
rect 49176 4864 49192 4928
rect 49256 4864 49272 4928
rect 49336 4864 49352 4928
rect 49416 4864 49424 4928
rect 49104 4863 49424 4864
rect 14365 4722 14431 4725
rect 44398 4722 44404 4724
rect 14365 4720 44404 4722
rect 14365 4664 14370 4720
rect 14426 4664 44404 4720
rect 14365 4662 44404 4664
rect 14365 4659 14431 4662
rect 44398 4660 44404 4662
rect 44468 4660 44474 4724
rect 15101 4586 15167 4589
rect 34462 4586 34468 4588
rect 15101 4584 34468 4586
rect 15101 4528 15106 4584
rect 15162 4528 34468 4584
rect 15101 4526 34468 4528
rect 15101 4523 15167 4526
rect 34462 4524 34468 4526
rect 34532 4524 34538 4588
rect 58157 4450 58223 4453
rect 59200 4450 60000 4480
rect 58157 4448 60000 4450
rect 58157 4392 58162 4448
rect 58218 4392 60000 4448
rect 58157 4390 60000 4392
rect 58157 4387 58223 4390
rect 20208 4384 20528 4385
rect 20208 4320 20216 4384
rect 20280 4320 20296 4384
rect 20360 4320 20376 4384
rect 20440 4320 20456 4384
rect 20520 4320 20528 4384
rect 20208 4319 20528 4320
rect 39472 4384 39792 4385
rect 39472 4320 39480 4384
rect 39544 4320 39560 4384
rect 39624 4320 39640 4384
rect 39704 4320 39720 4384
rect 39784 4320 39792 4384
rect 59200 4360 60000 4390
rect 39472 4319 39792 4320
rect 25773 4178 25839 4181
rect 41638 4178 41644 4180
rect 25773 4176 41644 4178
rect 25773 4120 25778 4176
rect 25834 4120 41644 4176
rect 25773 4118 41644 4120
rect 25773 4115 25839 4118
rect 41638 4116 41644 4118
rect 41708 4116 41714 4180
rect 18822 3980 18828 4044
rect 18892 4042 18898 4044
rect 47025 4042 47091 4045
rect 18892 4040 47091 4042
rect 18892 3984 47030 4040
rect 47086 3984 47091 4040
rect 18892 3982 47091 3984
rect 18892 3980 18898 3982
rect 47025 3979 47091 3982
rect 0 3906 800 3936
rect 1485 3906 1551 3909
rect 0 3904 1551 3906
rect 0 3848 1490 3904
rect 1546 3848 1551 3904
rect 0 3846 1551 3848
rect 0 3816 800 3846
rect 1485 3843 1551 3846
rect 10576 3840 10896 3841
rect 10576 3776 10584 3840
rect 10648 3776 10664 3840
rect 10728 3776 10744 3840
rect 10808 3776 10824 3840
rect 10888 3776 10896 3840
rect 10576 3775 10896 3776
rect 29840 3840 30160 3841
rect 29840 3776 29848 3840
rect 29912 3776 29928 3840
rect 29992 3776 30008 3840
rect 30072 3776 30088 3840
rect 30152 3776 30160 3840
rect 29840 3775 30160 3776
rect 49104 3840 49424 3841
rect 49104 3776 49112 3840
rect 49176 3776 49192 3840
rect 49256 3776 49272 3840
rect 49336 3776 49352 3840
rect 49416 3776 49424 3840
rect 49104 3775 49424 3776
rect 26918 3572 26924 3636
rect 26988 3634 26994 3636
rect 47209 3634 47275 3637
rect 26988 3632 47275 3634
rect 26988 3576 47214 3632
rect 47270 3576 47275 3632
rect 26988 3574 47275 3576
rect 26988 3572 26994 3574
rect 47209 3571 47275 3574
rect 15377 3498 15443 3501
rect 42926 3498 42932 3500
rect 15377 3496 42932 3498
rect 15377 3440 15382 3496
rect 15438 3440 42932 3496
rect 15377 3438 42932 3440
rect 15377 3435 15443 3438
rect 42926 3436 42932 3438
rect 42996 3436 43002 3500
rect 24853 3362 24919 3365
rect 29310 3362 29316 3364
rect 24853 3360 29316 3362
rect 24853 3304 24858 3360
rect 24914 3304 29316 3360
rect 24853 3302 29316 3304
rect 24853 3299 24919 3302
rect 29310 3300 29316 3302
rect 29380 3362 29386 3364
rect 37733 3362 37799 3365
rect 29380 3360 37799 3362
rect 29380 3304 37738 3360
rect 37794 3304 37799 3360
rect 29380 3302 37799 3304
rect 29380 3300 29386 3302
rect 37733 3299 37799 3302
rect 20208 3296 20528 3297
rect 20208 3232 20216 3296
rect 20280 3232 20296 3296
rect 20360 3232 20376 3296
rect 20440 3232 20456 3296
rect 20520 3232 20528 3296
rect 20208 3231 20528 3232
rect 39472 3296 39792 3297
rect 39472 3232 39480 3296
rect 39544 3232 39560 3296
rect 39624 3232 39640 3296
rect 39704 3232 39720 3296
rect 39784 3232 39792 3296
rect 39472 3231 39792 3232
rect 21173 2954 21239 2957
rect 46054 2954 46060 2956
rect 21173 2952 46060 2954
rect 21173 2896 21178 2952
rect 21234 2896 46060 2952
rect 21173 2894 46060 2896
rect 21173 2891 21239 2894
rect 46054 2892 46060 2894
rect 46124 2892 46130 2956
rect 10576 2752 10896 2753
rect 10576 2688 10584 2752
rect 10648 2688 10664 2752
rect 10728 2688 10744 2752
rect 10808 2688 10824 2752
rect 10888 2688 10896 2752
rect 10576 2687 10896 2688
rect 29840 2752 30160 2753
rect 29840 2688 29848 2752
rect 29912 2688 29928 2752
rect 29992 2688 30008 2752
rect 30072 2688 30088 2752
rect 30152 2688 30160 2752
rect 29840 2687 30160 2688
rect 49104 2752 49424 2753
rect 49104 2688 49112 2752
rect 49176 2688 49192 2752
rect 49256 2688 49272 2752
rect 49336 2688 49352 2752
rect 49416 2688 49424 2752
rect 49104 2687 49424 2688
rect 56501 2682 56567 2685
rect 59200 2682 60000 2712
rect 56501 2680 60000 2682
rect 56501 2624 56506 2680
rect 56562 2624 60000 2680
rect 56501 2622 60000 2624
rect 56501 2619 56567 2622
rect 59200 2592 60000 2622
rect 24577 2546 24643 2549
rect 46606 2546 46612 2548
rect 24577 2544 46612 2546
rect 24577 2488 24582 2544
rect 24638 2488 46612 2544
rect 24577 2486 46612 2488
rect 24577 2483 24643 2486
rect 46606 2484 46612 2486
rect 46676 2484 46682 2548
rect 21909 2410 21975 2413
rect 42742 2410 42748 2412
rect 21909 2408 42748 2410
rect 21909 2352 21914 2408
rect 21970 2352 42748 2408
rect 21909 2350 42748 2352
rect 21909 2347 21975 2350
rect 42742 2348 42748 2350
rect 42812 2348 42818 2412
rect 0 2274 800 2304
rect 1393 2274 1459 2277
rect 0 2272 1459 2274
rect 0 2216 1398 2272
rect 1454 2216 1459 2272
rect 0 2214 1459 2216
rect 0 2184 800 2214
rect 1393 2211 1459 2214
rect 20208 2208 20528 2209
rect 20208 2144 20216 2208
rect 20280 2144 20296 2208
rect 20360 2144 20376 2208
rect 20440 2144 20456 2208
rect 20520 2144 20528 2208
rect 20208 2143 20528 2144
rect 39472 2208 39792 2209
rect 39472 2144 39480 2208
rect 39544 2144 39560 2208
rect 39624 2144 39640 2208
rect 39704 2144 39720 2208
rect 39784 2144 39792 2208
rect 39472 2143 39792 2144
rect 14549 2002 14615 2005
rect 44214 2002 44220 2004
rect 14549 2000 44220 2002
rect 14549 1944 14554 2000
rect 14610 1944 44220 2000
rect 14549 1942 44220 1944
rect 14549 1939 14615 1942
rect 44214 1940 44220 1942
rect 44284 1940 44290 2004
rect 16430 1804 16436 1868
rect 16500 1866 16506 1868
rect 35014 1866 35020 1868
rect 16500 1806 35020 1866
rect 16500 1804 16506 1806
rect 35014 1804 35020 1806
rect 35084 1804 35090 1868
rect 18086 1668 18092 1732
rect 18156 1730 18162 1732
rect 38009 1730 38075 1733
rect 18156 1728 38075 1730
rect 18156 1672 38014 1728
rect 38070 1672 38075 1728
rect 18156 1670 38075 1672
rect 18156 1668 18162 1670
rect 38009 1667 38075 1670
rect 28441 1594 28507 1597
rect 44950 1594 44956 1596
rect 28441 1592 44956 1594
rect 28441 1536 28446 1592
rect 28502 1536 44956 1592
rect 28441 1534 44956 1536
rect 28441 1531 28507 1534
rect 44950 1532 44956 1534
rect 45020 1532 45026 1596
rect 57881 914 57947 917
rect 59200 914 60000 944
rect 57881 912 60000 914
rect 57881 856 57886 912
rect 57942 856 60000 912
rect 57881 854 60000 856
rect 57881 851 57947 854
rect 59200 824 60000 854
rect 0 778 800 808
rect 1485 778 1551 781
rect 0 776 1551 778
rect 0 720 1490 776
rect 1546 720 1551 776
rect 0 718 1551 720
rect 0 688 800 718
rect 1485 715 1551 718
<< via3 >>
rect 24348 29820 24412 29884
rect 19196 29684 19260 29748
rect 40172 29276 40236 29340
rect 16804 29140 16868 29204
rect 17540 29004 17604 29068
rect 21220 28868 21284 28932
rect 42748 28732 42812 28796
rect 45140 28596 45204 28660
rect 40356 28460 40420 28524
rect 37596 28324 37660 28388
rect 19012 28188 19076 28252
rect 42012 28188 42076 28252
rect 21772 28052 21836 28116
rect 38332 27916 38396 27980
rect 40908 27780 40972 27844
rect 10584 27772 10648 27776
rect 10584 27716 10588 27772
rect 10588 27716 10644 27772
rect 10644 27716 10648 27772
rect 10584 27712 10648 27716
rect 10664 27772 10728 27776
rect 10664 27716 10668 27772
rect 10668 27716 10724 27772
rect 10724 27716 10728 27772
rect 10664 27712 10728 27716
rect 10744 27772 10808 27776
rect 10744 27716 10748 27772
rect 10748 27716 10804 27772
rect 10804 27716 10808 27772
rect 10744 27712 10808 27716
rect 10824 27772 10888 27776
rect 10824 27716 10828 27772
rect 10828 27716 10884 27772
rect 10884 27716 10888 27772
rect 10824 27712 10888 27716
rect 29848 27772 29912 27776
rect 29848 27716 29852 27772
rect 29852 27716 29908 27772
rect 29908 27716 29912 27772
rect 29848 27712 29912 27716
rect 29928 27772 29992 27776
rect 29928 27716 29932 27772
rect 29932 27716 29988 27772
rect 29988 27716 29992 27772
rect 29928 27712 29992 27716
rect 30008 27772 30072 27776
rect 30008 27716 30012 27772
rect 30012 27716 30068 27772
rect 30068 27716 30072 27772
rect 30008 27712 30072 27716
rect 30088 27772 30152 27776
rect 30088 27716 30092 27772
rect 30092 27716 30148 27772
rect 30148 27716 30152 27772
rect 30088 27712 30152 27716
rect 49112 27772 49176 27776
rect 49112 27716 49116 27772
rect 49116 27716 49172 27772
rect 49172 27716 49176 27772
rect 49112 27712 49176 27716
rect 49192 27772 49256 27776
rect 49192 27716 49196 27772
rect 49196 27716 49252 27772
rect 49252 27716 49256 27772
rect 49192 27712 49256 27716
rect 49272 27772 49336 27776
rect 49272 27716 49276 27772
rect 49276 27716 49332 27772
rect 49332 27716 49336 27772
rect 49272 27712 49336 27716
rect 49352 27772 49416 27776
rect 49352 27716 49356 27772
rect 49356 27716 49412 27772
rect 49412 27716 49416 27772
rect 49352 27712 49416 27716
rect 19748 27508 19812 27572
rect 39252 27508 39316 27572
rect 20216 27228 20280 27232
rect 20216 27172 20220 27228
rect 20220 27172 20276 27228
rect 20276 27172 20280 27228
rect 20216 27168 20280 27172
rect 20296 27228 20360 27232
rect 20296 27172 20300 27228
rect 20300 27172 20356 27228
rect 20356 27172 20360 27228
rect 20296 27168 20360 27172
rect 20376 27228 20440 27232
rect 20376 27172 20380 27228
rect 20380 27172 20436 27228
rect 20436 27172 20440 27228
rect 20376 27168 20440 27172
rect 20456 27228 20520 27232
rect 20456 27172 20460 27228
rect 20460 27172 20516 27228
rect 20516 27172 20520 27228
rect 20456 27168 20520 27172
rect 39480 27228 39544 27232
rect 39480 27172 39484 27228
rect 39484 27172 39540 27228
rect 39540 27172 39544 27228
rect 39480 27168 39544 27172
rect 39560 27228 39624 27232
rect 39560 27172 39564 27228
rect 39564 27172 39620 27228
rect 39620 27172 39624 27228
rect 39560 27168 39624 27172
rect 39640 27228 39704 27232
rect 39640 27172 39644 27228
rect 39644 27172 39700 27228
rect 39700 27172 39704 27228
rect 39640 27168 39704 27172
rect 39720 27228 39784 27232
rect 39720 27172 39724 27228
rect 39724 27172 39780 27228
rect 39780 27172 39784 27228
rect 39720 27168 39784 27172
rect 10584 26684 10648 26688
rect 10584 26628 10588 26684
rect 10588 26628 10644 26684
rect 10644 26628 10648 26684
rect 10584 26624 10648 26628
rect 10664 26684 10728 26688
rect 10664 26628 10668 26684
rect 10668 26628 10724 26684
rect 10724 26628 10728 26684
rect 10664 26624 10728 26628
rect 10744 26684 10808 26688
rect 10744 26628 10748 26684
rect 10748 26628 10804 26684
rect 10804 26628 10808 26684
rect 10744 26624 10808 26628
rect 10824 26684 10888 26688
rect 10824 26628 10828 26684
rect 10828 26628 10884 26684
rect 10884 26628 10888 26684
rect 10824 26624 10888 26628
rect 29848 26684 29912 26688
rect 29848 26628 29852 26684
rect 29852 26628 29908 26684
rect 29908 26628 29912 26684
rect 29848 26624 29912 26628
rect 29928 26684 29992 26688
rect 29928 26628 29932 26684
rect 29932 26628 29988 26684
rect 29988 26628 29992 26684
rect 29928 26624 29992 26628
rect 30008 26684 30072 26688
rect 30008 26628 30012 26684
rect 30012 26628 30068 26684
rect 30068 26628 30072 26684
rect 30008 26624 30072 26628
rect 30088 26684 30152 26688
rect 30088 26628 30092 26684
rect 30092 26628 30148 26684
rect 30148 26628 30152 26684
rect 30088 26624 30152 26628
rect 38700 26692 38764 26756
rect 49112 26684 49176 26688
rect 49112 26628 49116 26684
rect 49116 26628 49172 26684
rect 49172 26628 49176 26684
rect 49112 26624 49176 26628
rect 49192 26684 49256 26688
rect 49192 26628 49196 26684
rect 49196 26628 49252 26684
rect 49252 26628 49256 26684
rect 49192 26624 49256 26628
rect 49272 26684 49336 26688
rect 49272 26628 49276 26684
rect 49276 26628 49332 26684
rect 49332 26628 49336 26684
rect 49272 26624 49336 26628
rect 49352 26684 49416 26688
rect 49352 26628 49356 26684
rect 49356 26628 49412 26684
rect 49412 26628 49416 26684
rect 49352 26624 49416 26628
rect 37412 26556 37476 26620
rect 21956 26284 22020 26348
rect 30788 26284 30852 26348
rect 32628 26284 32692 26348
rect 20216 26140 20280 26144
rect 20216 26084 20220 26140
rect 20220 26084 20276 26140
rect 20276 26084 20280 26140
rect 20216 26080 20280 26084
rect 20296 26140 20360 26144
rect 20296 26084 20300 26140
rect 20300 26084 20356 26140
rect 20356 26084 20360 26140
rect 20296 26080 20360 26084
rect 20376 26140 20440 26144
rect 20376 26084 20380 26140
rect 20380 26084 20436 26140
rect 20436 26084 20440 26140
rect 20376 26080 20440 26084
rect 20456 26140 20520 26144
rect 20456 26084 20460 26140
rect 20460 26084 20516 26140
rect 20516 26084 20520 26140
rect 20456 26080 20520 26084
rect 39480 26140 39544 26144
rect 39480 26084 39484 26140
rect 39484 26084 39540 26140
rect 39540 26084 39544 26140
rect 39480 26080 39544 26084
rect 39560 26140 39624 26144
rect 39560 26084 39564 26140
rect 39564 26084 39620 26140
rect 39620 26084 39624 26140
rect 39560 26080 39624 26084
rect 39640 26140 39704 26144
rect 39640 26084 39644 26140
rect 39644 26084 39700 26140
rect 39700 26084 39704 26140
rect 39640 26080 39704 26084
rect 39720 26140 39784 26144
rect 39720 26084 39724 26140
rect 39724 26084 39780 26140
rect 39780 26084 39784 26140
rect 39720 26080 39784 26084
rect 17908 25876 17972 25940
rect 19012 25604 19076 25668
rect 10584 25596 10648 25600
rect 10584 25540 10588 25596
rect 10588 25540 10644 25596
rect 10644 25540 10648 25596
rect 10584 25536 10648 25540
rect 10664 25596 10728 25600
rect 10664 25540 10668 25596
rect 10668 25540 10724 25596
rect 10724 25540 10728 25596
rect 10664 25536 10728 25540
rect 10744 25596 10808 25600
rect 10744 25540 10748 25596
rect 10748 25540 10804 25596
rect 10804 25540 10808 25596
rect 10744 25536 10808 25540
rect 10824 25596 10888 25600
rect 10824 25540 10828 25596
rect 10828 25540 10884 25596
rect 10884 25540 10888 25596
rect 10824 25536 10888 25540
rect 29848 25596 29912 25600
rect 29848 25540 29852 25596
rect 29852 25540 29908 25596
rect 29908 25540 29912 25596
rect 29848 25536 29912 25540
rect 29928 25596 29992 25600
rect 29928 25540 29932 25596
rect 29932 25540 29988 25596
rect 29988 25540 29992 25596
rect 29928 25536 29992 25540
rect 30008 25596 30072 25600
rect 30008 25540 30012 25596
rect 30012 25540 30068 25596
rect 30068 25540 30072 25596
rect 30008 25536 30072 25540
rect 30088 25596 30152 25600
rect 30088 25540 30092 25596
rect 30092 25540 30148 25596
rect 30148 25540 30152 25596
rect 30088 25536 30152 25540
rect 49112 25596 49176 25600
rect 49112 25540 49116 25596
rect 49116 25540 49172 25596
rect 49172 25540 49176 25596
rect 49112 25536 49176 25540
rect 49192 25596 49256 25600
rect 49192 25540 49196 25596
rect 49196 25540 49252 25596
rect 49252 25540 49256 25596
rect 49192 25536 49256 25540
rect 49272 25596 49336 25600
rect 49272 25540 49276 25596
rect 49276 25540 49332 25596
rect 49332 25540 49336 25596
rect 49272 25536 49336 25540
rect 49352 25596 49416 25600
rect 49352 25540 49356 25596
rect 49356 25540 49412 25596
rect 49412 25540 49416 25596
rect 49352 25536 49416 25540
rect 27476 25468 27540 25532
rect 28212 25332 28276 25396
rect 25268 25256 25332 25260
rect 25268 25200 25282 25256
rect 25282 25200 25332 25256
rect 25268 25196 25332 25200
rect 28396 25196 28460 25260
rect 29684 25196 29748 25260
rect 29316 25060 29380 25124
rect 20216 25052 20280 25056
rect 20216 24996 20220 25052
rect 20220 24996 20276 25052
rect 20276 24996 20280 25052
rect 20216 24992 20280 24996
rect 20296 25052 20360 25056
rect 20296 24996 20300 25052
rect 20300 24996 20356 25052
rect 20356 24996 20360 25052
rect 20296 24992 20360 24996
rect 20376 25052 20440 25056
rect 20376 24996 20380 25052
rect 20380 24996 20436 25052
rect 20436 24996 20440 25052
rect 20376 24992 20440 24996
rect 20456 25052 20520 25056
rect 20456 24996 20460 25052
rect 20460 24996 20516 25052
rect 20516 24996 20520 25052
rect 20456 24992 20520 24996
rect 39480 25052 39544 25056
rect 39480 24996 39484 25052
rect 39484 24996 39540 25052
rect 39540 24996 39544 25052
rect 39480 24992 39544 24996
rect 39560 25052 39624 25056
rect 39560 24996 39564 25052
rect 39564 24996 39620 25052
rect 39620 24996 39624 25052
rect 39560 24992 39624 24996
rect 39640 25052 39704 25056
rect 39640 24996 39644 25052
rect 39644 24996 39700 25052
rect 39700 24996 39704 25052
rect 39640 24992 39704 24996
rect 39720 25052 39784 25056
rect 39720 24996 39724 25052
rect 39724 24996 39780 25052
rect 39780 24996 39784 25052
rect 39720 24992 39784 24996
rect 34284 24984 34348 24988
rect 34284 24928 34334 24984
rect 34334 24928 34348 24984
rect 34284 24924 34348 24928
rect 28764 24516 28828 24580
rect 10584 24508 10648 24512
rect 10584 24452 10588 24508
rect 10588 24452 10644 24508
rect 10644 24452 10648 24508
rect 10584 24448 10648 24452
rect 10664 24508 10728 24512
rect 10664 24452 10668 24508
rect 10668 24452 10724 24508
rect 10724 24452 10728 24508
rect 10664 24448 10728 24452
rect 10744 24508 10808 24512
rect 10744 24452 10748 24508
rect 10748 24452 10804 24508
rect 10804 24452 10808 24508
rect 10744 24448 10808 24452
rect 10824 24508 10888 24512
rect 10824 24452 10828 24508
rect 10828 24452 10884 24508
rect 10884 24452 10888 24508
rect 10824 24448 10888 24452
rect 29848 24508 29912 24512
rect 29848 24452 29852 24508
rect 29852 24452 29908 24508
rect 29908 24452 29912 24508
rect 29848 24448 29912 24452
rect 29928 24508 29992 24512
rect 29928 24452 29932 24508
rect 29932 24452 29988 24508
rect 29988 24452 29992 24508
rect 29928 24448 29992 24452
rect 30008 24508 30072 24512
rect 30008 24452 30012 24508
rect 30012 24452 30068 24508
rect 30068 24452 30072 24508
rect 30008 24448 30072 24452
rect 30088 24508 30152 24512
rect 30088 24452 30092 24508
rect 30092 24452 30148 24508
rect 30148 24452 30152 24508
rect 30088 24448 30152 24452
rect 29316 24380 29380 24444
rect 37964 24652 38028 24716
rect 33364 24516 33428 24580
rect 36676 24516 36740 24580
rect 49112 24508 49176 24512
rect 49112 24452 49116 24508
rect 49116 24452 49172 24508
rect 49172 24452 49176 24508
rect 49112 24448 49176 24452
rect 49192 24508 49256 24512
rect 49192 24452 49196 24508
rect 49196 24452 49252 24508
rect 49252 24452 49256 24508
rect 49192 24448 49256 24452
rect 49272 24508 49336 24512
rect 49272 24452 49276 24508
rect 49276 24452 49332 24508
rect 49332 24452 49336 24508
rect 49272 24448 49336 24452
rect 49352 24508 49416 24512
rect 49352 24452 49356 24508
rect 49356 24452 49412 24508
rect 49412 24452 49416 24508
rect 49352 24448 49416 24452
rect 28580 24108 28644 24172
rect 41092 24108 41156 24172
rect 25820 23972 25884 24036
rect 27292 24032 27356 24036
rect 27292 23976 27342 24032
rect 27342 23976 27356 24032
rect 27292 23972 27356 23976
rect 20216 23964 20280 23968
rect 20216 23908 20220 23964
rect 20220 23908 20276 23964
rect 20276 23908 20280 23964
rect 20216 23904 20280 23908
rect 20296 23964 20360 23968
rect 20296 23908 20300 23964
rect 20300 23908 20356 23964
rect 20356 23908 20360 23964
rect 20296 23904 20360 23908
rect 20376 23964 20440 23968
rect 20376 23908 20380 23964
rect 20380 23908 20436 23964
rect 20436 23908 20440 23964
rect 20376 23904 20440 23908
rect 20456 23964 20520 23968
rect 20456 23908 20460 23964
rect 20460 23908 20516 23964
rect 20516 23908 20520 23964
rect 20456 23904 20520 23908
rect 39480 23964 39544 23968
rect 39480 23908 39484 23964
rect 39484 23908 39540 23964
rect 39540 23908 39544 23964
rect 39480 23904 39544 23908
rect 39560 23964 39624 23968
rect 39560 23908 39564 23964
rect 39564 23908 39620 23964
rect 39620 23908 39624 23964
rect 39560 23904 39624 23908
rect 39640 23964 39704 23968
rect 39640 23908 39644 23964
rect 39644 23908 39700 23964
rect 39700 23908 39704 23964
rect 39640 23904 39704 23908
rect 39720 23964 39784 23968
rect 39720 23908 39724 23964
rect 39724 23908 39780 23964
rect 39780 23908 39784 23964
rect 39720 23904 39784 23908
rect 28028 23836 28092 23900
rect 32996 23896 33060 23900
rect 32996 23840 33010 23896
rect 33010 23840 33060 23896
rect 32996 23836 33060 23840
rect 34836 23836 34900 23900
rect 24900 23700 24964 23764
rect 27108 23700 27172 23764
rect 30420 23564 30484 23628
rect 30972 23564 31036 23628
rect 35756 23624 35820 23628
rect 35756 23568 35770 23624
rect 35770 23568 35820 23624
rect 22324 23428 22388 23492
rect 24716 23428 24780 23492
rect 35756 23564 35820 23568
rect 33180 23488 33244 23492
rect 33180 23432 33194 23488
rect 33194 23432 33244 23488
rect 33180 23428 33244 23432
rect 37228 23428 37292 23492
rect 10584 23420 10648 23424
rect 10584 23364 10588 23420
rect 10588 23364 10644 23420
rect 10644 23364 10648 23420
rect 10584 23360 10648 23364
rect 10664 23420 10728 23424
rect 10664 23364 10668 23420
rect 10668 23364 10724 23420
rect 10724 23364 10728 23420
rect 10664 23360 10728 23364
rect 10744 23420 10808 23424
rect 10744 23364 10748 23420
rect 10748 23364 10804 23420
rect 10804 23364 10808 23420
rect 10744 23360 10808 23364
rect 10824 23420 10888 23424
rect 10824 23364 10828 23420
rect 10828 23364 10884 23420
rect 10884 23364 10888 23420
rect 10824 23360 10888 23364
rect 29848 23420 29912 23424
rect 29848 23364 29852 23420
rect 29852 23364 29908 23420
rect 29908 23364 29912 23420
rect 29848 23360 29912 23364
rect 29928 23420 29992 23424
rect 29928 23364 29932 23420
rect 29932 23364 29988 23420
rect 29988 23364 29992 23420
rect 29928 23360 29992 23364
rect 30008 23420 30072 23424
rect 30008 23364 30012 23420
rect 30012 23364 30068 23420
rect 30068 23364 30072 23420
rect 30008 23360 30072 23364
rect 30088 23420 30152 23424
rect 30088 23364 30092 23420
rect 30092 23364 30148 23420
rect 30148 23364 30152 23420
rect 30088 23360 30152 23364
rect 49112 23420 49176 23424
rect 49112 23364 49116 23420
rect 49116 23364 49172 23420
rect 49172 23364 49176 23420
rect 49112 23360 49176 23364
rect 49192 23420 49256 23424
rect 49192 23364 49196 23420
rect 49196 23364 49252 23420
rect 49252 23364 49256 23420
rect 49192 23360 49256 23364
rect 49272 23420 49336 23424
rect 49272 23364 49276 23420
rect 49276 23364 49332 23420
rect 49332 23364 49336 23420
rect 49272 23360 49336 23364
rect 49352 23420 49416 23424
rect 49352 23364 49356 23420
rect 49356 23364 49412 23420
rect 49412 23364 49416 23420
rect 49352 23360 49416 23364
rect 19564 23156 19628 23220
rect 21404 23020 21468 23084
rect 27844 23020 27908 23084
rect 30604 23020 30668 23084
rect 38884 22884 38948 22948
rect 20216 22876 20280 22880
rect 20216 22820 20220 22876
rect 20220 22820 20276 22876
rect 20276 22820 20280 22876
rect 20216 22816 20280 22820
rect 20296 22876 20360 22880
rect 20296 22820 20300 22876
rect 20300 22820 20356 22876
rect 20356 22820 20360 22876
rect 20296 22816 20360 22820
rect 20376 22876 20440 22880
rect 20376 22820 20380 22876
rect 20380 22820 20436 22876
rect 20436 22820 20440 22876
rect 20376 22816 20440 22820
rect 20456 22876 20520 22880
rect 20456 22820 20460 22876
rect 20460 22820 20516 22876
rect 20516 22820 20520 22876
rect 20456 22816 20520 22820
rect 39480 22876 39544 22880
rect 39480 22820 39484 22876
rect 39484 22820 39540 22876
rect 39540 22820 39544 22876
rect 39480 22816 39544 22820
rect 39560 22876 39624 22880
rect 39560 22820 39564 22876
rect 39564 22820 39620 22876
rect 39620 22820 39624 22876
rect 39560 22816 39624 22820
rect 39640 22876 39704 22880
rect 39640 22820 39644 22876
rect 39644 22820 39700 22876
rect 39700 22820 39704 22876
rect 39640 22816 39704 22820
rect 39720 22876 39784 22880
rect 39720 22820 39724 22876
rect 39724 22820 39780 22876
rect 39780 22820 39784 22876
rect 39720 22816 39784 22820
rect 28396 22748 28460 22812
rect 25820 22672 25884 22676
rect 25820 22616 25834 22672
rect 25834 22616 25884 22672
rect 25820 22612 25884 22616
rect 28580 22612 28644 22676
rect 29132 22612 29196 22676
rect 24164 22536 24228 22540
rect 24164 22480 24178 22536
rect 24178 22480 24228 22536
rect 24164 22476 24228 22480
rect 25084 22476 25148 22540
rect 21588 22340 21652 22404
rect 24348 22340 24412 22404
rect 34652 22476 34716 22540
rect 29316 22400 29380 22404
rect 29316 22344 29330 22400
rect 29330 22344 29380 22400
rect 10584 22332 10648 22336
rect 10584 22276 10588 22332
rect 10588 22276 10644 22332
rect 10644 22276 10648 22332
rect 10584 22272 10648 22276
rect 10664 22332 10728 22336
rect 10664 22276 10668 22332
rect 10668 22276 10724 22332
rect 10724 22276 10728 22332
rect 10664 22272 10728 22276
rect 10744 22332 10808 22336
rect 10744 22276 10748 22332
rect 10748 22276 10804 22332
rect 10804 22276 10808 22332
rect 10744 22272 10808 22276
rect 10824 22332 10888 22336
rect 10824 22276 10828 22332
rect 10828 22276 10884 22332
rect 10884 22276 10888 22332
rect 10824 22272 10888 22276
rect 20668 22204 20732 22268
rect 19932 22128 19996 22132
rect 29316 22340 29380 22344
rect 34468 22340 34532 22404
rect 29848 22332 29912 22336
rect 29848 22276 29852 22332
rect 29852 22276 29908 22332
rect 29908 22276 29912 22332
rect 29848 22272 29912 22276
rect 29928 22332 29992 22336
rect 29928 22276 29932 22332
rect 29932 22276 29988 22332
rect 29988 22276 29992 22332
rect 29928 22272 29992 22276
rect 30008 22332 30072 22336
rect 30008 22276 30012 22332
rect 30012 22276 30068 22332
rect 30068 22276 30072 22332
rect 30008 22272 30072 22276
rect 30088 22332 30152 22336
rect 30088 22276 30092 22332
rect 30092 22276 30148 22332
rect 30148 22276 30152 22332
rect 30088 22272 30152 22276
rect 29500 22204 29564 22268
rect 37044 22204 37108 22268
rect 49112 22332 49176 22336
rect 49112 22276 49116 22332
rect 49116 22276 49172 22332
rect 49172 22276 49176 22332
rect 49112 22272 49176 22276
rect 49192 22332 49256 22336
rect 49192 22276 49196 22332
rect 49196 22276 49252 22332
rect 49252 22276 49256 22332
rect 49192 22272 49256 22276
rect 49272 22332 49336 22336
rect 49272 22276 49276 22332
rect 49276 22276 49332 22332
rect 49332 22276 49336 22332
rect 49272 22272 49336 22276
rect 49352 22332 49416 22336
rect 49352 22276 49356 22332
rect 49356 22276 49412 22332
rect 49412 22276 49416 22332
rect 49352 22272 49416 22276
rect 19932 22072 19946 22128
rect 19946 22072 19996 22128
rect 19932 22068 19996 22072
rect 29132 21932 29196 21996
rect 33732 21992 33796 21996
rect 33732 21936 33746 21992
rect 33746 21936 33796 21992
rect 33732 21932 33796 21936
rect 37780 22068 37844 22132
rect 37596 21932 37660 21996
rect 21772 21796 21836 21860
rect 20216 21788 20280 21792
rect 20216 21732 20220 21788
rect 20220 21732 20276 21788
rect 20276 21732 20280 21788
rect 20216 21728 20280 21732
rect 20296 21788 20360 21792
rect 20296 21732 20300 21788
rect 20300 21732 20356 21788
rect 20356 21732 20360 21788
rect 20296 21728 20360 21732
rect 20376 21788 20440 21792
rect 20376 21732 20380 21788
rect 20380 21732 20436 21788
rect 20436 21732 20440 21788
rect 20376 21728 20440 21732
rect 20456 21788 20520 21792
rect 20456 21732 20460 21788
rect 20460 21732 20516 21788
rect 20516 21732 20520 21788
rect 20456 21728 20520 21732
rect 24348 21660 24412 21724
rect 24900 21796 24964 21860
rect 39480 21788 39544 21792
rect 39480 21732 39484 21788
rect 39484 21732 39540 21788
rect 39540 21732 39544 21788
rect 39480 21728 39544 21732
rect 39560 21788 39624 21792
rect 39560 21732 39564 21788
rect 39564 21732 39620 21788
rect 39620 21732 39624 21788
rect 39560 21728 39624 21732
rect 39640 21788 39704 21792
rect 39640 21732 39644 21788
rect 39644 21732 39700 21788
rect 39700 21732 39704 21788
rect 39640 21728 39704 21732
rect 39720 21788 39784 21792
rect 39720 21732 39724 21788
rect 39724 21732 39780 21788
rect 39780 21732 39784 21788
rect 39720 21728 39784 21732
rect 27844 21720 27908 21724
rect 27844 21664 27894 21720
rect 27894 21664 27908 21720
rect 27844 21660 27908 21664
rect 30972 21660 31036 21724
rect 33364 21660 33428 21724
rect 22692 21524 22756 21588
rect 26556 21524 26620 21588
rect 27476 21524 27540 21588
rect 18276 21388 18340 21452
rect 29500 21388 29564 21452
rect 30788 21252 30852 21316
rect 35572 21388 35636 21452
rect 37964 21252 38028 21316
rect 10584 21244 10648 21248
rect 10584 21188 10588 21244
rect 10588 21188 10644 21244
rect 10644 21188 10648 21244
rect 10584 21184 10648 21188
rect 10664 21244 10728 21248
rect 10664 21188 10668 21244
rect 10668 21188 10724 21244
rect 10724 21188 10728 21244
rect 10664 21184 10728 21188
rect 10744 21244 10808 21248
rect 10744 21188 10748 21244
rect 10748 21188 10804 21244
rect 10804 21188 10808 21244
rect 10744 21184 10808 21188
rect 10824 21244 10888 21248
rect 10824 21188 10828 21244
rect 10828 21188 10884 21244
rect 10884 21188 10888 21244
rect 10824 21184 10888 21188
rect 29848 21244 29912 21248
rect 29848 21188 29852 21244
rect 29852 21188 29908 21244
rect 29908 21188 29912 21244
rect 29848 21184 29912 21188
rect 29928 21244 29992 21248
rect 29928 21188 29932 21244
rect 29932 21188 29988 21244
rect 29988 21188 29992 21244
rect 29928 21184 29992 21188
rect 30008 21244 30072 21248
rect 30008 21188 30012 21244
rect 30012 21188 30068 21244
rect 30068 21188 30072 21244
rect 30008 21184 30072 21188
rect 30088 21244 30152 21248
rect 30088 21188 30092 21244
rect 30092 21188 30148 21244
rect 30148 21188 30152 21244
rect 30088 21184 30152 21188
rect 49112 21244 49176 21248
rect 49112 21188 49116 21244
rect 49116 21188 49172 21244
rect 49172 21188 49176 21244
rect 49112 21184 49176 21188
rect 49192 21244 49256 21248
rect 49192 21188 49196 21244
rect 49196 21188 49252 21244
rect 49252 21188 49256 21244
rect 49192 21184 49256 21188
rect 49272 21244 49336 21248
rect 49272 21188 49276 21244
rect 49276 21188 49332 21244
rect 49332 21188 49336 21244
rect 49272 21184 49336 21188
rect 49352 21244 49416 21248
rect 49352 21188 49356 21244
rect 49356 21188 49412 21244
rect 49412 21188 49416 21244
rect 49352 21184 49416 21188
rect 42012 21176 42076 21180
rect 42012 21120 42062 21176
rect 42062 21120 42076 21176
rect 42012 21116 42076 21120
rect 22692 20708 22756 20772
rect 30788 20708 30852 20772
rect 32260 20768 32324 20772
rect 32260 20712 32310 20768
rect 32310 20712 32324 20768
rect 32260 20708 32324 20712
rect 36860 20708 36924 20772
rect 20216 20700 20280 20704
rect 20216 20644 20220 20700
rect 20220 20644 20276 20700
rect 20276 20644 20280 20700
rect 20216 20640 20280 20644
rect 20296 20700 20360 20704
rect 20296 20644 20300 20700
rect 20300 20644 20356 20700
rect 20356 20644 20360 20700
rect 20296 20640 20360 20644
rect 20376 20700 20440 20704
rect 20376 20644 20380 20700
rect 20380 20644 20436 20700
rect 20436 20644 20440 20700
rect 20376 20640 20440 20644
rect 20456 20700 20520 20704
rect 20456 20644 20460 20700
rect 20460 20644 20516 20700
rect 20516 20644 20520 20700
rect 20456 20640 20520 20644
rect 39480 20700 39544 20704
rect 39480 20644 39484 20700
rect 39484 20644 39540 20700
rect 39540 20644 39544 20700
rect 39480 20640 39544 20644
rect 39560 20700 39624 20704
rect 39560 20644 39564 20700
rect 39564 20644 39620 20700
rect 39620 20644 39624 20700
rect 39560 20640 39624 20644
rect 39640 20700 39704 20704
rect 39640 20644 39644 20700
rect 39644 20644 39700 20700
rect 39700 20644 39704 20700
rect 39640 20640 39704 20644
rect 39720 20700 39784 20704
rect 39720 20644 39724 20700
rect 39724 20644 39780 20700
rect 39780 20644 39784 20700
rect 39720 20640 39784 20644
rect 19196 20436 19260 20500
rect 20668 20436 20732 20500
rect 27108 20436 27172 20500
rect 28396 20300 28460 20364
rect 10584 20156 10648 20160
rect 10584 20100 10588 20156
rect 10588 20100 10644 20156
rect 10644 20100 10648 20156
rect 10584 20096 10648 20100
rect 10664 20156 10728 20160
rect 10664 20100 10668 20156
rect 10668 20100 10724 20156
rect 10724 20100 10728 20156
rect 10664 20096 10728 20100
rect 10744 20156 10808 20160
rect 10744 20100 10748 20156
rect 10748 20100 10804 20156
rect 10804 20100 10808 20156
rect 10744 20096 10808 20100
rect 10824 20156 10888 20160
rect 10824 20100 10828 20156
rect 10828 20100 10884 20156
rect 10884 20100 10888 20156
rect 10824 20096 10888 20100
rect 29848 20156 29912 20160
rect 29848 20100 29852 20156
rect 29852 20100 29908 20156
rect 29908 20100 29912 20156
rect 29848 20096 29912 20100
rect 29928 20156 29992 20160
rect 29928 20100 29932 20156
rect 29932 20100 29988 20156
rect 29988 20100 29992 20156
rect 29928 20096 29992 20100
rect 30008 20156 30072 20160
rect 30008 20100 30012 20156
rect 30012 20100 30068 20156
rect 30068 20100 30072 20156
rect 30008 20096 30072 20100
rect 30088 20156 30152 20160
rect 30088 20100 30092 20156
rect 30092 20100 30148 20156
rect 30148 20100 30152 20156
rect 30088 20096 30152 20100
rect 20852 20028 20916 20092
rect 21220 20088 21284 20092
rect 21220 20032 21234 20088
rect 21234 20032 21284 20088
rect 21220 20028 21284 20032
rect 35940 20164 36004 20228
rect 49112 20156 49176 20160
rect 49112 20100 49116 20156
rect 49116 20100 49172 20156
rect 49172 20100 49176 20156
rect 49112 20096 49176 20100
rect 49192 20156 49256 20160
rect 49192 20100 49196 20156
rect 49196 20100 49252 20156
rect 49252 20100 49256 20156
rect 49192 20096 49256 20100
rect 49272 20156 49336 20160
rect 49272 20100 49276 20156
rect 49276 20100 49332 20156
rect 49332 20100 49336 20156
rect 49272 20096 49336 20100
rect 49352 20156 49416 20160
rect 49352 20100 49356 20156
rect 49356 20100 49412 20156
rect 49412 20100 49416 20156
rect 49352 20096 49416 20100
rect 34284 20028 34348 20092
rect 21036 19892 21100 19956
rect 22508 19892 22572 19956
rect 28764 19892 28828 19956
rect 18644 19756 18708 19820
rect 18828 19484 18892 19548
rect 18644 19348 18708 19412
rect 27844 19756 27908 19820
rect 27108 19680 27172 19684
rect 27108 19624 27158 19680
rect 27158 19624 27172 19680
rect 27108 19620 27172 19624
rect 34652 19620 34716 19684
rect 20216 19612 20280 19616
rect 20216 19556 20220 19612
rect 20220 19556 20276 19612
rect 20276 19556 20280 19612
rect 20216 19552 20280 19556
rect 20296 19612 20360 19616
rect 20296 19556 20300 19612
rect 20300 19556 20356 19612
rect 20356 19556 20360 19612
rect 20296 19552 20360 19556
rect 20376 19612 20440 19616
rect 20376 19556 20380 19612
rect 20380 19556 20436 19612
rect 20436 19556 20440 19612
rect 20376 19552 20440 19556
rect 20456 19612 20520 19616
rect 20456 19556 20460 19612
rect 20460 19556 20516 19612
rect 20516 19556 20520 19612
rect 20456 19552 20520 19556
rect 39480 19612 39544 19616
rect 39480 19556 39484 19612
rect 39484 19556 39540 19612
rect 39540 19556 39544 19612
rect 39480 19552 39544 19556
rect 39560 19612 39624 19616
rect 39560 19556 39564 19612
rect 39564 19556 39620 19612
rect 39620 19556 39624 19612
rect 39560 19552 39624 19556
rect 39640 19612 39704 19616
rect 39640 19556 39644 19612
rect 39644 19556 39700 19612
rect 39700 19556 39704 19612
rect 39640 19552 39704 19556
rect 39720 19612 39784 19616
rect 39720 19556 39724 19612
rect 39724 19556 39780 19612
rect 39780 19556 39784 19612
rect 39720 19552 39784 19556
rect 20668 19484 20732 19548
rect 22140 19408 22204 19412
rect 27108 19484 27172 19548
rect 29500 19484 29564 19548
rect 22140 19352 22190 19408
rect 22190 19352 22204 19408
rect 22140 19348 22204 19352
rect 27292 19348 27356 19412
rect 28028 19348 28092 19412
rect 36676 19484 36740 19548
rect 40908 19408 40972 19412
rect 40908 19352 40958 19408
rect 40958 19352 40972 19408
rect 40908 19348 40972 19352
rect 41644 19408 41708 19412
rect 41644 19352 41658 19408
rect 41658 19352 41708 19408
rect 41644 19348 41708 19352
rect 42748 19408 42812 19412
rect 42748 19352 42762 19408
rect 42762 19352 42812 19408
rect 42748 19348 42812 19352
rect 16804 19272 16868 19276
rect 16804 19216 16818 19272
rect 16818 19216 16868 19272
rect 16804 19212 16868 19216
rect 17172 19212 17236 19276
rect 18092 19212 18156 19276
rect 19932 19212 19996 19276
rect 20852 19212 20916 19276
rect 25268 19212 25332 19276
rect 19012 19076 19076 19140
rect 19196 19076 19260 19140
rect 10584 19068 10648 19072
rect 10584 19012 10588 19068
rect 10588 19012 10644 19068
rect 10644 19012 10648 19068
rect 10584 19008 10648 19012
rect 10664 19068 10728 19072
rect 10664 19012 10668 19068
rect 10668 19012 10724 19068
rect 10724 19012 10728 19068
rect 10664 19008 10728 19012
rect 10744 19068 10808 19072
rect 10744 19012 10748 19068
rect 10748 19012 10804 19068
rect 10804 19012 10808 19068
rect 10744 19008 10808 19012
rect 10824 19068 10888 19072
rect 10824 19012 10828 19068
rect 10828 19012 10884 19068
rect 10884 19012 10888 19068
rect 10824 19008 10888 19012
rect 17908 18940 17972 19004
rect 18276 18940 18340 19004
rect 25084 19076 25148 19140
rect 29500 19076 29564 19140
rect 33732 19212 33796 19276
rect 37412 19212 37476 19276
rect 38700 19272 38764 19276
rect 38700 19216 38714 19272
rect 38714 19216 38764 19272
rect 38700 19212 38764 19216
rect 29848 19068 29912 19072
rect 29848 19012 29852 19068
rect 29852 19012 29908 19068
rect 29908 19012 29912 19068
rect 29848 19008 29912 19012
rect 29928 19068 29992 19072
rect 29928 19012 29932 19068
rect 29932 19012 29988 19068
rect 29988 19012 29992 19068
rect 29928 19008 29992 19012
rect 30008 19068 30072 19072
rect 30008 19012 30012 19068
rect 30012 19012 30068 19068
rect 30068 19012 30072 19068
rect 30008 19008 30072 19012
rect 30088 19068 30152 19072
rect 30088 19012 30092 19068
rect 30092 19012 30148 19068
rect 30148 19012 30152 19068
rect 30088 19008 30152 19012
rect 49112 19068 49176 19072
rect 49112 19012 49116 19068
rect 49116 19012 49172 19068
rect 49172 19012 49176 19068
rect 49112 19008 49176 19012
rect 49192 19068 49256 19072
rect 49192 19012 49196 19068
rect 49196 19012 49252 19068
rect 49252 19012 49256 19068
rect 49192 19008 49256 19012
rect 49272 19068 49336 19072
rect 49272 19012 49276 19068
rect 49276 19012 49332 19068
rect 49332 19012 49336 19068
rect 49272 19008 49336 19012
rect 49352 19068 49416 19072
rect 49352 19012 49356 19068
rect 49356 19012 49412 19068
rect 49412 19012 49416 19068
rect 49352 19008 49416 19012
rect 30604 18940 30668 19004
rect 29684 18804 29748 18868
rect 16436 18532 16500 18596
rect 19380 18592 19444 18596
rect 19380 18536 19430 18592
rect 19430 18536 19444 18592
rect 19380 18532 19444 18536
rect 20852 18532 20916 18596
rect 34100 18668 34164 18732
rect 20216 18524 20280 18528
rect 20216 18468 20220 18524
rect 20220 18468 20276 18524
rect 20276 18468 20280 18524
rect 20216 18464 20280 18468
rect 20296 18524 20360 18528
rect 20296 18468 20300 18524
rect 20300 18468 20356 18524
rect 20356 18468 20360 18524
rect 20296 18464 20360 18468
rect 20376 18524 20440 18528
rect 20376 18468 20380 18524
rect 20380 18468 20436 18524
rect 20436 18468 20440 18524
rect 20376 18464 20440 18468
rect 20456 18524 20520 18528
rect 20456 18468 20460 18524
rect 20460 18468 20516 18524
rect 20516 18468 20520 18524
rect 20456 18464 20520 18468
rect 39480 18524 39544 18528
rect 39480 18468 39484 18524
rect 39484 18468 39540 18524
rect 39540 18468 39544 18524
rect 39480 18464 39544 18468
rect 39560 18524 39624 18528
rect 39560 18468 39564 18524
rect 39564 18468 39620 18524
rect 39620 18468 39624 18524
rect 39560 18464 39624 18468
rect 39640 18524 39704 18528
rect 39640 18468 39644 18524
rect 39644 18468 39700 18524
rect 39700 18468 39704 18524
rect 39640 18464 39704 18468
rect 39720 18524 39784 18528
rect 39720 18468 39724 18524
rect 39724 18468 39780 18524
rect 39780 18468 39784 18524
rect 39720 18464 39784 18468
rect 32628 18396 32692 18460
rect 34652 18456 34716 18460
rect 34652 18400 34702 18456
rect 34702 18400 34716 18456
rect 34652 18396 34716 18400
rect 33180 18260 33244 18324
rect 35572 18124 35636 18188
rect 10584 17980 10648 17984
rect 10584 17924 10588 17980
rect 10588 17924 10644 17980
rect 10644 17924 10648 17980
rect 10584 17920 10648 17924
rect 10664 17980 10728 17984
rect 10664 17924 10668 17980
rect 10668 17924 10724 17980
rect 10724 17924 10728 17980
rect 10664 17920 10728 17924
rect 10744 17980 10808 17984
rect 10744 17924 10748 17980
rect 10748 17924 10804 17980
rect 10804 17924 10808 17980
rect 10744 17920 10808 17924
rect 10824 17980 10888 17984
rect 10824 17924 10828 17980
rect 10828 17924 10884 17980
rect 10884 17924 10888 17980
rect 10824 17920 10888 17924
rect 17540 17852 17604 17916
rect 21956 17852 22020 17916
rect 29684 17988 29748 18052
rect 29848 17980 29912 17984
rect 29848 17924 29852 17980
rect 29852 17924 29908 17980
rect 29908 17924 29912 17980
rect 29848 17920 29912 17924
rect 29928 17980 29992 17984
rect 29928 17924 29932 17980
rect 29932 17924 29988 17980
rect 29988 17924 29992 17980
rect 29928 17920 29992 17924
rect 30008 17980 30072 17984
rect 30008 17924 30012 17980
rect 30012 17924 30068 17980
rect 30068 17924 30072 17980
rect 30008 17920 30072 17924
rect 30088 17980 30152 17984
rect 30088 17924 30092 17980
rect 30092 17924 30148 17980
rect 30148 17924 30152 17980
rect 30088 17920 30152 17924
rect 49112 17980 49176 17984
rect 49112 17924 49116 17980
rect 49116 17924 49172 17980
rect 49172 17924 49176 17980
rect 49112 17920 49176 17924
rect 49192 17980 49256 17984
rect 49192 17924 49196 17980
rect 49196 17924 49252 17980
rect 49252 17924 49256 17980
rect 49192 17920 49256 17924
rect 49272 17980 49336 17984
rect 49272 17924 49276 17980
rect 49276 17924 49332 17980
rect 49332 17924 49336 17980
rect 49272 17920 49336 17924
rect 49352 17980 49416 17984
rect 49352 17924 49356 17980
rect 49356 17924 49412 17980
rect 49412 17924 49416 17980
rect 49352 17920 49416 17924
rect 24716 17912 24780 17916
rect 24716 17856 24730 17912
rect 24730 17856 24780 17912
rect 24716 17852 24780 17856
rect 21220 17716 21284 17780
rect 45140 17912 45204 17916
rect 45140 17856 45154 17912
rect 45154 17856 45204 17912
rect 45140 17852 45204 17856
rect 18092 17580 18156 17644
rect 20216 17436 20280 17440
rect 20216 17380 20220 17436
rect 20220 17380 20276 17436
rect 20276 17380 20280 17436
rect 20216 17376 20280 17380
rect 20296 17436 20360 17440
rect 20296 17380 20300 17436
rect 20300 17380 20356 17436
rect 20356 17380 20360 17436
rect 20296 17376 20360 17380
rect 20376 17436 20440 17440
rect 20376 17380 20380 17436
rect 20380 17380 20436 17436
rect 20436 17380 20440 17436
rect 20376 17376 20440 17380
rect 20456 17436 20520 17440
rect 20456 17380 20460 17436
rect 20460 17380 20516 17436
rect 20516 17380 20520 17436
rect 20456 17376 20520 17380
rect 39480 17436 39544 17440
rect 39480 17380 39484 17436
rect 39484 17380 39540 17436
rect 39540 17380 39544 17436
rect 39480 17376 39544 17380
rect 39560 17436 39624 17440
rect 39560 17380 39564 17436
rect 39564 17380 39620 17436
rect 39620 17380 39624 17436
rect 39560 17376 39624 17380
rect 39640 17436 39704 17440
rect 39640 17380 39644 17436
rect 39644 17380 39700 17436
rect 39700 17380 39704 17436
rect 39640 17376 39704 17380
rect 39720 17436 39784 17440
rect 39720 17380 39724 17436
rect 39724 17380 39780 17436
rect 39780 17380 39784 17436
rect 39720 17376 39784 17380
rect 41092 17368 41156 17372
rect 41092 17312 41142 17368
rect 41142 17312 41156 17368
rect 20852 17172 20916 17236
rect 41092 17308 41156 17312
rect 46060 17308 46124 17372
rect 36860 17172 36924 17236
rect 37228 17172 37292 17236
rect 37780 17172 37844 17236
rect 32444 16900 32508 16964
rect 37044 16900 37108 16964
rect 10584 16892 10648 16896
rect 10584 16836 10588 16892
rect 10588 16836 10644 16892
rect 10644 16836 10648 16892
rect 10584 16832 10648 16836
rect 10664 16892 10728 16896
rect 10664 16836 10668 16892
rect 10668 16836 10724 16892
rect 10724 16836 10728 16892
rect 10664 16832 10728 16836
rect 10744 16892 10808 16896
rect 10744 16836 10748 16892
rect 10748 16836 10804 16892
rect 10804 16836 10808 16892
rect 10744 16832 10808 16836
rect 10824 16892 10888 16896
rect 10824 16836 10828 16892
rect 10828 16836 10884 16892
rect 10884 16836 10888 16892
rect 10824 16832 10888 16836
rect 29848 16892 29912 16896
rect 29848 16836 29852 16892
rect 29852 16836 29908 16892
rect 29908 16836 29912 16892
rect 29848 16832 29912 16836
rect 29928 16892 29992 16896
rect 29928 16836 29932 16892
rect 29932 16836 29988 16892
rect 29988 16836 29992 16892
rect 29928 16832 29992 16836
rect 30008 16892 30072 16896
rect 30008 16836 30012 16892
rect 30012 16836 30068 16892
rect 30068 16836 30072 16892
rect 30008 16832 30072 16836
rect 30088 16892 30152 16896
rect 30088 16836 30092 16892
rect 30092 16836 30148 16892
rect 30148 16836 30152 16892
rect 30088 16832 30152 16836
rect 15332 16688 15396 16692
rect 15332 16632 15346 16688
rect 15346 16632 15396 16688
rect 15332 16628 15396 16632
rect 17540 16688 17604 16692
rect 17540 16632 17554 16688
rect 17554 16632 17604 16688
rect 17540 16628 17604 16632
rect 18828 16628 18892 16692
rect 19748 16628 19812 16692
rect 18460 16492 18524 16556
rect 19012 16492 19076 16556
rect 19932 16492 19996 16556
rect 26372 16628 26436 16692
rect 31892 16764 31956 16828
rect 34468 16764 34532 16828
rect 49112 16892 49176 16896
rect 49112 16836 49116 16892
rect 49116 16836 49172 16892
rect 49172 16836 49176 16892
rect 49112 16832 49176 16836
rect 49192 16892 49256 16896
rect 49192 16836 49196 16892
rect 49196 16836 49252 16892
rect 49252 16836 49256 16892
rect 49192 16832 49256 16836
rect 49272 16892 49336 16896
rect 49272 16836 49276 16892
rect 49276 16836 49332 16892
rect 49332 16836 49336 16892
rect 49272 16832 49336 16836
rect 49352 16892 49416 16896
rect 49352 16836 49356 16892
rect 49356 16836 49412 16892
rect 49412 16836 49416 16892
rect 49352 16832 49416 16836
rect 25452 16492 25516 16556
rect 26556 16492 26620 16556
rect 42196 16628 42260 16692
rect 46612 16628 46676 16692
rect 20216 16348 20280 16352
rect 20216 16292 20220 16348
rect 20220 16292 20276 16348
rect 20276 16292 20280 16348
rect 20216 16288 20280 16292
rect 20296 16348 20360 16352
rect 20296 16292 20300 16348
rect 20300 16292 20356 16348
rect 20356 16292 20360 16348
rect 20296 16288 20360 16292
rect 20376 16348 20440 16352
rect 20376 16292 20380 16348
rect 20380 16292 20436 16348
rect 20436 16292 20440 16348
rect 20376 16288 20440 16292
rect 20456 16348 20520 16352
rect 20456 16292 20460 16348
rect 20460 16292 20516 16348
rect 20516 16292 20520 16348
rect 20456 16288 20520 16292
rect 20852 16356 20916 16420
rect 22140 16220 22204 16284
rect 21036 16144 21100 16148
rect 21036 16088 21086 16144
rect 21086 16088 21100 16144
rect 21036 16084 21100 16088
rect 21588 16144 21652 16148
rect 21588 16088 21602 16144
rect 21602 16088 21652 16144
rect 21588 16084 21652 16088
rect 24532 16084 24596 16148
rect 28212 16356 28276 16420
rect 36124 16356 36188 16420
rect 39480 16348 39544 16352
rect 39480 16292 39484 16348
rect 39484 16292 39540 16348
rect 39540 16292 39544 16348
rect 39480 16288 39544 16292
rect 39560 16348 39624 16352
rect 39560 16292 39564 16348
rect 39564 16292 39620 16348
rect 39620 16292 39624 16348
rect 39560 16288 39624 16292
rect 39640 16348 39704 16352
rect 39640 16292 39644 16348
rect 39644 16292 39700 16348
rect 39700 16292 39704 16348
rect 39640 16288 39704 16292
rect 39720 16348 39784 16352
rect 39720 16292 39724 16348
rect 39724 16292 39780 16348
rect 39780 16292 39784 16348
rect 39720 16288 39784 16292
rect 38884 16220 38948 16284
rect 30972 16084 31036 16148
rect 32076 15948 32140 16012
rect 10584 15804 10648 15808
rect 10584 15748 10588 15804
rect 10588 15748 10644 15804
rect 10644 15748 10648 15804
rect 10584 15744 10648 15748
rect 10664 15804 10728 15808
rect 10664 15748 10668 15804
rect 10668 15748 10724 15804
rect 10724 15748 10728 15804
rect 10664 15744 10728 15748
rect 10744 15804 10808 15808
rect 10744 15748 10748 15804
rect 10748 15748 10804 15804
rect 10804 15748 10808 15804
rect 10744 15744 10808 15748
rect 10824 15804 10888 15808
rect 10824 15748 10828 15804
rect 10828 15748 10884 15804
rect 10884 15748 10888 15804
rect 10824 15744 10888 15748
rect 29500 15872 29564 15876
rect 29500 15816 29550 15872
rect 29550 15816 29564 15872
rect 29500 15812 29564 15816
rect 46060 15872 46124 15876
rect 46060 15816 46074 15872
rect 46074 15816 46124 15872
rect 29848 15804 29912 15808
rect 29848 15748 29852 15804
rect 29852 15748 29908 15804
rect 29908 15748 29912 15804
rect 29848 15744 29912 15748
rect 29928 15804 29992 15808
rect 29928 15748 29932 15804
rect 29932 15748 29988 15804
rect 29988 15748 29992 15804
rect 29928 15744 29992 15748
rect 30008 15804 30072 15808
rect 30008 15748 30012 15804
rect 30012 15748 30068 15804
rect 30068 15748 30072 15804
rect 30008 15744 30072 15748
rect 30088 15804 30152 15808
rect 30088 15748 30092 15804
rect 30092 15748 30148 15804
rect 30148 15748 30152 15804
rect 30088 15744 30152 15748
rect 23428 15540 23492 15604
rect 28948 15540 29012 15604
rect 46060 15812 46124 15816
rect 49112 15804 49176 15808
rect 49112 15748 49116 15804
rect 49116 15748 49172 15804
rect 49172 15748 49176 15804
rect 49112 15744 49176 15748
rect 49192 15804 49256 15808
rect 49192 15748 49196 15804
rect 49196 15748 49252 15804
rect 49252 15748 49256 15804
rect 49192 15744 49256 15748
rect 49272 15804 49336 15808
rect 49272 15748 49276 15804
rect 49276 15748 49332 15804
rect 49332 15748 49336 15804
rect 49272 15744 49336 15748
rect 49352 15804 49416 15808
rect 49352 15748 49356 15804
rect 49356 15748 49412 15804
rect 49412 15748 49416 15804
rect 49352 15744 49416 15748
rect 38700 15464 38764 15468
rect 38700 15408 38750 15464
rect 38750 15408 38764 15464
rect 38700 15404 38764 15408
rect 17356 15328 17420 15332
rect 17356 15272 17370 15328
rect 17370 15272 17420 15328
rect 17356 15268 17420 15272
rect 18092 15328 18156 15332
rect 18092 15272 18142 15328
rect 18142 15272 18156 15328
rect 18092 15268 18156 15272
rect 20216 15260 20280 15264
rect 20216 15204 20220 15260
rect 20220 15204 20276 15260
rect 20276 15204 20280 15260
rect 20216 15200 20280 15204
rect 20296 15260 20360 15264
rect 20296 15204 20300 15260
rect 20300 15204 20356 15260
rect 20356 15204 20360 15260
rect 20296 15200 20360 15204
rect 20376 15260 20440 15264
rect 20376 15204 20380 15260
rect 20380 15204 20436 15260
rect 20436 15204 20440 15260
rect 20376 15200 20440 15204
rect 20456 15260 20520 15264
rect 20456 15204 20460 15260
rect 20460 15204 20516 15260
rect 20516 15204 20520 15260
rect 20456 15200 20520 15204
rect 17172 14996 17236 15060
rect 21772 15328 21836 15332
rect 21772 15272 21786 15328
rect 21786 15272 21836 15328
rect 21772 15268 21836 15272
rect 22140 15268 22204 15332
rect 28764 15328 28828 15332
rect 28764 15272 28778 15328
rect 28778 15272 28828 15328
rect 28764 15268 28828 15272
rect 30604 15268 30668 15332
rect 38884 15268 38948 15332
rect 44404 15404 44468 15468
rect 42564 15268 42628 15332
rect 44220 15268 44284 15332
rect 44956 15328 45020 15332
rect 44956 15272 44970 15328
rect 44970 15272 45020 15328
rect 44956 15268 45020 15272
rect 39480 15260 39544 15264
rect 39480 15204 39484 15260
rect 39484 15204 39540 15260
rect 39540 15204 39544 15260
rect 39480 15200 39544 15204
rect 39560 15260 39624 15264
rect 39560 15204 39564 15260
rect 39564 15204 39620 15260
rect 39620 15204 39624 15260
rect 39560 15200 39624 15204
rect 39640 15260 39704 15264
rect 39640 15204 39644 15260
rect 39644 15204 39700 15260
rect 39700 15204 39704 15260
rect 39640 15200 39704 15204
rect 39720 15260 39784 15264
rect 39720 15204 39724 15260
rect 39724 15204 39780 15260
rect 39780 15204 39784 15260
rect 39720 15200 39784 15204
rect 19564 14860 19628 14924
rect 20668 14860 20732 14924
rect 23980 14860 24044 14924
rect 27476 14860 27540 14924
rect 30236 14724 30300 14788
rect 30788 14724 30852 14788
rect 36308 14724 36372 14788
rect 10584 14716 10648 14720
rect 10584 14660 10588 14716
rect 10588 14660 10644 14716
rect 10644 14660 10648 14716
rect 10584 14656 10648 14660
rect 10664 14716 10728 14720
rect 10664 14660 10668 14716
rect 10668 14660 10724 14716
rect 10724 14660 10728 14716
rect 10664 14656 10728 14660
rect 10744 14716 10808 14720
rect 10744 14660 10748 14716
rect 10748 14660 10804 14716
rect 10804 14660 10808 14716
rect 10744 14656 10808 14660
rect 10824 14716 10888 14720
rect 10824 14660 10828 14716
rect 10828 14660 10884 14716
rect 10884 14660 10888 14716
rect 10824 14656 10888 14660
rect 29848 14716 29912 14720
rect 29848 14660 29852 14716
rect 29852 14660 29908 14716
rect 29908 14660 29912 14716
rect 29848 14656 29912 14660
rect 29928 14716 29992 14720
rect 29928 14660 29932 14716
rect 29932 14660 29988 14716
rect 29988 14660 29992 14716
rect 29928 14656 29992 14660
rect 30008 14716 30072 14720
rect 30008 14660 30012 14716
rect 30012 14660 30068 14716
rect 30068 14660 30072 14716
rect 30008 14656 30072 14660
rect 30088 14716 30152 14720
rect 30088 14660 30092 14716
rect 30092 14660 30148 14716
rect 30148 14660 30152 14716
rect 30088 14656 30152 14660
rect 49112 14716 49176 14720
rect 49112 14660 49116 14716
rect 49116 14660 49172 14716
rect 49172 14660 49176 14716
rect 49112 14656 49176 14660
rect 49192 14716 49256 14720
rect 49192 14660 49196 14716
rect 49196 14660 49252 14716
rect 49252 14660 49256 14716
rect 49192 14656 49256 14660
rect 49272 14716 49336 14720
rect 49272 14660 49276 14716
rect 49276 14660 49332 14716
rect 49332 14660 49336 14716
rect 49272 14656 49336 14660
rect 49352 14716 49416 14720
rect 49352 14660 49356 14716
rect 49356 14660 49412 14716
rect 49412 14660 49416 14716
rect 49352 14656 49416 14660
rect 33180 14588 33244 14652
rect 35940 14588 36004 14652
rect 36492 14648 36556 14652
rect 36492 14592 36506 14648
rect 36506 14592 36556 14648
rect 36492 14588 36556 14592
rect 30788 14512 30852 14516
rect 30788 14456 30802 14512
rect 30802 14456 30852 14512
rect 30788 14452 30852 14456
rect 20216 14172 20280 14176
rect 20216 14116 20220 14172
rect 20220 14116 20276 14172
rect 20276 14116 20280 14172
rect 20216 14112 20280 14116
rect 20296 14172 20360 14176
rect 20296 14116 20300 14172
rect 20300 14116 20356 14172
rect 20356 14116 20360 14172
rect 20296 14112 20360 14116
rect 20376 14172 20440 14176
rect 20376 14116 20380 14172
rect 20380 14116 20436 14172
rect 20436 14116 20440 14172
rect 20376 14112 20440 14116
rect 20456 14172 20520 14176
rect 20456 14116 20460 14172
rect 20460 14116 20516 14172
rect 20516 14116 20520 14172
rect 20456 14112 20520 14116
rect 28028 14180 28092 14244
rect 28396 14180 28460 14244
rect 21772 14044 21836 14108
rect 22324 14044 22388 14108
rect 21404 13908 21468 13972
rect 21956 13908 22020 13972
rect 39480 14172 39544 14176
rect 39480 14116 39484 14172
rect 39484 14116 39540 14172
rect 39540 14116 39544 14172
rect 39480 14112 39544 14116
rect 39560 14172 39624 14176
rect 39560 14116 39564 14172
rect 39564 14116 39620 14172
rect 39620 14116 39624 14172
rect 39560 14112 39624 14116
rect 39640 14172 39704 14176
rect 39640 14116 39644 14172
rect 39644 14116 39700 14172
rect 39700 14116 39704 14172
rect 39640 14112 39704 14116
rect 39720 14172 39784 14176
rect 39720 14116 39724 14172
rect 39724 14116 39780 14172
rect 39780 14116 39784 14172
rect 39720 14112 39784 14116
rect 40172 14104 40236 14108
rect 40172 14048 40186 14104
rect 40186 14048 40236 14104
rect 40172 14044 40236 14048
rect 34836 13908 34900 13972
rect 39252 13968 39316 13972
rect 39252 13912 39266 13968
rect 39266 13912 39316 13968
rect 39252 13908 39316 13912
rect 39988 13908 40052 13972
rect 40356 13908 40420 13972
rect 24716 13832 24780 13836
rect 24716 13776 24730 13832
rect 24730 13776 24780 13832
rect 24716 13772 24780 13776
rect 24900 13832 24964 13836
rect 24900 13776 24950 13832
rect 24950 13776 24964 13832
rect 24900 13772 24964 13776
rect 28948 13772 29012 13836
rect 35204 13772 35268 13836
rect 35940 13832 36004 13836
rect 42932 13908 42996 13972
rect 35940 13776 35990 13832
rect 35990 13776 36004 13832
rect 35940 13772 36004 13776
rect 42748 13772 42812 13836
rect 21036 13636 21100 13700
rect 10584 13628 10648 13632
rect 10584 13572 10588 13628
rect 10588 13572 10644 13628
rect 10644 13572 10648 13628
rect 10584 13568 10648 13572
rect 10664 13628 10728 13632
rect 10664 13572 10668 13628
rect 10668 13572 10724 13628
rect 10724 13572 10728 13628
rect 10664 13568 10728 13572
rect 10744 13628 10808 13632
rect 10744 13572 10748 13628
rect 10748 13572 10804 13628
rect 10804 13572 10808 13628
rect 10744 13568 10808 13572
rect 10824 13628 10888 13632
rect 10824 13572 10828 13628
rect 10828 13572 10884 13628
rect 10884 13572 10888 13628
rect 10824 13568 10888 13572
rect 29848 13628 29912 13632
rect 29848 13572 29852 13628
rect 29852 13572 29908 13628
rect 29908 13572 29912 13628
rect 29848 13568 29912 13572
rect 29928 13628 29992 13632
rect 29928 13572 29932 13628
rect 29932 13572 29988 13628
rect 29988 13572 29992 13628
rect 29928 13568 29992 13572
rect 30008 13628 30072 13632
rect 30008 13572 30012 13628
rect 30012 13572 30068 13628
rect 30068 13572 30072 13628
rect 30008 13568 30072 13572
rect 30088 13628 30152 13632
rect 30088 13572 30092 13628
rect 30092 13572 30148 13628
rect 30148 13572 30152 13628
rect 30088 13568 30152 13572
rect 49112 13628 49176 13632
rect 49112 13572 49116 13628
rect 49116 13572 49172 13628
rect 49172 13572 49176 13628
rect 49112 13568 49176 13572
rect 49192 13628 49256 13632
rect 49192 13572 49196 13628
rect 49196 13572 49252 13628
rect 49252 13572 49256 13628
rect 49192 13568 49256 13572
rect 49272 13628 49336 13632
rect 49272 13572 49276 13628
rect 49276 13572 49332 13628
rect 49332 13572 49336 13628
rect 49272 13568 49336 13572
rect 49352 13628 49416 13632
rect 49352 13572 49356 13628
rect 49356 13572 49412 13628
rect 49412 13572 49416 13628
rect 49352 13568 49416 13572
rect 19380 13500 19444 13564
rect 25268 13228 25332 13292
rect 33732 13364 33796 13428
rect 38332 13560 38396 13564
rect 38332 13504 38346 13560
rect 38346 13504 38396 13560
rect 38332 13500 38396 13504
rect 20216 13084 20280 13088
rect 20216 13028 20220 13084
rect 20220 13028 20276 13084
rect 20276 13028 20280 13084
rect 20216 13024 20280 13028
rect 20296 13084 20360 13088
rect 20296 13028 20300 13084
rect 20300 13028 20356 13084
rect 20356 13028 20360 13084
rect 20296 13024 20360 13028
rect 20376 13084 20440 13088
rect 20376 13028 20380 13084
rect 20380 13028 20436 13084
rect 20436 13028 20440 13084
rect 20376 13024 20440 13028
rect 20456 13084 20520 13088
rect 20456 13028 20460 13084
rect 20460 13028 20516 13084
rect 20516 13028 20520 13084
rect 20456 13024 20520 13028
rect 21220 12956 21284 13020
rect 26372 13016 26436 13020
rect 26372 12960 26422 13016
rect 26422 12960 26436 13016
rect 26372 12956 26436 12960
rect 27660 12956 27724 13020
rect 38700 12880 38764 12884
rect 39480 13084 39544 13088
rect 39480 13028 39484 13084
rect 39484 13028 39540 13084
rect 39540 13028 39544 13084
rect 39480 13024 39544 13028
rect 39560 13084 39624 13088
rect 39560 13028 39564 13084
rect 39564 13028 39620 13084
rect 39620 13028 39624 13084
rect 39560 13024 39624 13028
rect 39640 13084 39704 13088
rect 39640 13028 39644 13084
rect 39644 13028 39700 13084
rect 39700 13028 39704 13084
rect 39640 13024 39704 13028
rect 39720 13084 39784 13088
rect 39720 13028 39724 13084
rect 39724 13028 39780 13084
rect 39780 13028 39784 13084
rect 39720 13024 39784 13028
rect 38700 12824 38750 12880
rect 38750 12824 38764 12880
rect 38700 12820 38764 12824
rect 20668 12684 20732 12748
rect 25820 12684 25884 12748
rect 27844 12684 27908 12748
rect 10584 12540 10648 12544
rect 10584 12484 10588 12540
rect 10588 12484 10644 12540
rect 10644 12484 10648 12540
rect 10584 12480 10648 12484
rect 10664 12540 10728 12544
rect 10664 12484 10668 12540
rect 10668 12484 10724 12540
rect 10724 12484 10728 12540
rect 10664 12480 10728 12484
rect 10744 12540 10808 12544
rect 10744 12484 10748 12540
rect 10748 12484 10804 12540
rect 10804 12484 10808 12540
rect 10744 12480 10808 12484
rect 10824 12540 10888 12544
rect 10824 12484 10828 12540
rect 10828 12484 10884 12540
rect 10884 12484 10888 12540
rect 10824 12480 10888 12484
rect 21588 12412 21652 12476
rect 24532 12276 24596 12340
rect 28028 12548 28092 12612
rect 29500 12608 29564 12612
rect 29500 12552 29550 12608
rect 29550 12552 29564 12608
rect 29500 12548 29564 12552
rect 30972 12684 31036 12748
rect 38884 12744 38948 12748
rect 38884 12688 38934 12744
rect 38934 12688 38948 12744
rect 38884 12684 38948 12688
rect 29848 12540 29912 12544
rect 29848 12484 29852 12540
rect 29852 12484 29908 12540
rect 29908 12484 29912 12540
rect 29848 12480 29912 12484
rect 29928 12540 29992 12544
rect 29928 12484 29932 12540
rect 29932 12484 29988 12540
rect 29988 12484 29992 12540
rect 29928 12480 29992 12484
rect 30008 12540 30072 12544
rect 30008 12484 30012 12540
rect 30012 12484 30068 12540
rect 30068 12484 30072 12540
rect 30008 12480 30072 12484
rect 30088 12540 30152 12544
rect 30088 12484 30092 12540
rect 30092 12484 30148 12540
rect 30148 12484 30152 12540
rect 30088 12480 30152 12484
rect 31892 12276 31956 12340
rect 33732 12548 33796 12612
rect 49112 12540 49176 12544
rect 49112 12484 49116 12540
rect 49116 12484 49172 12540
rect 49172 12484 49176 12540
rect 49112 12480 49176 12484
rect 49192 12540 49256 12544
rect 49192 12484 49196 12540
rect 49196 12484 49252 12540
rect 49252 12484 49256 12540
rect 49192 12480 49256 12484
rect 49272 12540 49336 12544
rect 49272 12484 49276 12540
rect 49276 12484 49332 12540
rect 49332 12484 49336 12540
rect 49272 12480 49336 12484
rect 49352 12540 49416 12544
rect 49352 12484 49356 12540
rect 49356 12484 49412 12540
rect 49412 12484 49416 12540
rect 49352 12480 49416 12484
rect 40356 12336 40420 12340
rect 40356 12280 40406 12336
rect 40406 12280 40420 12336
rect 40356 12276 40420 12280
rect 20852 12064 20916 12068
rect 20852 12008 20902 12064
rect 20902 12008 20916 12064
rect 20852 12004 20916 12008
rect 28580 12004 28644 12068
rect 30236 12004 30300 12068
rect 34652 12004 34716 12068
rect 20216 11996 20280 12000
rect 20216 11940 20220 11996
rect 20220 11940 20276 11996
rect 20276 11940 20280 11996
rect 20216 11936 20280 11940
rect 20296 11996 20360 12000
rect 20296 11940 20300 11996
rect 20300 11940 20356 11996
rect 20356 11940 20360 11996
rect 20296 11936 20360 11940
rect 20376 11996 20440 12000
rect 20376 11940 20380 11996
rect 20380 11940 20436 11996
rect 20436 11940 20440 11996
rect 20376 11936 20440 11940
rect 20456 11996 20520 12000
rect 20456 11940 20460 11996
rect 20460 11940 20516 11996
rect 20516 11940 20520 11996
rect 20456 11936 20520 11940
rect 39988 12004 40052 12068
rect 39480 11996 39544 12000
rect 39480 11940 39484 11996
rect 39484 11940 39540 11996
rect 39540 11940 39544 11996
rect 39480 11936 39544 11940
rect 39560 11996 39624 12000
rect 39560 11940 39564 11996
rect 39564 11940 39620 11996
rect 39620 11940 39624 11996
rect 39560 11936 39624 11940
rect 39640 11996 39704 12000
rect 39640 11940 39644 11996
rect 39644 11940 39700 11996
rect 39700 11940 39704 11996
rect 39640 11936 39704 11940
rect 39720 11996 39784 12000
rect 39720 11940 39724 11996
rect 39724 11940 39780 11996
rect 39780 11940 39784 11996
rect 39720 11936 39784 11940
rect 29316 11732 29380 11796
rect 30420 11596 30484 11660
rect 36308 11596 36372 11660
rect 21220 11460 21284 11524
rect 29316 11520 29380 11524
rect 29316 11464 29330 11520
rect 29330 11464 29380 11520
rect 29316 11460 29380 11464
rect 30236 11460 30300 11524
rect 35756 11520 35820 11524
rect 35756 11464 35806 11520
rect 35806 11464 35820 11520
rect 35756 11460 35820 11464
rect 37596 11520 37660 11524
rect 37596 11464 37646 11520
rect 37646 11464 37660 11520
rect 37596 11460 37660 11464
rect 10584 11452 10648 11456
rect 10584 11396 10588 11452
rect 10588 11396 10644 11452
rect 10644 11396 10648 11452
rect 10584 11392 10648 11396
rect 10664 11452 10728 11456
rect 10664 11396 10668 11452
rect 10668 11396 10724 11452
rect 10724 11396 10728 11452
rect 10664 11392 10728 11396
rect 10744 11452 10808 11456
rect 10744 11396 10748 11452
rect 10748 11396 10804 11452
rect 10804 11396 10808 11452
rect 10744 11392 10808 11396
rect 10824 11452 10888 11456
rect 10824 11396 10828 11452
rect 10828 11396 10884 11452
rect 10884 11396 10888 11452
rect 10824 11392 10888 11396
rect 29848 11452 29912 11456
rect 29848 11396 29852 11452
rect 29852 11396 29908 11452
rect 29908 11396 29912 11452
rect 29848 11392 29912 11396
rect 29928 11452 29992 11456
rect 29928 11396 29932 11452
rect 29932 11396 29988 11452
rect 29988 11396 29992 11452
rect 29928 11392 29992 11396
rect 30008 11452 30072 11456
rect 30008 11396 30012 11452
rect 30012 11396 30068 11452
rect 30068 11396 30072 11452
rect 30008 11392 30072 11396
rect 30088 11452 30152 11456
rect 30088 11396 30092 11452
rect 30092 11396 30148 11452
rect 30148 11396 30152 11452
rect 30088 11392 30152 11396
rect 49112 11452 49176 11456
rect 49112 11396 49116 11452
rect 49116 11396 49172 11452
rect 49172 11396 49176 11452
rect 49112 11392 49176 11396
rect 49192 11452 49256 11456
rect 49192 11396 49196 11452
rect 49196 11396 49252 11452
rect 49252 11396 49256 11452
rect 49192 11392 49256 11396
rect 49272 11452 49336 11456
rect 49272 11396 49276 11452
rect 49276 11396 49332 11452
rect 49332 11396 49336 11452
rect 49272 11392 49336 11396
rect 49352 11452 49416 11456
rect 49352 11396 49356 11452
rect 49356 11396 49412 11452
rect 49412 11396 49416 11452
rect 49352 11392 49416 11396
rect 20668 11324 20732 11388
rect 22140 11324 22204 11388
rect 24164 11324 24228 11388
rect 25452 11324 25516 11388
rect 27108 11324 27172 11388
rect 28580 11324 28644 11388
rect 23980 11052 24044 11116
rect 26924 11052 26988 11116
rect 28948 11052 29012 11116
rect 32812 11052 32876 11116
rect 33548 11188 33612 11252
rect 35940 11188 36004 11252
rect 20216 10908 20280 10912
rect 20216 10852 20220 10908
rect 20220 10852 20276 10908
rect 20276 10852 20280 10908
rect 20216 10848 20280 10852
rect 20296 10908 20360 10912
rect 20296 10852 20300 10908
rect 20300 10852 20356 10908
rect 20356 10852 20360 10908
rect 20296 10848 20360 10852
rect 20376 10908 20440 10912
rect 20376 10852 20380 10908
rect 20380 10852 20436 10908
rect 20436 10852 20440 10908
rect 20376 10848 20440 10852
rect 20456 10908 20520 10912
rect 20456 10852 20460 10908
rect 20460 10852 20516 10908
rect 20516 10852 20520 10908
rect 20456 10848 20520 10852
rect 33180 10916 33244 10980
rect 39480 10908 39544 10912
rect 39480 10852 39484 10908
rect 39484 10852 39540 10908
rect 39540 10852 39544 10908
rect 39480 10848 39544 10852
rect 39560 10908 39624 10912
rect 39560 10852 39564 10908
rect 39564 10852 39620 10908
rect 39620 10852 39624 10908
rect 39560 10848 39624 10852
rect 39640 10908 39704 10912
rect 39640 10852 39644 10908
rect 39644 10852 39700 10908
rect 39700 10852 39704 10908
rect 39640 10848 39704 10852
rect 39720 10908 39784 10912
rect 39720 10852 39724 10908
rect 39724 10852 39780 10908
rect 39780 10852 39784 10908
rect 39720 10848 39784 10852
rect 36124 10780 36188 10844
rect 29132 10644 29196 10708
rect 33732 10704 33796 10708
rect 33732 10648 33782 10704
rect 33782 10648 33796 10704
rect 33732 10644 33796 10648
rect 37228 10372 37292 10436
rect 10584 10364 10648 10368
rect 10584 10308 10588 10364
rect 10588 10308 10644 10364
rect 10644 10308 10648 10364
rect 10584 10304 10648 10308
rect 10664 10364 10728 10368
rect 10664 10308 10668 10364
rect 10668 10308 10724 10364
rect 10724 10308 10728 10364
rect 10664 10304 10728 10308
rect 10744 10364 10808 10368
rect 10744 10308 10748 10364
rect 10748 10308 10804 10364
rect 10804 10308 10808 10364
rect 10744 10304 10808 10308
rect 10824 10364 10888 10368
rect 10824 10308 10828 10364
rect 10828 10308 10884 10364
rect 10884 10308 10888 10364
rect 10824 10304 10888 10308
rect 29848 10364 29912 10368
rect 29848 10308 29852 10364
rect 29852 10308 29908 10364
rect 29908 10308 29912 10364
rect 29848 10304 29912 10308
rect 29928 10364 29992 10368
rect 29928 10308 29932 10364
rect 29932 10308 29988 10364
rect 29988 10308 29992 10364
rect 29928 10304 29992 10308
rect 30008 10364 30072 10368
rect 30008 10308 30012 10364
rect 30012 10308 30068 10364
rect 30068 10308 30072 10364
rect 30008 10304 30072 10308
rect 30088 10364 30152 10368
rect 30088 10308 30092 10364
rect 30092 10308 30148 10364
rect 30148 10308 30152 10364
rect 30088 10304 30152 10308
rect 49112 10364 49176 10368
rect 49112 10308 49116 10364
rect 49116 10308 49172 10364
rect 49172 10308 49176 10364
rect 49112 10304 49176 10308
rect 49192 10364 49256 10368
rect 49192 10308 49196 10364
rect 49196 10308 49252 10364
rect 49252 10308 49256 10364
rect 49192 10304 49256 10308
rect 49272 10364 49336 10368
rect 49272 10308 49276 10364
rect 49276 10308 49332 10364
rect 49332 10308 49336 10364
rect 49272 10304 49336 10308
rect 49352 10364 49416 10368
rect 49352 10308 49356 10364
rect 49356 10308 49412 10364
rect 49412 10308 49416 10364
rect 49352 10304 49416 10308
rect 25268 9964 25332 10028
rect 35756 10100 35820 10164
rect 20216 9820 20280 9824
rect 20216 9764 20220 9820
rect 20220 9764 20276 9820
rect 20276 9764 20280 9820
rect 20216 9760 20280 9764
rect 20296 9820 20360 9824
rect 20296 9764 20300 9820
rect 20300 9764 20356 9820
rect 20356 9764 20360 9820
rect 20296 9760 20360 9764
rect 20376 9820 20440 9824
rect 20376 9764 20380 9820
rect 20380 9764 20436 9820
rect 20436 9764 20440 9820
rect 20376 9760 20440 9764
rect 20456 9820 20520 9824
rect 20456 9764 20460 9820
rect 20460 9764 20516 9820
rect 20516 9764 20520 9820
rect 20456 9760 20520 9764
rect 21956 9692 22020 9756
rect 30236 9692 30300 9756
rect 32076 9752 32140 9756
rect 32076 9696 32126 9752
rect 32126 9696 32140 9752
rect 32076 9692 32140 9696
rect 29684 9556 29748 9620
rect 32996 9692 33060 9756
rect 34468 9752 34532 9756
rect 34468 9696 34518 9752
rect 34518 9696 34532 9752
rect 34468 9692 34532 9696
rect 39480 9820 39544 9824
rect 39480 9764 39484 9820
rect 39484 9764 39540 9820
rect 39540 9764 39544 9820
rect 39480 9760 39544 9764
rect 39560 9820 39624 9824
rect 39560 9764 39564 9820
rect 39564 9764 39620 9820
rect 39620 9764 39624 9820
rect 39560 9760 39624 9764
rect 39640 9820 39704 9824
rect 39640 9764 39644 9820
rect 39644 9764 39700 9820
rect 39700 9764 39704 9820
rect 39640 9760 39704 9764
rect 39720 9820 39784 9824
rect 39720 9764 39724 9820
rect 39724 9764 39780 9820
rect 39780 9764 39784 9820
rect 39720 9760 39784 9764
rect 32444 9556 32508 9620
rect 34100 9556 34164 9620
rect 35020 9556 35084 9620
rect 10584 9276 10648 9280
rect 10584 9220 10588 9276
rect 10588 9220 10644 9276
rect 10644 9220 10648 9276
rect 10584 9216 10648 9220
rect 10664 9276 10728 9280
rect 10664 9220 10668 9276
rect 10668 9220 10724 9276
rect 10724 9220 10728 9276
rect 10664 9216 10728 9220
rect 10744 9276 10808 9280
rect 10744 9220 10748 9276
rect 10748 9220 10804 9276
rect 10804 9220 10808 9276
rect 10744 9216 10808 9220
rect 10824 9276 10888 9280
rect 10824 9220 10828 9276
rect 10828 9220 10884 9276
rect 10884 9220 10888 9276
rect 10824 9216 10888 9220
rect 24900 9420 24964 9484
rect 30972 9420 31036 9484
rect 32260 9420 32324 9484
rect 29848 9276 29912 9280
rect 29848 9220 29852 9276
rect 29852 9220 29908 9276
rect 29908 9220 29912 9276
rect 29848 9216 29912 9220
rect 29928 9276 29992 9280
rect 29928 9220 29932 9276
rect 29932 9220 29988 9276
rect 29988 9220 29992 9276
rect 29928 9216 29992 9220
rect 30008 9276 30072 9280
rect 30008 9220 30012 9276
rect 30012 9220 30068 9276
rect 30068 9220 30072 9276
rect 30008 9216 30072 9220
rect 30088 9276 30152 9280
rect 30088 9220 30092 9276
rect 30092 9220 30148 9276
rect 30148 9220 30152 9276
rect 30088 9216 30152 9220
rect 49112 9276 49176 9280
rect 49112 9220 49116 9276
rect 49116 9220 49172 9276
rect 49172 9220 49176 9276
rect 49112 9216 49176 9220
rect 49192 9276 49256 9280
rect 49192 9220 49196 9276
rect 49196 9220 49252 9276
rect 49252 9220 49256 9276
rect 49192 9216 49256 9220
rect 49272 9276 49336 9280
rect 49272 9220 49276 9276
rect 49276 9220 49332 9276
rect 49332 9220 49336 9276
rect 49272 9216 49336 9220
rect 49352 9276 49416 9280
rect 49352 9220 49356 9276
rect 49356 9220 49412 9276
rect 49412 9220 49416 9276
rect 49352 9216 49416 9220
rect 26556 9148 26620 9212
rect 27476 9012 27540 9076
rect 37412 9012 37476 9076
rect 30604 8740 30668 8804
rect 20216 8732 20280 8736
rect 20216 8676 20220 8732
rect 20220 8676 20276 8732
rect 20276 8676 20280 8732
rect 20216 8672 20280 8676
rect 20296 8732 20360 8736
rect 20296 8676 20300 8732
rect 20300 8676 20356 8732
rect 20356 8676 20360 8732
rect 20296 8672 20360 8676
rect 20376 8732 20440 8736
rect 20376 8676 20380 8732
rect 20380 8676 20436 8732
rect 20436 8676 20440 8732
rect 20376 8672 20440 8676
rect 20456 8732 20520 8736
rect 20456 8676 20460 8732
rect 20460 8676 20516 8732
rect 20516 8676 20520 8732
rect 20456 8672 20520 8676
rect 39480 8732 39544 8736
rect 39480 8676 39484 8732
rect 39484 8676 39540 8732
rect 39540 8676 39544 8732
rect 39480 8672 39544 8676
rect 39560 8732 39624 8736
rect 39560 8676 39564 8732
rect 39564 8676 39620 8732
rect 39620 8676 39624 8732
rect 39560 8672 39624 8676
rect 39640 8732 39704 8736
rect 39640 8676 39644 8732
rect 39644 8676 39700 8732
rect 39700 8676 39704 8732
rect 39640 8672 39704 8676
rect 39720 8732 39784 8736
rect 39720 8676 39724 8732
rect 39724 8676 39780 8732
rect 39780 8676 39784 8732
rect 39720 8672 39784 8676
rect 23428 8604 23492 8668
rect 27660 8332 27724 8396
rect 28948 8332 29012 8396
rect 15332 8196 15396 8260
rect 29500 8196 29564 8260
rect 10584 8188 10648 8192
rect 10584 8132 10588 8188
rect 10588 8132 10644 8188
rect 10644 8132 10648 8188
rect 10584 8128 10648 8132
rect 10664 8188 10728 8192
rect 10664 8132 10668 8188
rect 10668 8132 10724 8188
rect 10724 8132 10728 8188
rect 10664 8128 10728 8132
rect 10744 8188 10808 8192
rect 10744 8132 10748 8188
rect 10748 8132 10804 8188
rect 10804 8132 10808 8188
rect 10744 8128 10808 8132
rect 10824 8188 10888 8192
rect 10824 8132 10828 8188
rect 10828 8132 10884 8188
rect 10884 8132 10888 8188
rect 10824 8128 10888 8132
rect 29848 8188 29912 8192
rect 29848 8132 29852 8188
rect 29852 8132 29908 8188
rect 29908 8132 29912 8188
rect 29848 8128 29912 8132
rect 29928 8188 29992 8192
rect 29928 8132 29932 8188
rect 29932 8132 29988 8188
rect 29988 8132 29992 8188
rect 29928 8128 29992 8132
rect 30008 8188 30072 8192
rect 30008 8132 30012 8188
rect 30012 8132 30068 8188
rect 30068 8132 30072 8188
rect 30008 8128 30072 8132
rect 30088 8188 30152 8192
rect 30088 8132 30092 8188
rect 30092 8132 30148 8188
rect 30148 8132 30152 8188
rect 30088 8128 30152 8132
rect 49112 8188 49176 8192
rect 49112 8132 49116 8188
rect 49116 8132 49172 8188
rect 49172 8132 49176 8188
rect 49112 8128 49176 8132
rect 49192 8188 49256 8192
rect 49192 8132 49196 8188
rect 49196 8132 49252 8188
rect 49252 8132 49256 8188
rect 49192 8128 49256 8132
rect 49272 8188 49336 8192
rect 49272 8132 49276 8188
rect 49276 8132 49332 8188
rect 49332 8132 49336 8188
rect 49272 8128 49336 8132
rect 49352 8188 49416 8192
rect 49352 8132 49356 8188
rect 49356 8132 49412 8188
rect 49412 8132 49416 8188
rect 49352 8128 49416 8132
rect 19748 8060 19812 8124
rect 24716 8120 24780 8124
rect 24716 8064 24766 8120
rect 24766 8064 24780 8120
rect 24716 8060 24780 8064
rect 25820 8060 25884 8124
rect 21772 7788 21836 7852
rect 20216 7644 20280 7648
rect 20216 7588 20220 7644
rect 20220 7588 20276 7644
rect 20276 7588 20280 7644
rect 20216 7584 20280 7588
rect 20296 7644 20360 7648
rect 20296 7588 20300 7644
rect 20300 7588 20356 7644
rect 20356 7588 20360 7644
rect 20296 7584 20360 7588
rect 20376 7644 20440 7648
rect 20376 7588 20380 7644
rect 20380 7588 20436 7644
rect 20436 7588 20440 7644
rect 20376 7584 20440 7588
rect 20456 7644 20520 7648
rect 20456 7588 20460 7644
rect 20460 7588 20516 7644
rect 20516 7588 20520 7644
rect 20456 7584 20520 7588
rect 39480 7644 39544 7648
rect 39480 7588 39484 7644
rect 39484 7588 39540 7644
rect 39540 7588 39544 7644
rect 39480 7584 39544 7588
rect 39560 7644 39624 7648
rect 39560 7588 39564 7644
rect 39564 7588 39620 7644
rect 39620 7588 39624 7644
rect 39560 7584 39624 7588
rect 39640 7644 39704 7648
rect 39640 7588 39644 7644
rect 39644 7588 39700 7644
rect 39700 7588 39704 7644
rect 39640 7584 39704 7588
rect 39720 7644 39784 7648
rect 39720 7588 39724 7644
rect 39724 7588 39780 7644
rect 39780 7588 39784 7644
rect 39720 7584 39784 7588
rect 30236 7576 30300 7580
rect 30236 7520 30286 7576
rect 30286 7520 30300 7576
rect 30236 7516 30300 7520
rect 28764 7380 28828 7444
rect 33548 7380 33612 7444
rect 10584 7100 10648 7104
rect 10584 7044 10588 7100
rect 10588 7044 10644 7100
rect 10644 7044 10648 7100
rect 10584 7040 10648 7044
rect 10664 7100 10728 7104
rect 10664 7044 10668 7100
rect 10668 7044 10724 7100
rect 10724 7044 10728 7100
rect 10664 7040 10728 7044
rect 10744 7100 10808 7104
rect 10744 7044 10748 7100
rect 10748 7044 10804 7100
rect 10804 7044 10808 7100
rect 10744 7040 10808 7044
rect 10824 7100 10888 7104
rect 10824 7044 10828 7100
rect 10828 7044 10884 7100
rect 10884 7044 10888 7100
rect 10824 7040 10888 7044
rect 29848 7100 29912 7104
rect 29848 7044 29852 7100
rect 29852 7044 29908 7100
rect 29908 7044 29912 7100
rect 29848 7040 29912 7044
rect 29928 7100 29992 7104
rect 29928 7044 29932 7100
rect 29932 7044 29988 7100
rect 29988 7044 29992 7100
rect 29928 7040 29992 7044
rect 30008 7100 30072 7104
rect 30008 7044 30012 7100
rect 30012 7044 30068 7100
rect 30068 7044 30072 7100
rect 30008 7040 30072 7044
rect 30088 7100 30152 7104
rect 30088 7044 30092 7100
rect 30092 7044 30148 7100
rect 30148 7044 30152 7100
rect 30088 7040 30152 7044
rect 49112 7100 49176 7104
rect 49112 7044 49116 7100
rect 49116 7044 49172 7100
rect 49172 7044 49176 7100
rect 49112 7040 49176 7044
rect 49192 7100 49256 7104
rect 49192 7044 49196 7100
rect 49196 7044 49252 7100
rect 49252 7044 49256 7100
rect 49192 7040 49256 7044
rect 49272 7100 49336 7104
rect 49272 7044 49276 7100
rect 49276 7044 49332 7100
rect 49332 7044 49336 7100
rect 49272 7040 49336 7044
rect 49352 7100 49416 7104
rect 49352 7044 49356 7100
rect 49356 7044 49412 7100
rect 49412 7044 49416 7100
rect 49352 7040 49416 7044
rect 17540 6836 17604 6900
rect 32812 6836 32876 6900
rect 18460 6700 18524 6764
rect 36492 6700 36556 6764
rect 20216 6556 20280 6560
rect 20216 6500 20220 6556
rect 20220 6500 20276 6556
rect 20276 6500 20280 6556
rect 20216 6496 20280 6500
rect 20296 6556 20360 6560
rect 20296 6500 20300 6556
rect 20300 6500 20356 6556
rect 20356 6500 20360 6556
rect 20296 6496 20360 6500
rect 20376 6556 20440 6560
rect 20376 6500 20380 6556
rect 20380 6500 20436 6556
rect 20436 6500 20440 6556
rect 20376 6496 20440 6500
rect 20456 6556 20520 6560
rect 20456 6500 20460 6556
rect 20460 6500 20516 6556
rect 20516 6500 20520 6556
rect 20456 6496 20520 6500
rect 28396 6488 28460 6492
rect 39480 6556 39544 6560
rect 39480 6500 39484 6556
rect 39484 6500 39540 6556
rect 39540 6500 39544 6556
rect 39480 6496 39544 6500
rect 39560 6556 39624 6560
rect 39560 6500 39564 6556
rect 39564 6500 39620 6556
rect 39620 6500 39624 6556
rect 39560 6496 39624 6500
rect 39640 6556 39704 6560
rect 39640 6500 39644 6556
rect 39644 6500 39700 6556
rect 39700 6500 39704 6556
rect 39640 6496 39704 6500
rect 39720 6556 39784 6560
rect 39720 6500 39724 6556
rect 39724 6500 39780 6556
rect 39780 6500 39784 6556
rect 39720 6496 39784 6500
rect 28396 6432 28446 6488
rect 28446 6432 28460 6488
rect 28396 6428 28460 6432
rect 17356 6292 17420 6356
rect 42564 6292 42628 6356
rect 30236 6156 30300 6220
rect 10584 6012 10648 6016
rect 10584 5956 10588 6012
rect 10588 5956 10644 6012
rect 10644 5956 10648 6012
rect 10584 5952 10648 5956
rect 10664 6012 10728 6016
rect 10664 5956 10668 6012
rect 10668 5956 10724 6012
rect 10724 5956 10728 6012
rect 10664 5952 10728 5956
rect 10744 6012 10808 6016
rect 10744 5956 10748 6012
rect 10748 5956 10804 6012
rect 10804 5956 10808 6012
rect 10744 5952 10808 5956
rect 10824 6012 10888 6016
rect 10824 5956 10828 6012
rect 10828 5956 10884 6012
rect 10884 5956 10888 6012
rect 10824 5952 10888 5956
rect 29848 6012 29912 6016
rect 29848 5956 29852 6012
rect 29852 5956 29908 6012
rect 29908 5956 29912 6012
rect 29848 5952 29912 5956
rect 29928 6012 29992 6016
rect 29928 5956 29932 6012
rect 29932 5956 29988 6012
rect 29988 5956 29992 6012
rect 29928 5952 29992 5956
rect 30008 6012 30072 6016
rect 30008 5956 30012 6012
rect 30012 5956 30068 6012
rect 30068 5956 30072 6012
rect 30008 5952 30072 5956
rect 30088 6012 30152 6016
rect 30088 5956 30092 6012
rect 30092 5956 30148 6012
rect 30148 5956 30152 6012
rect 30088 5952 30152 5956
rect 49112 6012 49176 6016
rect 49112 5956 49116 6012
rect 49116 5956 49172 6012
rect 49172 5956 49176 6012
rect 49112 5952 49176 5956
rect 49192 6012 49256 6016
rect 49192 5956 49196 6012
rect 49196 5956 49252 6012
rect 49252 5956 49256 6012
rect 49192 5952 49256 5956
rect 49272 6012 49336 6016
rect 49272 5956 49276 6012
rect 49276 5956 49332 6012
rect 49332 5956 49336 6012
rect 49272 5952 49336 5956
rect 49352 6012 49416 6016
rect 49352 5956 49356 6012
rect 49356 5956 49412 6012
rect 49412 5956 49416 6012
rect 49352 5952 49416 5956
rect 32812 5944 32876 5948
rect 32812 5888 32862 5944
rect 32862 5888 32876 5944
rect 32812 5884 32876 5888
rect 20216 5468 20280 5472
rect 20216 5412 20220 5468
rect 20220 5412 20276 5468
rect 20276 5412 20280 5468
rect 20216 5408 20280 5412
rect 20296 5468 20360 5472
rect 20296 5412 20300 5468
rect 20300 5412 20356 5468
rect 20356 5412 20360 5468
rect 20296 5408 20360 5412
rect 20376 5468 20440 5472
rect 20376 5412 20380 5468
rect 20380 5412 20436 5468
rect 20436 5412 20440 5468
rect 20376 5408 20440 5412
rect 20456 5468 20520 5472
rect 20456 5412 20460 5468
rect 20460 5412 20516 5468
rect 20516 5412 20520 5468
rect 20456 5408 20520 5412
rect 29500 5400 29564 5404
rect 29500 5344 29514 5400
rect 29514 5344 29564 5400
rect 29500 5340 29564 5344
rect 39480 5468 39544 5472
rect 39480 5412 39484 5468
rect 39484 5412 39540 5468
rect 39540 5412 39544 5468
rect 39480 5408 39544 5412
rect 39560 5468 39624 5472
rect 39560 5412 39564 5468
rect 39564 5412 39620 5468
rect 39620 5412 39624 5468
rect 39560 5408 39624 5412
rect 39640 5468 39704 5472
rect 39640 5412 39644 5468
rect 39644 5412 39700 5468
rect 39700 5412 39704 5468
rect 39640 5408 39704 5412
rect 39720 5468 39784 5472
rect 39720 5412 39724 5468
rect 39724 5412 39780 5468
rect 39780 5412 39784 5468
rect 39720 5408 39784 5412
rect 35940 5204 36004 5268
rect 42196 5204 42260 5268
rect 33548 5068 33612 5132
rect 37596 5068 37660 5132
rect 10584 4924 10648 4928
rect 10584 4868 10588 4924
rect 10588 4868 10644 4924
rect 10644 4868 10648 4924
rect 10584 4864 10648 4868
rect 10664 4924 10728 4928
rect 10664 4868 10668 4924
rect 10668 4868 10724 4924
rect 10724 4868 10728 4924
rect 10664 4864 10728 4868
rect 10744 4924 10808 4928
rect 10744 4868 10748 4924
rect 10748 4868 10804 4924
rect 10804 4868 10808 4924
rect 10744 4864 10808 4868
rect 10824 4924 10888 4928
rect 10824 4868 10828 4924
rect 10828 4868 10884 4924
rect 10884 4868 10888 4924
rect 10824 4864 10888 4868
rect 29848 4924 29912 4928
rect 29848 4868 29852 4924
rect 29852 4868 29908 4924
rect 29908 4868 29912 4924
rect 29848 4864 29912 4868
rect 29928 4924 29992 4928
rect 29928 4868 29932 4924
rect 29932 4868 29988 4924
rect 29988 4868 29992 4924
rect 29928 4864 29992 4868
rect 30008 4924 30072 4928
rect 30008 4868 30012 4924
rect 30012 4868 30068 4924
rect 30068 4868 30072 4924
rect 30008 4864 30072 4868
rect 30088 4924 30152 4928
rect 30088 4868 30092 4924
rect 30092 4868 30148 4924
rect 30148 4868 30152 4924
rect 30088 4864 30152 4868
rect 49112 4924 49176 4928
rect 49112 4868 49116 4924
rect 49116 4868 49172 4924
rect 49172 4868 49176 4924
rect 49112 4864 49176 4868
rect 49192 4924 49256 4928
rect 49192 4868 49196 4924
rect 49196 4868 49252 4924
rect 49252 4868 49256 4924
rect 49192 4864 49256 4868
rect 49272 4924 49336 4928
rect 49272 4868 49276 4924
rect 49276 4868 49332 4924
rect 49332 4868 49336 4924
rect 49272 4864 49336 4868
rect 49352 4924 49416 4928
rect 49352 4868 49356 4924
rect 49356 4868 49412 4924
rect 49412 4868 49416 4924
rect 49352 4864 49416 4868
rect 44404 4660 44468 4724
rect 34468 4524 34532 4588
rect 20216 4380 20280 4384
rect 20216 4324 20220 4380
rect 20220 4324 20276 4380
rect 20276 4324 20280 4380
rect 20216 4320 20280 4324
rect 20296 4380 20360 4384
rect 20296 4324 20300 4380
rect 20300 4324 20356 4380
rect 20356 4324 20360 4380
rect 20296 4320 20360 4324
rect 20376 4380 20440 4384
rect 20376 4324 20380 4380
rect 20380 4324 20436 4380
rect 20436 4324 20440 4380
rect 20376 4320 20440 4324
rect 20456 4380 20520 4384
rect 20456 4324 20460 4380
rect 20460 4324 20516 4380
rect 20516 4324 20520 4380
rect 20456 4320 20520 4324
rect 39480 4380 39544 4384
rect 39480 4324 39484 4380
rect 39484 4324 39540 4380
rect 39540 4324 39544 4380
rect 39480 4320 39544 4324
rect 39560 4380 39624 4384
rect 39560 4324 39564 4380
rect 39564 4324 39620 4380
rect 39620 4324 39624 4380
rect 39560 4320 39624 4324
rect 39640 4380 39704 4384
rect 39640 4324 39644 4380
rect 39644 4324 39700 4380
rect 39700 4324 39704 4380
rect 39640 4320 39704 4324
rect 39720 4380 39784 4384
rect 39720 4324 39724 4380
rect 39724 4324 39780 4380
rect 39780 4324 39784 4380
rect 39720 4320 39784 4324
rect 41644 4116 41708 4180
rect 18828 3980 18892 4044
rect 10584 3836 10648 3840
rect 10584 3780 10588 3836
rect 10588 3780 10644 3836
rect 10644 3780 10648 3836
rect 10584 3776 10648 3780
rect 10664 3836 10728 3840
rect 10664 3780 10668 3836
rect 10668 3780 10724 3836
rect 10724 3780 10728 3836
rect 10664 3776 10728 3780
rect 10744 3836 10808 3840
rect 10744 3780 10748 3836
rect 10748 3780 10804 3836
rect 10804 3780 10808 3836
rect 10744 3776 10808 3780
rect 10824 3836 10888 3840
rect 10824 3780 10828 3836
rect 10828 3780 10884 3836
rect 10884 3780 10888 3836
rect 10824 3776 10888 3780
rect 29848 3836 29912 3840
rect 29848 3780 29852 3836
rect 29852 3780 29908 3836
rect 29908 3780 29912 3836
rect 29848 3776 29912 3780
rect 29928 3836 29992 3840
rect 29928 3780 29932 3836
rect 29932 3780 29988 3836
rect 29988 3780 29992 3836
rect 29928 3776 29992 3780
rect 30008 3836 30072 3840
rect 30008 3780 30012 3836
rect 30012 3780 30068 3836
rect 30068 3780 30072 3836
rect 30008 3776 30072 3780
rect 30088 3836 30152 3840
rect 30088 3780 30092 3836
rect 30092 3780 30148 3836
rect 30148 3780 30152 3836
rect 30088 3776 30152 3780
rect 49112 3836 49176 3840
rect 49112 3780 49116 3836
rect 49116 3780 49172 3836
rect 49172 3780 49176 3836
rect 49112 3776 49176 3780
rect 49192 3836 49256 3840
rect 49192 3780 49196 3836
rect 49196 3780 49252 3836
rect 49252 3780 49256 3836
rect 49192 3776 49256 3780
rect 49272 3836 49336 3840
rect 49272 3780 49276 3836
rect 49276 3780 49332 3836
rect 49332 3780 49336 3836
rect 49272 3776 49336 3780
rect 49352 3836 49416 3840
rect 49352 3780 49356 3836
rect 49356 3780 49412 3836
rect 49412 3780 49416 3836
rect 49352 3776 49416 3780
rect 26924 3572 26988 3636
rect 42932 3436 42996 3500
rect 29316 3300 29380 3364
rect 20216 3292 20280 3296
rect 20216 3236 20220 3292
rect 20220 3236 20276 3292
rect 20276 3236 20280 3292
rect 20216 3232 20280 3236
rect 20296 3292 20360 3296
rect 20296 3236 20300 3292
rect 20300 3236 20356 3292
rect 20356 3236 20360 3292
rect 20296 3232 20360 3236
rect 20376 3292 20440 3296
rect 20376 3236 20380 3292
rect 20380 3236 20436 3292
rect 20436 3236 20440 3292
rect 20376 3232 20440 3236
rect 20456 3292 20520 3296
rect 20456 3236 20460 3292
rect 20460 3236 20516 3292
rect 20516 3236 20520 3292
rect 20456 3232 20520 3236
rect 39480 3292 39544 3296
rect 39480 3236 39484 3292
rect 39484 3236 39540 3292
rect 39540 3236 39544 3292
rect 39480 3232 39544 3236
rect 39560 3292 39624 3296
rect 39560 3236 39564 3292
rect 39564 3236 39620 3292
rect 39620 3236 39624 3292
rect 39560 3232 39624 3236
rect 39640 3292 39704 3296
rect 39640 3236 39644 3292
rect 39644 3236 39700 3292
rect 39700 3236 39704 3292
rect 39640 3232 39704 3236
rect 39720 3292 39784 3296
rect 39720 3236 39724 3292
rect 39724 3236 39780 3292
rect 39780 3236 39784 3292
rect 39720 3232 39784 3236
rect 46060 2892 46124 2956
rect 10584 2748 10648 2752
rect 10584 2692 10588 2748
rect 10588 2692 10644 2748
rect 10644 2692 10648 2748
rect 10584 2688 10648 2692
rect 10664 2748 10728 2752
rect 10664 2692 10668 2748
rect 10668 2692 10724 2748
rect 10724 2692 10728 2748
rect 10664 2688 10728 2692
rect 10744 2748 10808 2752
rect 10744 2692 10748 2748
rect 10748 2692 10804 2748
rect 10804 2692 10808 2748
rect 10744 2688 10808 2692
rect 10824 2748 10888 2752
rect 10824 2692 10828 2748
rect 10828 2692 10884 2748
rect 10884 2692 10888 2748
rect 10824 2688 10888 2692
rect 29848 2748 29912 2752
rect 29848 2692 29852 2748
rect 29852 2692 29908 2748
rect 29908 2692 29912 2748
rect 29848 2688 29912 2692
rect 29928 2748 29992 2752
rect 29928 2692 29932 2748
rect 29932 2692 29988 2748
rect 29988 2692 29992 2748
rect 29928 2688 29992 2692
rect 30008 2748 30072 2752
rect 30008 2692 30012 2748
rect 30012 2692 30068 2748
rect 30068 2692 30072 2748
rect 30008 2688 30072 2692
rect 30088 2748 30152 2752
rect 30088 2692 30092 2748
rect 30092 2692 30148 2748
rect 30148 2692 30152 2748
rect 30088 2688 30152 2692
rect 49112 2748 49176 2752
rect 49112 2692 49116 2748
rect 49116 2692 49172 2748
rect 49172 2692 49176 2748
rect 49112 2688 49176 2692
rect 49192 2748 49256 2752
rect 49192 2692 49196 2748
rect 49196 2692 49252 2748
rect 49252 2692 49256 2748
rect 49192 2688 49256 2692
rect 49272 2748 49336 2752
rect 49272 2692 49276 2748
rect 49276 2692 49332 2748
rect 49332 2692 49336 2748
rect 49272 2688 49336 2692
rect 49352 2748 49416 2752
rect 49352 2692 49356 2748
rect 49356 2692 49412 2748
rect 49412 2692 49416 2748
rect 49352 2688 49416 2692
rect 46612 2484 46676 2548
rect 42748 2348 42812 2412
rect 20216 2204 20280 2208
rect 20216 2148 20220 2204
rect 20220 2148 20276 2204
rect 20276 2148 20280 2204
rect 20216 2144 20280 2148
rect 20296 2204 20360 2208
rect 20296 2148 20300 2204
rect 20300 2148 20356 2204
rect 20356 2148 20360 2204
rect 20296 2144 20360 2148
rect 20376 2204 20440 2208
rect 20376 2148 20380 2204
rect 20380 2148 20436 2204
rect 20436 2148 20440 2204
rect 20376 2144 20440 2148
rect 20456 2204 20520 2208
rect 20456 2148 20460 2204
rect 20460 2148 20516 2204
rect 20516 2148 20520 2204
rect 20456 2144 20520 2148
rect 39480 2204 39544 2208
rect 39480 2148 39484 2204
rect 39484 2148 39540 2204
rect 39540 2148 39544 2204
rect 39480 2144 39544 2148
rect 39560 2204 39624 2208
rect 39560 2148 39564 2204
rect 39564 2148 39620 2204
rect 39620 2148 39624 2204
rect 39560 2144 39624 2148
rect 39640 2204 39704 2208
rect 39640 2148 39644 2204
rect 39644 2148 39700 2204
rect 39700 2148 39704 2204
rect 39640 2144 39704 2148
rect 39720 2204 39784 2208
rect 39720 2148 39724 2204
rect 39724 2148 39780 2204
rect 39780 2148 39784 2204
rect 39720 2144 39784 2148
rect 44220 1940 44284 2004
rect 16436 1804 16500 1868
rect 35020 1804 35084 1868
rect 18092 1668 18156 1732
rect 44956 1532 45020 1596
<< metal4 >>
rect 24347 29884 24413 29885
rect 24347 29820 24348 29884
rect 24412 29820 24413 29884
rect 24347 29819 24413 29820
rect 19195 29748 19261 29749
rect 19195 29684 19196 29748
rect 19260 29684 19261 29748
rect 19195 29683 19261 29684
rect 16803 29204 16869 29205
rect 16803 29140 16804 29204
rect 16868 29140 16869 29204
rect 16803 29139 16869 29140
rect 10576 27776 10896 27792
rect 10576 27712 10584 27776
rect 10648 27712 10664 27776
rect 10728 27712 10744 27776
rect 10808 27712 10824 27776
rect 10888 27712 10896 27776
rect 10576 26688 10896 27712
rect 10576 26624 10584 26688
rect 10648 26624 10664 26688
rect 10728 26624 10744 26688
rect 10808 26624 10824 26688
rect 10888 26624 10896 26688
rect 10576 25600 10896 26624
rect 10576 25536 10584 25600
rect 10648 25536 10664 25600
rect 10728 25536 10744 25600
rect 10808 25536 10824 25600
rect 10888 25536 10896 25600
rect 10576 24512 10896 25536
rect 10576 24448 10584 24512
rect 10648 24448 10664 24512
rect 10728 24448 10744 24512
rect 10808 24448 10824 24512
rect 10888 24448 10896 24512
rect 10576 23424 10896 24448
rect 10576 23360 10584 23424
rect 10648 23360 10664 23424
rect 10728 23360 10744 23424
rect 10808 23360 10824 23424
rect 10888 23360 10896 23424
rect 10576 22336 10896 23360
rect 10576 22272 10584 22336
rect 10648 22272 10664 22336
rect 10728 22272 10744 22336
rect 10808 22272 10824 22336
rect 10888 22272 10896 22336
rect 10576 21248 10896 22272
rect 10576 21184 10584 21248
rect 10648 21184 10664 21248
rect 10728 21184 10744 21248
rect 10808 21184 10824 21248
rect 10888 21184 10896 21248
rect 10576 20160 10896 21184
rect 10576 20096 10584 20160
rect 10648 20096 10664 20160
rect 10728 20096 10744 20160
rect 10808 20096 10824 20160
rect 10888 20096 10896 20160
rect 10576 19072 10896 20096
rect 16806 19277 16866 29139
rect 17539 29068 17605 29069
rect 17539 29004 17540 29068
rect 17604 29004 17605 29068
rect 17539 29003 17605 29004
rect 16803 19276 16869 19277
rect 16803 19212 16804 19276
rect 16868 19212 16869 19276
rect 16803 19211 16869 19212
rect 17171 19276 17237 19277
rect 17171 19212 17172 19276
rect 17236 19212 17237 19276
rect 17171 19211 17237 19212
rect 10576 19008 10584 19072
rect 10648 19008 10664 19072
rect 10728 19008 10744 19072
rect 10808 19008 10824 19072
rect 10888 19008 10896 19072
rect 10576 17984 10896 19008
rect 16435 18596 16501 18597
rect 16435 18532 16436 18596
rect 16500 18532 16501 18596
rect 16435 18531 16501 18532
rect 10576 17920 10584 17984
rect 10648 17920 10664 17984
rect 10728 17920 10744 17984
rect 10808 17920 10824 17984
rect 10888 17920 10896 17984
rect 10576 16896 10896 17920
rect 10576 16832 10584 16896
rect 10648 16832 10664 16896
rect 10728 16832 10744 16896
rect 10808 16832 10824 16896
rect 10888 16832 10896 16896
rect 10576 15808 10896 16832
rect 15331 16692 15397 16693
rect 15331 16628 15332 16692
rect 15396 16628 15397 16692
rect 15331 16627 15397 16628
rect 10576 15744 10584 15808
rect 10648 15744 10664 15808
rect 10728 15744 10744 15808
rect 10808 15744 10824 15808
rect 10888 15744 10896 15808
rect 10576 14720 10896 15744
rect 10576 14656 10584 14720
rect 10648 14656 10664 14720
rect 10728 14656 10744 14720
rect 10808 14656 10824 14720
rect 10888 14656 10896 14720
rect 10576 13632 10896 14656
rect 10576 13568 10584 13632
rect 10648 13568 10664 13632
rect 10728 13568 10744 13632
rect 10808 13568 10824 13632
rect 10888 13568 10896 13632
rect 10576 12544 10896 13568
rect 10576 12480 10584 12544
rect 10648 12480 10664 12544
rect 10728 12480 10744 12544
rect 10808 12480 10824 12544
rect 10888 12480 10896 12544
rect 10576 11456 10896 12480
rect 10576 11392 10584 11456
rect 10648 11392 10664 11456
rect 10728 11392 10744 11456
rect 10808 11392 10824 11456
rect 10888 11392 10896 11456
rect 10576 10368 10896 11392
rect 10576 10304 10584 10368
rect 10648 10304 10664 10368
rect 10728 10304 10744 10368
rect 10808 10304 10824 10368
rect 10888 10304 10896 10368
rect 10576 9280 10896 10304
rect 10576 9216 10584 9280
rect 10648 9216 10664 9280
rect 10728 9216 10744 9280
rect 10808 9216 10824 9280
rect 10888 9216 10896 9280
rect 10576 8192 10896 9216
rect 15334 8261 15394 16627
rect 15331 8260 15397 8261
rect 15331 8196 15332 8260
rect 15396 8196 15397 8260
rect 15331 8195 15397 8196
rect 10576 8128 10584 8192
rect 10648 8128 10664 8192
rect 10728 8128 10744 8192
rect 10808 8128 10824 8192
rect 10888 8128 10896 8192
rect 10576 7104 10896 8128
rect 10576 7040 10584 7104
rect 10648 7040 10664 7104
rect 10728 7040 10744 7104
rect 10808 7040 10824 7104
rect 10888 7040 10896 7104
rect 10576 6016 10896 7040
rect 10576 5952 10584 6016
rect 10648 5952 10664 6016
rect 10728 5952 10744 6016
rect 10808 5952 10824 6016
rect 10888 5952 10896 6016
rect 10576 4928 10896 5952
rect 10576 4864 10584 4928
rect 10648 4864 10664 4928
rect 10728 4864 10744 4928
rect 10808 4864 10824 4928
rect 10888 4864 10896 4928
rect 10576 3840 10896 4864
rect 10576 3776 10584 3840
rect 10648 3776 10664 3840
rect 10728 3776 10744 3840
rect 10808 3776 10824 3840
rect 10888 3776 10896 3840
rect 10576 2752 10896 3776
rect 10576 2688 10584 2752
rect 10648 2688 10664 2752
rect 10728 2688 10744 2752
rect 10808 2688 10824 2752
rect 10888 2688 10896 2752
rect 10576 2128 10896 2688
rect 16438 1869 16498 18531
rect 17174 15061 17234 19211
rect 17542 17917 17602 29003
rect 19011 28252 19077 28253
rect 19011 28188 19012 28252
rect 19076 28188 19077 28252
rect 19011 28187 19077 28188
rect 19014 27630 19074 28187
rect 18646 27570 19074 27630
rect 17907 25940 17973 25941
rect 17907 25876 17908 25940
rect 17972 25876 17973 25940
rect 17907 25875 17973 25876
rect 17910 19005 17970 25875
rect 18275 21452 18341 21453
rect 18275 21388 18276 21452
rect 18340 21388 18341 21452
rect 18275 21387 18341 21388
rect 18091 19276 18157 19277
rect 18091 19212 18092 19276
rect 18156 19212 18157 19276
rect 18091 19211 18157 19212
rect 17907 19004 17973 19005
rect 17907 18940 17908 19004
rect 17972 18940 17973 19004
rect 17907 18939 17973 18940
rect 17539 17916 17605 17917
rect 17539 17852 17540 17916
rect 17604 17852 17605 17916
rect 17539 17851 17605 17852
rect 18094 17645 18154 19211
rect 18278 19005 18338 21387
rect 18646 19821 18706 27570
rect 19011 25668 19077 25669
rect 19011 25604 19012 25668
rect 19076 25604 19077 25668
rect 19011 25603 19077 25604
rect 18643 19820 18709 19821
rect 18643 19756 18644 19820
rect 18708 19756 18709 19820
rect 18643 19755 18709 19756
rect 18646 19413 18706 19755
rect 18827 19548 18893 19549
rect 18827 19484 18828 19548
rect 18892 19484 18893 19548
rect 18827 19483 18893 19484
rect 18643 19412 18709 19413
rect 18643 19348 18644 19412
rect 18708 19348 18709 19412
rect 18643 19347 18709 19348
rect 18275 19004 18341 19005
rect 18275 18940 18276 19004
rect 18340 18940 18341 19004
rect 18275 18939 18341 18940
rect 18830 17970 18890 19483
rect 19014 19141 19074 25603
rect 19198 20501 19258 29683
rect 21219 28932 21285 28933
rect 21219 28868 21220 28932
rect 21284 28868 21285 28932
rect 21219 28867 21285 28868
rect 19747 27572 19813 27573
rect 19747 27508 19748 27572
rect 19812 27508 19813 27572
rect 19747 27507 19813 27508
rect 19563 23220 19629 23221
rect 19563 23156 19564 23220
rect 19628 23156 19629 23220
rect 19563 23155 19629 23156
rect 19195 20500 19261 20501
rect 19195 20436 19196 20500
rect 19260 20436 19261 20500
rect 19195 20435 19261 20436
rect 19198 19141 19258 20435
rect 19011 19140 19077 19141
rect 19011 19076 19012 19140
rect 19076 19076 19077 19140
rect 19011 19075 19077 19076
rect 19195 19140 19261 19141
rect 19195 19076 19196 19140
rect 19260 19076 19261 19140
rect 19195 19075 19261 19076
rect 19379 18596 19445 18597
rect 19379 18532 19380 18596
rect 19444 18532 19445 18596
rect 19379 18531 19445 18532
rect 18830 17910 19074 17970
rect 18091 17644 18157 17645
rect 18091 17580 18092 17644
rect 18156 17580 18157 17644
rect 18091 17579 18157 17580
rect 17539 16692 17605 16693
rect 17539 16628 17540 16692
rect 17604 16628 17605 16692
rect 17539 16627 17605 16628
rect 18827 16692 18893 16693
rect 18827 16628 18828 16692
rect 18892 16628 18893 16692
rect 18827 16627 18893 16628
rect 17355 15332 17421 15333
rect 17355 15268 17356 15332
rect 17420 15268 17421 15332
rect 17355 15267 17421 15268
rect 17171 15060 17237 15061
rect 17171 14996 17172 15060
rect 17236 14996 17237 15060
rect 17171 14995 17237 14996
rect 17358 6357 17418 15267
rect 17542 6901 17602 16627
rect 18459 16556 18525 16557
rect 18459 16492 18460 16556
rect 18524 16492 18525 16556
rect 18459 16491 18525 16492
rect 18091 15332 18157 15333
rect 18091 15268 18092 15332
rect 18156 15268 18157 15332
rect 18091 15267 18157 15268
rect 17539 6900 17605 6901
rect 17539 6836 17540 6900
rect 17604 6836 17605 6900
rect 17539 6835 17605 6836
rect 17355 6356 17421 6357
rect 17355 6292 17356 6356
rect 17420 6292 17421 6356
rect 17355 6291 17421 6292
rect 16435 1868 16501 1869
rect 16435 1804 16436 1868
rect 16500 1804 16501 1868
rect 16435 1803 16501 1804
rect 18094 1733 18154 15267
rect 18462 6765 18522 16491
rect 18459 6764 18525 6765
rect 18459 6700 18460 6764
rect 18524 6700 18525 6764
rect 18459 6699 18525 6700
rect 18830 4045 18890 16627
rect 19014 16557 19074 17910
rect 19011 16556 19077 16557
rect 19011 16492 19012 16556
rect 19076 16492 19077 16556
rect 19011 16491 19077 16492
rect 19382 13565 19442 18531
rect 19566 14925 19626 23155
rect 19750 17370 19810 27507
rect 20208 27232 20528 27792
rect 20208 27168 20216 27232
rect 20280 27168 20296 27232
rect 20360 27168 20376 27232
rect 20440 27168 20456 27232
rect 20520 27168 20528 27232
rect 20208 26144 20528 27168
rect 20208 26080 20216 26144
rect 20280 26080 20296 26144
rect 20360 26080 20376 26144
rect 20440 26080 20456 26144
rect 20520 26080 20528 26144
rect 20208 25056 20528 26080
rect 20208 24992 20216 25056
rect 20280 24992 20296 25056
rect 20360 24992 20376 25056
rect 20440 24992 20456 25056
rect 20520 24992 20528 25056
rect 20208 23968 20528 24992
rect 20208 23904 20216 23968
rect 20280 23904 20296 23968
rect 20360 23904 20376 23968
rect 20440 23904 20456 23968
rect 20520 23904 20528 23968
rect 20208 22880 20528 23904
rect 20208 22816 20216 22880
rect 20280 22816 20296 22880
rect 20360 22816 20376 22880
rect 20440 22816 20456 22880
rect 20520 22816 20528 22880
rect 19931 22132 19997 22133
rect 19931 22068 19932 22132
rect 19996 22068 19997 22132
rect 19931 22067 19997 22068
rect 19934 19277 19994 22067
rect 20208 21792 20528 22816
rect 20667 22268 20733 22269
rect 20667 22204 20668 22268
rect 20732 22204 20733 22268
rect 20667 22203 20733 22204
rect 20208 21728 20216 21792
rect 20280 21728 20296 21792
rect 20360 21728 20376 21792
rect 20440 21728 20456 21792
rect 20520 21728 20528 21792
rect 20208 20704 20528 21728
rect 20208 20640 20216 20704
rect 20280 20640 20296 20704
rect 20360 20640 20376 20704
rect 20440 20640 20456 20704
rect 20520 20640 20528 20704
rect 20208 19616 20528 20640
rect 20670 20501 20730 22203
rect 20667 20500 20733 20501
rect 20667 20436 20668 20500
rect 20732 20436 20733 20500
rect 20667 20435 20733 20436
rect 21222 20093 21282 28867
rect 21771 28116 21837 28117
rect 21771 28052 21772 28116
rect 21836 28052 21837 28116
rect 21771 28051 21837 28052
rect 21403 23084 21469 23085
rect 21403 23020 21404 23084
rect 21468 23020 21469 23084
rect 21403 23019 21469 23020
rect 20851 20092 20917 20093
rect 20851 20028 20852 20092
rect 20916 20028 20917 20092
rect 20851 20027 20917 20028
rect 21219 20092 21285 20093
rect 21219 20028 21220 20092
rect 21284 20028 21285 20092
rect 21219 20027 21285 20028
rect 20208 19552 20216 19616
rect 20280 19552 20296 19616
rect 20360 19552 20376 19616
rect 20440 19552 20456 19616
rect 20520 19552 20528 19616
rect 19931 19276 19997 19277
rect 19931 19212 19932 19276
rect 19996 19212 19997 19276
rect 19931 19211 19997 19212
rect 20208 18528 20528 19552
rect 20667 19548 20733 19549
rect 20667 19484 20668 19548
rect 20732 19484 20733 19548
rect 20667 19483 20733 19484
rect 20208 18464 20216 18528
rect 20280 18464 20296 18528
rect 20360 18464 20376 18528
rect 20440 18464 20456 18528
rect 20520 18464 20528 18528
rect 20208 17440 20528 18464
rect 20208 17376 20216 17440
rect 20280 17376 20296 17440
rect 20360 17376 20376 17440
rect 20440 17376 20456 17440
rect 20520 17376 20528 17440
rect 19750 17310 19994 17370
rect 19747 16692 19813 16693
rect 19747 16628 19748 16692
rect 19812 16628 19813 16692
rect 19747 16627 19813 16628
rect 19563 14924 19629 14925
rect 19563 14860 19564 14924
rect 19628 14860 19629 14924
rect 19563 14859 19629 14860
rect 19379 13564 19445 13565
rect 19379 13500 19380 13564
rect 19444 13500 19445 13564
rect 19379 13499 19445 13500
rect 19750 8125 19810 16627
rect 19934 16557 19994 17310
rect 19931 16556 19997 16557
rect 19931 16492 19932 16556
rect 19996 16492 19997 16556
rect 19931 16491 19997 16492
rect 20208 16352 20528 17376
rect 20208 16288 20216 16352
rect 20280 16288 20296 16352
rect 20360 16288 20376 16352
rect 20440 16288 20456 16352
rect 20520 16288 20528 16352
rect 20208 15264 20528 16288
rect 20208 15200 20216 15264
rect 20280 15200 20296 15264
rect 20360 15200 20376 15264
rect 20440 15200 20456 15264
rect 20520 15200 20528 15264
rect 20208 14176 20528 15200
rect 20670 14925 20730 19483
rect 20854 19277 20914 20027
rect 21035 19956 21101 19957
rect 21035 19892 21036 19956
rect 21100 19892 21101 19956
rect 21035 19891 21101 19892
rect 20851 19276 20917 19277
rect 20851 19212 20852 19276
rect 20916 19212 20917 19276
rect 20851 19211 20917 19212
rect 20851 18596 20917 18597
rect 20851 18532 20852 18596
rect 20916 18532 20917 18596
rect 20851 18531 20917 18532
rect 20854 17237 20914 18531
rect 20851 17236 20917 17237
rect 20851 17172 20852 17236
rect 20916 17172 20917 17236
rect 20851 17171 20917 17172
rect 20851 16420 20917 16421
rect 20851 16356 20852 16420
rect 20916 16356 20917 16420
rect 20851 16355 20917 16356
rect 20667 14924 20733 14925
rect 20667 14860 20668 14924
rect 20732 14860 20733 14924
rect 20667 14859 20733 14860
rect 20208 14112 20216 14176
rect 20280 14112 20296 14176
rect 20360 14112 20376 14176
rect 20440 14112 20456 14176
rect 20520 14112 20528 14176
rect 20208 13088 20528 14112
rect 20208 13024 20216 13088
rect 20280 13024 20296 13088
rect 20360 13024 20376 13088
rect 20440 13024 20456 13088
rect 20520 13024 20528 13088
rect 20208 12000 20528 13024
rect 20670 12749 20730 14859
rect 20667 12748 20733 12749
rect 20667 12684 20668 12748
rect 20732 12684 20733 12748
rect 20667 12683 20733 12684
rect 20208 11936 20216 12000
rect 20280 11936 20296 12000
rect 20360 11936 20376 12000
rect 20440 11936 20456 12000
rect 20520 11936 20528 12000
rect 20208 10912 20528 11936
rect 20670 11389 20730 12683
rect 20854 12069 20914 16355
rect 21038 16149 21098 19891
rect 21219 17780 21285 17781
rect 21219 17716 21220 17780
rect 21284 17716 21285 17780
rect 21219 17715 21285 17716
rect 21035 16148 21101 16149
rect 21035 16084 21036 16148
rect 21100 16084 21101 16148
rect 21035 16083 21101 16084
rect 21038 13701 21098 16083
rect 21035 13700 21101 13701
rect 21035 13636 21036 13700
rect 21100 13636 21101 13700
rect 21035 13635 21101 13636
rect 21222 13021 21282 17715
rect 21406 13973 21466 23019
rect 21587 22404 21653 22405
rect 21587 22340 21588 22404
rect 21652 22340 21653 22404
rect 21587 22339 21653 22340
rect 21590 16149 21650 22339
rect 21774 21861 21834 28051
rect 21955 26348 22021 26349
rect 21955 26284 21956 26348
rect 22020 26284 22021 26348
rect 21955 26283 22021 26284
rect 21771 21860 21837 21861
rect 21771 21796 21772 21860
rect 21836 21796 21837 21860
rect 21771 21795 21837 21796
rect 21958 17917 22018 26283
rect 22323 23492 22389 23493
rect 22323 23428 22324 23492
rect 22388 23428 22389 23492
rect 22323 23427 22389 23428
rect 22326 20090 22386 23427
rect 24163 22540 24229 22541
rect 24163 22476 24164 22540
rect 24228 22476 24229 22540
rect 24163 22475 24229 22476
rect 22691 21588 22757 21589
rect 22691 21524 22692 21588
rect 22756 21524 22757 21588
rect 22691 21523 22757 21524
rect 22694 20773 22754 21523
rect 22691 20772 22757 20773
rect 22691 20708 22692 20772
rect 22756 20708 22757 20772
rect 22691 20707 22757 20708
rect 22326 20030 22570 20090
rect 22139 19412 22205 19413
rect 22139 19348 22140 19412
rect 22204 19348 22205 19412
rect 22139 19347 22205 19348
rect 21955 17916 22021 17917
rect 21955 17852 21956 17916
rect 22020 17852 22021 17916
rect 21955 17851 22021 17852
rect 22142 16285 22202 19347
rect 22139 16284 22205 16285
rect 22139 16220 22140 16284
rect 22204 16220 22205 16284
rect 22139 16219 22205 16220
rect 21587 16148 21653 16149
rect 21587 16084 21588 16148
rect 21652 16084 21653 16148
rect 21587 16083 21653 16084
rect 21771 15332 21837 15333
rect 21771 15330 21772 15332
rect 21590 15270 21772 15330
rect 21403 13972 21469 13973
rect 21403 13908 21404 13972
rect 21468 13908 21469 13972
rect 21403 13907 21469 13908
rect 21219 13020 21285 13021
rect 21219 12956 21220 13020
rect 21284 12956 21285 13020
rect 21219 12955 21285 12956
rect 20851 12068 20917 12069
rect 20851 12004 20852 12068
rect 20916 12004 20917 12068
rect 20851 12003 20917 12004
rect 21222 11525 21282 12955
rect 21590 12477 21650 15270
rect 21771 15268 21772 15270
rect 21836 15268 21837 15332
rect 21771 15267 21837 15268
rect 22139 15332 22205 15333
rect 22139 15268 22140 15332
rect 22204 15268 22205 15332
rect 22139 15267 22205 15268
rect 21771 14108 21837 14109
rect 21771 14044 21772 14108
rect 21836 14044 21837 14108
rect 21771 14043 21837 14044
rect 21587 12476 21653 12477
rect 21587 12412 21588 12476
rect 21652 12412 21653 12476
rect 21587 12411 21653 12412
rect 21219 11524 21285 11525
rect 21219 11460 21220 11524
rect 21284 11460 21285 11524
rect 21219 11459 21285 11460
rect 20667 11388 20733 11389
rect 20667 11324 20668 11388
rect 20732 11324 20733 11388
rect 20667 11323 20733 11324
rect 20208 10848 20216 10912
rect 20280 10848 20296 10912
rect 20360 10848 20376 10912
rect 20440 10848 20456 10912
rect 20520 10848 20528 10912
rect 20208 9824 20528 10848
rect 20208 9760 20216 9824
rect 20280 9760 20296 9824
rect 20360 9760 20376 9824
rect 20440 9760 20456 9824
rect 20520 9760 20528 9824
rect 20208 8736 20528 9760
rect 20208 8672 20216 8736
rect 20280 8672 20296 8736
rect 20360 8672 20376 8736
rect 20440 8672 20456 8736
rect 20520 8672 20528 8736
rect 19747 8124 19813 8125
rect 19747 8060 19748 8124
rect 19812 8060 19813 8124
rect 19747 8059 19813 8060
rect 20208 7648 20528 8672
rect 21774 7853 21834 14043
rect 21955 13972 22021 13973
rect 21955 13908 21956 13972
rect 22020 13908 22021 13972
rect 21955 13907 22021 13908
rect 21958 9757 22018 13907
rect 22142 11389 22202 15267
rect 22326 14109 22386 20030
rect 22510 19957 22570 20030
rect 22507 19956 22573 19957
rect 22507 19892 22508 19956
rect 22572 19892 22573 19956
rect 22507 19891 22573 19892
rect 23427 15604 23493 15605
rect 23427 15540 23428 15604
rect 23492 15540 23493 15604
rect 23427 15539 23493 15540
rect 22323 14108 22389 14109
rect 22323 14044 22324 14108
rect 22388 14044 22389 14108
rect 22323 14043 22389 14044
rect 22139 11388 22205 11389
rect 22139 11324 22140 11388
rect 22204 11324 22205 11388
rect 22139 11323 22205 11324
rect 21955 9756 22021 9757
rect 21955 9692 21956 9756
rect 22020 9692 22021 9756
rect 21955 9691 22021 9692
rect 23430 8669 23490 15539
rect 23979 14924 24045 14925
rect 23979 14860 23980 14924
rect 24044 14860 24045 14924
rect 23979 14859 24045 14860
rect 23982 11117 24042 14859
rect 24166 11389 24226 22475
rect 24350 22405 24410 29819
rect 40171 29340 40237 29341
rect 40171 29276 40172 29340
rect 40236 29276 40237 29340
rect 40171 29275 40237 29276
rect 37595 28388 37661 28389
rect 37595 28324 37596 28388
rect 37660 28324 37661 28388
rect 37595 28323 37661 28324
rect 29840 27776 30160 27792
rect 29840 27712 29848 27776
rect 29912 27712 29928 27776
rect 29992 27712 30008 27776
rect 30072 27712 30088 27776
rect 30152 27712 30160 27776
rect 29840 26688 30160 27712
rect 29840 26624 29848 26688
rect 29912 26624 29928 26688
rect 29992 26624 30008 26688
rect 30072 26624 30088 26688
rect 30152 26624 30160 26688
rect 29840 25600 30160 26624
rect 37411 26620 37477 26621
rect 37411 26556 37412 26620
rect 37476 26556 37477 26620
rect 37411 26555 37477 26556
rect 30787 26348 30853 26349
rect 30787 26284 30788 26348
rect 30852 26284 30853 26348
rect 30787 26283 30853 26284
rect 32627 26348 32693 26349
rect 32627 26284 32628 26348
rect 32692 26284 32693 26348
rect 32627 26283 32693 26284
rect 29840 25536 29848 25600
rect 29912 25536 29928 25600
rect 29992 25536 30008 25600
rect 30072 25536 30088 25600
rect 30152 25536 30160 25600
rect 27475 25532 27541 25533
rect 27475 25468 27476 25532
rect 27540 25468 27541 25532
rect 27475 25467 27541 25468
rect 25267 25260 25333 25261
rect 25267 25196 25268 25260
rect 25332 25196 25333 25260
rect 25267 25195 25333 25196
rect 24899 23764 24965 23765
rect 24899 23700 24900 23764
rect 24964 23700 24965 23764
rect 24899 23699 24965 23700
rect 24715 23492 24781 23493
rect 24715 23428 24716 23492
rect 24780 23428 24781 23492
rect 24715 23427 24781 23428
rect 24347 22404 24413 22405
rect 24347 22340 24348 22404
rect 24412 22340 24413 22404
rect 24347 22339 24413 22340
rect 24350 21725 24410 22339
rect 24347 21724 24413 21725
rect 24347 21660 24348 21724
rect 24412 21660 24413 21724
rect 24347 21659 24413 21660
rect 24718 17917 24778 23427
rect 24902 21861 24962 23699
rect 25083 22540 25149 22541
rect 25083 22476 25084 22540
rect 25148 22476 25149 22540
rect 25083 22475 25149 22476
rect 24899 21860 24965 21861
rect 24899 21796 24900 21860
rect 24964 21796 24965 21860
rect 24899 21795 24965 21796
rect 25086 19141 25146 22475
rect 25270 19277 25330 25195
rect 25819 24036 25885 24037
rect 25819 23972 25820 24036
rect 25884 23972 25885 24036
rect 25819 23971 25885 23972
rect 27291 24036 27357 24037
rect 27291 23972 27292 24036
rect 27356 23972 27357 24036
rect 27291 23971 27357 23972
rect 25822 22677 25882 23971
rect 27107 23764 27173 23765
rect 27107 23700 27108 23764
rect 27172 23700 27173 23764
rect 27107 23699 27173 23700
rect 25819 22676 25885 22677
rect 25819 22612 25820 22676
rect 25884 22612 25885 22676
rect 25819 22611 25885 22612
rect 26555 21588 26621 21589
rect 26555 21524 26556 21588
rect 26620 21524 26621 21588
rect 26555 21523 26621 21524
rect 25267 19276 25333 19277
rect 25267 19212 25268 19276
rect 25332 19212 25333 19276
rect 25267 19211 25333 19212
rect 25083 19140 25149 19141
rect 25083 19076 25084 19140
rect 25148 19076 25149 19140
rect 25083 19075 25149 19076
rect 24715 17916 24781 17917
rect 24715 17852 24716 17916
rect 24780 17852 24781 17916
rect 24715 17851 24781 17852
rect 26371 16692 26437 16693
rect 26371 16628 26372 16692
rect 26436 16628 26437 16692
rect 26371 16627 26437 16628
rect 25451 16556 25517 16557
rect 25451 16492 25452 16556
rect 25516 16492 25517 16556
rect 25451 16491 25517 16492
rect 24531 16148 24597 16149
rect 24531 16084 24532 16148
rect 24596 16084 24597 16148
rect 24531 16083 24597 16084
rect 24534 12341 24594 16083
rect 24715 13836 24781 13837
rect 24715 13772 24716 13836
rect 24780 13772 24781 13836
rect 24715 13771 24781 13772
rect 24899 13836 24965 13837
rect 24899 13772 24900 13836
rect 24964 13772 24965 13836
rect 24899 13771 24965 13772
rect 24531 12340 24597 12341
rect 24531 12276 24532 12340
rect 24596 12276 24597 12340
rect 24531 12275 24597 12276
rect 24163 11388 24229 11389
rect 24163 11324 24164 11388
rect 24228 11324 24229 11388
rect 24163 11323 24229 11324
rect 23979 11116 24045 11117
rect 23979 11052 23980 11116
rect 24044 11052 24045 11116
rect 23979 11051 24045 11052
rect 23427 8668 23493 8669
rect 23427 8604 23428 8668
rect 23492 8604 23493 8668
rect 23427 8603 23493 8604
rect 24718 8125 24778 13771
rect 24902 9485 24962 13771
rect 25267 13292 25333 13293
rect 25267 13228 25268 13292
rect 25332 13228 25333 13292
rect 25267 13227 25333 13228
rect 25270 10029 25330 13227
rect 25454 11389 25514 16491
rect 26374 13021 26434 16627
rect 26558 16557 26618 21523
rect 27110 20501 27170 23699
rect 27107 20500 27173 20501
rect 27107 20436 27108 20500
rect 27172 20436 27173 20500
rect 27107 20435 27173 20436
rect 27110 19685 27170 20435
rect 27107 19684 27173 19685
rect 27107 19620 27108 19684
rect 27172 19620 27173 19684
rect 27107 19619 27173 19620
rect 27107 19548 27173 19549
rect 27107 19484 27108 19548
rect 27172 19484 27173 19548
rect 27107 19483 27173 19484
rect 26555 16556 26621 16557
rect 26555 16492 26556 16556
rect 26620 16492 26621 16556
rect 26555 16491 26621 16492
rect 26371 13020 26437 13021
rect 26371 12956 26372 13020
rect 26436 12956 26437 13020
rect 26371 12955 26437 12956
rect 25819 12748 25885 12749
rect 25819 12684 25820 12748
rect 25884 12684 25885 12748
rect 25819 12683 25885 12684
rect 25451 11388 25517 11389
rect 25451 11324 25452 11388
rect 25516 11324 25517 11388
rect 25451 11323 25517 11324
rect 25267 10028 25333 10029
rect 25267 9964 25268 10028
rect 25332 9964 25333 10028
rect 25267 9963 25333 9964
rect 24899 9484 24965 9485
rect 24899 9420 24900 9484
rect 24964 9420 24965 9484
rect 24899 9419 24965 9420
rect 25822 8125 25882 12683
rect 26558 9213 26618 16491
rect 27110 11389 27170 19483
rect 27294 19413 27354 23971
rect 27478 21589 27538 25467
rect 28211 25396 28277 25397
rect 28211 25332 28212 25396
rect 28276 25332 28277 25396
rect 28211 25331 28277 25332
rect 28027 23900 28093 23901
rect 28027 23836 28028 23900
rect 28092 23836 28093 23900
rect 28027 23835 28093 23836
rect 27843 23084 27909 23085
rect 27843 23020 27844 23084
rect 27908 23020 27909 23084
rect 27843 23019 27909 23020
rect 27846 21725 27906 23019
rect 27843 21724 27909 21725
rect 27843 21660 27844 21724
rect 27908 21660 27909 21724
rect 27843 21659 27909 21660
rect 27475 21588 27541 21589
rect 27475 21524 27476 21588
rect 27540 21524 27541 21588
rect 27475 21523 27541 21524
rect 27843 19820 27909 19821
rect 27843 19756 27844 19820
rect 27908 19756 27909 19820
rect 27843 19755 27909 19756
rect 27291 19412 27357 19413
rect 27291 19348 27292 19412
rect 27356 19348 27357 19412
rect 27291 19347 27357 19348
rect 27475 14924 27541 14925
rect 27475 14860 27476 14924
rect 27540 14860 27541 14924
rect 27475 14859 27541 14860
rect 27107 11388 27173 11389
rect 27107 11324 27108 11388
rect 27172 11324 27173 11388
rect 27107 11323 27173 11324
rect 26923 11116 26989 11117
rect 26923 11052 26924 11116
rect 26988 11052 26989 11116
rect 26923 11051 26989 11052
rect 26555 9212 26621 9213
rect 26555 9148 26556 9212
rect 26620 9148 26621 9212
rect 26555 9147 26621 9148
rect 24715 8124 24781 8125
rect 24715 8060 24716 8124
rect 24780 8060 24781 8124
rect 24715 8059 24781 8060
rect 25819 8124 25885 8125
rect 25819 8060 25820 8124
rect 25884 8060 25885 8124
rect 25819 8059 25885 8060
rect 21771 7852 21837 7853
rect 21771 7788 21772 7852
rect 21836 7788 21837 7852
rect 21771 7787 21837 7788
rect 20208 7584 20216 7648
rect 20280 7584 20296 7648
rect 20360 7584 20376 7648
rect 20440 7584 20456 7648
rect 20520 7584 20528 7648
rect 20208 6560 20528 7584
rect 20208 6496 20216 6560
rect 20280 6496 20296 6560
rect 20360 6496 20376 6560
rect 20440 6496 20456 6560
rect 20520 6496 20528 6560
rect 20208 5472 20528 6496
rect 20208 5408 20216 5472
rect 20280 5408 20296 5472
rect 20360 5408 20376 5472
rect 20440 5408 20456 5472
rect 20520 5408 20528 5472
rect 20208 4384 20528 5408
rect 20208 4320 20216 4384
rect 20280 4320 20296 4384
rect 20360 4320 20376 4384
rect 20440 4320 20456 4384
rect 20520 4320 20528 4384
rect 18827 4044 18893 4045
rect 18827 3980 18828 4044
rect 18892 3980 18893 4044
rect 18827 3979 18893 3980
rect 20208 3296 20528 4320
rect 26926 3637 26986 11051
rect 27478 9077 27538 14859
rect 27659 13020 27725 13021
rect 27659 12956 27660 13020
rect 27724 12956 27725 13020
rect 27659 12955 27725 12956
rect 27475 9076 27541 9077
rect 27475 9012 27476 9076
rect 27540 9012 27541 9076
rect 27475 9011 27541 9012
rect 27662 8397 27722 12955
rect 27846 12749 27906 19755
rect 28030 19413 28090 23835
rect 28027 19412 28093 19413
rect 28027 19348 28028 19412
rect 28092 19348 28093 19412
rect 28027 19347 28093 19348
rect 28214 16421 28274 25331
rect 28395 25260 28461 25261
rect 28395 25196 28396 25260
rect 28460 25196 28461 25260
rect 28395 25195 28461 25196
rect 29683 25260 29749 25261
rect 29683 25196 29684 25260
rect 29748 25196 29749 25260
rect 29683 25195 29749 25196
rect 28398 22813 28458 25195
rect 29315 25124 29381 25125
rect 29315 25060 29316 25124
rect 29380 25060 29381 25124
rect 29315 25059 29381 25060
rect 28763 24580 28829 24581
rect 28763 24516 28764 24580
rect 28828 24516 28829 24580
rect 28763 24515 28829 24516
rect 28579 24172 28645 24173
rect 28579 24108 28580 24172
rect 28644 24108 28645 24172
rect 28579 24107 28645 24108
rect 28395 22812 28461 22813
rect 28395 22748 28396 22812
rect 28460 22748 28461 22812
rect 28395 22747 28461 22748
rect 28582 22677 28642 24107
rect 28579 22676 28645 22677
rect 28579 22612 28580 22676
rect 28644 22612 28645 22676
rect 28579 22611 28645 22612
rect 28395 20364 28461 20365
rect 28395 20300 28396 20364
rect 28460 20300 28461 20364
rect 28395 20299 28461 20300
rect 28398 19350 28458 20299
rect 28766 19957 28826 24515
rect 29318 24445 29378 25059
rect 29315 24444 29381 24445
rect 29315 24380 29316 24444
rect 29380 24380 29381 24444
rect 29315 24379 29381 24380
rect 29131 22676 29197 22677
rect 29131 22612 29132 22676
rect 29196 22612 29197 22676
rect 29131 22611 29197 22612
rect 29134 22266 29194 22611
rect 29318 22405 29378 24379
rect 29315 22404 29381 22405
rect 29315 22340 29316 22404
rect 29380 22340 29381 22404
rect 29315 22339 29381 22340
rect 29499 22268 29565 22269
rect 29134 22206 29378 22266
rect 29131 21996 29197 21997
rect 29131 21932 29132 21996
rect 29196 21932 29197 21996
rect 29131 21931 29197 21932
rect 28763 19956 28829 19957
rect 28763 19892 28764 19956
rect 28828 19892 28829 19956
rect 28763 19891 28829 19892
rect 28398 19290 28642 19350
rect 28211 16420 28277 16421
rect 28211 16356 28212 16420
rect 28276 16356 28277 16420
rect 28211 16355 28277 16356
rect 28027 14244 28093 14245
rect 28027 14180 28028 14244
rect 28092 14180 28093 14244
rect 28027 14179 28093 14180
rect 28395 14244 28461 14245
rect 28395 14180 28396 14244
rect 28460 14180 28461 14244
rect 28395 14179 28461 14180
rect 27843 12748 27909 12749
rect 27843 12684 27844 12748
rect 27908 12684 27909 12748
rect 27843 12683 27909 12684
rect 28030 12613 28090 14179
rect 28027 12612 28093 12613
rect 28027 12548 28028 12612
rect 28092 12548 28093 12612
rect 28027 12547 28093 12548
rect 27659 8396 27725 8397
rect 27659 8332 27660 8396
rect 27724 8332 27725 8396
rect 27659 8331 27725 8332
rect 28398 6493 28458 14179
rect 28582 12069 28642 19290
rect 28947 15604 29013 15605
rect 28947 15540 28948 15604
rect 29012 15540 29013 15604
rect 28947 15539 29013 15540
rect 28763 15332 28829 15333
rect 28763 15268 28764 15332
rect 28828 15268 28829 15332
rect 28763 15267 28829 15268
rect 28579 12068 28645 12069
rect 28579 12004 28580 12068
rect 28644 12004 28645 12068
rect 28579 12003 28645 12004
rect 28582 11389 28642 12003
rect 28579 11388 28645 11389
rect 28579 11324 28580 11388
rect 28644 11324 28645 11388
rect 28579 11323 28645 11324
rect 28766 7445 28826 15267
rect 28950 13837 29010 15539
rect 28947 13836 29013 13837
rect 28947 13772 28948 13836
rect 29012 13772 29013 13836
rect 28947 13771 29013 13772
rect 28947 11116 29013 11117
rect 28947 11052 28948 11116
rect 29012 11052 29013 11116
rect 28947 11051 29013 11052
rect 28950 8397 29010 11051
rect 29134 10709 29194 21931
rect 29318 11797 29378 22206
rect 29499 22204 29500 22268
rect 29564 22204 29565 22268
rect 29499 22203 29565 22204
rect 29502 21453 29562 22203
rect 29499 21452 29565 21453
rect 29499 21388 29500 21452
rect 29564 21388 29565 21452
rect 29499 21387 29565 21388
rect 29499 19548 29565 19549
rect 29499 19484 29500 19548
rect 29564 19484 29565 19548
rect 29499 19483 29565 19484
rect 29502 19141 29562 19483
rect 29499 19140 29565 19141
rect 29499 19076 29500 19140
rect 29564 19076 29565 19140
rect 29499 19075 29565 19076
rect 29502 15877 29562 19075
rect 29686 18869 29746 25195
rect 29840 24512 30160 25536
rect 29840 24448 29848 24512
rect 29912 24448 29928 24512
rect 29992 24448 30008 24512
rect 30072 24448 30088 24512
rect 30152 24448 30160 24512
rect 29840 23424 30160 24448
rect 30419 23628 30485 23629
rect 30419 23564 30420 23628
rect 30484 23564 30485 23628
rect 30419 23563 30485 23564
rect 29840 23360 29848 23424
rect 29912 23360 29928 23424
rect 29992 23360 30008 23424
rect 30072 23360 30088 23424
rect 30152 23360 30160 23424
rect 29840 22336 30160 23360
rect 29840 22272 29848 22336
rect 29912 22272 29928 22336
rect 29992 22272 30008 22336
rect 30072 22272 30088 22336
rect 30152 22272 30160 22336
rect 29840 21248 30160 22272
rect 29840 21184 29848 21248
rect 29912 21184 29928 21248
rect 29992 21184 30008 21248
rect 30072 21184 30088 21248
rect 30152 21184 30160 21248
rect 29840 20160 30160 21184
rect 29840 20096 29848 20160
rect 29912 20096 29928 20160
rect 29992 20096 30008 20160
rect 30072 20096 30088 20160
rect 30152 20096 30160 20160
rect 29840 19072 30160 20096
rect 29840 19008 29848 19072
rect 29912 19008 29928 19072
rect 29992 19008 30008 19072
rect 30072 19008 30088 19072
rect 30152 19008 30160 19072
rect 29683 18868 29749 18869
rect 29683 18804 29684 18868
rect 29748 18804 29749 18868
rect 29683 18803 29749 18804
rect 29683 18052 29749 18053
rect 29683 17988 29684 18052
rect 29748 17988 29749 18052
rect 29683 17987 29749 17988
rect 29499 15876 29565 15877
rect 29499 15812 29500 15876
rect 29564 15812 29565 15876
rect 29499 15811 29565 15812
rect 29499 12612 29565 12613
rect 29499 12548 29500 12612
rect 29564 12548 29565 12612
rect 29499 12547 29565 12548
rect 29315 11796 29381 11797
rect 29315 11732 29316 11796
rect 29380 11732 29381 11796
rect 29315 11731 29381 11732
rect 29315 11524 29381 11525
rect 29315 11460 29316 11524
rect 29380 11460 29381 11524
rect 29315 11459 29381 11460
rect 29131 10708 29197 10709
rect 29131 10644 29132 10708
rect 29196 10644 29197 10708
rect 29131 10643 29197 10644
rect 28947 8396 29013 8397
rect 28947 8332 28948 8396
rect 29012 8332 29013 8396
rect 28947 8331 29013 8332
rect 28763 7444 28829 7445
rect 28763 7380 28764 7444
rect 28828 7380 28829 7444
rect 28763 7379 28829 7380
rect 28395 6492 28461 6493
rect 28395 6428 28396 6492
rect 28460 6428 28461 6492
rect 28395 6427 28461 6428
rect 26923 3636 26989 3637
rect 26923 3572 26924 3636
rect 26988 3572 26989 3636
rect 26923 3571 26989 3572
rect 29318 3365 29378 11459
rect 29502 8261 29562 12547
rect 29686 9621 29746 17987
rect 29840 17984 30160 19008
rect 29840 17920 29848 17984
rect 29912 17920 29928 17984
rect 29992 17920 30008 17984
rect 30072 17920 30088 17984
rect 30152 17920 30160 17984
rect 29840 16896 30160 17920
rect 29840 16832 29848 16896
rect 29912 16832 29928 16896
rect 29992 16832 30008 16896
rect 30072 16832 30088 16896
rect 30152 16832 30160 16896
rect 29840 15808 30160 16832
rect 29840 15744 29848 15808
rect 29912 15744 29928 15808
rect 29992 15744 30008 15808
rect 30072 15744 30088 15808
rect 30152 15744 30160 15808
rect 29840 14720 30160 15744
rect 30235 14788 30301 14789
rect 30235 14724 30236 14788
rect 30300 14724 30301 14788
rect 30235 14723 30301 14724
rect 29840 14656 29848 14720
rect 29912 14656 29928 14720
rect 29992 14656 30008 14720
rect 30072 14656 30088 14720
rect 30152 14656 30160 14720
rect 29840 13632 30160 14656
rect 29840 13568 29848 13632
rect 29912 13568 29928 13632
rect 29992 13568 30008 13632
rect 30072 13568 30088 13632
rect 30152 13568 30160 13632
rect 29840 12544 30160 13568
rect 29840 12480 29848 12544
rect 29912 12480 29928 12544
rect 29992 12480 30008 12544
rect 30072 12480 30088 12544
rect 30152 12480 30160 12544
rect 29840 11456 30160 12480
rect 30238 12069 30298 14723
rect 30235 12068 30301 12069
rect 30235 12004 30236 12068
rect 30300 12004 30301 12068
rect 30235 12003 30301 12004
rect 30422 11661 30482 23563
rect 30603 23084 30669 23085
rect 30603 23020 30604 23084
rect 30668 23020 30669 23084
rect 30603 23019 30669 23020
rect 30606 19005 30666 23019
rect 30790 21317 30850 26283
rect 30971 23628 31037 23629
rect 30971 23564 30972 23628
rect 31036 23564 31037 23628
rect 30971 23563 31037 23564
rect 30974 21725 31034 23563
rect 30971 21724 31037 21725
rect 30971 21660 30972 21724
rect 31036 21660 31037 21724
rect 30971 21659 31037 21660
rect 30787 21316 30853 21317
rect 30787 21252 30788 21316
rect 30852 21252 30853 21316
rect 30787 21251 30853 21252
rect 30787 20772 30853 20773
rect 30787 20708 30788 20772
rect 30852 20708 30853 20772
rect 30787 20707 30853 20708
rect 30603 19004 30669 19005
rect 30603 18940 30604 19004
rect 30668 18940 30669 19004
rect 30603 18939 30669 18940
rect 30603 15332 30669 15333
rect 30603 15268 30604 15332
rect 30668 15268 30669 15332
rect 30603 15267 30669 15268
rect 30419 11660 30485 11661
rect 30419 11596 30420 11660
rect 30484 11596 30485 11660
rect 30419 11595 30485 11596
rect 30235 11524 30301 11525
rect 30235 11460 30236 11524
rect 30300 11460 30301 11524
rect 30235 11459 30301 11460
rect 29840 11392 29848 11456
rect 29912 11392 29928 11456
rect 29992 11392 30008 11456
rect 30072 11392 30088 11456
rect 30152 11392 30160 11456
rect 29840 10368 30160 11392
rect 29840 10304 29848 10368
rect 29912 10304 29928 10368
rect 29992 10304 30008 10368
rect 30072 10304 30088 10368
rect 30152 10304 30160 10368
rect 29683 9620 29749 9621
rect 29683 9556 29684 9620
rect 29748 9556 29749 9620
rect 29683 9555 29749 9556
rect 29840 9280 30160 10304
rect 30238 9757 30298 11459
rect 30235 9756 30301 9757
rect 30235 9692 30236 9756
rect 30300 9692 30301 9756
rect 30235 9691 30301 9692
rect 29840 9216 29848 9280
rect 29912 9216 29928 9280
rect 29992 9216 30008 9280
rect 30072 9216 30088 9280
rect 30152 9216 30160 9280
rect 29499 8260 29565 8261
rect 29499 8196 29500 8260
rect 29564 8196 29565 8260
rect 29499 8195 29565 8196
rect 29502 5405 29562 8195
rect 29840 8192 30160 9216
rect 30606 8805 30666 15267
rect 30790 14789 30850 20707
rect 30974 16149 31034 21659
rect 32259 20772 32325 20773
rect 32259 20708 32260 20772
rect 32324 20708 32325 20772
rect 32259 20707 32325 20708
rect 31891 16828 31957 16829
rect 31891 16764 31892 16828
rect 31956 16764 31957 16828
rect 31891 16763 31957 16764
rect 30971 16148 31037 16149
rect 30971 16084 30972 16148
rect 31036 16084 31037 16148
rect 30971 16083 31037 16084
rect 30787 14788 30853 14789
rect 30787 14724 30788 14788
rect 30852 14724 30853 14788
rect 30787 14723 30853 14724
rect 30790 14517 30850 14723
rect 30787 14516 30853 14517
rect 30787 14452 30788 14516
rect 30852 14452 30853 14516
rect 30787 14451 30853 14452
rect 30971 12748 31037 12749
rect 30971 12684 30972 12748
rect 31036 12684 31037 12748
rect 30971 12683 31037 12684
rect 30974 9485 31034 12683
rect 31894 12341 31954 16763
rect 32075 16012 32141 16013
rect 32075 15948 32076 16012
rect 32140 15948 32141 16012
rect 32075 15947 32141 15948
rect 31891 12340 31957 12341
rect 31891 12276 31892 12340
rect 31956 12276 31957 12340
rect 31891 12275 31957 12276
rect 32078 9757 32138 15947
rect 32075 9756 32141 9757
rect 32075 9692 32076 9756
rect 32140 9692 32141 9756
rect 32075 9691 32141 9692
rect 32262 9485 32322 20707
rect 32630 18461 32690 26283
rect 34283 24988 34349 24989
rect 34283 24924 34284 24988
rect 34348 24924 34349 24988
rect 34283 24923 34349 24924
rect 33363 24580 33429 24581
rect 33363 24516 33364 24580
rect 33428 24516 33429 24580
rect 33363 24515 33429 24516
rect 32995 23900 33061 23901
rect 32995 23836 32996 23900
rect 33060 23836 33061 23900
rect 32995 23835 33061 23836
rect 32627 18460 32693 18461
rect 32627 18396 32628 18460
rect 32692 18396 32693 18460
rect 32627 18395 32693 18396
rect 32443 16964 32509 16965
rect 32443 16900 32444 16964
rect 32508 16900 32509 16964
rect 32443 16899 32509 16900
rect 32446 9621 32506 16899
rect 32811 11116 32877 11117
rect 32811 11052 32812 11116
rect 32876 11052 32877 11116
rect 32811 11051 32877 11052
rect 32443 9620 32509 9621
rect 32443 9556 32444 9620
rect 32508 9556 32509 9620
rect 32443 9555 32509 9556
rect 30971 9484 31037 9485
rect 30971 9420 30972 9484
rect 31036 9420 31037 9484
rect 30971 9419 31037 9420
rect 32259 9484 32325 9485
rect 32259 9420 32260 9484
rect 32324 9420 32325 9484
rect 32259 9419 32325 9420
rect 30603 8804 30669 8805
rect 30603 8740 30604 8804
rect 30668 8740 30669 8804
rect 30603 8739 30669 8740
rect 29840 8128 29848 8192
rect 29912 8128 29928 8192
rect 29992 8128 30008 8192
rect 30072 8128 30088 8192
rect 30152 8128 30160 8192
rect 29840 7104 30160 8128
rect 30235 7580 30301 7581
rect 30235 7516 30236 7580
rect 30300 7516 30301 7580
rect 30235 7515 30301 7516
rect 29840 7040 29848 7104
rect 29912 7040 29928 7104
rect 29992 7040 30008 7104
rect 30072 7040 30088 7104
rect 30152 7040 30160 7104
rect 29840 6016 30160 7040
rect 30238 6221 30298 7515
rect 32814 6901 32874 11051
rect 32998 9757 33058 23835
rect 33179 23492 33245 23493
rect 33179 23428 33180 23492
rect 33244 23428 33245 23492
rect 33179 23427 33245 23428
rect 33182 18325 33242 23427
rect 33366 21725 33426 24515
rect 33731 21996 33797 21997
rect 33731 21932 33732 21996
rect 33796 21932 33797 21996
rect 33731 21931 33797 21932
rect 33363 21724 33429 21725
rect 33363 21660 33364 21724
rect 33428 21660 33429 21724
rect 33363 21659 33429 21660
rect 33734 19277 33794 21931
rect 34286 20093 34346 24923
rect 36675 24580 36741 24581
rect 36675 24516 36676 24580
rect 36740 24516 36741 24580
rect 36675 24515 36741 24516
rect 34835 23900 34901 23901
rect 34835 23836 34836 23900
rect 34900 23836 34901 23900
rect 34835 23835 34901 23836
rect 34651 22540 34717 22541
rect 34651 22476 34652 22540
rect 34716 22476 34717 22540
rect 34651 22475 34717 22476
rect 34467 22404 34533 22405
rect 34467 22340 34468 22404
rect 34532 22340 34533 22404
rect 34467 22339 34533 22340
rect 34283 20092 34349 20093
rect 34283 20028 34284 20092
rect 34348 20028 34349 20092
rect 34283 20027 34349 20028
rect 33731 19276 33797 19277
rect 33731 19212 33732 19276
rect 33796 19212 33797 19276
rect 33731 19211 33797 19212
rect 34099 18732 34165 18733
rect 34099 18668 34100 18732
rect 34164 18668 34165 18732
rect 34099 18667 34165 18668
rect 33179 18324 33245 18325
rect 33179 18260 33180 18324
rect 33244 18260 33245 18324
rect 33179 18259 33245 18260
rect 33179 14652 33245 14653
rect 33179 14588 33180 14652
rect 33244 14588 33245 14652
rect 33179 14587 33245 14588
rect 33182 10981 33242 14587
rect 33731 13428 33797 13429
rect 33731 13364 33732 13428
rect 33796 13364 33797 13428
rect 33731 13363 33797 13364
rect 33734 12613 33794 13363
rect 33731 12612 33797 12613
rect 33731 12548 33732 12612
rect 33796 12548 33797 12612
rect 33731 12547 33797 12548
rect 33547 11252 33613 11253
rect 33547 11188 33548 11252
rect 33612 11188 33613 11252
rect 33547 11187 33613 11188
rect 33179 10980 33245 10981
rect 33179 10916 33180 10980
rect 33244 10916 33245 10980
rect 33179 10915 33245 10916
rect 32995 9756 33061 9757
rect 32995 9692 32996 9756
rect 33060 9692 33061 9756
rect 32995 9691 33061 9692
rect 33550 7445 33610 11187
rect 33734 10709 33794 12547
rect 33731 10708 33797 10709
rect 33731 10644 33732 10708
rect 33796 10644 33797 10708
rect 33731 10643 33797 10644
rect 34102 9621 34162 18667
rect 34470 16829 34530 22339
rect 34654 19685 34714 22475
rect 34651 19684 34717 19685
rect 34651 19620 34652 19684
rect 34716 19620 34717 19684
rect 34651 19619 34717 19620
rect 34651 18460 34717 18461
rect 34651 18396 34652 18460
rect 34716 18396 34717 18460
rect 34651 18395 34717 18396
rect 34467 16828 34533 16829
rect 34467 16764 34468 16828
rect 34532 16764 34533 16828
rect 34467 16763 34533 16764
rect 34654 12069 34714 18395
rect 34838 13973 34898 23835
rect 35755 23628 35821 23629
rect 35755 23564 35756 23628
rect 35820 23564 35821 23628
rect 35755 23563 35821 23564
rect 35571 21452 35637 21453
rect 35571 21388 35572 21452
rect 35636 21388 35637 21452
rect 35571 21387 35637 21388
rect 35574 18189 35634 21387
rect 35571 18188 35637 18189
rect 35571 18124 35572 18188
rect 35636 18124 35637 18188
rect 35571 18123 35637 18124
rect 34835 13972 34901 13973
rect 34835 13908 34836 13972
rect 34900 13908 34901 13972
rect 34835 13907 34901 13908
rect 35203 13836 35269 13837
rect 35203 13772 35204 13836
rect 35268 13772 35269 13836
rect 35203 13771 35269 13772
rect 35206 12450 35266 13771
rect 35022 12390 35266 12450
rect 34651 12068 34717 12069
rect 34651 12004 34652 12068
rect 34716 12004 34717 12068
rect 34651 12003 34717 12004
rect 34467 9756 34533 9757
rect 34467 9692 34468 9756
rect 34532 9692 34533 9756
rect 34467 9691 34533 9692
rect 34099 9620 34165 9621
rect 34099 9556 34100 9620
rect 34164 9556 34165 9620
rect 34099 9555 34165 9556
rect 33547 7444 33613 7445
rect 33547 7380 33548 7444
rect 33612 7380 33613 7444
rect 33547 7379 33613 7380
rect 32811 6900 32877 6901
rect 32811 6836 32812 6900
rect 32876 6836 32877 6900
rect 32811 6835 32877 6836
rect 30235 6220 30301 6221
rect 30235 6156 30236 6220
rect 30300 6156 30301 6220
rect 30235 6155 30301 6156
rect 29840 5952 29848 6016
rect 29912 5952 29928 6016
rect 29992 5952 30008 6016
rect 30072 5952 30088 6016
rect 30152 5952 30160 6016
rect 29499 5404 29565 5405
rect 29499 5340 29500 5404
rect 29564 5340 29565 5404
rect 29499 5339 29565 5340
rect 29840 4928 30160 5952
rect 32814 5949 32874 6835
rect 32811 5948 32877 5949
rect 32811 5884 32812 5948
rect 32876 5884 32877 5948
rect 32811 5883 32877 5884
rect 33550 5133 33610 7379
rect 33547 5132 33613 5133
rect 33547 5068 33548 5132
rect 33612 5068 33613 5132
rect 33547 5067 33613 5068
rect 29840 4864 29848 4928
rect 29912 4864 29928 4928
rect 29992 4864 30008 4928
rect 30072 4864 30088 4928
rect 30152 4864 30160 4928
rect 29840 3840 30160 4864
rect 34470 4589 34530 9691
rect 35022 9621 35082 12390
rect 35758 11525 35818 23563
rect 35939 20228 36005 20229
rect 35939 20164 35940 20228
rect 36004 20164 36005 20228
rect 35939 20163 36005 20164
rect 35942 14653 36002 20163
rect 36678 19549 36738 24515
rect 37227 23492 37293 23493
rect 37227 23428 37228 23492
rect 37292 23428 37293 23492
rect 37227 23427 37293 23428
rect 37043 22268 37109 22269
rect 37043 22204 37044 22268
rect 37108 22204 37109 22268
rect 37043 22203 37109 22204
rect 36859 20772 36925 20773
rect 36859 20708 36860 20772
rect 36924 20708 36925 20772
rect 36859 20707 36925 20708
rect 36675 19548 36741 19549
rect 36675 19484 36676 19548
rect 36740 19484 36741 19548
rect 36675 19483 36741 19484
rect 36862 17237 36922 20707
rect 36859 17236 36925 17237
rect 36859 17172 36860 17236
rect 36924 17172 36925 17236
rect 36859 17171 36925 17172
rect 37046 16965 37106 22203
rect 37230 17370 37290 23427
rect 37414 19277 37474 26555
rect 37598 21997 37658 28323
rect 38331 27980 38397 27981
rect 38331 27916 38332 27980
rect 38396 27916 38397 27980
rect 38331 27915 38397 27916
rect 37963 24716 38029 24717
rect 37963 24652 37964 24716
rect 38028 24652 38029 24716
rect 37963 24651 38029 24652
rect 37779 22132 37845 22133
rect 37779 22068 37780 22132
rect 37844 22068 37845 22132
rect 37779 22067 37845 22068
rect 37595 21996 37661 21997
rect 37595 21932 37596 21996
rect 37660 21932 37661 21996
rect 37595 21931 37661 21932
rect 37411 19276 37477 19277
rect 37411 19212 37412 19276
rect 37476 19212 37477 19276
rect 37411 19211 37477 19212
rect 37230 17310 37474 17370
rect 37227 17236 37293 17237
rect 37227 17172 37228 17236
rect 37292 17172 37293 17236
rect 37227 17171 37293 17172
rect 37043 16964 37109 16965
rect 37043 16900 37044 16964
rect 37108 16900 37109 16964
rect 37043 16899 37109 16900
rect 36123 16420 36189 16421
rect 36123 16356 36124 16420
rect 36188 16356 36189 16420
rect 36123 16355 36189 16356
rect 35939 14652 36005 14653
rect 35939 14588 35940 14652
rect 36004 14588 36005 14652
rect 35939 14587 36005 14588
rect 35942 13837 36002 14587
rect 35939 13836 36005 13837
rect 35939 13772 35940 13836
rect 36004 13772 36005 13836
rect 35939 13771 36005 13772
rect 35755 11524 35821 11525
rect 35755 11460 35756 11524
rect 35820 11460 35821 11524
rect 35755 11459 35821 11460
rect 35758 10165 35818 11459
rect 35939 11252 36005 11253
rect 35939 11188 35940 11252
rect 36004 11188 36005 11252
rect 35939 11187 36005 11188
rect 35755 10164 35821 10165
rect 35755 10100 35756 10164
rect 35820 10100 35821 10164
rect 35755 10099 35821 10100
rect 35019 9620 35085 9621
rect 35019 9556 35020 9620
rect 35084 9556 35085 9620
rect 35019 9555 35085 9556
rect 34467 4588 34533 4589
rect 34467 4524 34468 4588
rect 34532 4524 34533 4588
rect 34467 4523 34533 4524
rect 29840 3776 29848 3840
rect 29912 3776 29928 3840
rect 29992 3776 30008 3840
rect 30072 3776 30088 3840
rect 30152 3776 30160 3840
rect 29315 3364 29381 3365
rect 29315 3300 29316 3364
rect 29380 3300 29381 3364
rect 29315 3299 29381 3300
rect 20208 3232 20216 3296
rect 20280 3232 20296 3296
rect 20360 3232 20376 3296
rect 20440 3232 20456 3296
rect 20520 3232 20528 3296
rect 20208 2208 20528 3232
rect 20208 2144 20216 2208
rect 20280 2144 20296 2208
rect 20360 2144 20376 2208
rect 20440 2144 20456 2208
rect 20520 2144 20528 2208
rect 20208 2128 20528 2144
rect 29840 2752 30160 3776
rect 29840 2688 29848 2752
rect 29912 2688 29928 2752
rect 29992 2688 30008 2752
rect 30072 2688 30088 2752
rect 30152 2688 30160 2752
rect 29840 2128 30160 2688
rect 35022 1869 35082 9555
rect 35942 5269 36002 11187
rect 36126 10845 36186 16355
rect 36307 14788 36373 14789
rect 36307 14724 36308 14788
rect 36372 14724 36373 14788
rect 36307 14723 36373 14724
rect 36310 11661 36370 14723
rect 36491 14652 36557 14653
rect 36491 14588 36492 14652
rect 36556 14588 36557 14652
rect 36491 14587 36557 14588
rect 36307 11660 36373 11661
rect 36307 11596 36308 11660
rect 36372 11596 36373 11660
rect 36307 11595 36373 11596
rect 36123 10844 36189 10845
rect 36123 10780 36124 10844
rect 36188 10780 36189 10844
rect 36123 10779 36189 10780
rect 36494 6765 36554 14587
rect 37230 10437 37290 17171
rect 37227 10436 37293 10437
rect 37227 10372 37228 10436
rect 37292 10372 37293 10436
rect 37227 10371 37293 10372
rect 37414 9077 37474 17310
rect 37782 17237 37842 22067
rect 37966 21317 38026 24651
rect 37963 21316 38029 21317
rect 37963 21252 37964 21316
rect 38028 21252 38029 21316
rect 37963 21251 38029 21252
rect 37779 17236 37845 17237
rect 37779 17172 37780 17236
rect 37844 17172 37845 17236
rect 37779 17171 37845 17172
rect 38334 13565 38394 27915
rect 39251 27572 39317 27573
rect 39251 27508 39252 27572
rect 39316 27508 39317 27572
rect 39251 27507 39317 27508
rect 38699 26756 38765 26757
rect 38699 26692 38700 26756
rect 38764 26692 38765 26756
rect 38699 26691 38765 26692
rect 38702 19277 38762 26691
rect 38883 22948 38949 22949
rect 38883 22884 38884 22948
rect 38948 22884 38949 22948
rect 38883 22883 38949 22884
rect 38699 19276 38765 19277
rect 38699 19212 38700 19276
rect 38764 19212 38765 19276
rect 38699 19211 38765 19212
rect 38886 16285 38946 22883
rect 38883 16284 38949 16285
rect 38883 16220 38884 16284
rect 38948 16220 38949 16284
rect 38883 16219 38949 16220
rect 38699 15468 38765 15469
rect 38699 15404 38700 15468
rect 38764 15404 38765 15468
rect 38699 15403 38765 15404
rect 38331 13564 38397 13565
rect 38331 13500 38332 13564
rect 38396 13500 38397 13564
rect 38331 13499 38397 13500
rect 38702 12885 38762 15403
rect 38886 15333 38946 16219
rect 38883 15332 38949 15333
rect 38883 15268 38884 15332
rect 38948 15268 38949 15332
rect 38883 15267 38949 15268
rect 38699 12884 38765 12885
rect 38699 12820 38700 12884
rect 38764 12820 38765 12884
rect 38699 12819 38765 12820
rect 38886 12749 38946 15267
rect 39254 13973 39314 27507
rect 39472 27232 39792 27792
rect 39472 27168 39480 27232
rect 39544 27168 39560 27232
rect 39624 27168 39640 27232
rect 39704 27168 39720 27232
rect 39784 27168 39792 27232
rect 39472 26144 39792 27168
rect 39472 26080 39480 26144
rect 39544 26080 39560 26144
rect 39624 26080 39640 26144
rect 39704 26080 39720 26144
rect 39784 26080 39792 26144
rect 39472 25056 39792 26080
rect 39472 24992 39480 25056
rect 39544 24992 39560 25056
rect 39624 24992 39640 25056
rect 39704 24992 39720 25056
rect 39784 24992 39792 25056
rect 39472 23968 39792 24992
rect 39472 23904 39480 23968
rect 39544 23904 39560 23968
rect 39624 23904 39640 23968
rect 39704 23904 39720 23968
rect 39784 23904 39792 23968
rect 39472 22880 39792 23904
rect 39472 22816 39480 22880
rect 39544 22816 39560 22880
rect 39624 22816 39640 22880
rect 39704 22816 39720 22880
rect 39784 22816 39792 22880
rect 39472 21792 39792 22816
rect 39472 21728 39480 21792
rect 39544 21728 39560 21792
rect 39624 21728 39640 21792
rect 39704 21728 39720 21792
rect 39784 21728 39792 21792
rect 39472 20704 39792 21728
rect 39472 20640 39480 20704
rect 39544 20640 39560 20704
rect 39624 20640 39640 20704
rect 39704 20640 39720 20704
rect 39784 20640 39792 20704
rect 39472 19616 39792 20640
rect 39472 19552 39480 19616
rect 39544 19552 39560 19616
rect 39624 19552 39640 19616
rect 39704 19552 39720 19616
rect 39784 19552 39792 19616
rect 39472 18528 39792 19552
rect 39472 18464 39480 18528
rect 39544 18464 39560 18528
rect 39624 18464 39640 18528
rect 39704 18464 39720 18528
rect 39784 18464 39792 18528
rect 39472 17440 39792 18464
rect 39472 17376 39480 17440
rect 39544 17376 39560 17440
rect 39624 17376 39640 17440
rect 39704 17376 39720 17440
rect 39784 17376 39792 17440
rect 39472 16352 39792 17376
rect 39472 16288 39480 16352
rect 39544 16288 39560 16352
rect 39624 16288 39640 16352
rect 39704 16288 39720 16352
rect 39784 16288 39792 16352
rect 39472 15264 39792 16288
rect 39472 15200 39480 15264
rect 39544 15200 39560 15264
rect 39624 15200 39640 15264
rect 39704 15200 39720 15264
rect 39784 15200 39792 15264
rect 39472 14176 39792 15200
rect 39472 14112 39480 14176
rect 39544 14112 39560 14176
rect 39624 14112 39640 14176
rect 39704 14112 39720 14176
rect 39784 14112 39792 14176
rect 39251 13972 39317 13973
rect 39251 13908 39252 13972
rect 39316 13908 39317 13972
rect 39251 13907 39317 13908
rect 39472 13088 39792 14112
rect 40174 14109 40234 29275
rect 42747 28796 42813 28797
rect 42747 28732 42748 28796
rect 42812 28732 42813 28796
rect 42747 28731 42813 28732
rect 40355 28524 40421 28525
rect 40355 28460 40356 28524
rect 40420 28460 40421 28524
rect 40355 28459 40421 28460
rect 40171 14108 40237 14109
rect 40171 14044 40172 14108
rect 40236 14044 40237 14108
rect 40171 14043 40237 14044
rect 40358 13973 40418 28459
rect 42011 28252 42077 28253
rect 42011 28188 42012 28252
rect 42076 28188 42077 28252
rect 42011 28187 42077 28188
rect 40907 27844 40973 27845
rect 40907 27780 40908 27844
rect 40972 27780 40973 27844
rect 40907 27779 40973 27780
rect 40910 19413 40970 27779
rect 41091 24172 41157 24173
rect 41091 24108 41092 24172
rect 41156 24108 41157 24172
rect 41091 24107 41157 24108
rect 40907 19412 40973 19413
rect 40907 19348 40908 19412
rect 40972 19348 40973 19412
rect 40907 19347 40973 19348
rect 41094 17373 41154 24107
rect 42014 21181 42074 28187
rect 42011 21180 42077 21181
rect 42011 21116 42012 21180
rect 42076 21116 42077 21180
rect 42011 21115 42077 21116
rect 42750 19413 42810 28731
rect 45139 28660 45205 28661
rect 45139 28596 45140 28660
rect 45204 28596 45205 28660
rect 45139 28595 45205 28596
rect 41643 19412 41709 19413
rect 41643 19348 41644 19412
rect 41708 19348 41709 19412
rect 41643 19347 41709 19348
rect 42747 19412 42813 19413
rect 42747 19348 42748 19412
rect 42812 19348 42813 19412
rect 42747 19347 42813 19348
rect 41091 17372 41157 17373
rect 41091 17308 41092 17372
rect 41156 17308 41157 17372
rect 41091 17307 41157 17308
rect 39987 13972 40053 13973
rect 39987 13908 39988 13972
rect 40052 13908 40053 13972
rect 39987 13907 40053 13908
rect 40355 13972 40421 13973
rect 40355 13908 40356 13972
rect 40420 13908 40421 13972
rect 40355 13907 40421 13908
rect 39472 13024 39480 13088
rect 39544 13024 39560 13088
rect 39624 13024 39640 13088
rect 39704 13024 39720 13088
rect 39784 13024 39792 13088
rect 38883 12748 38949 12749
rect 38883 12684 38884 12748
rect 38948 12684 38949 12748
rect 38883 12683 38949 12684
rect 39472 12000 39792 13024
rect 39990 12069 40050 13907
rect 40358 12341 40418 13907
rect 40355 12340 40421 12341
rect 40355 12276 40356 12340
rect 40420 12276 40421 12340
rect 40355 12275 40421 12276
rect 39987 12068 40053 12069
rect 39987 12004 39988 12068
rect 40052 12004 40053 12068
rect 39987 12003 40053 12004
rect 39472 11936 39480 12000
rect 39544 11936 39560 12000
rect 39624 11936 39640 12000
rect 39704 11936 39720 12000
rect 39784 11936 39792 12000
rect 37595 11524 37661 11525
rect 37595 11460 37596 11524
rect 37660 11460 37661 11524
rect 37595 11459 37661 11460
rect 37411 9076 37477 9077
rect 37411 9012 37412 9076
rect 37476 9012 37477 9076
rect 37411 9011 37477 9012
rect 36491 6764 36557 6765
rect 36491 6700 36492 6764
rect 36556 6700 36557 6764
rect 36491 6699 36557 6700
rect 35939 5268 36005 5269
rect 35939 5204 35940 5268
rect 36004 5204 36005 5268
rect 35939 5203 36005 5204
rect 37598 5133 37658 11459
rect 39472 10912 39792 11936
rect 39472 10848 39480 10912
rect 39544 10848 39560 10912
rect 39624 10848 39640 10912
rect 39704 10848 39720 10912
rect 39784 10848 39792 10912
rect 39472 9824 39792 10848
rect 39472 9760 39480 9824
rect 39544 9760 39560 9824
rect 39624 9760 39640 9824
rect 39704 9760 39720 9824
rect 39784 9760 39792 9824
rect 39472 8736 39792 9760
rect 39472 8672 39480 8736
rect 39544 8672 39560 8736
rect 39624 8672 39640 8736
rect 39704 8672 39720 8736
rect 39784 8672 39792 8736
rect 39472 7648 39792 8672
rect 39472 7584 39480 7648
rect 39544 7584 39560 7648
rect 39624 7584 39640 7648
rect 39704 7584 39720 7648
rect 39784 7584 39792 7648
rect 39472 6560 39792 7584
rect 39472 6496 39480 6560
rect 39544 6496 39560 6560
rect 39624 6496 39640 6560
rect 39704 6496 39720 6560
rect 39784 6496 39792 6560
rect 39472 5472 39792 6496
rect 39472 5408 39480 5472
rect 39544 5408 39560 5472
rect 39624 5408 39640 5472
rect 39704 5408 39720 5472
rect 39784 5408 39792 5472
rect 37595 5132 37661 5133
rect 37595 5068 37596 5132
rect 37660 5068 37661 5132
rect 37595 5067 37661 5068
rect 39472 4384 39792 5408
rect 39472 4320 39480 4384
rect 39544 4320 39560 4384
rect 39624 4320 39640 4384
rect 39704 4320 39720 4384
rect 39784 4320 39792 4384
rect 39472 3296 39792 4320
rect 41646 4181 41706 19347
rect 45142 17917 45202 28595
rect 49104 27776 49424 27792
rect 49104 27712 49112 27776
rect 49176 27712 49192 27776
rect 49256 27712 49272 27776
rect 49336 27712 49352 27776
rect 49416 27712 49424 27776
rect 49104 26688 49424 27712
rect 49104 26624 49112 26688
rect 49176 26624 49192 26688
rect 49256 26624 49272 26688
rect 49336 26624 49352 26688
rect 49416 26624 49424 26688
rect 49104 25600 49424 26624
rect 49104 25536 49112 25600
rect 49176 25536 49192 25600
rect 49256 25536 49272 25600
rect 49336 25536 49352 25600
rect 49416 25536 49424 25600
rect 49104 24512 49424 25536
rect 49104 24448 49112 24512
rect 49176 24448 49192 24512
rect 49256 24448 49272 24512
rect 49336 24448 49352 24512
rect 49416 24448 49424 24512
rect 49104 23424 49424 24448
rect 49104 23360 49112 23424
rect 49176 23360 49192 23424
rect 49256 23360 49272 23424
rect 49336 23360 49352 23424
rect 49416 23360 49424 23424
rect 49104 22336 49424 23360
rect 49104 22272 49112 22336
rect 49176 22272 49192 22336
rect 49256 22272 49272 22336
rect 49336 22272 49352 22336
rect 49416 22272 49424 22336
rect 49104 21248 49424 22272
rect 49104 21184 49112 21248
rect 49176 21184 49192 21248
rect 49256 21184 49272 21248
rect 49336 21184 49352 21248
rect 49416 21184 49424 21248
rect 49104 20160 49424 21184
rect 49104 20096 49112 20160
rect 49176 20096 49192 20160
rect 49256 20096 49272 20160
rect 49336 20096 49352 20160
rect 49416 20096 49424 20160
rect 49104 19072 49424 20096
rect 49104 19008 49112 19072
rect 49176 19008 49192 19072
rect 49256 19008 49272 19072
rect 49336 19008 49352 19072
rect 49416 19008 49424 19072
rect 49104 17984 49424 19008
rect 49104 17920 49112 17984
rect 49176 17920 49192 17984
rect 49256 17920 49272 17984
rect 49336 17920 49352 17984
rect 49416 17920 49424 17984
rect 45139 17916 45205 17917
rect 45139 17852 45140 17916
rect 45204 17852 45205 17916
rect 45139 17851 45205 17852
rect 46059 17372 46125 17373
rect 46059 17308 46060 17372
rect 46124 17308 46125 17372
rect 46059 17307 46125 17308
rect 42195 16692 42261 16693
rect 42195 16628 42196 16692
rect 42260 16628 42261 16692
rect 42195 16627 42261 16628
rect 42198 5269 42258 16627
rect 46062 15877 46122 17307
rect 49104 16896 49424 17920
rect 49104 16832 49112 16896
rect 49176 16832 49192 16896
rect 49256 16832 49272 16896
rect 49336 16832 49352 16896
rect 49416 16832 49424 16896
rect 46611 16692 46677 16693
rect 46611 16628 46612 16692
rect 46676 16628 46677 16692
rect 46611 16627 46677 16628
rect 46059 15876 46125 15877
rect 46059 15812 46060 15876
rect 46124 15812 46125 15876
rect 46059 15811 46125 15812
rect 44403 15468 44469 15469
rect 44403 15404 44404 15468
rect 44468 15404 44469 15468
rect 44403 15403 44469 15404
rect 42563 15332 42629 15333
rect 42563 15268 42564 15332
rect 42628 15268 42629 15332
rect 42563 15267 42629 15268
rect 44219 15332 44285 15333
rect 44219 15268 44220 15332
rect 44284 15268 44285 15332
rect 44219 15267 44285 15268
rect 42566 6357 42626 15267
rect 42931 13972 42997 13973
rect 42931 13908 42932 13972
rect 42996 13908 42997 13972
rect 42931 13907 42997 13908
rect 42747 13836 42813 13837
rect 42747 13772 42748 13836
rect 42812 13772 42813 13836
rect 42747 13771 42813 13772
rect 42563 6356 42629 6357
rect 42563 6292 42564 6356
rect 42628 6292 42629 6356
rect 42563 6291 42629 6292
rect 42195 5268 42261 5269
rect 42195 5204 42196 5268
rect 42260 5204 42261 5268
rect 42195 5203 42261 5204
rect 41643 4180 41709 4181
rect 41643 4116 41644 4180
rect 41708 4116 41709 4180
rect 41643 4115 41709 4116
rect 39472 3232 39480 3296
rect 39544 3232 39560 3296
rect 39624 3232 39640 3296
rect 39704 3232 39720 3296
rect 39784 3232 39792 3296
rect 39472 2208 39792 3232
rect 42750 2413 42810 13771
rect 42934 3501 42994 13907
rect 42931 3500 42997 3501
rect 42931 3436 42932 3500
rect 42996 3436 42997 3500
rect 42931 3435 42997 3436
rect 42747 2412 42813 2413
rect 42747 2348 42748 2412
rect 42812 2348 42813 2412
rect 42747 2347 42813 2348
rect 39472 2144 39480 2208
rect 39544 2144 39560 2208
rect 39624 2144 39640 2208
rect 39704 2144 39720 2208
rect 39784 2144 39792 2208
rect 39472 2128 39792 2144
rect 44222 2005 44282 15267
rect 44406 4725 44466 15403
rect 44955 15332 45021 15333
rect 44955 15268 44956 15332
rect 45020 15268 45021 15332
rect 44955 15267 45021 15268
rect 44403 4724 44469 4725
rect 44403 4660 44404 4724
rect 44468 4660 44469 4724
rect 44403 4659 44469 4660
rect 44219 2004 44285 2005
rect 44219 1940 44220 2004
rect 44284 1940 44285 2004
rect 44219 1939 44285 1940
rect 35019 1868 35085 1869
rect 35019 1804 35020 1868
rect 35084 1804 35085 1868
rect 35019 1803 35085 1804
rect 18091 1732 18157 1733
rect 18091 1668 18092 1732
rect 18156 1668 18157 1732
rect 18091 1667 18157 1668
rect 44958 1597 45018 15267
rect 46062 2957 46122 15811
rect 46059 2956 46125 2957
rect 46059 2892 46060 2956
rect 46124 2892 46125 2956
rect 46059 2891 46125 2892
rect 46614 2549 46674 16627
rect 49104 15808 49424 16832
rect 49104 15744 49112 15808
rect 49176 15744 49192 15808
rect 49256 15744 49272 15808
rect 49336 15744 49352 15808
rect 49416 15744 49424 15808
rect 49104 14720 49424 15744
rect 49104 14656 49112 14720
rect 49176 14656 49192 14720
rect 49256 14656 49272 14720
rect 49336 14656 49352 14720
rect 49416 14656 49424 14720
rect 49104 13632 49424 14656
rect 49104 13568 49112 13632
rect 49176 13568 49192 13632
rect 49256 13568 49272 13632
rect 49336 13568 49352 13632
rect 49416 13568 49424 13632
rect 49104 12544 49424 13568
rect 49104 12480 49112 12544
rect 49176 12480 49192 12544
rect 49256 12480 49272 12544
rect 49336 12480 49352 12544
rect 49416 12480 49424 12544
rect 49104 11456 49424 12480
rect 49104 11392 49112 11456
rect 49176 11392 49192 11456
rect 49256 11392 49272 11456
rect 49336 11392 49352 11456
rect 49416 11392 49424 11456
rect 49104 10368 49424 11392
rect 49104 10304 49112 10368
rect 49176 10304 49192 10368
rect 49256 10304 49272 10368
rect 49336 10304 49352 10368
rect 49416 10304 49424 10368
rect 49104 9280 49424 10304
rect 49104 9216 49112 9280
rect 49176 9216 49192 9280
rect 49256 9216 49272 9280
rect 49336 9216 49352 9280
rect 49416 9216 49424 9280
rect 49104 8192 49424 9216
rect 49104 8128 49112 8192
rect 49176 8128 49192 8192
rect 49256 8128 49272 8192
rect 49336 8128 49352 8192
rect 49416 8128 49424 8192
rect 49104 7104 49424 8128
rect 49104 7040 49112 7104
rect 49176 7040 49192 7104
rect 49256 7040 49272 7104
rect 49336 7040 49352 7104
rect 49416 7040 49424 7104
rect 49104 6016 49424 7040
rect 49104 5952 49112 6016
rect 49176 5952 49192 6016
rect 49256 5952 49272 6016
rect 49336 5952 49352 6016
rect 49416 5952 49424 6016
rect 49104 4928 49424 5952
rect 49104 4864 49112 4928
rect 49176 4864 49192 4928
rect 49256 4864 49272 4928
rect 49336 4864 49352 4928
rect 49416 4864 49424 4928
rect 49104 3840 49424 4864
rect 49104 3776 49112 3840
rect 49176 3776 49192 3840
rect 49256 3776 49272 3840
rect 49336 3776 49352 3840
rect 49416 3776 49424 3840
rect 49104 2752 49424 3776
rect 49104 2688 49112 2752
rect 49176 2688 49192 2752
rect 49256 2688 49272 2752
rect 49336 2688 49352 2752
rect 49416 2688 49424 2752
rect 46611 2548 46677 2549
rect 46611 2484 46612 2548
rect 46676 2484 46677 2548
rect 46611 2483 46677 2484
rect 49104 2128 49424 2688
rect 44955 1596 45021 1597
rect 44955 1532 44956 1596
rect 45020 1532 45021 1596
rect 44955 1531 45021 1532
use sky130_fd_sc_hd__diode_2  ANTENNA__225__1_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 32292 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__2_A
timestamp 1644511149
transform -1 0 24564 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A
timestamp 1644511149
transform 1 0 30728 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__A
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A
timestamp 1644511149
transform -1 0 21344 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A
timestamp 1644511149
transform -1 0 39376 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1644511149
transform -1 0 31372 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A
timestamp 1644511149
transform 1 0 36616 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A
timestamp 1644511149
transform -1 0 39376 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1644511149
transform 1 0 41768 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A
timestamp 1644511149
transform -1 0 23920 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1644511149
transform -1 0 20608 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A
timestamp 1644511149
transform -1 0 44528 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A
timestamp 1644511149
transform 1 0 37720 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__A
timestamp 1644511149
transform -1 0 39836 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A
timestamp 1644511149
transform 1 0 18584 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A
timestamp 1644511149
transform -1 0 16192 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__A
timestamp 1644511149
transform 1 0 19136 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A
timestamp 1644511149
transform 1 0 45540 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A
timestamp 1644511149
transform 1 0 41124 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1644511149
transform -1 0 35880 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A
timestamp 1644511149
transform 1 0 42872 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__B_N
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A_N
timestamp 1644511149
transform 1 0 40388 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__B
timestamp 1644511149
transform 1 0 40940 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__C
timestamp 1644511149
transform 1 0 43424 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__B1
timestamp 1644511149
transform -1 0 38824 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A1
timestamp 1644511149
transform 1 0 23000 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A2
timestamp 1644511149
transform 1 0 22356 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A3
timestamp 1644511149
transform 1 0 25208 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A
timestamp 1644511149
transform -1 0 34224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A
timestamp 1644511149
transform 1 0 41676 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A1
timestamp 1644511149
transform -1 0 27140 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__S
timestamp 1644511149
transform -1 0 27140 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A
timestamp 1644511149
transform 1 0 19320 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__B
timestamp 1644511149
transform -1 0 18768 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A
timestamp 1644511149
transform 1 0 21804 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__B
timestamp 1644511149
transform 1 0 20608 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__C
timestamp 1644511149
transform -1 0 22632 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__B1
timestamp 1644511149
transform -1 0 15456 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__C1
timestamp 1644511149
transform -1 0 14904 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A1
timestamp 1644511149
transform -1 0 29072 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A
timestamp 1644511149
transform 1 0 22632 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__A1
timestamp 1644511149
transform -1 0 45632 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__A2
timestamp 1644511149
transform -1 0 44344 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__B1
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__A
timestamp 1644511149
transform 1 0 35880 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__B
timestamp 1644511149
transform -1 0 36800 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__C
timestamp 1644511149
transform -1 0 37444 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__A2
timestamp 1644511149
transform -1 0 23920 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__B1
timestamp 1644511149
transform 1 0 21160 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__C1
timestamp 1644511149
transform 1 0 20056 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A1
timestamp 1644511149
transform 1 0 17848 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__B1
timestamp 1644511149
transform -1 0 17388 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__B
timestamp 1644511149
transform -1 0 28336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A
timestamp 1644511149
transform 1 0 20976 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__A
timestamp 1644511149
transform -1 0 36800 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__A
timestamp 1644511149
transform 1 0 46368 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__B
timestamp 1644511149
transform -1 0 46184 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A
timestamp 1644511149
transform -1 0 29072 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__B
timestamp 1644511149
transform -1 0 27784 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__B
timestamp 1644511149
transform -1 0 32568 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__B
timestamp 1644511149
transform -1 0 29532 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A
timestamp 1644511149
transform -1 0 30360 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__B
timestamp 1644511149
transform -1 0 34868 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__B
timestamp 1644511149
transform -1 0 38732 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__B
timestamp 1644511149
transform -1 0 40664 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A
timestamp 1644511149
transform 1 0 23184 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__301__A
timestamp 1644511149
transform 1 0 36708 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__A
timestamp 1644511149
transform -1 0 30636 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__A
timestamp 1644511149
transform -1 0 28244 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__B
timestamp 1644511149
transform -1 0 29256 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__304__A
timestamp 1644511149
transform 1 0 26312 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__304__D
timestamp 1644511149
transform 1 0 27232 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__B
timestamp 1644511149
transform -1 0 33672 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__C
timestamp 1644511149
transform -1 0 37444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__D
timestamp 1644511149
transform -1 0 35420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__B
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__C
timestamp 1644511149
transform -1 0 38456 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__D
timestamp 1644511149
transform 1 0 39192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__A
timestamp 1644511149
transform 1 0 41032 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__A1
timestamp 1644511149
transform 1 0 27048 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__A2
timestamp 1644511149
transform -1 0 24380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__A3
timestamp 1644511149
transform 1 0 23184 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__A4
timestamp 1644511149
transform -1 0 28520 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__B1
timestamp 1644511149
transform -1 0 27692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__A
timestamp 1644511149
transform 1 0 21528 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__D
timestamp 1644511149
transform -1 0 20792 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A
timestamp 1644511149
transform 1 0 28244 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__B
timestamp 1644511149
transform -1 0 25668 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__C
timestamp 1644511149
transform 1 0 27692 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__D
timestamp 1644511149
transform -1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__A
timestamp 1644511149
transform 1 0 26680 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__B
timestamp 1644511149
transform 1 0 27140 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__C
timestamp 1644511149
transform -1 0 25944 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__D
timestamp 1644511149
transform 1 0 24932 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__A1
timestamp 1644511149
transform -1 0 34316 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__A2
timestamp 1644511149
transform -1 0 20056 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__A3
timestamp 1644511149
transform -1 0 28980 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__A4
timestamp 1644511149
transform 1 0 22080 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__B1
timestamp 1644511149
transform 1 0 19320 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__A
timestamp 1644511149
transform 1 0 20608 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__B
timestamp 1644511149
transform 1 0 23644 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__C
timestamp 1644511149
transform 1 0 22632 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__A
timestamp 1644511149
transform -1 0 30084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__B
timestamp 1644511149
transform -1 0 31188 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__C
timestamp 1644511149
transform -1 0 30268 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__A
timestamp 1644511149
transform 1 0 36248 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__B
timestamp 1644511149
transform 1 0 18032 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__C
timestamp 1644511149
transform -1 0 21160 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__D
timestamp 1644511149
transform 1 0 18584 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__A
timestamp 1644511149
transform -1 0 17388 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A
timestamp 1644511149
transform 1 0 27508 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__A
timestamp 1644511149
transform -1 0 26128 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__A
timestamp 1644511149
transform 1 0 25208 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__A
timestamp 1644511149
transform -1 0 37996 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__B1
timestamp 1644511149
transform -1 0 40388 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__A
timestamp 1644511149
transform 1 0 22632 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__A_N
timestamp 1644511149
transform -1 0 32844 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__A1
timestamp 1644511149
transform -1 0 18952 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__A2
timestamp 1644511149
transform -1 0 20976 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__B1
timestamp 1644511149
transform -1 0 19688 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A
timestamp 1644511149
transform 1 0 20056 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__A0
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__A1
timestamp 1644511149
transform 1 0 20424 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__S
timestamp 1644511149
transform -1 0 27048 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A
timestamp 1644511149
transform -1 0 28428 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__A
timestamp 1644511149
transform -1 0 16468 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A
timestamp 1644511149
transform -1 0 41216 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__B
timestamp 1644511149
transform -1 0 41768 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__C
timestamp 1644511149
transform -1 0 40020 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__A1
timestamp 1644511149
transform -1 0 15640 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__A2
timestamp 1644511149
transform 1 0 17480 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__A3
timestamp 1644511149
transform -1 0 18216 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__B1
timestamp 1644511149
transform -1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A
timestamp 1644511149
transform 1 0 25392 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__A
timestamp 1644511149
transform -1 0 28704 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A
timestamp 1644511149
transform -1 0 22264 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__A2
timestamp 1644511149
transform -1 0 19688 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__B1
timestamp 1644511149
transform 1 0 21160 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A
timestamp 1644511149
transform -1 0 26496 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A
timestamp 1644511149
transform 1 0 24472 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A1
timestamp 1644511149
transform -1 0 24840 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__S
timestamp 1644511149
transform -1 0 23920 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__344__A
timestamp 1644511149
transform -1 0 22632 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A
timestamp 1644511149
transform -1 0 18768 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__A
timestamp 1644511149
transform -1 0 42780 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__B
timestamp 1644511149
transform -1 0 43884 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__C
timestamp 1644511149
transform -1 0 41768 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__A
timestamp 1644511149
transform 1 0 26496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__B
timestamp 1644511149
transform -1 0 30820 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__C
timestamp 1644511149
transform -1 0 28704 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A2
timestamp 1644511149
transform -1 0 36616 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__B1
timestamp 1644511149
transform -1 0 38272 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A
timestamp 1644511149
transform 1 0 40756 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__A2
timestamp 1644511149
transform -1 0 18216 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__B1
timestamp 1644511149
transform 1 0 20056 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A
timestamp 1644511149
transform -1 0 17112 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A
timestamp 1644511149
transform -1 0 17480 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A
timestamp 1644511149
transform -1 0 24288 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__B
timestamp 1644511149
transform -1 0 21712 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A
timestamp 1644511149
transform -1 0 27968 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__B
timestamp 1644511149
transform -1 0 29072 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A
timestamp 1644511149
transform 1 0 34592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A1
timestamp 1644511149
transform -1 0 40572 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__B1
timestamp 1644511149
transform 1 0 42228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A
timestamp 1644511149
transform -1 0 16192 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__B
timestamp 1644511149
transform -1 0 20700 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A
timestamp 1644511149
transform -1 0 43148 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__B
timestamp 1644511149
transform -1 0 41124 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__C
timestamp 1644511149
transform -1 0 44160 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1644511149
transform -1 0 32292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__B
timestamp 1644511149
transform -1 0 31740 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__C
timestamp 1644511149
transform -1 0 33120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__B1
timestamp 1644511149
transform 1 0 44712 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A
timestamp 1644511149
transform -1 0 16192 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__B
timestamp 1644511149
transform -1 0 15456 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A
timestamp 1644511149
transform 1 0 25944 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__B
timestamp 1644511149
transform 1 0 27232 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__C
timestamp 1644511149
transform -1 0 24748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__D
timestamp 1644511149
transform 1 0 26312 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__A
timestamp 1644511149
transform -1 0 16836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__B
timestamp 1644511149
transform 1 0 17480 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__C
timestamp 1644511149
transform 1 0 16744 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__D
timestamp 1644511149
transform 1 0 18216 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A
timestamp 1644511149
transform 1 0 37260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__A2
timestamp 1644511149
transform -1 0 39008 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__B1
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1644511149
transform -1 0 16284 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__B
timestamp 1644511149
transform -1 0 15640 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__B
timestamp 1644511149
transform -1 0 28060 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__C
timestamp 1644511149
transform -1 0 25576 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1644511149
transform 1 0 23092 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__A
timestamp 1644511149
transform 1 0 21896 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__B
timestamp 1644511149
transform 1 0 23736 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__B
timestamp 1644511149
transform -1 0 15088 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__D
timestamp 1644511149
transform -1 0 17112 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__A
timestamp 1644511149
transform -1 0 22264 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A
timestamp 1644511149
transform -1 0 45172 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__B
timestamp 1644511149
transform -1 0 46276 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__376__A
timestamp 1644511149
transform -1 0 32844 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__376__B
timestamp 1644511149
transform -1 0 33672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A
timestamp 1644511149
transform -1 0 43792 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__B
timestamp 1644511149
transform -1 0 44620 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__B
timestamp 1644511149
transform -1 0 22724 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__379__A
timestamp 1644511149
transform -1 0 45724 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A
timestamp 1644511149
transform -1 0 14904 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__B
timestamp 1644511149
transform -1 0 15732 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A
timestamp 1644511149
transform 1 0 44160 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1644511149
transform -1 0 16192 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__385__A
timestamp 1644511149
transform -1 0 20424 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__385__B
timestamp 1644511149
transform 1 0 19504 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__B
timestamp 1644511149
transform 1 0 39744 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__C
timestamp 1644511149
transform 1 0 37812 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__D
timestamp 1644511149
transform 1 0 40296 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__B
timestamp 1644511149
transform -1 0 32292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__C
timestamp 1644511149
transform -1 0 32844 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__B
timestamp 1644511149
transform 1 0 36340 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__D
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__A
timestamp 1644511149
transform -1 0 42596 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A1
timestamp 1644511149
transform 1 0 18952 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A2
timestamp 1644511149
transform -1 0 21712 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A3
timestamp 1644511149
transform -1 0 23368 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A4
timestamp 1644511149
transform -1 0 26680 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__B1
timestamp 1644511149
transform -1 0 25944 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__A
timestamp 1644511149
transform -1 0 28060 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__B
timestamp 1644511149
transform -1 0 28888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__C
timestamp 1644511149
transform -1 0 29440 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__D
timestamp 1644511149
transform -1 0 27508 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A
timestamp 1644511149
transform -1 0 35328 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__B
timestamp 1644511149
transform 1 0 34040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__C
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__D
timestamp 1644511149
transform -1 0 33948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__A
timestamp 1644511149
transform -1 0 33396 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__B
timestamp 1644511149
transform -1 0 34868 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__D
timestamp 1644511149
transform -1 0 33948 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A1
timestamp 1644511149
transform -1 0 15916 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A2
timestamp 1644511149
transform -1 0 15364 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A3
timestamp 1644511149
transform 1 0 17480 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A4
timestamp 1644511149
transform -1 0 16560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__B1
timestamp 1644511149
transform -1 0 20056 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__A
timestamp 1644511149
transform 1 0 18216 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__B
timestamp 1644511149
transform 1 0 17664 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__C
timestamp 1644511149
transform 1 0 14996 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A
timestamp 1644511149
transform -1 0 47104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__B
timestamp 1644511149
transform 1 0 45264 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__C
timestamp 1644511149
transform -1 0 46736 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A
timestamp 1644511149
transform -1 0 37996 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A_N
timestamp 1644511149
transform 1 0 14628 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__B
timestamp 1644511149
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__C
timestamp 1644511149
transform -1 0 15088 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__D
timestamp 1644511149
transform -1 0 14352 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__B
timestamp 1644511149
transform -1 0 28336 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__A
timestamp 1644511149
transform 1 0 19688 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__B
timestamp 1644511149
transform -1 0 17848 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__403__A
timestamp 1644511149
transform 1 0 23184 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A
timestamp 1644511149
transform -1 0 14536 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__A
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__B
timestamp 1644511149
transform -1 0 42964 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__C
timestamp 1644511149
transform -1 0 46276 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A
timestamp 1644511149
transform -1 0 33856 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__B
timestamp 1644511149
transform -1 0 34868 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__C
timestamp 1644511149
transform -1 0 34868 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__B1
timestamp 1644511149
transform -1 0 46000 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A
timestamp 1644511149
transform -1 0 14352 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__B
timestamp 1644511149
transform -1 0 14536 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A_N
timestamp 1644511149
transform -1 0 45172 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A1
timestamp 1644511149
transform -1 0 45724 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A2
timestamp 1644511149
transform -1 0 46276 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__B1
timestamp 1644511149
transform -1 0 43332 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A
timestamp 1644511149
transform 1 0 24840 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__B
timestamp 1644511149
transform -1 0 24196 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A0
timestamp 1644511149
transform -1 0 26128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A1
timestamp 1644511149
transform -1 0 18584 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__S
timestamp 1644511149
transform -1 0 22172 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__413__A
timestamp 1644511149
transform -1 0 13984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__A
timestamp 1644511149
transform 1 0 18676 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__A
timestamp 1644511149
transform 1 0 43332 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__B
timestamp 1644511149
transform -1 0 44252 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A1
timestamp 1644511149
transform -1 0 33580 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A2
timestamp 1644511149
transform -1 0 32568 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A3
timestamp 1644511149
transform -1 0 35420 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__B1
timestamp 1644511149
transform -1 0 34132 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__A
timestamp 1644511149
transform -1 0 24748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__B
timestamp 1644511149
transform -1 0 25300 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A
timestamp 1644511149
transform -1 0 22816 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__A
timestamp 1644511149
transform -1 0 21160 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__A2
timestamp 1644511149
transform 1 0 16376 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__B1
timestamp 1644511149
transform -1 0 13616 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__A
timestamp 1644511149
transform 1 0 19688 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A1
timestamp 1644511149
transform 1 0 17112 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__S
timestamp 1644511149
transform -1 0 15640 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__A
timestamp 1644511149
transform 1 0 22080 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__A
timestamp 1644511149
transform -1 0 13616 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__A
timestamp 1644511149
transform -1 0 47196 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__B
timestamp 1644511149
transform -1 0 47748 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__C
timestamp 1644511149
transform -1 0 48300 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__A
timestamp 1644511149
transform 1 0 35696 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__B
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__C
timestamp 1644511149
transform -1 0 39100 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__A1
timestamp 1644511149
transform -1 0 34500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__B1
timestamp 1644511149
transform 1 0 35236 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__A
timestamp 1644511149
transform 1 0 15824 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__A
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A2
timestamp 1644511149
transform -1 0 31372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__B1
timestamp 1644511149
transform -1 0 30820 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__A
timestamp 1644511149
transform -1 0 17296 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__A
timestamp 1644511149
transform 1 0 41492 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__A
timestamp 1644511149
transform 1 0 23184 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__B
timestamp 1644511149
transform -1 0 23368 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__A
timestamp 1644511149
transform -1 0 35972 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__B
timestamp 1644511149
transform 1 0 36984 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__B1
timestamp 1644511149
transform -1 0 33120 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__A
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__B
timestamp 1644511149
transform -1 0 38548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__A
timestamp 1644511149
transform 1 0 17848 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__B
timestamp 1644511149
transform -1 0 15640 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__C
timestamp 1644511149
transform -1 0 17112 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__A
timestamp 1644511149
transform -1 0 40572 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__B
timestamp 1644511149
transform -1 0 36432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__C
timestamp 1644511149
transform -1 0 39100 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__A1
timestamp 1644511149
transform -1 0 45172 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__B1
timestamp 1644511149
transform -1 0 44804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__441__A
timestamp 1644511149
transform -1 0 14628 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__441__B
timestamp 1644511149
transform -1 0 15088 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__A
timestamp 1644511149
transform -1 0 37996 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__B
timestamp 1644511149
transform 1 0 39100 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__C
timestamp 1644511149
transform 1 0 38640 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__D
timestamp 1644511149
transform -1 0 40572 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__A
timestamp 1644511149
transform -1 0 33672 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__B
timestamp 1644511149
transform -1 0 34684 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__C
timestamp 1644511149
transform -1 0 35420 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__D
timestamp 1644511149
transform -1 0 36524 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__A2
timestamp 1644511149
transform -1 0 46828 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__B1
timestamp 1644511149
transform -1 0 47656 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__A
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__B
timestamp 1644511149
transform -1 0 18032 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__A_N
timestamp 1644511149
transform -1 0 41492 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__B
timestamp 1644511149
transform -1 0 37720 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__C
timestamp 1644511149
transform -1 0 39836 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__A
timestamp 1644511149
transform -1 0 13432 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__B
timestamp 1644511149
transform -1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__A
timestamp 1644511149
transform -1 0 41032 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__B
timestamp 1644511149
transform -1 0 41676 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__A_N
timestamp 1644511149
transform -1 0 13064 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__B
timestamp 1644511149
transform -1 0 12512 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__C
timestamp 1644511149
transform -1 0 15456 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__D
timestamp 1644511149
transform 1 0 16560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__A
timestamp 1644511149
transform -1 0 42596 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__B
timestamp 1644511149
transform -1 0 41584 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__A
timestamp 1644511149
transform -1 0 27416 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__A
timestamp 1644511149
transform 1 0 42136 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__B
timestamp 1644511149
transform 1 0 42964 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__456__A
timestamp 1644511149
transform -1 0 39376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__457__S
timestamp 1644511149
transform -1 0 47748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__458__B
timestamp 1644511149
transform -1 0 23920 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__459__B
timestamp 1644511149
transform -1 0 16192 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__A
timestamp 1644511149
transform -1 0 25024 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__B
timestamp 1644511149
transform 1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__462__A
timestamp 1644511149
transform 1 0 43700 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__463__A
timestamp 1644511149
transform 1 0 26312 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__463__B
timestamp 1644511149
transform -1 0 28152 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__A
timestamp 1644511149
transform 1 0 34040 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__B
timestamp 1644511149
transform 1 0 35052 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__C
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__A
timestamp 1644511149
transform -1 0 25944 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__B
timestamp 1644511149
transform -1 0 27600 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__A
timestamp 1644511149
transform -1 0 45724 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__B
timestamp 1644511149
transform -1 0 46828 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__A
timestamp 1644511149
transform -1 0 20792 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__A
timestamp 1644511149
transform -1 0 21344 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__471__A
timestamp 1644511149
transform -1 0 48208 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__A
timestamp 1644511149
transform -1 0 20792 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__473__A
timestamp 1644511149
transform -1 0 48300 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__A
timestamp 1644511149
transform -1 0 19320 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__A
timestamp 1644511149
transform 1 0 19320 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__A
timestamp 1644511149
transform -1 0 47748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__A
timestamp 1644511149
transform -1 0 18308 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__A
timestamp 1644511149
transform -1 0 14812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__A
timestamp 1644511149
transform -1 0 13984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__A
timestamp 1644511149
transform -1 0 40388 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__A
timestamp 1644511149
transform -1 0 14536 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__A
timestamp 1644511149
transform -1 0 18216 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__A
timestamp 1644511149
transform -1 0 42228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__A
timestamp 1644511149
transform -1 0 13616 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__A
timestamp 1644511149
transform -1 0 31372 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__A
timestamp 1644511149
transform -1 0 44436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__A
timestamp 1644511149
transform -1 0 32292 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__500__A
timestamp 1644511149
transform -1 0 38548 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__501__A
timestamp 1644511149
transform -1 0 45172 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__505__A
timestamp 1644511149
transform -1 0 44988 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__513__A
timestamp 1644511149
transform -1 0 39100 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__5_A
timestamp 1644511149
transform -1 0 43700 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__A
timestamp 1644511149
transform -1 0 25576 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__A
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__A
timestamp 1644511149
transform 1 0 42964 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__A
timestamp 1644511149
transform -1 0 27416 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__A
timestamp 1644511149
transform -1 0 37628 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__A
timestamp 1644511149
transform -1 0 22816 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__A
timestamp 1644511149
transform -1 0 46828 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__527__A
timestamp 1644511149
transform 1 0 12512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__528__A
timestamp 1644511149
transform 1 0 46368 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__529__A
timestamp 1644511149
transform 1 0 42596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__530__A
timestamp 1644511149
transform 1 0 45540 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__531__A
timestamp 1644511149
transform -1 0 46276 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__532__A
timestamp 1644511149
transform 1 0 35604 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__533__A
timestamp 1644511149
transform 1 0 36156 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__534__A
timestamp 1644511149
transform 1 0 36340 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__535__A
timestamp 1644511149
transform -1 0 17480 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__536__A
timestamp 1644511149
transform -1 0 30268 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__537__A
timestamp 1644511149
transform 1 0 43884 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__538__A
timestamp 1644511149
transform 1 0 40020 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__539__A
timestamp 1644511149
transform -1 0 29716 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__540__A
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__541__A
timestamp 1644511149
transform 1 0 26312 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__542__A
timestamp 1644511149
transform -1 0 47748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__543__A
timestamp 1644511149
transform 1 0 21896 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__544__A
timestamp 1644511149
transform -1 0 31924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__545__A
timestamp 1644511149
transform 1 0 48668 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__A
timestamp 1644511149
transform 1 0 32660 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__547__A
timestamp 1644511149
transform -1 0 29072 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__548__A
timestamp 1644511149
transform 1 0 45540 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__549__A
timestamp 1644511149
transform -1 0 35052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__550__A
timestamp 1644511149
transform -1 0 37444 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__551__A
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__552__A
timestamp 1644511149
transform 1 0 38088 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__553__A
timestamp 1644511149
transform -1 0 37076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__554__A
timestamp 1644511149
transform 1 0 37812 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__A
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__556__A
timestamp 1644511149
transform -1 0 16008 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__556__B
timestamp 1644511149
transform -1 0 15088 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__557__A
timestamp 1644511149
transform -1 0 15456 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__558__A
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__560__A
timestamp 1644511149
transform -1 0 38824 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__562__A
timestamp 1644511149
transform 1 0 42688 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__564__A
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__RESET_B
timestamp 1644511149
transform 1 0 48576 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__567__RESET_B
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__568__RESET_B
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__569__CLK
timestamp 1644511149
transform 1 0 22632 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__569__RESET_B
timestamp 1644511149
transform 1 0 17296 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__570__RESET_B
timestamp 1644511149
transform 1 0 23920 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__571__CLK
timestamp 1644511149
transform 1 0 41492 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__571__RESET_B
timestamp 1644511149
transform 1 0 40756 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__572__CLK
timestamp 1644511149
transform -1 0 45540 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__572__RESET_B
timestamp 1644511149
transform 1 0 43240 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__CLK
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__RESET_B
timestamp 1644511149
transform 1 0 44068 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__574__CLK
timestamp 1644511149
transform 1 0 24840 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__574__RESET_B
timestamp 1644511149
transform 1 0 25116 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__575__CLK
timestamp 1644511149
transform -1 0 47380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__575__RESET_B
timestamp 1644511149
transform 1 0 46644 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__576__CLK
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__576__RESET_B
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__577__CLK
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__577__D
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__577__RESET_B
timestamp 1644511149
transform 1 0 40388 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__578__CLK
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__578__RESET_B
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__579__CLK
timestamp 1644511149
transform 1 0 45172 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__580__CLK
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__582__CLK
timestamp 1644511149
transform 1 0 14720 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__584__CLK
timestamp 1644511149
transform 1 0 12696 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__584__D
timestamp 1644511149
transform -1 0 11960 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__586__CLK
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__586__RESET_B
timestamp 1644511149
transform -1 0 13064 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__587__CLK
timestamp 1644511149
transform -1 0 29532 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__588__CLK
timestamp 1644511149
transform 1 0 15456 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__588__RESET_B
timestamp 1644511149
transform -1 0 28520 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__589__CLK
timestamp 1644511149
transform -1 0 22264 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__589__RESET_B
timestamp 1644511149
transform -1 0 23920 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__590__CLK
timestamp 1644511149
transform -1 0 21344 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__590__D
timestamp 1644511149
transform -1 0 20148 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__590__RESET_B
timestamp 1644511149
transform -1 0 26496 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__591__CLK
timestamp 1644511149
transform 1 0 19412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__592__CLK
timestamp 1644511149
transform 1 0 48116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__593__CLK
timestamp 1644511149
transform 1 0 41308 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__594__CLK
timestamp 1644511149
transform 1 0 47748 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__596__CLK
timestamp 1644511149
transform 1 0 22632 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__599__CLK
timestamp 1644511149
transform 1 0 13800 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__599__RESET_B
timestamp 1644511149
transform 1 0 23184 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__600__CLK
timestamp 1644511149
transform -1 0 30084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__600__SET_B
timestamp 1644511149
transform 1 0 48116 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__601__CLK
timestamp 1644511149
transform 1 0 25760 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__601__RESET_B
timestamp 1644511149
transform 1 0 42964 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__602__CLK
timestamp 1644511149
transform 1 0 32292 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__602__RESET_B
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__603__CLK
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__603__D
timestamp 1644511149
transform -1 0 47104 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__603__RESET_B
timestamp 1644511149
transform 1 0 47748 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__604__CLK
timestamp 1644511149
transform 1 0 18584 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__604__RESET_B
timestamp 1644511149
transform 1 0 16744 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__605__CLK
timestamp 1644511149
transform -1 0 12144 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__605__RESET_B
timestamp 1644511149
transform 1 0 12328 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__606__CLK
timestamp 1644511149
transform 1 0 45908 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__606__RESET_B
timestamp 1644511149
transform 1 0 43792 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__607__CLK
timestamp 1644511149
transform 1 0 17572 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__607__RESET_B
timestamp 1644511149
transform 1 0 48668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__608__CLK
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__608__RESET_B
timestamp 1644511149
transform 1 0 44344 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__609__CLK
timestamp 1644511149
transform 1 0 49128 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__609__D
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__609__RESET_B
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__610__CLK
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__610__D
timestamp 1644511149
transform -1 0 41676 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__610__RESET_B
timestamp 1644511149
transform 1 0 38916 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__611__CLK
timestamp 1644511149
transform 1 0 49220 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__611__RESET_B
timestamp 1644511149
transform 1 0 49220 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__612__CLK
timestamp 1644511149
transform 1 0 21528 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__612__RESET_B
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__613__CLK
timestamp 1644511149
transform 1 0 16008 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__613__RESET_B
timestamp 1644511149
transform 1 0 46644 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__614__CLK
timestamp 1644511149
transform 1 0 27232 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__614__RESET_B
timestamp 1644511149
transform 1 0 26680 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__616__CLK
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__617__D
timestamp 1644511149
transform -1 0 25944 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__618__CLK
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__620__CLK
timestamp 1644511149
transform 1 0 44068 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__622__CLK
timestamp 1644511149
transform -1 0 37444 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__623__CLK
timestamp 1644511149
transform -1 0 25024 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__623__D
timestamp 1644511149
transform -1 0 22264 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__CLK
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__625__D
timestamp 1644511149
transform -1 0 19964 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__626__CLK
timestamp 1644511149
transform 1 0 46644 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__628__CLK
timestamp 1644511149
transform 1 0 39192 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__630__CLK
timestamp 1644511149
transform -1 0 24472 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__631__CLK
timestamp 1644511149
transform -1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__631__D
timestamp 1644511149
transform -1 0 13616 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__632__CLK
timestamp 1644511149
transform -1 0 47748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__635__CLK
timestamp 1644511149
transform 1 0 18584 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__635__RESET_B
timestamp 1644511149
transform 1 0 16744 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__636__CLK
timestamp 1644511149
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__636__SET_B
timestamp 1644511149
transform 1 0 48300 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__637__CLK
timestamp 1644511149
transform 1 0 49772 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__637__D
timestamp 1644511149
transform -1 0 50508 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__637__RESET_B
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__638__CLK
timestamp 1644511149
transform -1 0 32292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__638__D
timestamp 1644511149
transform -1 0 33028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__638__RESET_B
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__639__CLK
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__639__D
timestamp 1644511149
transform -1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__639__RESET_B
timestamp 1644511149
transform 1 0 48852 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__640__CLK
timestamp 1644511149
transform -1 0 28980 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__640__D
timestamp 1644511149
transform -1 0 29716 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__640__RESET_B
timestamp 1644511149
transform 1 0 33764 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__641__CLK
timestamp 1644511149
transform 1 0 23184 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__641__RESET_B
timestamp 1644511149
transform 1 0 37444 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__642__CLK
timestamp 1644511149
transform 1 0 49220 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__642__D
timestamp 1644511149
transform -1 0 50324 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__642__RESET_B
timestamp 1644511149
transform 1 0 48852 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__643__CLK
timestamp 1644511149
transform 1 0 45540 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__643__RESET_B
timestamp 1644511149
transform 1 0 46460 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__644__CLK
timestamp 1644511149
transform 1 0 26128 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__644__RESET_B
timestamp 1644511149
transform 1 0 22632 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__645__CLK
timestamp 1644511149
transform 1 0 36340 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__645__RESET_B
timestamp 1644511149
transform 1 0 41124 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__646__CLK
timestamp 1644511149
transform 1 0 40020 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__646__RESET_B
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__647__CLK
timestamp 1644511149
transform -1 0 50324 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__647__RESET_B
timestamp 1644511149
transform 1 0 38548 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__648__CLK
timestamp 1644511149
transform 1 0 20976 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__648__RESET_B
timestamp 1644511149
transform 1 0 20056 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__649__CLK
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__649__RESET_B
timestamp 1644511149
transform 1 0 11776 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__650__CLK
timestamp 1644511149
transform 1 0 20056 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__650__D
timestamp 1644511149
transform -1 0 15640 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__650__RESET_B
timestamp 1644511149
transform 1 0 22080 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__652__CLK
timestamp 1644511149
transform 1 0 47196 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__654__CLK
timestamp 1644511149
transform 1 0 45172 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__655__CLK
timestamp 1644511149
transform -1 0 14904 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__656__CLK
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__658__CLK
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__659__A
timestamp 1644511149
transform -1 0 36340 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__660__A
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__661__A
timestamp 1644511149
transform -1 0 20792 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__662__A
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__663__A
timestamp 1644511149
transform 1 0 40480 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__664__A
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__665__A
timestamp 1644511149
transform 1 0 12144 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__666__A
timestamp 1644511149
transform 1 0 12788 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__667__A
timestamp 1644511149
transform 1 0 11960 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__668__A
timestamp 1644511149
transform 1 0 11224 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__669__A
timestamp 1644511149
transform 1 0 11868 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__670__A
timestamp 1644511149
transform -1 0 11040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__671__A
timestamp 1644511149
transform 1 0 13432 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__672__A
timestamp 1644511149
transform -1 0 12880 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__674__A
timestamp 1644511149
transform -1 0 26496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__675__A
timestamp 1644511149
transform 1 0 17296 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__681__A
timestamp 1644511149
transform 1 0 4416 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__682__A
timestamp 1644511149
transform 1 0 37444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__683__A
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_master_A
timestamp 1644511149
transform 1 0 30452 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
timestamp 1644511149
transform -1 0 42780 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
timestamp 1644511149
transform 1 0 20608 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 24564 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 19504 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf_A
timestamp 1644511149
transform -1 0 48300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 18032 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 16192 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_A
timestamp 1644511149
transform -1 0 49588 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
timestamp 1644511149
transform 1 0 17020 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 23736 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 20976 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_A
timestamp 1644511149
transform -1 0 49956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
timestamp 1644511149
transform 1 0 12880 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 12052 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 11224 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_A
timestamp 1644511149
transform -1 0 42228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
timestamp 1644511149
transform 1 0 20056 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 17480 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_RESET_B
timestamp 1644511149
transform -1 0 25392 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_A
timestamp 1644511149
transform -1 0 43884 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
timestamp 1644511149
transform 1 0 15640 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 14904 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 14168 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_A
timestamp 1644511149
transform -1 0 47932 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
timestamp 1644511149
transform -1 0 12328 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 16008 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 12880 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_A
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
timestamp 1644511149
transform 1 0 12328 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_GATE_N
timestamp 1644511149
transform -1 0 11684 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 18308 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_A
timestamp 1644511149
transform -1 0 38180 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
timestamp 1644511149
transform -1 0 23368 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_GATE_N
timestamp 1644511149
transform -1 0 37444 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 38916 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
timestamp 1644511149
transform 1 0 42964 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 40388 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 37812 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf_A
timestamp 1644511149
transform -1 0 14352 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
timestamp 1644511149
transform 1 0 35972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 37444 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_A
timestamp 1644511149
transform -1 0 46460 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 45540 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_A
timestamp 1644511149
transform -1 0 49956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 40020 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_A
timestamp 1644511149
transform -1 0 45356 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_A
timestamp 1644511149
transform -1 0 50508 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
timestamp 1644511149
transform -1 0 48300 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 42596 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_A
timestamp 1644511149
transform -1 0 33580 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
timestamp 1644511149
transform 1 0 47748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
timestamp 1644511149
transform -1 0 34500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 35236 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_A
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
timestamp 1644511149
transform -1 0 35052 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_GATE_N
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_RESET_B
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1644511149
transform -1 0 58236 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1644511149
transform -1 0 14904 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1644511149
transform -1 0 30820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1644511149
transform -1 0 58236 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1644511149
transform -1 0 58236 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1644511149
transform -1 0 58236 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1644511149
transform -1 0 58236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1644511149
transform -1 0 58236 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1644511149
transform -1 0 58236 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1644511149
transform -1 0 58236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1644511149
transform -1 0 58236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1644511149
transform -1 0 58236 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1644511149
transform -1 0 58236 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1644511149
transform -1 0 58236 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1644511149
transform -1 0 58236 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1644511149
transform -1 0 57408 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1644511149
transform -1 0 40480 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1644511149
transform -1 0 46000 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1644511149
transform -1 0 58052 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1644511149
transform -1 0 58236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output21_A
timestamp 1644511149
transform -1 0 25944 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output24_A
timestamp 1644511149
transform -1 0 3956 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output26_A
timestamp 1644511149
transform -1 0 2300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output27_A
timestamp 1644511149
transform -1 0 9844 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output28_A
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output41_A
timestamp 1644511149
transform 1 0 2116 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output49_A
timestamp 1644511149
transform 1 0 7084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_38
timestamp 1644511149
transform 1 0 4600 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61
timestamp 1644511149
transform 1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_67
timestamp 1644511149
transform 1 0 7268 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79
timestamp 1644511149
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1644511149
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp 1644511149
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1644511149
transform 1 0 19412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_211
timestamp 1644511149
transform 1 0 20516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_237
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1644511149
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1644511149
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1644511149
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_313
timestamp 1644511149
transform 1 0 29900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_317
timestamp 1644511149
transform 1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_323
timestamp 1644511149
transform 1 0 30820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1644511149
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1644511149
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_397
timestamp 1644511149
transform 1 0 37628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_409
timestamp 1644511149
transform 1 0 38732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1644511149
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_433
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1644511149
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_453
timestamp 1644511149
transform 1 0 42780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_465
timestamp 1644511149
transform 1 0 43884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1644511149
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_489
timestamp 1644511149
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1644511149
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_517
timestamp 1644511149
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1644511149
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_533
timestamp 1644511149
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_545
timestamp 1644511149
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1644511149
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_561
timestamp 1644511149
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_573
timestamp 1644511149
transform 1 0 53820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_579
timestamp 1644511149
transform 1 0 54372 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_587
timestamp 1644511149
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_589
timestamp 1644511149
transform 1 0 55292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_595
timestamp 1644511149
transform 1 0 55844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_612
timestamp 1644511149
transform 1 0 57408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_619
timestamp 1644511149
transform 1 0 58052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_6
timestamp 1644511149
transform 1 0 1656 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_18
timestamp 1644511149
transform 1 0 2760 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_30
timestamp 1644511149
transform 1 0 3864 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_42
timestamp 1644511149
transform 1 0 4968 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1644511149
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_137
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_193
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_205
timestamp 1644511149
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_261
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_317
timestamp 1644511149
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_349
timestamp 1644511149
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_373
timestamp 1644511149
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1644511149
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_401
timestamp 1644511149
transform 1 0 37996 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_413
timestamp 1644511149
transform 1 0 39100 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_425
timestamp 1644511149
transform 1 0 40204 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_437
timestamp 1644511149
transform 1 0 41308 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_445
timestamp 1644511149
transform 1 0 42044 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_461
timestamp 1644511149
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_473
timestamp 1644511149
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_485
timestamp 1644511149
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1644511149
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1644511149
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_517
timestamp 1644511149
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_529
timestamp 1644511149
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_541
timestamp 1644511149
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1644511149
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1644511149
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_561
timestamp 1644511149
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_573
timestamp 1644511149
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_585
timestamp 1644511149
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_597
timestamp 1644511149
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1644511149
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1644511149
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_617
timestamp 1644511149
transform 1 0 57868 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_121
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1644511149
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_424
timestamp 1644511149
transform 1 0 40112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_430
timestamp 1644511149
transform 1 0 40664 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_442
timestamp 1644511149
transform 1 0 41768 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_454
timestamp 1644511149
transform 1 0 42872 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_466
timestamp 1644511149
transform 1 0 43976 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_474
timestamp 1644511149
transform 1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_477
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_489
timestamp 1644511149
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_501
timestamp 1644511149
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_513
timestamp 1644511149
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1644511149
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1644511149
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_533
timestamp 1644511149
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_545
timestamp 1644511149
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_557
timestamp 1644511149
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_569
timestamp 1644511149
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1644511149
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1644511149
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_589
timestamp 1644511149
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_601
timestamp 1644511149
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_613
timestamp 1644511149
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1644511149
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_13
timestamp 1644511149
transform 1 0 2300 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_25
timestamp 1644511149
transform 1 0 3404 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_37
timestamp 1644511149
transform 1 0 4508 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp 1644511149
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_417
timestamp 1644511149
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_429
timestamp 1644511149
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1644511149
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_461
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_473
timestamp 1644511149
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_485
timestamp 1644511149
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1644511149
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1644511149
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_517
timestamp 1644511149
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_529
timestamp 1644511149
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_541
timestamp 1644511149
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1644511149
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1644511149
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_561
timestamp 1644511149
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_573
timestamp 1644511149
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_585
timestamp 1644511149
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_597
timestamp 1644511149
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1644511149
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1644511149
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_617
timestamp 1644511149
transform 1 0 57868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_621
timestamp 1644511149
transform 1 0 58236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_311
timestamp 1644511149
transform 1 0 29716 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_323
timestamp 1644511149
transform 1 0 30820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_335
timestamp 1644511149
transform 1 0 31924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_347
timestamp 1644511149
transform 1 0 33028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_359
timestamp 1644511149
transform 1 0 34132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_457
timestamp 1644511149
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1644511149
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_501
timestamp 1644511149
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_513
timestamp 1644511149
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1644511149
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1644511149
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_533
timestamp 1644511149
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_545
timestamp 1644511149
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_557
timestamp 1644511149
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_569
timestamp 1644511149
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1644511149
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1644511149
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_589
timestamp 1644511149
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_601
timestamp 1644511149
transform 1 0 56396 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_609
timestamp 1644511149
transform 1 0 57132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_621
timestamp 1644511149
transform 1 0 58236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_303
timestamp 1644511149
transform 1 0 28980 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_309
timestamp 1644511149
transform 1 0 29532 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_315
timestamp 1644511149
transform 1 0 30084 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_321
timestamp 1644511149
transform 1 0 30636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_333
timestamp 1644511149
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_339
timestamp 1644511149
transform 1 0 32292 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_351
timestamp 1644511149
transform 1 0 33396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_363
timestamp 1644511149
transform 1 0 34500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_375
timestamp 1644511149
transform 1 0 35604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_387
timestamp 1644511149
transform 1 0 36708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1644511149
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_517
timestamp 1644511149
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_529
timestamp 1644511149
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_541
timestamp 1644511149
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1644511149
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1644511149
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_561
timestamp 1644511149
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_573
timestamp 1644511149
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_585
timestamp 1644511149
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_597
timestamp 1644511149
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1644511149
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1644511149
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_617
timestamp 1644511149
transform 1 0 57868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_621
timestamp 1644511149
transform 1 0 58236 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_7
timestamp 1644511149
transform 1 0 1748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_19
timestamp 1644511149
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_129
timestamp 1644511149
transform 1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1644511149
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_143
timestamp 1644511149
transform 1 0 14260 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_155
timestamp 1644511149
transform 1 0 15364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_167
timestamp 1644511149
transform 1 0 16468 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_179
timestamp 1644511149
transform 1 0 17572 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_191
timestamp 1644511149
transform 1 0 18676 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_295
timestamp 1644511149
transform 1 0 28244 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_298
timestamp 1644511149
transform 1 0 28520 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_304
timestamp 1644511149
transform 1 0 29072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_311
timestamp 1644511149
transform 1 0 29716 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_317
timestamp 1644511149
transform 1 0 30268 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_323
timestamp 1644511149
transform 1 0 30820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_329
timestamp 1644511149
transform 1 0 31372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_335
timestamp 1644511149
transform 1 0 31924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_341
timestamp 1644511149
transform 1 0 32476 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_347
timestamp 1644511149
transform 1 0 33028 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_353
timestamp 1644511149
transform 1 0 33580 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_359
timestamp 1644511149
transform 1 0 34132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1644511149
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1644511149
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_533
timestamp 1644511149
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_545
timestamp 1644511149
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_557
timestamp 1644511149
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_569
timestamp 1644511149
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1644511149
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1644511149
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_589
timestamp 1644511149
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_601
timestamp 1644511149
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_613
timestamp 1644511149
transform 1 0 57500 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_621
timestamp 1644511149
transform 1 0 58236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_286
timestamp 1644511149
transform 1 0 27416 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_296
timestamp 1644511149
transform 1 0 28336 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_302
timestamp 1644511149
transform 1 0 28888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_308
timestamp 1644511149
transform 1 0 29440 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_314
timestamp 1644511149
transform 1 0 29992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_323
timestamp 1644511149
transform 1 0 30820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_339
timestamp 1644511149
transform 1 0 32292 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_345
timestamp 1644511149
transform 1 0 32844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_351
timestamp 1644511149
transform 1 0 33396 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_357
timestamp 1644511149
transform 1 0 33948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_363
timestamp 1644511149
transform 1 0 34500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_369
timestamp 1644511149
transform 1 0 35052 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_375
timestamp 1644511149
transform 1 0 35604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_387
timestamp 1644511149
transform 1 0 36708 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_517
timestamp 1644511149
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_529
timestamp 1644511149
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_541
timestamp 1644511149
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1644511149
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1644511149
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_561
timestamp 1644511149
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_573
timestamp 1644511149
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_585
timestamp 1644511149
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_597
timestamp 1644511149
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1644511149
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1644511149
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_617
timestamp 1644511149
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_271
timestamp 1644511149
transform 1 0 26036 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_274
timestamp 1644511149
transform 1 0 26312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_280
timestamp 1644511149
transform 1 0 26864 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_286
timestamp 1644511149
transform 1 0 27416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_290
timestamp 1644511149
transform 1 0 27784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_293
timestamp 1644511149
transform 1 0 28060 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_304
timestamp 1644511149
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_315
timestamp 1644511149
transform 1 0 30084 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_327
timestamp 1644511149
transform 1 0 31188 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_339
timestamp 1644511149
transform 1 0 32292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_351
timestamp 1644511149
transform 1 0 33396 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_367
timestamp 1644511149
transform 1 0 34868 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_373
timestamp 1644511149
transform 1 0 35420 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_379
timestamp 1644511149
transform 1 0 35972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_391
timestamp 1644511149
transform 1 0 37076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_403
timestamp 1644511149
transform 1 0 38180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_415
timestamp 1644511149
transform 1 0 39284 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1644511149
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1644511149
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_533
timestamp 1644511149
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_545
timestamp 1644511149
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_557
timestamp 1644511149
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_569
timestamp 1644511149
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1644511149
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1644511149
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_589
timestamp 1644511149
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_601
timestamp 1644511149
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_613
timestamp 1644511149
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_7
timestamp 1644511149
transform 1 0 1748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_19
timestamp 1644511149
transform 1 0 2852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_31
timestamp 1644511149
transform 1 0 3956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_43
timestamp 1644511149
transform 1 0 5060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_267
timestamp 1644511149
transform 1 0 25668 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_270
timestamp 1644511149
transform 1 0 25944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1644511149
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_287
timestamp 1644511149
transform 1 0 27508 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_297
timestamp 1644511149
transform 1 0 28428 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_300
timestamp 1644511149
transform 1 0 28704 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_306
timestamp 1644511149
transform 1 0 29256 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_313
timestamp 1644511149
transform 1 0 29900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_320
timestamp 1644511149
transform 1 0 30544 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_327
timestamp 1644511149
transform 1 0 31188 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_339
timestamp 1644511149
transform 1 0 32292 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_345
timestamp 1644511149
transform 1 0 32844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_351
timestamp 1644511149
transform 1 0 33396 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_357
timestamp 1644511149
transform 1 0 33948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_363
timestamp 1644511149
transform 1 0 34500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_369
timestamp 1644511149
transform 1 0 35052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_375
timestamp 1644511149
transform 1 0 35604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_381
timestamp 1644511149
transform 1 0 36156 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_387
timestamp 1644511149
transform 1 0 36708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_517
timestamp 1644511149
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_529
timestamp 1644511149
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_541
timestamp 1644511149
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1644511149
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1644511149
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_561
timestamp 1644511149
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_573
timestamp 1644511149
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_585
timestamp 1644511149
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_597
timestamp 1644511149
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1644511149
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1644511149
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_617
timestamp 1644511149
transform 1 0 57868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_621
timestamp 1644511149
transform 1 0 58236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1644511149
transform 1 0 14812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_155
timestamp 1644511149
transform 1 0 15364 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_167
timestamp 1644511149
transform 1 0 16468 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_179
timestamp 1644511149
transform 1 0 17572 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_191
timestamp 1644511149
transform 1 0 18676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_257
timestamp 1644511149
transform 1 0 24748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_260
timestamp 1644511149
transform 1 0 25024 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_266
timestamp 1644511149
transform 1 0 25576 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_272
timestamp 1644511149
transform 1 0 26128 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_278
timestamp 1644511149
transform 1 0 26680 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_286
timestamp 1644511149
transform 1 0 27416 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_292
timestamp 1644511149
transform 1 0 27968 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_298
timestamp 1644511149
transform 1 0 28520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1644511149
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_313
timestamp 1644511149
transform 1 0 29900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_329
timestamp 1644511149
transform 1 0 31372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_336
timestamp 1644511149
transform 1 0 32016 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_342
timestamp 1644511149
transform 1 0 32568 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_348
timestamp 1644511149
transform 1 0 33120 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_354
timestamp 1644511149
transform 1 0 33672 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_360
timestamp 1644511149
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_367
timestamp 1644511149
transform 1 0 34868 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_373
timestamp 1644511149
transform 1 0 35420 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_379
timestamp 1644511149
transform 1 0 35972 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_385
timestamp 1644511149
transform 1 0 36524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_391
timestamp 1644511149
transform 1 0 37076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_397
timestamp 1644511149
transform 1 0 37628 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_409
timestamp 1644511149
transform 1 0 38732 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_417
timestamp 1644511149
transform 1 0 39468 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_501
timestamp 1644511149
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_513
timestamp 1644511149
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1644511149
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1644511149
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_533
timestamp 1644511149
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_545
timestamp 1644511149
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_557
timestamp 1644511149
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_569
timestamp 1644511149
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1644511149
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1644511149
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_589
timestamp 1644511149
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_601
timestamp 1644511149
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_613
timestamp 1644511149
transform 1 0 57500 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_621
timestamp 1644511149
transform 1 0 58236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_245
timestamp 1644511149
transform 1 0 23644 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_250
timestamp 1644511149
transform 1 0 24104 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_254
timestamp 1644511149
transform 1 0 24472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_257
timestamp 1644511149
transform 1 0 24748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_263
timestamp 1644511149
transform 1 0 25300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_267
timestamp 1644511149
transform 1 0 25668 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_270
timestamp 1644511149
transform 1 0 25944 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1644511149
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_283
timestamp 1644511149
transform 1 0 27140 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_289
timestamp 1644511149
transform 1 0 27692 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_295
timestamp 1644511149
transform 1 0 28244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_302
timestamp 1644511149
transform 1 0 28888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_313
timestamp 1644511149
transform 1 0 29900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_322
timestamp 1644511149
transform 1 0 30728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_331
timestamp 1644511149
transform 1 0 31556 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_341
timestamp 1644511149
transform 1 0 32476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_348
timestamp 1644511149
transform 1 0 33120 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_354
timestamp 1644511149
transform 1 0 33672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_360
timestamp 1644511149
transform 1 0 34224 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_366
timestamp 1644511149
transform 1 0 34776 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_372
timestamp 1644511149
transform 1 0 35328 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_378
timestamp 1644511149
transform 1 0 35880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_384
timestamp 1644511149
transform 1 0 36432 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_395
timestamp 1644511149
transform 1 0 37444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_401
timestamp 1644511149
transform 1 0 37996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_407
timestamp 1644511149
transform 1 0 38548 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_419
timestamp 1644511149
transform 1 0 39652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_431
timestamp 1644511149
transform 1 0 40756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_443
timestamp 1644511149
transform 1 0 41860 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_517
timestamp 1644511149
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_529
timestamp 1644511149
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_541
timestamp 1644511149
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1644511149
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1644511149
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_561
timestamp 1644511149
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_573
timestamp 1644511149
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_585
timestamp 1644511149
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_597
timestamp 1644511149
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1644511149
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1644511149
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1644511149
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_7
timestamp 1644511149
transform 1 0 1748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_19
timestamp 1644511149
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_236
timestamp 1644511149
transform 1 0 22816 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_242
timestamp 1644511149
transform 1 0 23368 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1644511149
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_257
timestamp 1644511149
transform 1 0 24748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_260
timestamp 1644511149
transform 1 0 25024 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_266
timestamp 1644511149
transform 1 0 25576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_272
timestamp 1644511149
transform 1 0 26128 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_278
timestamp 1644511149
transform 1 0 26680 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_284
timestamp 1644511149
transform 1 0 27232 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_290
timestamp 1644511149
transform 1 0 27784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_296
timestamp 1644511149
transform 1 0 28336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1644511149
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_314
timestamp 1644511149
transform 1 0 29992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_325
timestamp 1644511149
transform 1 0 31004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_335
timestamp 1644511149
transform 1 0 31924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_343
timestamp 1644511149
transform 1 0 32660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_347
timestamp 1644511149
transform 1 0 33028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_352
timestamp 1644511149
transform 1 0 33488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_359
timestamp 1644511149
transform 1 0 34132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_367
timestamp 1644511149
transform 1 0 34868 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_373
timestamp 1644511149
transform 1 0 35420 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_379
timestamp 1644511149
transform 1 0 35972 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_385
timestamp 1644511149
transform 1 0 36524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_391
timestamp 1644511149
transform 1 0 37076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_397
timestamp 1644511149
transform 1 0 37628 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_403
timestamp 1644511149
transform 1 0 38180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_409
timestamp 1644511149
transform 1 0 38732 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_415
timestamp 1644511149
transform 1 0 39284 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_513
timestamp 1644511149
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1644511149
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1644511149
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_533
timestamp 1644511149
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_545
timestamp 1644511149
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_557
timestamp 1644511149
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_569
timestamp 1644511149
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1644511149
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1644511149
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_589
timestamp 1644511149
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_601
timestamp 1644511149
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_613
timestamp 1644511149
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_104
timestamp 1644511149
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_115
timestamp 1644511149
transform 1 0 11684 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_127
timestamp 1644511149
transform 1 0 12788 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_139
timestamp 1644511149
transform 1 0 13892 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_151
timestamp 1644511149
transform 1 0 14996 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_163
timestamp 1644511149
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_230
timestamp 1644511149
transform 1 0 22264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_236
timestamp 1644511149
transform 1 0 22816 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_242
timestamp 1644511149
transform 1 0 23368 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_248
timestamp 1644511149
transform 1 0 23920 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_251
timestamp 1644511149
transform 1 0 24196 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_257
timestamp 1644511149
transform 1 0 24748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_263
timestamp 1644511149
transform 1 0 25300 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_274
timestamp 1644511149
transform 1 0 26312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_289
timestamp 1644511149
transform 1 0 27692 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_300
timestamp 1644511149
transform 1 0 28704 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_309
timestamp 1644511149
transform 1 0 29532 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_320
timestamp 1644511149
transform 1 0 30544 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_331
timestamp 1644511149
transform 1 0 31556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_344
timestamp 1644511149
transform 1 0 32752 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_352
timestamp 1644511149
transform 1 0 33488 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_358
timestamp 1644511149
transform 1 0 34040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_365
timestamp 1644511149
transform 1 0 34684 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_372
timestamp 1644511149
transform 1 0 35328 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_378
timestamp 1644511149
transform 1 0 35880 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_384
timestamp 1644511149
transform 1 0 36432 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_395
timestamp 1644511149
transform 1 0 37444 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_401
timestamp 1644511149
transform 1 0 37996 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_407
timestamp 1644511149
transform 1 0 38548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_413
timestamp 1644511149
transform 1 0 39100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_419
timestamp 1644511149
transform 1 0 39652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_425
timestamp 1644511149
transform 1 0 40204 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_437
timestamp 1644511149
transform 1 0 41308 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_445
timestamp 1644511149
transform 1 0 42044 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_517
timestamp 1644511149
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_529
timestamp 1644511149
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_541
timestamp 1644511149
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1644511149
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1644511149
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_561
timestamp 1644511149
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_573
timestamp 1644511149
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_585
timestamp 1644511149
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_597
timestamp 1644511149
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1644511149
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1644511149
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_617
timestamp 1644511149
transform 1 0 57868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_621
timestamp 1644511149
transform 1 0 58236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_215
timestamp 1644511149
transform 1 0 20884 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_218
timestamp 1644511149
transform 1 0 21160 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_224
timestamp 1644511149
transform 1 0 21712 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_230
timestamp 1644511149
transform 1 0 22264 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_236
timestamp 1644511149
transform 1 0 22816 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_242
timestamp 1644511149
transform 1 0 23368 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1644511149
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_256
timestamp 1644511149
transform 1 0 24656 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_264
timestamp 1644511149
transform 1 0 25392 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_276
timestamp 1644511149
transform 1 0 26496 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_284
timestamp 1644511149
transform 1 0 27232 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_293
timestamp 1644511149
transform 1 0 28060 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1644511149
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_331
timestamp 1644511149
transform 1 0 31556 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_349
timestamp 1644511149
transform 1 0 33212 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_360
timestamp 1644511149
transform 1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_369
timestamp 1644511149
transform 1 0 35052 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_376
timestamp 1644511149
transform 1 0 35696 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_383
timestamp 1644511149
transform 1 0 36340 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_395
timestamp 1644511149
transform 1 0 37444 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_407
timestamp 1644511149
transform 1 0 38548 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_423
timestamp 1644511149
transform 1 0 40020 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_429
timestamp 1644511149
transform 1 0 40572 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_435
timestamp 1644511149
transform 1 0 41124 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_447
timestamp 1644511149
transform 1 0 42228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_459
timestamp 1644511149
transform 1 0 43332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_471
timestamp 1644511149
transform 1 0 44436 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_501
timestamp 1644511149
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_513
timestamp 1644511149
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1644511149
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1644511149
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_533
timestamp 1644511149
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_545
timestamp 1644511149
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_557
timestamp 1644511149
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_569
timestamp 1644511149
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1644511149
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1644511149
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_589
timestamp 1644511149
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_601
timestamp 1644511149
transform 1 0 56396 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_609
timestamp 1644511149
transform 1 0 57132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_621
timestamp 1644511149
transform 1 0 58236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_7
timestamp 1644511149
transform 1 0 1748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_19
timestamp 1644511149
transform 1 0 2852 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_31
timestamp 1644511149
transform 1 0 3956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_43
timestamp 1644511149
transform 1 0 5060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_116
timestamp 1644511149
transform 1 0 11776 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_122
timestamp 1644511149
transform 1 0 12328 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_134
timestamp 1644511149
transform 1 0 13432 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_146
timestamp 1644511149
transform 1 0 14536 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_158
timestamp 1644511149
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1644511149
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_208
timestamp 1644511149
transform 1 0 20240 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_214
timestamp 1644511149
transform 1 0 20792 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1644511149
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_229
timestamp 1644511149
transform 1 0 22172 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_235
timestamp 1644511149
transform 1 0 22724 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_241
timestamp 1644511149
transform 1 0 23276 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_247
timestamp 1644511149
transform 1 0 23828 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_253
timestamp 1644511149
transform 1 0 24380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_260
timestamp 1644511149
transform 1 0 25024 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_268
timestamp 1644511149
transform 1 0 25760 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1644511149
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_285
timestamp 1644511149
transform 1 0 27324 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_321
timestamp 1644511149
transform 1 0 30636 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_324
timestamp 1644511149
transform 1 0 30912 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_332
timestamp 1644511149
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_351
timestamp 1644511149
transform 1 0 33396 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_370
timestamp 1644511149
transform 1 0 35144 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_377
timestamp 1644511149
transform 1 0 35788 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_384
timestamp 1644511149
transform 1 0 36432 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_395
timestamp 1644511149
transform 1 0 37444 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_401
timestamp 1644511149
transform 1 0 37996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_407
timestamp 1644511149
transform 1 0 38548 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_413
timestamp 1644511149
transform 1 0 39100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_419
timestamp 1644511149
transform 1 0 39652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_425
timestamp 1644511149
transform 1 0 40204 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_431
timestamp 1644511149
transform 1 0 40756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_437
timestamp 1644511149
transform 1 0 41308 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_443
timestamp 1644511149
transform 1 0 41860 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_517
timestamp 1644511149
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_529
timestamp 1644511149
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_541
timestamp 1644511149
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1644511149
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1644511149
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_561
timestamp 1644511149
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_573
timestamp 1644511149
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_585
timestamp 1644511149
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_597
timestamp 1644511149
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1644511149
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1644511149
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_617
timestamp 1644511149
transform 1 0 57868 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_621
timestamp 1644511149
transform 1 0 58236 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_199
timestamp 1644511149
transform 1 0 19412 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_205
timestamp 1644511149
transform 1 0 19964 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_211
timestamp 1644511149
transform 1 0 20516 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_215
timestamp 1644511149
transform 1 0 20884 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_218
timestamp 1644511149
transform 1 0 21160 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_224
timestamp 1644511149
transform 1 0 21712 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_230
timestamp 1644511149
transform 1 0 22264 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_236
timestamp 1644511149
transform 1 0 22816 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_242
timestamp 1644511149
transform 1 0 23368 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1644511149
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_257
timestamp 1644511149
transform 1 0 24748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_261
timestamp 1644511149
transform 1 0 25116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_269
timestamp 1644511149
transform 1 0 25852 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_280
timestamp 1644511149
transform 1 0 26864 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_291
timestamp 1644511149
transform 1 0 27876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1644511149
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_346
timestamp 1644511149
transform 1 0 32936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_360
timestamp 1644511149
transform 1 0 34224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_371
timestamp 1644511149
transform 1 0 35236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_380
timestamp 1644511149
transform 1 0 36064 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_387
timestamp 1644511149
transform 1 0 36708 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_394
timestamp 1644511149
transform 1 0 37352 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_400
timestamp 1644511149
transform 1 0 37904 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_406
timestamp 1644511149
transform 1 0 38456 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_412
timestamp 1644511149
transform 1 0 39008 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_423
timestamp 1644511149
transform 1 0 40020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_429
timestamp 1644511149
transform 1 0 40572 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_435
timestamp 1644511149
transform 1 0 41124 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_441
timestamp 1644511149
transform 1 0 41676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_447
timestamp 1644511149
transform 1 0 42228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_453
timestamp 1644511149
transform 1 0 42780 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_465
timestamp 1644511149
transform 1 0 43884 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_473
timestamp 1644511149
transform 1 0 44620 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_501
timestamp 1644511149
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_513
timestamp 1644511149
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1644511149
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1644511149
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_533
timestamp 1644511149
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_545
timestamp 1644511149
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_557
timestamp 1644511149
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_569
timestamp 1644511149
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1644511149
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1644511149
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_589
timestamp 1644511149
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_601
timestamp 1644511149
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_613
timestamp 1644511149
transform 1 0 57500 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_621
timestamp 1644511149
transform 1 0 58236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 1644511149
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_192
timestamp 1644511149
transform 1 0 18768 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_198
timestamp 1644511149
transform 1 0 19320 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_204
timestamp 1644511149
transform 1 0 19872 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_212
timestamp 1644511149
transform 1 0 20608 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_218
timestamp 1644511149
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_228
timestamp 1644511149
transform 1 0 22080 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_234
timestamp 1644511149
transform 1 0 22632 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_240
timestamp 1644511149
transform 1 0 23184 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_247
timestamp 1644511149
transform 1 0 23828 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_254
timestamp 1644511149
transform 1 0 24472 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_265
timestamp 1644511149
transform 1 0 25484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_276
timestamp 1644511149
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_307
timestamp 1644511149
transform 1 0 29348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_311
timestamp 1644511149
transform 1 0 29716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1644511149
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_357
timestamp 1644511149
transform 1 0 33948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_371
timestamp 1644511149
transform 1 0 35236 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_381
timestamp 1644511149
transform 1 0 36156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_388
timestamp 1644511149
transform 1 0 36800 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_396
timestamp 1644511149
transform 1 0 37536 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_403
timestamp 1644511149
transform 1 0 38180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_407
timestamp 1644511149
transform 1 0 38548 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_410
timestamp 1644511149
transform 1 0 38824 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_416
timestamp 1644511149
transform 1 0 39376 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_422
timestamp 1644511149
transform 1 0 39928 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_428
timestamp 1644511149
transform 1 0 40480 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_434
timestamp 1644511149
transform 1 0 41032 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_440
timestamp 1644511149
transform 1 0 41584 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_451
timestamp 1644511149
transform 1 0 42596 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_457
timestamp 1644511149
transform 1 0 43148 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_463
timestamp 1644511149
transform 1 0 43700 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_475
timestamp 1644511149
transform 1 0 44804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_487
timestamp 1644511149
transform 1 0 45908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_499
timestamp 1644511149
transform 1 0 47012 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_517
timestamp 1644511149
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_529
timestamp 1644511149
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_541
timestamp 1644511149
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1644511149
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1644511149
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_561
timestamp 1644511149
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_573
timestamp 1644511149
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_585
timestamp 1644511149
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_597
timestamp 1644511149
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1644511149
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1644511149
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1644511149
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_7
timestamp 1644511149
transform 1 0 1748 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_19
timestamp 1644511149
transform 1 0 2852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_117
timestamp 1644511149
transform 1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_123
timestamp 1644511149
transform 1 0 12420 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_129
timestamp 1644511149
transform 1 0 12972 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1644511149
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_183
timestamp 1644511149
transform 1 0 17940 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1644511149
transform 1 0 18216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1644511149
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_201
timestamp 1644511149
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_204
timestamp 1644511149
transform 1 0 19872 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1644511149
transform 1 0 20424 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_216
timestamp 1644511149
transform 1 0 20976 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_224
timestamp 1644511149
transform 1 0 21712 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_227
timestamp 1644511149
transform 1 0 21988 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_240
timestamp 1644511149
transform 1 0 23184 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1644511149
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_258
timestamp 1644511149
transform 1 0 24840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_269
timestamp 1644511149
transform 1 0 25852 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_280
timestamp 1644511149
transform 1 0 26864 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1644511149
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_331
timestamp 1644511149
transform 1 0 31556 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_355
timestamp 1644511149
transform 1 0 33764 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_375
timestamp 1644511149
transform 1 0 35604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_386
timestamp 1644511149
transform 1 0 36616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_394
timestamp 1644511149
transform 1 0 37352 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_402
timestamp 1644511149
transform 1 0 38088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_409
timestamp 1644511149
transform 1 0 38732 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_415
timestamp 1644511149
transform 1 0 39284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_423
timestamp 1644511149
transform 1 0 40020 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_429
timestamp 1644511149
transform 1 0 40572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_435
timestamp 1644511149
transform 1 0 41124 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_441
timestamp 1644511149
transform 1 0 41676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_447
timestamp 1644511149
transform 1 0 42228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_453
timestamp 1644511149
transform 1 0 42780 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_459
timestamp 1644511149
transform 1 0 43332 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_465
timestamp 1644511149
transform 1 0 43884 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_471
timestamp 1644511149
transform 1 0 44436 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1644511149
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1644511149
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_533
timestamp 1644511149
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_545
timestamp 1644511149
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_557
timestamp 1644511149
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_569
timestamp 1644511149
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1644511149
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1644511149
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_589
timestamp 1644511149
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_601
timestamp 1644511149
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_613
timestamp 1644511149
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_172
timestamp 1644511149
transform 1 0 16928 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1644511149
transform 1 0 17480 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_184
timestamp 1644511149
transform 1 0 18032 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_190
timestamp 1644511149
transform 1 0 18584 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_196
timestamp 1644511149
transform 1 0 19136 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_202
timestamp 1644511149
transform 1 0 19688 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_208
timestamp 1644511149
transform 1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_214
timestamp 1644511149
transform 1 0 20792 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1644511149
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_229
timestamp 1644511149
transform 1 0 22172 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_233
timestamp 1644511149
transform 1 0 22540 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_241
timestamp 1644511149
transform 1 0 23276 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_252
timestamp 1644511149
transform 1 0 24288 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_263
timestamp 1644511149
transform 1 0 25300 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1644511149
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_357
timestamp 1644511149
transform 1 0 33948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_375
timestamp 1644511149
transform 1 0 35604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_386
timestamp 1644511149
transform 1 0 36616 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_400
timestamp 1644511149
transform 1 0 37904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_408
timestamp 1644511149
transform 1 0 38640 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_415
timestamp 1644511149
transform 1 0 39284 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_422
timestamp 1644511149
transform 1 0 39928 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_426
timestamp 1644511149
transform 1 0 40296 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_435
timestamp 1644511149
transform 1 0 41124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_451
timestamp 1644511149
transform 1 0 42596 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_457
timestamp 1644511149
transform 1 0 43148 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_463
timestamp 1644511149
transform 1 0 43700 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_469
timestamp 1644511149
transform 1 0 44252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_475
timestamp 1644511149
transform 1 0 44804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_481
timestamp 1644511149
transform 1 0 45356 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_493
timestamp 1644511149
transform 1 0 46460 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_501
timestamp 1644511149
transform 1 0 47196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_517
timestamp 1644511149
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_529
timestamp 1644511149
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_541
timestamp 1644511149
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1644511149
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1644511149
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_561
timestamp 1644511149
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_573
timestamp 1644511149
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_585
timestamp 1644511149
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_597
timestamp 1644511149
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1644511149
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1644511149
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_617
timestamp 1644511149
transform 1 0 57868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_621
timestamp 1644511149
transform 1 0 58236 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_114
timestamp 1644511149
transform 1 0 11592 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_120
timestamp 1644511149
transform 1 0 12144 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_132
timestamp 1644511149
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_161
timestamp 1644511149
transform 1 0 15916 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_164
timestamp 1644511149
transform 1 0 16192 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_170
timestamp 1644511149
transform 1 0 16744 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_176
timestamp 1644511149
transform 1 0 17296 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_182
timestamp 1644511149
transform 1 0 17848 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_188
timestamp 1644511149
transform 1 0 18400 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_202
timestamp 1644511149
transform 1 0 19688 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_208
timestamp 1644511149
transform 1 0 20240 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_214
timestamp 1644511149
transform 1 0 20792 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1644511149
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_266
timestamp 1644511149
transform 1 0 25576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_280
timestamp 1644511149
transform 1 0 26864 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1644511149
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_332
timestamp 1644511149
transform 1 0 31648 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_356
timestamp 1644511149
transform 1 0 33856 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_379
timestamp 1644511149
transform 1 0 35972 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_397
timestamp 1644511149
transform 1 0 37628 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_408
timestamp 1644511149
transform 1 0 38640 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_416
timestamp 1644511149
transform 1 0 39376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_424
timestamp 1644511149
transform 1 0 40112 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_431
timestamp 1644511149
transform 1 0 40756 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_437
timestamp 1644511149
transform 1 0 41308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_443
timestamp 1644511149
transform 1 0 41860 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_449
timestamp 1644511149
transform 1 0 42412 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_455
timestamp 1644511149
transform 1 0 42964 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_461
timestamp 1644511149
transform 1 0 43516 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_467
timestamp 1644511149
transform 1 0 44068 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_479
timestamp 1644511149
transform 1 0 45172 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_485
timestamp 1644511149
transform 1 0 45724 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_491
timestamp 1644511149
transform 1 0 46276 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_503
timestamp 1644511149
transform 1 0 47380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_515
timestamp 1644511149
transform 1 0 48484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_527
timestamp 1644511149
transform 1 0 49588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1644511149
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_533
timestamp 1644511149
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_545
timestamp 1644511149
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_557
timestamp 1644511149
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_569
timestamp 1644511149
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1644511149
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1644511149
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_589
timestamp 1644511149
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_601
timestamp 1644511149
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_613
timestamp 1644511149
transform 1 0 57500 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_621
timestamp 1644511149
transform 1 0 58236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_7
timestamp 1644511149
transform 1 0 1748 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_19
timestamp 1644511149
transform 1 0 2852 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_31
timestamp 1644511149
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_43
timestamp 1644511149
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_155
timestamp 1644511149
transform 1 0 15364 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_158
timestamp 1644511149
transform 1 0 15640 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1644511149
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_173
timestamp 1644511149
transform 1 0 17020 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_176
timestamp 1644511149
transform 1 0 17296 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_182
timestamp 1644511149
transform 1 0 17848 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_188
timestamp 1644511149
transform 1 0 18400 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_194
timestamp 1644511149
transform 1 0 18952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_200
timestamp 1644511149
transform 1 0 19504 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_208
timestamp 1644511149
transform 1 0 20240 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_212
timestamp 1644511149
transform 1 0 20608 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1644511149
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_230
timestamp 1644511149
transform 1 0 22264 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_241
timestamp 1644511149
transform 1 0 23276 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_252
timestamp 1644511149
transform 1 0 24288 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1644511149
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_285
timestamp 1644511149
transform 1 0 27324 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_306
timestamp 1644511149
transform 1 0 29256 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_330
timestamp 1644511149
transform 1 0 31464 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_357
timestamp 1644511149
transform 1 0 33948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_381
timestamp 1644511149
transform 1 0 36156 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_388
timestamp 1644511149
transform 1 0 36800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_407
timestamp 1644511149
transform 1 0 38548 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_418
timestamp 1644511149
transform 1 0 39560 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_426
timestamp 1644511149
transform 1 0 40296 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_434
timestamp 1644511149
transform 1 0 41032 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_451
timestamp 1644511149
transform 1 0 42596 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_457
timestamp 1644511149
transform 1 0 43148 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_463
timestamp 1644511149
transform 1 0 43700 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_469
timestamp 1644511149
transform 1 0 44252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_475
timestamp 1644511149
transform 1 0 44804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_481
timestamp 1644511149
transform 1 0 45356 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_487
timestamp 1644511149
transform 1 0 45908 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_493
timestamp 1644511149
transform 1 0 46460 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_499
timestamp 1644511149
transform 1 0 47012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_517
timestamp 1644511149
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_529
timestamp 1644511149
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_541
timestamp 1644511149
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1644511149
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1644511149
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_561
timestamp 1644511149
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_573
timestamp 1644511149
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_585
timestamp 1644511149
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_597
timestamp 1644511149
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1644511149
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1644511149
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1644511149
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_106
timestamp 1644511149
transform 1 0 10856 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_112
timestamp 1644511149
transform 1 0 11408 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_124
timestamp 1644511149
transform 1 0 12512 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1644511149
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_144
timestamp 1644511149
transform 1 0 14352 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_150
timestamp 1644511149
transform 1 0 14904 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_156
timestamp 1644511149
transform 1 0 15456 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_162
timestamp 1644511149
transform 1 0 16008 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_168
timestamp 1644511149
transform 1 0 16560 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_174
timestamp 1644511149
transform 1 0 17112 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_180
timestamp 1644511149
transform 1 0 17664 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_186
timestamp 1644511149
transform 1 0 18216 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1644511149
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_204
timestamp 1644511149
transform 1 0 19872 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_212
timestamp 1644511149
transform 1 0 20608 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_223
timestamp 1644511149
transform 1 0 21620 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_234
timestamp 1644511149
transform 1 0 22632 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1644511149
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_256
timestamp 1644511149
transform 1 0 24656 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_280
timestamp 1644511149
transform 1 0 26864 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1644511149
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_319
timestamp 1644511149
transform 1 0 30452 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_344
timestamp 1644511149
transform 1 0 32752 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_358
timestamp 1644511149
transform 1 0 34040 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_385
timestamp 1644511149
transform 1 0 36524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_403
timestamp 1644511149
transform 1 0 38180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_414
timestamp 1644511149
transform 1 0 39192 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_427
timestamp 1644511149
transform 1 0 40388 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_435
timestamp 1644511149
transform 1 0 41124 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_443
timestamp 1644511149
transform 1 0 41860 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_450
timestamp 1644511149
transform 1 0 42504 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_456
timestamp 1644511149
transform 1 0 43056 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_462
timestamp 1644511149
transform 1 0 43608 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_468
timestamp 1644511149
transform 1 0 44160 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_479
timestamp 1644511149
transform 1 0 45172 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_485
timestamp 1644511149
transform 1 0 45724 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_491
timestamp 1644511149
transform 1 0 46276 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_497
timestamp 1644511149
transform 1 0 46828 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_503
timestamp 1644511149
transform 1 0 47380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_509
timestamp 1644511149
transform 1 0 47932 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_521
timestamp 1644511149
transform 1 0 49036 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_529
timestamp 1644511149
transform 1 0 49772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_533
timestamp 1644511149
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_545
timestamp 1644511149
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_557
timestamp 1644511149
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_569
timestamp 1644511149
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1644511149
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1644511149
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_589
timestamp 1644511149
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_601
timestamp 1644511149
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_613
timestamp 1644511149
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_7
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_19
timestamp 1644511149
transform 1 0 2852 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_31
timestamp 1644511149
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_43
timestamp 1644511149
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_140
timestamp 1644511149
transform 1 0 13984 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_146
timestamp 1644511149
transform 1 0 14536 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_152
timestamp 1644511149
transform 1 0 15088 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_158
timestamp 1644511149
transform 1 0 15640 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1644511149
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_172
timestamp 1644511149
transform 1 0 16928 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_178
timestamp 1644511149
transform 1 0 17480 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1644511149
transform 1 0 18032 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_191
timestamp 1644511149
transform 1 0 18676 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_198
timestamp 1644511149
transform 1 0 19320 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_209
timestamp 1644511149
transform 1 0 20332 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1644511149
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_238
timestamp 1644511149
transform 1 0 23000 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_252
timestamp 1644511149
transform 1 0 24288 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1644511149
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_283
timestamp 1644511149
transform 1 0 27140 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_307
timestamp 1644511149
transform 1 0 29348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_332
timestamp 1644511149
transform 1 0 31648 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_358
timestamp 1644511149
transform 1 0 34040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_382
timestamp 1644511149
transform 1 0 36248 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1644511149
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_407
timestamp 1644511149
transform 1 0 38548 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_425
timestamp 1644511149
transform 1 0 40204 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_436
timestamp 1644511149
transform 1 0 41216 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_444
timestamp 1644511149
transform 1 0 41952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_457
timestamp 1644511149
transform 1 0 43148 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_464
timestamp 1644511149
transform 1 0 43792 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_470
timestamp 1644511149
transform 1 0 44344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_476
timestamp 1644511149
transform 1 0 44896 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_482
timestamp 1644511149
transform 1 0 45448 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_488
timestamp 1644511149
transform 1 0 46000 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_494
timestamp 1644511149
transform 1 0 46552 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_500
timestamp 1644511149
transform 1 0 47104 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_507
timestamp 1644511149
transform 1 0 47748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_513
timestamp 1644511149
transform 1 0 48300 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_525
timestamp 1644511149
transform 1 0 49404 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_537
timestamp 1644511149
transform 1 0 50508 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_549
timestamp 1644511149
transform 1 0 51612 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_557
timestamp 1644511149
transform 1 0 52348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_561
timestamp 1644511149
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_573
timestamp 1644511149
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_585
timestamp 1644511149
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_597
timestamp 1644511149
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1644511149
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1644511149
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_617
timestamp 1644511149
transform 1 0 57868 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_621
timestamp 1644511149
transform 1 0 58236 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_113
timestamp 1644511149
transform 1 0 11500 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_119
timestamp 1644511149
transform 1 0 12052 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_127
timestamp 1644511149
transform 1 0 12788 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_130
timestamp 1644511149
transform 1 0 13064 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1644511149
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_147
timestamp 1644511149
transform 1 0 14628 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1644511149
transform 1 0 15732 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_171
timestamp 1644511149
transform 1 0 16836 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_184
timestamp 1644511149
transform 1 0 18032 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_205
timestamp 1644511149
transform 1 0 19964 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_216
timestamp 1644511149
transform 1 0 20976 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_228
timestamp 1644511149
transform 1 0 22080 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1644511149
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_256
timestamp 1644511149
transform 1 0 24656 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_280
timestamp 1644511149
transform 1 0 26864 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1644511149
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_313
timestamp 1644511149
transform 1 0 29900 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_335
timestamp 1644511149
transform 1 0 31924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_360
timestamp 1644511149
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_385
timestamp 1644511149
transform 1 0 36524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_409
timestamp 1644511149
transform 1 0 38732 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_416
timestamp 1644511149
transform 1 0 39376 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_435
timestamp 1644511149
transform 1 0 41124 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_453
timestamp 1644511149
transform 1 0 42780 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_461
timestamp 1644511149
transform 1 0 43516 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_468
timestamp 1644511149
transform 1 0 44160 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_479
timestamp 1644511149
transform 1 0 45172 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_485
timestamp 1644511149
transform 1 0 45724 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_491
timestamp 1644511149
transform 1 0 46276 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_497
timestamp 1644511149
transform 1 0 46828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_503
timestamp 1644511149
transform 1 0 47380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_509
timestamp 1644511149
transform 1 0 47932 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_515
timestamp 1644511149
transform 1 0 48484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_521
timestamp 1644511149
transform 1 0 49036 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_527
timestamp 1644511149
transform 1 0 49588 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1644511149
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_533
timestamp 1644511149
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_545
timestamp 1644511149
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_557
timestamp 1644511149
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_569
timestamp 1644511149
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1644511149
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1644511149
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_589
timestamp 1644511149
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_601
timestamp 1644511149
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_613
timestamp 1644511149
transform 1 0 57500 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_621
timestamp 1644511149
transform 1 0 58236 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1644511149
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_122
timestamp 1644511149
transform 1 0 12328 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_128
timestamp 1644511149
transform 1 0 12880 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_134
timestamp 1644511149
transform 1 0 13432 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_140
timestamp 1644511149
transform 1 0 13984 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_146
timestamp 1644511149
transform 1 0 14536 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_152
timestamp 1644511149
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_158
timestamp 1644511149
transform 1 0 15640 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1644511149
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_171
timestamp 1644511149
transform 1 0 16836 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1644511149
transform 1 0 17480 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_186
timestamp 1644511149
transform 1 0 18216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_197
timestamp 1644511149
transform 1 0 19228 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1644511149
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1644511149
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_228
timestamp 1644511149
transform 1 0 22080 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_252
timestamp 1644511149
transform 1 0 24288 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1644511149
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_331
timestamp 1644511149
transform 1 0 31556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_358
timestamp 1644511149
transform 1 0 34040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_383
timestamp 1644511149
transform 1 0 36340 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_413
timestamp 1644511149
transform 1 0 39100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_430
timestamp 1644511149
transform 1 0 40664 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_444
timestamp 1644511149
transform 1 0 41952 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_455
timestamp 1644511149
transform 1 0 42964 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_463
timestamp 1644511149
transform 1 0 43700 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_471
timestamp 1644511149
transform 1 0 44436 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_478
timestamp 1644511149
transform 1 0 45080 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_484
timestamp 1644511149
transform 1 0 45632 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_490
timestamp 1644511149
transform 1 0 46184 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_496
timestamp 1644511149
transform 1 0 46736 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_507
timestamp 1644511149
transform 1 0 47748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_513
timestamp 1644511149
transform 1 0 48300 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_519
timestamp 1644511149
transform 1 0 48852 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_525
timestamp 1644511149
transform 1 0 49404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_531
timestamp 1644511149
transform 1 0 49956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_543
timestamp 1644511149
transform 1 0 51060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_555
timestamp 1644511149
transform 1 0 52164 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1644511149
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_561
timestamp 1644511149
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_573
timestamp 1644511149
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_585
timestamp 1644511149
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_597
timestamp 1644511149
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1644511149
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1644511149
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_617
timestamp 1644511149
transform 1 0 57868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_621
timestamp 1644511149
transform 1 0 58236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_7
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1644511149
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_115
timestamp 1644511149
transform 1 0 11684 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_118
timestamp 1644511149
transform 1 0 11960 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_124
timestamp 1644511149
transform 1 0 12512 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_130
timestamp 1644511149
transform 1 0 13064 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_144
timestamp 1644511149
transform 1 0 14352 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_150
timestamp 1644511149
transform 1 0 14904 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_156
timestamp 1644511149
transform 1 0 15456 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1644511149
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1644511149
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_181
timestamp 1644511149
transform 1 0 17756 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_207
timestamp 1644511149
transform 1 0 20148 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_224
timestamp 1644511149
transform 1 0 21712 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1644511149
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_255
timestamp 1644511149
transform 1 0 24564 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_279
timestamp 1644511149
transform 1 0 26772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1644511149
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_334
timestamp 1644511149
transform 1 0 31832 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1644511149
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_386
timestamp 1644511149
transform 1 0 36616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_410
timestamp 1644511149
transform 1 0 38824 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_416
timestamp 1644511149
transform 1 0 39376 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_441
timestamp 1644511149
transform 1 0 41676 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_452
timestamp 1644511149
transform 1 0 42688 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_463
timestamp 1644511149
transform 1 0 43700 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_472
timestamp 1644511149
transform 1 0 44528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_481
timestamp 1644511149
transform 1 0 45356 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_488
timestamp 1644511149
transform 1 0 46000 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_494
timestamp 1644511149
transform 1 0 46552 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_500
timestamp 1644511149
transform 1 0 47104 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_506
timestamp 1644511149
transform 1 0 47656 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_518
timestamp 1644511149
transform 1 0 48760 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_524
timestamp 1644511149
transform 1 0 49312 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_535
timestamp 1644511149
transform 1 0 50324 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_547
timestamp 1644511149
transform 1 0 51428 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_559
timestamp 1644511149
transform 1 0 52532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_571
timestamp 1644511149
transform 1 0 53636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_583
timestamp 1644511149
transform 1 0 54740 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1644511149
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_589
timestamp 1644511149
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_601
timestamp 1644511149
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_613
timestamp 1644511149
transform 1 0 57500 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_621
timestamp 1644511149
transform 1 0 58236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1644511149
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_117
timestamp 1644511149
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_120
timestamp 1644511149
transform 1 0 12144 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_126
timestamp 1644511149
transform 1 0 12696 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_133
timestamp 1644511149
transform 1 0 13340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_143
timestamp 1644511149
transform 1 0 14260 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_156
timestamp 1644511149
transform 1 0 15456 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1644511149
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_179
timestamp 1644511149
transform 1 0 17572 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_190
timestamp 1644511149
transform 1 0 18584 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_202
timestamp 1644511149
transform 1 0 19688 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1644511149
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_228
timestamp 1644511149
transform 1 0 22080 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_252
timestamp 1644511149
transform 1 0 24288 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1644511149
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_303
timestamp 1644511149
transform 1 0 28980 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_328
timestamp 1644511149
transform 1 0 31280 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_358
timestamp 1644511149
transform 1 0 34040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_383
timestamp 1644511149
transform 1 0 36340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_414
timestamp 1644511149
transform 1 0 39192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_438
timestamp 1644511149
transform 1 0 41400 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_444
timestamp 1644511149
transform 1 0 41952 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_459
timestamp 1644511149
transform 1 0 43332 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_470
timestamp 1644511149
transform 1 0 44344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_480
timestamp 1644511149
transform 1 0 45264 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_488
timestamp 1644511149
transform 1 0 46000 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_495
timestamp 1644511149
transform 1 0 46644 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_507
timestamp 1644511149
transform 1 0 47748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_513
timestamp 1644511149
transform 1 0 48300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_519
timestamp 1644511149
transform 1 0 48852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_525
timestamp 1644511149
transform 1 0 49404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_531
timestamp 1644511149
transform 1 0 49956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_537
timestamp 1644511149
transform 1 0 50508 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_549
timestamp 1644511149
transform 1 0 51612 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_557
timestamp 1644511149
transform 1 0 52348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_561
timestamp 1644511149
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_573
timestamp 1644511149
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_585
timestamp 1644511149
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_597
timestamp 1644511149
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1644511149
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1644511149
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1644511149
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_112
timestamp 1644511149
transform 1 0 11408 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_118
timestamp 1644511149
transform 1 0 11960 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_124
timestamp 1644511149
transform 1 0 12512 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_130
timestamp 1644511149
transform 1 0 13064 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1644511149
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_144
timestamp 1644511149
transform 1 0 14352 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_150
timestamp 1644511149
transform 1 0 14904 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_156
timestamp 1644511149
transform 1 0 15456 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_163
timestamp 1644511149
transform 1 0 16100 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1644511149
transform 1 0 16744 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_181
timestamp 1644511149
transform 1 0 17756 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1644511149
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_206
timestamp 1644511149
transform 1 0 20056 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_224
timestamp 1644511149
transform 1 0 21712 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1644511149
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_255
timestamp 1644511149
transform 1 0 24564 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_279
timestamp 1644511149
transform 1 0 26772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1644511149
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_332
timestamp 1644511149
transform 1 0 31648 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_386
timestamp 1644511149
transform 1 0 36616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_410
timestamp 1644511149
transform 1 0 38824 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_416
timestamp 1644511149
transform 1 0 39376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_441
timestamp 1644511149
transform 1 0 41676 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_454
timestamp 1644511149
transform 1 0 42872 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_465
timestamp 1644511149
transform 1 0 43884 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_472
timestamp 1644511149
transform 1 0 44528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_481
timestamp 1644511149
transform 1 0 45356 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_488
timestamp 1644511149
transform 1 0 46000 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_495
timestamp 1644511149
transform 1 0 46644 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_501
timestamp 1644511149
transform 1 0 47196 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_507
timestamp 1644511149
transform 1 0 47748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_513
timestamp 1644511149
transform 1 0 48300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_519
timestamp 1644511149
transform 1 0 48852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1644511149
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1644511149
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_535
timestamp 1644511149
transform 1 0 50324 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_547
timestamp 1644511149
transform 1 0 51428 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_559
timestamp 1644511149
transform 1 0 52532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_571
timestamp 1644511149
transform 1 0 53636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_583
timestamp 1644511149
transform 1 0 54740 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1644511149
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_589
timestamp 1644511149
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_601
timestamp 1644511149
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_613
timestamp 1644511149
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_7
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_19
timestamp 1644511149
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_31
timestamp 1644511149
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_43
timestamp 1644511149
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_115
timestamp 1644511149
transform 1 0 11684 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_121
timestamp 1644511149
transform 1 0 12236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_127
timestamp 1644511149
transform 1 0 12788 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_134
timestamp 1644511149
transform 1 0 13432 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_140
timestamp 1644511149
transform 1 0 13984 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_146
timestamp 1644511149
transform 1 0 14536 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_152
timestamp 1644511149
transform 1 0 15088 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_158
timestamp 1644511149
transform 1 0 15640 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1644511149
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_172
timestamp 1644511149
transform 1 0 16928 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1644511149
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_191
timestamp 1644511149
transform 1 0 18676 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_202
timestamp 1644511149
transform 1 0 19688 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_228
timestamp 1644511149
transform 1 0 22080 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_252
timestamp 1644511149
transform 1 0 24288 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1644511149
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_285
timestamp 1644511149
transform 1 0 27324 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_307
timestamp 1644511149
transform 1 0 29348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1644511149
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_358
timestamp 1644511149
transform 1 0 34040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_383
timestamp 1644511149
transform 1 0 36340 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_413
timestamp 1644511149
transform 1 0 39100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_437
timestamp 1644511149
transform 1 0 41308 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_444
timestamp 1644511149
transform 1 0 41952 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_456
timestamp 1644511149
transform 1 0 43056 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_464
timestamp 1644511149
transform 1 0 43792 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_472
timestamp 1644511149
transform 1 0 44528 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_479
timestamp 1644511149
transform 1 0 45172 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_491
timestamp 1644511149
transform 1 0 46276 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_507
timestamp 1644511149
transform 1 0 47748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_513
timestamp 1644511149
transform 1 0 48300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_519
timestamp 1644511149
transform 1 0 48852 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_525
timestamp 1644511149
transform 1 0 49404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_531
timestamp 1644511149
transform 1 0 49956 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_537
timestamp 1644511149
transform 1 0 50508 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_549
timestamp 1644511149
transform 1 0 51612 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_557
timestamp 1644511149
transform 1 0 52348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_561
timestamp 1644511149
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_573
timestamp 1644511149
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_585
timestamp 1644511149
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_597
timestamp 1644511149
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1644511149
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1644511149
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_617
timestamp 1644511149
transform 1 0 57868 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_621
timestamp 1644511149
transform 1 0 58236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_124
timestamp 1644511149
transform 1 0 12512 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_130
timestamp 1644511149
transform 1 0 13064 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_143
timestamp 1644511149
transform 1 0 14260 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1644511149
transform 1 0 14812 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_155
timestamp 1644511149
transform 1 0 15364 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_161
timestamp 1644511149
transform 1 0 15916 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_167
timestamp 1644511149
transform 1 0 16468 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_174
timestamp 1644511149
transform 1 0 17112 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1644511149
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1644511149
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_201
timestamp 1644511149
transform 1 0 19596 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_212
timestamp 1644511149
transform 1 0 20608 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_224
timestamp 1644511149
transform 1 0 21712 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1644511149
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_256
timestamp 1644511149
transform 1 0 24656 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_280
timestamp 1644511149
transform 1 0 26864 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_334
timestamp 1644511149
transform 1 0 31832 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_359
timestamp 1644511149
transform 1 0 34132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_385
timestamp 1644511149
transform 1 0 36524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_409
timestamp 1644511149
transform 1 0 38732 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_416
timestamp 1644511149
transform 1 0 39376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_441
timestamp 1644511149
transform 1 0 41676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_451
timestamp 1644511149
transform 1 0 42596 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_459
timestamp 1644511149
transform 1 0 43332 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_466
timestamp 1644511149
transform 1 0 43976 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_472
timestamp 1644511149
transform 1 0 44528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_479
timestamp 1644511149
transform 1 0 45172 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_485
timestamp 1644511149
transform 1 0 45724 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_491
timestamp 1644511149
transform 1 0 46276 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_497
timestamp 1644511149
transform 1 0 46828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_503
timestamp 1644511149
transform 1 0 47380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_509
timestamp 1644511149
transform 1 0 47932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_515
timestamp 1644511149
transform 1 0 48484 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_521
timestamp 1644511149
transform 1 0 49036 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_527
timestamp 1644511149
transform 1 0 49588 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1644511149
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_533
timestamp 1644511149
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_545
timestamp 1644511149
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_557
timestamp 1644511149
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_569
timestamp 1644511149
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1644511149
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1644511149
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_589
timestamp 1644511149
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_601
timestamp 1644511149
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_613
timestamp 1644511149
transform 1 0 57500 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_621
timestamp 1644511149
transform 1 0 58236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1644511149
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_128
timestamp 1644511149
transform 1 0 12880 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_136
timestamp 1644511149
transform 1 0 13616 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_146
timestamp 1644511149
transform 1 0 14536 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_152
timestamp 1644511149
transform 1 0 15088 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_158
timestamp 1644511149
transform 1 0 15640 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1644511149
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_171
timestamp 1644511149
transform 1 0 16836 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_177
timestamp 1644511149
transform 1 0 17388 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_184
timestamp 1644511149
transform 1 0 18032 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_191
timestamp 1644511149
transform 1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_198
timestamp 1644511149
transform 1 0 19320 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_209
timestamp 1644511149
transform 1 0 20332 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1644511149
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_234
timestamp 1644511149
transform 1 0 22632 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_252
timestamp 1644511149
transform 1 0 24288 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1644511149
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_283
timestamp 1644511149
transform 1 0 27140 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_307
timestamp 1644511149
transform 1 0 29348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1644511149
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_358
timestamp 1644511149
transform 1 0 34040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_382
timestamp 1644511149
transform 1 0 36248 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_388
timestamp 1644511149
transform 1 0 36800 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_413
timestamp 1644511149
transform 1 0 39100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_430
timestamp 1644511149
transform 1 0 40664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_440
timestamp 1644511149
transform 1 0 41584 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_453
timestamp 1644511149
transform 1 0 42780 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_460
timestamp 1644511149
transform 1 0 43424 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_467
timestamp 1644511149
transform 1 0 44068 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_479
timestamp 1644511149
transform 1 0 45172 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_491
timestamp 1644511149
transform 1 0 46276 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_507
timestamp 1644511149
transform 1 0 47748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_513
timestamp 1644511149
transform 1 0 48300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_519
timestamp 1644511149
transform 1 0 48852 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_531
timestamp 1644511149
transform 1 0 49956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_543
timestamp 1644511149
transform 1 0 51060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_555
timestamp 1644511149
transform 1 0 52164 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1644511149
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_561
timestamp 1644511149
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_573
timestamp 1644511149
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_585
timestamp 1644511149
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_597
timestamp 1644511149
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1644511149
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1644511149
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_617
timestamp 1644511149
transform 1 0 57868 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_621
timestamp 1644511149
transform 1 0 58236 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_19
timestamp 1644511149
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1644511149
transform 1 0 12604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 1644511149
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_144
timestamp 1644511149
transform 1 0 14352 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_150
timestamp 1644511149
transform 1 0 14904 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_156
timestamp 1644511149
transform 1 0 15456 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_162
timestamp 1644511149
transform 1 0 16008 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_168
timestamp 1644511149
transform 1 0 16560 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_174
timestamp 1644511149
transform 1 0 17112 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1644511149
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_186
timestamp 1644511149
transform 1 0 18216 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1644511149
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_201
timestamp 1644511149
transform 1 0 19596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_208
timestamp 1644511149
transform 1 0 20240 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_219
timestamp 1644511149
transform 1 0 21252 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_230
timestamp 1644511149
transform 1 0 22264 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1644511149
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_256
timestamp 1644511149
transform 1 0 24656 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_280
timestamp 1644511149
transform 1 0 26864 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1644511149
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_318
timestamp 1644511149
transform 1 0 30360 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_343
timestamp 1644511149
transform 1 0 32660 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_360
timestamp 1644511149
transform 1 0 34224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_385
timestamp 1644511149
transform 1 0 36524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_409
timestamp 1644511149
transform 1 0 38732 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_416
timestamp 1644511149
transform 1 0 39376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_427
timestamp 1644511149
transform 1 0 40388 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_437
timestamp 1644511149
transform 1 0 41308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_444
timestamp 1644511149
transform 1 0 41952 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_451
timestamp 1644511149
transform 1 0 42596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_458
timestamp 1644511149
transform 1 0 43240 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_464
timestamp 1644511149
transform 1 0 43792 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_470
timestamp 1644511149
transform 1 0 44344 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_479
timestamp 1644511149
transform 1 0 45172 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_485
timestamp 1644511149
transform 1 0 45724 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_491
timestamp 1644511149
transform 1 0 46276 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_497
timestamp 1644511149
transform 1 0 46828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_503
timestamp 1644511149
transform 1 0 47380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_509
timestamp 1644511149
transform 1 0 47932 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_521
timestamp 1644511149
transform 1 0 49036 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_529
timestamp 1644511149
transform 1 0 49772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_533
timestamp 1644511149
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_545
timestamp 1644511149
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_557
timestamp 1644511149
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_569
timestamp 1644511149
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1644511149
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1644511149
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_589
timestamp 1644511149
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_601
timestamp 1644511149
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_613
timestamp 1644511149
transform 1 0 57500 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_621
timestamp 1644511149
transform 1 0 58236 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_152
timestamp 1644511149
transform 1 0 15088 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_158
timestamp 1644511149
transform 1 0 15640 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_174
timestamp 1644511149
transform 1 0 17112 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_180
timestamp 1644511149
transform 1 0 17664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_186
timestamp 1644511149
transform 1 0 18216 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1644511149
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_198
timestamp 1644511149
transform 1 0 19320 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_212
timestamp 1644511149
transform 1 0 20608 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1644511149
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_228
timestamp 1644511149
transform 1 0 22080 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_239
timestamp 1644511149
transform 1 0 23092 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_252
timestamp 1644511149
transform 1 0 24288 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1644511149
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_301
timestamp 1644511149
transform 1 0 28796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_325
timestamp 1644511149
transform 1 0 31004 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_332
timestamp 1644511149
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_357
timestamp 1644511149
transform 1 0 33948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_381
timestamp 1644511149
transform 1 0 36156 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_388
timestamp 1644511149
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_406
timestamp 1644511149
transform 1 0 38456 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_419
timestamp 1644511149
transform 1 0 39652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_427
timestamp 1644511149
transform 1 0 40388 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_435
timestamp 1644511149
transform 1 0 41124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_442
timestamp 1644511149
transform 1 0 41768 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_452
timestamp 1644511149
transform 1 0 42688 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_459
timestamp 1644511149
transform 1 0 43332 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_465
timestamp 1644511149
transform 1 0 43884 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_471
timestamp 1644511149
transform 1 0 44436 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_477
timestamp 1644511149
transform 1 0 44988 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_483
timestamp 1644511149
transform 1 0 45540 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_489
timestamp 1644511149
transform 1 0 46092 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_495
timestamp 1644511149
transform 1 0 46644 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_517
timestamp 1644511149
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_529
timestamp 1644511149
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_541
timestamp 1644511149
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1644511149
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1644511149
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_561
timestamp 1644511149
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_573
timestamp 1644511149
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_585
timestamp 1644511149
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_597
timestamp 1644511149
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1644511149
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1644511149
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1644511149
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_157
timestamp 1644511149
transform 1 0 15548 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_160
timestamp 1644511149
transform 1 0 15824 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_166
timestamp 1644511149
transform 1 0 16376 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_172
timestamp 1644511149
transform 1 0 16928 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_178
timestamp 1644511149
transform 1 0 17480 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_184
timestamp 1644511149
transform 1 0 18032 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1644511149
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_200
timestamp 1644511149
transform 1 0 19504 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_206
timestamp 1644511149
transform 1 0 20056 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_212
timestamp 1644511149
transform 1 0 20608 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_219
timestamp 1644511149
transform 1 0 21252 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_226
timestamp 1644511149
transform 1 0 21896 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_237
timestamp 1644511149
transform 1 0 22908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1644511149
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_262
timestamp 1644511149
transform 1 0 25208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_280
timestamp 1644511149
transform 1 0 26864 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1644511149
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_317
timestamp 1644511149
transform 1 0 30268 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_341
timestamp 1644511149
transform 1 0 32476 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_359
timestamp 1644511149
transform 1 0 34132 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_385
timestamp 1644511149
transform 1 0 36524 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_409
timestamp 1644511149
transform 1 0 38732 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_416
timestamp 1644511149
transform 1 0 39376 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_425
timestamp 1644511149
transform 1 0 40204 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_440
timestamp 1644511149
transform 1 0 41584 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_447
timestamp 1644511149
transform 1 0 42228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_453
timestamp 1644511149
transform 1 0 42780 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_459
timestamp 1644511149
transform 1 0 43332 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_465
timestamp 1644511149
transform 1 0 43884 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_471
timestamp 1644511149
transform 1 0 44436 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_479
timestamp 1644511149
transform 1 0 45172 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_485
timestamp 1644511149
transform 1 0 45724 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_491
timestamp 1644511149
transform 1 0 46276 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_503
timestamp 1644511149
transform 1 0 47380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_515
timestamp 1644511149
transform 1 0 48484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_527
timestamp 1644511149
transform 1 0 49588 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1644511149
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_533
timestamp 1644511149
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_545
timestamp 1644511149
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_557
timestamp 1644511149
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_569
timestamp 1644511149
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1644511149
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1644511149
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_589
timestamp 1644511149
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_601
timestamp 1644511149
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_613
timestamp 1644511149
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_7
timestamp 1644511149
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_19
timestamp 1644511149
transform 1 0 2852 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_31
timestamp 1644511149
transform 1 0 3956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_43
timestamp 1644511149
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_175
timestamp 1644511149
transform 1 0 17204 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_187
timestamp 1644511149
transform 1 0 18308 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_199
timestamp 1644511149
transform 1 0 19412 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_202
timestamp 1644511149
transform 1 0 19688 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_208
timestamp 1644511149
transform 1 0 20240 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_214
timestamp 1644511149
transform 1 0 20792 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_232
timestamp 1644511149
transform 1 0 22448 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_258
timestamp 1644511149
transform 1 0 24840 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_284
timestamp 1644511149
transform 1 0 27232 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_308
timestamp 1644511149
transform 1 0 29440 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1644511149
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_357
timestamp 1644511149
transform 1 0 33948 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_381
timestamp 1644511149
transform 1 0 36156 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_388
timestamp 1644511149
transform 1 0 36800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_403
timestamp 1644511149
transform 1 0 38180 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_415
timestamp 1644511149
transform 1 0 39284 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_423
timestamp 1644511149
transform 1 0 40020 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_430
timestamp 1644511149
transform 1 0 40664 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_436
timestamp 1644511149
transform 1 0 41216 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_442
timestamp 1644511149
transform 1 0 41768 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_451
timestamp 1644511149
transform 1 0 42596 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_457
timestamp 1644511149
transform 1 0 43148 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_463
timestamp 1644511149
transform 1 0 43700 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_469
timestamp 1644511149
transform 1 0 44252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_475
timestamp 1644511149
transform 1 0 44804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_481
timestamp 1644511149
transform 1 0 45356 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_493
timestamp 1644511149
transform 1 0 46460 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_501
timestamp 1644511149
transform 1 0 47196 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_517
timestamp 1644511149
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_529
timestamp 1644511149
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_541
timestamp 1644511149
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1644511149
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1644511149
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_561
timestamp 1644511149
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_573
timestamp 1644511149
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_585
timestamp 1644511149
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_597
timestamp 1644511149
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1644511149
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1644511149
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_617
timestamp 1644511149
transform 1 0 57868 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_621
timestamp 1644511149
transform 1 0 58236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_180
timestamp 1644511149
transform 1 0 17664 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_186
timestamp 1644511149
transform 1 0 18216 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1644511149
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_200
timestamp 1644511149
transform 1 0 19504 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_206
timestamp 1644511149
transform 1 0 20056 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_212
timestamp 1644511149
transform 1 0 20608 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_218
timestamp 1644511149
transform 1 0 21160 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_224
timestamp 1644511149
transform 1 0 21712 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_231
timestamp 1644511149
transform 1 0 22356 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_240
timestamp 1644511149
transform 1 0 23184 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1644511149
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_256
timestamp 1644511149
transform 1 0 24656 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_267
timestamp 1644511149
transform 1 0 25668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_280
timestamp 1644511149
transform 1 0 26864 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1644511149
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_331
timestamp 1644511149
transform 1 0 31556 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_355
timestamp 1644511149
transform 1 0 33764 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_369
timestamp 1644511149
transform 1 0 35052 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_390
timestamp 1644511149
transform 1 0 36984 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_409
timestamp 1644511149
transform 1 0 38732 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1644511149
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_424
timestamp 1644511149
transform 1 0 40112 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_430
timestamp 1644511149
transform 1 0 40664 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_436
timestamp 1644511149
transform 1 0 41216 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_442
timestamp 1644511149
transform 1 0 41768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_448
timestamp 1644511149
transform 1 0 42320 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_454
timestamp 1644511149
transform 1 0 42872 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_460
timestamp 1644511149
transform 1 0 43424 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_466
timestamp 1644511149
transform 1 0 43976 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_472
timestamp 1644511149
transform 1 0 44528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_489
timestamp 1644511149
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_501
timestamp 1644511149
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_513
timestamp 1644511149
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1644511149
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1644511149
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_533
timestamp 1644511149
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_545
timestamp 1644511149
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_557
timestamp 1644511149
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_569
timestamp 1644511149
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1644511149
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1644511149
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_589
timestamp 1644511149
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_601
timestamp 1644511149
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_613
timestamp 1644511149
transform 1 0 57500 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_621
timestamp 1644511149
transform 1 0 58236 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_189
timestamp 1644511149
transform 1 0 18492 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_195
timestamp 1644511149
transform 1 0 19044 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_201
timestamp 1644511149
transform 1 0 19596 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_207
timestamp 1644511149
transform 1 0 20148 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_213
timestamp 1644511149
transform 1 0 20700 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1644511149
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_230
timestamp 1644511149
transform 1 0 22264 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_236
timestamp 1644511149
transform 1 0 22816 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_240
timestamp 1644511149
transform 1 0 23184 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_244
timestamp 1644511149
transform 1 0 23552 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_251
timestamp 1644511149
transform 1 0 24196 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_262
timestamp 1644511149
transform 1 0 25208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1644511149
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_287
timestamp 1644511149
transform 1 0 27508 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_357
timestamp 1644511149
transform 1 0 33948 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_378
timestamp 1644511149
transform 1 0 35880 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_382
timestamp 1644511149
transform 1 0 36248 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_388
timestamp 1644511149
transform 1 0 36800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_400
timestamp 1644511149
transform 1 0 37904 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_408
timestamp 1644511149
transform 1 0 38640 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_415
timestamp 1644511149
transform 1 0 39284 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_421
timestamp 1644511149
transform 1 0 39836 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_427
timestamp 1644511149
transform 1 0 40388 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_433
timestamp 1644511149
transform 1 0 40940 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_439
timestamp 1644511149
transform 1 0 41492 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_451
timestamp 1644511149
transform 1 0 42596 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_457
timestamp 1644511149
transform 1 0 43148 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_463
timestamp 1644511149
transform 1 0 43700 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_475
timestamp 1644511149
transform 1 0 44804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_487
timestamp 1644511149
transform 1 0 45908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_499
timestamp 1644511149
transform 1 0 47012 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_517
timestamp 1644511149
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_529
timestamp 1644511149
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_541
timestamp 1644511149
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1644511149
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1644511149
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_561
timestamp 1644511149
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_573
timestamp 1644511149
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_585
timestamp 1644511149
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_597
timestamp 1644511149
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1644511149
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1644511149
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_617
timestamp 1644511149
transform 1 0 57868 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_7
timestamp 1644511149
transform 1 0 1748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_13
timestamp 1644511149
transform 1 0 2300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_25
timestamp 1644511149
transform 1 0 3404 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_202
timestamp 1644511149
transform 1 0 19688 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_208
timestamp 1644511149
transform 1 0 20240 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_214
timestamp 1644511149
transform 1 0 20792 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_224
timestamp 1644511149
transform 1 0 21712 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_230
timestamp 1644511149
transform 1 0 22264 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_236
timestamp 1644511149
transform 1 0 22816 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_242
timestamp 1644511149
transform 1 0 23368 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_257
timestamp 1644511149
transform 1 0 24748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_276
timestamp 1644511149
transform 1 0 26496 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_287
timestamp 1644511149
transform 1 0 27508 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1644511149
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_313
timestamp 1644511149
transform 1 0 29900 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_334
timestamp 1644511149
transform 1 0 31832 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_358
timestamp 1644511149
transform 1 0 34040 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_372
timestamp 1644511149
transform 1 0 35328 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_387
timestamp 1644511149
transform 1 0 36708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_397
timestamp 1644511149
transform 1 0 37628 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_404
timestamp 1644511149
transform 1 0 38272 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_411
timestamp 1644511149
transform 1 0 38916 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_423
timestamp 1644511149
transform 1 0 40020 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_429
timestamp 1644511149
transform 1 0 40572 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_435
timestamp 1644511149
transform 1 0 41124 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_441
timestamp 1644511149
transform 1 0 41676 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_447
timestamp 1644511149
transform 1 0 42228 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_453
timestamp 1644511149
transform 1 0 42780 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_465
timestamp 1644511149
transform 1 0 43884 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_473
timestamp 1644511149
transform 1 0 44620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_513
timestamp 1644511149
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1644511149
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1644511149
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_533
timestamp 1644511149
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_545
timestamp 1644511149
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_557
timestamp 1644511149
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_569
timestamp 1644511149
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1644511149
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1644511149
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_589
timestamp 1644511149
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_601
timestamp 1644511149
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_613
timestamp 1644511149
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_208
timestamp 1644511149
transform 1 0 20240 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_214
timestamp 1644511149
transform 1 0 20792 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1644511149
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_228
timestamp 1644511149
transform 1 0 22080 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_234
timestamp 1644511149
transform 1 0 22632 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_259
timestamp 1644511149
transform 1 0 24932 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_268
timestamp 1644511149
transform 1 0 25760 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_291
timestamp 1644511149
transform 1 0 27876 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_302
timestamp 1644511149
transform 1 0 28888 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_310
timestamp 1644511149
transform 1 0 29624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_331
timestamp 1644511149
transform 1 0 31556 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_350
timestamp 1644511149
transform 1 0 33304 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_370
timestamp 1644511149
transform 1 0 35144 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_379
timestamp 1644511149
transform 1 0 35972 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_387
timestamp 1644511149
transform 1 0 36708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_396
timestamp 1644511149
transform 1 0 37536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_403
timestamp 1644511149
transform 1 0 38180 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_409
timestamp 1644511149
transform 1 0 38732 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_415
timestamp 1644511149
transform 1 0 39284 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_421
timestamp 1644511149
transform 1 0 39836 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_427
timestamp 1644511149
transform 1 0 40388 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_433
timestamp 1644511149
transform 1 0 40940 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_439
timestamp 1644511149
transform 1 0 41492 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_485
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_505
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_517
timestamp 1644511149
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_529
timestamp 1644511149
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_541
timestamp 1644511149
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1644511149
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1644511149
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_561
timestamp 1644511149
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_573
timestamp 1644511149
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_585
timestamp 1644511149
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_597
timestamp 1644511149
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1644511149
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1644511149
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_617
timestamp 1644511149
transform 1 0 57868 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_621
timestamp 1644511149
transform 1 0 58236 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_149
timestamp 1644511149
transform 1 0 14812 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_161
timestamp 1644511149
transform 1 0 15916 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_167
timestamp 1644511149
transform 1 0 16468 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_172
timestamp 1644511149
transform 1 0 16928 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_178
timestamp 1644511149
transform 1 0 17480 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_190
timestamp 1644511149
transform 1 0 18584 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_215
timestamp 1644511149
transform 1 0 20884 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_218
timestamp 1644511149
transform 1 0 21160 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_224
timestamp 1644511149
transform 1 0 21712 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_230
timestamp 1644511149
transform 1 0 22264 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_236
timestamp 1644511149
transform 1 0 22816 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_242
timestamp 1644511149
transform 1 0 23368 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1644511149
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_255
timestamp 1644511149
transform 1 0 24564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_261
timestamp 1644511149
transform 1 0 25116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_267
timestamp 1644511149
transform 1 0 25668 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_274
timestamp 1644511149
transform 1 0 26312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_282
timestamp 1644511149
transform 1 0 27048 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_293
timestamp 1644511149
transform 1 0 28060 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1644511149
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_316
timestamp 1644511149
transform 1 0 30176 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_340
timestamp 1644511149
transform 1 0 32384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_351
timestamp 1644511149
transform 1 0 33396 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1644511149
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_369
timestamp 1644511149
transform 1 0 35052 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_373
timestamp 1644511149
transform 1 0 35420 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_384
timestamp 1644511149
transform 1 0 36432 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_391
timestamp 1644511149
transform 1 0 37076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_398
timestamp 1644511149
transform 1 0 37720 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_404
timestamp 1644511149
transform 1 0 38272 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_410
timestamp 1644511149
transform 1 0 38824 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_416
timestamp 1644511149
transform 1 0 39376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_423
timestamp 1644511149
transform 1 0 40020 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_429
timestamp 1644511149
transform 1 0 40572 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_435
timestamp 1644511149
transform 1 0 41124 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_447
timestamp 1644511149
transform 1 0 42228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_459
timestamp 1644511149
transform 1 0 43332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_471
timestamp 1644511149
transform 1 0 44436 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_501
timestamp 1644511149
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_513
timestamp 1644511149
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1644511149
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1644511149
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_533
timestamp 1644511149
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_545
timestamp 1644511149
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_557
timestamp 1644511149
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_569
timestamp 1644511149
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1644511149
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1644511149
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_589
timestamp 1644511149
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_601
timestamp 1644511149
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_613
timestamp 1644511149
transform 1 0 57500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_621
timestamp 1644511149
transform 1 0 58236 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_7
timestamp 1644511149
transform 1 0 1748 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_19
timestamp 1644511149
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_31
timestamp 1644511149
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_43
timestamp 1644511149
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_116
timestamp 1644511149
transform 1 0 11776 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_128
timestamp 1644511149
transform 1 0 12880 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_140
timestamp 1644511149
transform 1 0 13984 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_152
timestamp 1644511149
transform 1 0 15088 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1644511149
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_230
timestamp 1644511149
transform 1 0 22264 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_236
timestamp 1644511149
transform 1 0 22816 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_242
timestamp 1644511149
transform 1 0 23368 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_252
timestamp 1644511149
transform 1 0 24288 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_258
timestamp 1644511149
transform 1 0 24840 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_264
timestamp 1644511149
transform 1 0 25392 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_270
timestamp 1644511149
transform 1 0 25944 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1644511149
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_287
timestamp 1644511149
transform 1 0 27508 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_296
timestamp 1644511149
transform 1 0 28336 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_307
timestamp 1644511149
transform 1 0 29348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_325
timestamp 1644511149
transform 1 0 31004 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_332
timestamp 1644511149
transform 1 0 31648 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_344
timestamp 1644511149
transform 1 0 32752 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_352
timestamp 1644511149
transform 1 0 33488 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_360
timestamp 1644511149
transform 1 0 34224 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_368
timestamp 1644511149
transform 1 0 34960 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_375
timestamp 1644511149
transform 1 0 35604 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_382
timestamp 1644511149
transform 1 0 36248 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_388
timestamp 1644511149
transform 1 0 36800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_395
timestamp 1644511149
transform 1 0 37444 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_401
timestamp 1644511149
transform 1 0 37996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_407
timestamp 1644511149
transform 1 0 38548 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_413
timestamp 1644511149
transform 1 0 39100 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_419
timestamp 1644511149
transform 1 0 39652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_425
timestamp 1644511149
transform 1 0 40204 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_431
timestamp 1644511149
transform 1 0 40756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_443
timestamp 1644511149
transform 1 0 41860 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1644511149
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_505
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_517
timestamp 1644511149
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_529
timestamp 1644511149
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_541
timestamp 1644511149
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1644511149
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1644511149
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_561
timestamp 1644511149
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_573
timestamp 1644511149
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_585
timestamp 1644511149
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_597
timestamp 1644511149
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1644511149
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1644511149
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_617
timestamp 1644511149
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_149
timestamp 1644511149
transform 1 0 14812 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_161
timestamp 1644511149
transform 1 0 15916 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_173
timestamp 1644511149
transform 1 0 17020 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_185
timestamp 1644511149
transform 1 0 18124 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_193
timestamp 1644511149
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_239
timestamp 1644511149
transform 1 0 23092 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_242
timestamp 1644511149
transform 1 0 23368 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_257
timestamp 1644511149
transform 1 0 24748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_260
timestamp 1644511149
transform 1 0 25024 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_266
timestamp 1644511149
transform 1 0 25576 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_272
timestamp 1644511149
transform 1 0 26128 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_280
timestamp 1644511149
transform 1 0 26864 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_286
timestamp 1644511149
transform 1 0 27416 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_293
timestamp 1644511149
transform 1 0 28060 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_302
timestamp 1644511149
transform 1 0 28888 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_314
timestamp 1644511149
transform 1 0 29992 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_325
timestamp 1644511149
transform 1 0 31004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_334
timestamp 1644511149
transform 1 0 31832 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_343
timestamp 1644511149
transform 1 0 32660 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_351
timestamp 1644511149
transform 1 0 33396 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_358
timestamp 1644511149
transform 1 0 34040 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_367
timestamp 1644511149
transform 1 0 34868 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_374
timestamp 1644511149
transform 1 0 35512 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_380
timestamp 1644511149
transform 1 0 36064 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_386
timestamp 1644511149
transform 1 0 36616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_392
timestamp 1644511149
transform 1 0 37168 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_398
timestamp 1644511149
transform 1 0 37720 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_404
timestamp 1644511149
transform 1 0 38272 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_410
timestamp 1644511149
transform 1 0 38824 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_416
timestamp 1644511149
transform 1 0 39376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_501
timestamp 1644511149
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_513
timestamp 1644511149
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1644511149
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1644511149
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_533
timestamp 1644511149
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_545
timestamp 1644511149
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_557
timestamp 1644511149
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_569
timestamp 1644511149
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1644511149
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1644511149
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_589
timestamp 1644511149
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_601
timestamp 1644511149
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_613
timestamp 1644511149
transform 1 0 57500 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_621
timestamp 1644511149
transform 1 0 58236 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_242
timestamp 1644511149
transform 1 0 23368 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_248
timestamp 1644511149
transform 1 0 23920 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_254
timestamp 1644511149
transform 1 0 24472 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_260
timestamp 1644511149
transform 1 0 25024 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_266
timestamp 1644511149
transform 1 0 25576 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1644511149
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_285
timestamp 1644511149
transform 1 0 27324 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_291
timestamp 1644511149
transform 1 0 27876 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_297
timestamp 1644511149
transform 1 0 28428 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_304
timestamp 1644511149
transform 1 0 29072 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_315
timestamp 1644511149
transform 1 0 30084 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_325
timestamp 1644511149
transform 1 0 31004 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1644511149
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_341
timestamp 1644511149
transform 1 0 32476 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_348
timestamp 1644511149
transform 1 0 33120 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_355
timestamp 1644511149
transform 1 0 33764 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_367
timestamp 1644511149
transform 1 0 34868 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_379
timestamp 1644511149
transform 1 0 35972 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_395
timestamp 1644511149
transform 1 0 37444 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_401
timestamp 1644511149
transform 1 0 37996 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_407
timestamp 1644511149
transform 1 0 38548 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_413
timestamp 1644511149
transform 1 0 39100 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_425
timestamp 1644511149
transform 1 0 40204 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_437
timestamp 1644511149
transform 1 0 41308 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_445
timestamp 1644511149
transform 1 0 42044 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_467
timestamp 1644511149
transform 1 0 44068 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_471
timestamp 1644511149
transform 1 0 44436 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_483
timestamp 1644511149
transform 1 0 45540 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_495
timestamp 1644511149
transform 1 0 46644 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_508
timestamp 1644511149
transform 1 0 47840 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_520
timestamp 1644511149
transform 1 0 48944 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_532
timestamp 1644511149
transform 1 0 50048 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_544
timestamp 1644511149
transform 1 0 51152 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_556
timestamp 1644511149
transform 1 0 52256 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_561
timestamp 1644511149
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_573
timestamp 1644511149
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_585
timestamp 1644511149
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_597
timestamp 1644511149
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1644511149
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1644511149
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_621
timestamp 1644511149
transform 1 0 58236 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_7
timestamp 1644511149
transform 1 0 1748 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_19
timestamp 1644511149
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_257
timestamp 1644511149
transform 1 0 24748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_263
timestamp 1644511149
transform 1 0 25300 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_267
timestamp 1644511149
transform 1 0 25668 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_270
timestamp 1644511149
transform 1 0 25944 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_276
timestamp 1644511149
transform 1 0 26496 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_282
timestamp 1644511149
transform 1 0 27048 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_286
timestamp 1644511149
transform 1 0 27416 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_297
timestamp 1644511149
transform 1 0 28428 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1644511149
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_313
timestamp 1644511149
transform 1 0 29900 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_329
timestamp 1644511149
transform 1 0 31372 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_336
timestamp 1644511149
transform 1 0 32016 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_343
timestamp 1644511149
transform 1 0 32660 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_350
timestamp 1644511149
transform 1 0 33304 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_356
timestamp 1644511149
transform 1 0 33856 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_367
timestamp 1644511149
transform 1 0 34868 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_373
timestamp 1644511149
transform 1 0 35420 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_379
timestamp 1644511149
transform 1 0 35972 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_385
timestamp 1644511149
transform 1 0 36524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_391
timestamp 1644511149
transform 1 0 37076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_397
timestamp 1644511149
transform 1 0 37628 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_403
timestamp 1644511149
transform 1 0 38180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_415
timestamp 1644511149
transform 1 0 39284 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1644511149
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1644511149
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_533
timestamp 1644511149
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_545
timestamp 1644511149
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_557
timestamp 1644511149
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_569
timestamp 1644511149
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1644511149
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1644511149
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_589
timestamp 1644511149
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_601
timestamp 1644511149
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_613
timestamp 1644511149
transform 1 0 57500 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_621
timestamp 1644511149
transform 1 0 58236 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_7
timestamp 1644511149
transform 1 0 1748 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_19
timestamp 1644511149
transform 1 0 2852 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_31
timestamp 1644511149
transform 1 0 3956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_43
timestamp 1644511149
transform 1 0 5060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_213
timestamp 1644511149
transform 1 0 20700 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_227
timestamp 1644511149
transform 1 0 21988 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_239
timestamp 1644511149
transform 1 0 23092 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_251
timestamp 1644511149
transform 1 0 24196 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_259
timestamp 1644511149
transform 1 0 24932 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_264
timestamp 1644511149
transform 1 0 25392 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_270
timestamp 1644511149
transform 1 0 25944 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1644511149
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_286
timestamp 1644511149
transform 1 0 27416 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_294
timestamp 1644511149
transform 1 0 28152 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_297
timestamp 1644511149
transform 1 0 28428 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_303
timestamp 1644511149
transform 1 0 28980 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_309
timestamp 1644511149
transform 1 0 29532 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_315
timestamp 1644511149
transform 1 0 30084 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_318
timestamp 1644511149
transform 1 0 30360 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_325
timestamp 1644511149
transform 1 0 31004 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1644511149
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_339
timestamp 1644511149
transform 1 0 32292 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_345
timestamp 1644511149
transform 1 0 32844 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_353
timestamp 1644511149
transform 1 0 33580 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_359
timestamp 1644511149
transform 1 0 34132 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_365
timestamp 1644511149
transform 1 0 34684 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_371
timestamp 1644511149
transform 1 0 35236 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_377
timestamp 1644511149
transform 1 0 35788 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_383
timestamp 1644511149
transform 1 0 36340 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_395
timestamp 1644511149
transform 1 0 37444 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_407
timestamp 1644511149
transform 1 0 38548 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_419
timestamp 1644511149
transform 1 0 39652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_431
timestamp 1644511149
transform 1 0 40756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_443
timestamp 1644511149
transform 1 0 41860 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_517
timestamp 1644511149
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_529
timestamp 1644511149
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_541
timestamp 1644511149
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1644511149
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1644511149
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_561
timestamp 1644511149
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_573
timestamp 1644511149
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_585
timestamp 1644511149
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_597
timestamp 1644511149
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_609
timestamp 1644511149
transform 1 0 57132 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_612
timestamp 1644511149
transform 1 0 57408 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_621
timestamp 1644511149
transform 1 0 58236 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_7
timestamp 1644511149
transform 1 0 1748 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_22
timestamp 1644511149
transform 1 0 3128 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_31
timestamp 1644511149
transform 1 0 3956 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_43
timestamp 1644511149
transform 1 0 5060 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_55
timestamp 1644511149
transform 1 0 6164 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_57
timestamp 1644511149
transform 1 0 6348 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_69
timestamp 1644511149
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1644511149
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_89
timestamp 1644511149
transform 1 0 9292 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_95
timestamp 1644511149
transform 1 0 9844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_107
timestamp 1644511149
transform 1 0 10948 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_111
timestamp 1644511149
transform 1 0 11316 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_113
timestamp 1644511149
transform 1 0 11500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_125
timestamp 1644511149
transform 1 0 12604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1644511149
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_144
timestamp 1644511149
transform 1 0 14352 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_150
timestamp 1644511149
transform 1 0 14904 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_162
timestamp 1644511149
transform 1 0 16008 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_169
timestamp 1644511149
transform 1 0 16652 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_181
timestamp 1644511149
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_193
timestamp 1644511149
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_201
timestamp 1644511149
transform 1 0 19596 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_208
timestamp 1644511149
transform 1 0 20240 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_214
timestamp 1644511149
transform 1 0 20792 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_222
timestamp 1644511149
transform 1 0 21528 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_225
timestamp 1644511149
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_237
timestamp 1644511149
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1644511149
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_259
timestamp 1644511149
transform 1 0 24932 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_267
timestamp 1644511149
transform 1 0 25668 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_270
timestamp 1644511149
transform 1 0 25944 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_276
timestamp 1644511149
transform 1 0 26496 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_281
timestamp 1644511149
transform 1 0 26956 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_285
timestamp 1644511149
transform 1 0 27324 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_288
timestamp 1644511149
transform 1 0 27600 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_294
timestamp 1644511149
transform 1 0 28152 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_300
timestamp 1644511149
transform 1 0 28704 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_313
timestamp 1644511149
transform 1 0 29900 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_318
timestamp 1644511149
transform 1 0 30360 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_326
timestamp 1644511149
transform 1 0 31096 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_329
timestamp 1644511149
transform 1 0 31372 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_335
timestamp 1644511149
transform 1 0 31924 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_337
timestamp 1644511149
transform 1 0 32108 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_342
timestamp 1644511149
transform 1 0 32568 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_348
timestamp 1644511149
transform 1 0 33120 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_354
timestamp 1644511149
transform 1 0 33672 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_360
timestamp 1644511149
transform 1 0 34224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_368
timestamp 1644511149
transform 1 0 34960 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_372
timestamp 1644511149
transform 1 0 35328 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_383
timestamp 1644511149
transform 1 0 36340 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_391
timestamp 1644511149
transform 1 0 37076 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_393
timestamp 1644511149
transform 1 0 37260 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_405
timestamp 1644511149
transform 1 0 38364 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_417
timestamp 1644511149
transform 1 0 39468 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_425
timestamp 1644511149
transform 1 0 40204 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_428
timestamp 1644511149
transform 1 0 40480 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_436
timestamp 1644511149
transform 1 0 41216 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_449
timestamp 1644511149
transform 1 0 42412 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_461
timestamp 1644511149
transform 1 0 43516 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_473
timestamp 1644511149
transform 1 0 44620 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_485
timestamp 1644511149
transform 1 0 45724 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_488
timestamp 1644511149
transform 1 0 46000 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_496
timestamp 1644511149
transform 1 0 46736 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_505
timestamp 1644511149
transform 1 0 47564 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_517
timestamp 1644511149
transform 1 0 48668 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_529
timestamp 1644511149
transform 1 0 49772 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_533
timestamp 1644511149
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_545
timestamp 1644511149
transform 1 0 51244 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_555
timestamp 1644511149
transform 1 0 52164 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_559
timestamp 1644511149
transform 1 0 52532 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_561
timestamp 1644511149
transform 1 0 52716 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_573
timestamp 1644511149
transform 1 0 53820 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_585
timestamp 1644511149
transform 1 0 54924 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_589
timestamp 1644511149
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_601
timestamp 1644511149
transform 1 0 56396 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_605
timestamp 1644511149
transform 1 0 56764 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_612
timestamp 1644511149
transform 1 0 57408 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_621
timestamp 1644511149
transform 1 0 58236 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1644511149
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1644511149
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1644511149
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1644511149
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1644511149
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1644511149
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 32016 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 37168 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 42320 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 47472 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 52624 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 57776 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _225__1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 31648 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _226__2
timestamp 1644511149
transform -1 0 24656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227__3
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228__4
timestamp 1644511149
transform -1 0 36800 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _229_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1644511149
transform -1 0 24656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _237_
timestamp 1644511149
transform -1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1644511149
transform -1 0 31648 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1644511149
transform -1 0 36800 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _243_
timestamp 1644511149
transform -1 0 25852 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1644511149
transform -1 0 41952 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1644511149
transform -1 0 36800 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23552 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1644511149
transform -1 0 39376 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1644511149
transform 1 0 19964 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1644511149
transform 1 0 16468 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1644511149
transform 1 0 16468 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1644511149
transform 1 0 19044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _255_
timestamp 1644511149
transform -1 0 43792 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _256_
timestamp 1644511149
transform -1 0 37352 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _257_
timestamp 1644511149
transform -1 0 39376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1644511149
transform -1 0 34132 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34408 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 42044 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 40388 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38272 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _263_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 34040 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1644511149
transform -1 0 40112 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _267_
timestamp 1644511149
transform 1 0 19044 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22264 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20056 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28244 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 24840 0 -1 21760
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_1  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _273_
timestamp 1644511149
transform -1 0 35144 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _274_
timestamp 1644511149
transform 1 0 23644 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21344 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_4  _276_
timestamp 1644511149
transform 1 0 29532 0 -1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _277_
timestamp 1644511149
transform 1 0 27324 0 -1 11968
box -38 -48 2062 592
use sky130_fd_sc_hd__clkinv_2  _278_
timestamp 1644511149
transform 1 0 20240 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_8  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23920 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__and2b_1  _280_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 39284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _281_
timestamp 1644511149
transform -1 0 21896 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _282_
timestamp 1644511149
transform -1 0 40388 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _283_
timestamp 1644511149
transform -1 0 29992 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _284_
timestamp 1644511149
transform -1 0 35788 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _285_
timestamp 1644511149
transform -1 0 41584 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _286_
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _287_
timestamp 1644511149
transform -1 0 41308 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _288_
timestamp 1644511149
transform -1 0 31832 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _289_
timestamp 1644511149
transform -1 0 37536 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _290_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 39192 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _291_
timestamp 1644511149
transform -1 0 42688 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _292_
timestamp 1644511149
transform 1 0 29900 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _293_
timestamp 1644511149
transform 1 0 30912 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _294_
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _295_
timestamp 1644511149
transform 1 0 30360 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _296_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 34224 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _297_
timestamp 1644511149
transform -1 0 35880 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _298_
timestamp 1644511149
transform -1 0 38456 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _299_
timestamp 1644511149
transform 1 0 21620 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _300_
timestamp 1644511149
transform 1 0 23552 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 34040 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _302_
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 29072 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _304_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _305_
timestamp 1644511149
transform -1 0 34316 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _306_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 36616 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1644511149
transform -1 0 40664 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28244 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _309_
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _310_
timestamp 1644511149
transform -1 0 30636 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 21344 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _312_
timestamp 1644511149
transform -1 0 29072 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _313_
timestamp 1644511149
transform -1 0 27508 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _316_
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _317_
timestamp 1644511149
transform -1 0 35696 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1644511149
transform 1 0 35512 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _319_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21896 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _320_
timestamp 1644511149
transform 1 0 26220 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _321_
timestamp 1644511149
transform 1 0 19964 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _322_
timestamp 1644511149
transform 1 0 27232 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _323_
timestamp 1644511149
transform 1 0 25024 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _324_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _325_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27876 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1644511149
transform -1 0 36708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _327_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38364 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _328_
timestamp 1644511149
transform 1 0 23276 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _329_
timestamp 1644511149
transform -1 0 31004 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _330_
timestamp 1644511149
transform 1 0 20976 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _331_
timestamp 1644511149
transform 1 0 22448 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _332_
timestamp 1644511149
transform -1 0 26864 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _333_
timestamp 1644511149
transform 1 0 28796 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _334_
timestamp 1644511149
transform 1 0 19044 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _335_
timestamp 1644511149
transform 1 0 39652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _336_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18768 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _337_
timestamp 1644511149
transform 1 0 25484 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _338_
timestamp 1644511149
transform -1 0 29348 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1644511149
transform -1 0 22448 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _340_
timestamp 1644511149
transform -1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _341_
timestamp 1644511149
transform 1 0 27232 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp 1644511149
transform 1 0 24196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _343_
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _344_
timestamp 1644511149
transform 1 0 24472 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _345_
timestamp 1644511149
transform 1 0 22264 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _346_
timestamp 1644511149
transform 1 0 40020 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _347_
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _348_
timestamp 1644511149
transform -1 0 36708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _349_
timestamp 1644511149
transform -1 0 37996 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _350_
timestamp 1644511149
transform 1 0 25944 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1644511149
transform -1 0 25116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _352_
timestamp 1644511149
transform -1 0 20608 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _353_
timestamp 1644511149
transform 1 0 20608 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _354_
timestamp 1644511149
transform 1 0 23368 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _355_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 24196 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _356_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29072 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _357_
timestamp 1644511149
transform -1 0 34224 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _358_
timestamp 1644511149
transform -1 0 40296 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _359_
timestamp 1644511149
transform 1 0 19688 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _360_
timestamp 1644511149
transform -1 0 41124 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _361_
timestamp 1644511149
transform 1 0 31096 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _362_
timestamp 1644511149
transform 1 0 41584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _363_
timestamp 1644511149
transform 1 0 17940 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _364_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 28060 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _365_
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _366_
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _367_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 35236 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _368_
timestamp 1644511149
transform 1 0 19596 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _369_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27876 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _370_
timestamp 1644511149
transform 1 0 25208 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _371_
timestamp 1644511149
transform -1 0 25300 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _372_
timestamp 1644511149
transform 1 0 20608 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _373_
timestamp 1644511149
transform 1 0 22632 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _374_
timestamp 1644511149
transform -1 0 43700 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _375_
timestamp 1644511149
transform -1 0 44344 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _376_
timestamp 1644511149
transform 1 0 30360 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _377_
timestamp 1644511149
transform -1 0 43884 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _378_
timestamp 1644511149
transform 1 0 27416 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _379_
timestamp 1644511149
transform -1 0 40664 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _380_
timestamp 1644511149
transform 1 0 20516 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _381_
timestamp 1644511149
transform -1 0 33304 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _382_
timestamp 1644511149
transform -1 0 40664 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _383_
timestamp 1644511149
transform 1 0 27876 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _384_
timestamp 1644511149
transform 1 0 18400 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _385_
timestamp 1644511149
transform 1 0 21988 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _386_
timestamp 1644511149
transform 1 0 35604 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _387_
timestamp 1644511149
transform -1 0 31924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _388_
timestamp 1644511149
transform 1 0 35972 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp 1644511149
transform -1 0 41768 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _390_
timestamp 1644511149
transform -1 0 26496 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _391_
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _392_
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _393_
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _394_
timestamp 1644511149
transform 1 0 33580 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _395_
timestamp 1644511149
transform -1 0 32752 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _396_
timestamp 1644511149
transform 1 0 20976 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _397_
timestamp 1644511149
transform 1 0 17848 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _398_
timestamp 1644511149
transform -1 0 44528 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _399_
timestamp 1644511149
transform -1 0 37536 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _400_
timestamp 1644511149
transform 1 0 18952 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _401_
timestamp 1644511149
transform 1 0 29256 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _402_
timestamp 1644511149
transform 1 0 20700 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _403_
timestamp 1644511149
transform 1 0 22908 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _404_
timestamp 1644511149
transform 1 0 18124 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _405_
timestamp 1644511149
transform -1 0 42780 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _406_
timestamp 1644511149
transform 1 0 33764 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _407_
timestamp 1644511149
transform 1 0 43332 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _408_
timestamp 1644511149
transform 1 0 16928 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _409_
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _410_
timestamp 1644511149
transform -1 0 43332 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _411_
timestamp 1644511149
transform 1 0 25852 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp 1644511149
transform 1 0 24748 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _413_
timestamp 1644511149
transform -1 0 17480 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _414_
timestamp 1644511149
transform 1 0 18032 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _415_
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _416_
timestamp 1644511149
transform 1 0 32752 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _417_
timestamp 1644511149
transform -1 0 25024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _418_
timestamp 1644511149
transform 1 0 26220 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 1644511149
transform -1 0 22540 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _420_
timestamp 1644511149
transform -1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _421_
timestamp 1644511149
transform 1 0 23644 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _422_
timestamp 1644511149
transform -1 0 23000 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _423_
timestamp 1644511149
transform 1 0 23552 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _424_
timestamp 1644511149
transform 1 0 17112 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _425_
timestamp 1644511149
transform 1 0 45632 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _426_
timestamp 1644511149
transform -1 0 35144 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _427_
timestamp 1644511149
transform -1 0 33488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _428_
timestamp 1644511149
transform -1 0 37904 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _429_
timestamp 1644511149
transform 1 0 23000 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1644511149
transform -1 0 38732 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _431_
timestamp 1644511149
transform -1 0 30636 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _432_
timestamp 1644511149
transform 1 0 20976 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _433_
timestamp 1644511149
transform 1 0 41032 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _434_
timestamp 1644511149
transform -1 0 23184 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _435_
timestamp 1644511149
transform -1 0 35972 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _436_
timestamp 1644511149
transform 1 0 30268 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _437_
timestamp 1644511149
transform -1 0 38640 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _438_
timestamp 1644511149
transform -1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _439_
timestamp 1644511149
transform 1 0 35604 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _440_
timestamp 1644511149
transform -1 0 44436 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _441_
timestamp 1644511149
transform 1 0 19320 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _442_
timestamp 1644511149
transform -1 0 36800 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _443_
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _444_
timestamp 1644511149
transform -1 0 45264 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _445_
timestamp 1644511149
transform 1 0 19688 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _446_
timestamp 1644511149
transform -1 0 37904 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _447_
timestamp 1644511149
transform 1 0 18584 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _448_
timestamp 1644511149
transform -1 0 41216 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _449_
timestamp 1644511149
transform 1 0 19412 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _450_
timestamp 1644511149
transform -1 0 39560 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _451_
timestamp 1644511149
transform -1 0 26496 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _452_
timestamp 1644511149
transform 1 0 33672 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _453_
timestamp 1644511149
transform -1 0 28060 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _454_
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _455_
timestamp 1644511149
transform -1 0 41584 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _456_
timestamp 1644511149
transform -1 0 39376 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _457_
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _458_
timestamp 1644511149
transform 1 0 24840 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _459_
timestamp 1644511149
transform 1 0 17112 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _460_
timestamp 1644511149
transform -1 0 25208 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _461_
timestamp 1644511149
transform -1 0 21252 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _462_
timestamp 1644511149
transform -1 0 41952 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _463_
timestamp 1644511149
transform -1 0 28888 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _464_
timestamp 1644511149
transform 1 0 22080 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _465_
timestamp 1644511149
transform 1 0 32200 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _466_
timestamp 1644511149
transform -1 0 30084 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _467_
timestamp 1644511149
transform -1 0 43056 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _468_
timestamp 1644511149
transform 1 0 39008 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 1644511149
transform -1 0 20608 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _470_
timestamp 1644511149
transform -1 0 21436 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _471_
timestamp 1644511149
transform -1 0 45356 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _472_
timestamp 1644511149
transform -1 0 20608 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _473_
timestamp 1644511149
transform -1 0 45356 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _474_
timestamp 1644511149
transform 1 0 19596 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _475_
timestamp 1644511149
transform -1 0 29900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _476_
timestamp 1644511149
transform -1 0 19596 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _477_
timestamp 1644511149
transform -1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _478_
timestamp 1644511149
transform 1 0 33120 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _479_
timestamp 1644511149
transform -1 0 44528 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _480_
timestamp 1644511149
transform 1 0 18400 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _481_
timestamp 1644511149
transform 1 0 31004 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _482_
timestamp 1644511149
transform 1 0 17480 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _483_
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _484_
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _485_
timestamp 1644511149
transform 1 0 43148 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _486_
timestamp 1644511149
transform 1 0 26036 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _487_
timestamp 1644511149
transform -1 0 16100 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _488_
timestamp 1644511149
transform -1 0 40756 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _489_
timestamp 1644511149
transform -1 0 41676 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _490_
timestamp 1644511149
transform -1 0 39284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _491_
timestamp 1644511149
transform 1 0 17756 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _492_
timestamp 1644511149
transform 1 0 18400 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _493_
timestamp 1644511149
transform 1 0 37720 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _494_
timestamp 1644511149
transform 1 0 15824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _495_
timestamp 1644511149
transform 1 0 31004 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _496_
timestamp 1644511149
transform -1 0 42688 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _497_
timestamp 1644511149
transform 1 0 32292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _498_
timestamp 1644511149
transform 1 0 42228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _499_
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _500_
timestamp 1644511149
transform 1 0 36156 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _501_
timestamp 1644511149
transform -1 0 42780 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _502_
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _503_
timestamp 1644511149
transform 1 0 33028 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _504_
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _505_
timestamp 1644511149
transform -1 0 42596 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _506_
timestamp 1644511149
transform -1 0 19964 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _507_
timestamp 1644511149
transform -1 0 28060 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _508_
timestamp 1644511149
transform 1 0 38640 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _509_
timestamp 1644511149
transform 1 0 37260 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _510_
timestamp 1644511149
transform 1 0 43700 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _511_
timestamp 1644511149
transform 1 0 33856 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _512_
timestamp 1644511149
transform 1 0 32384 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _513_
timestamp 1644511149
transform -1 0 38640 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _514_
timestamp 1644511149
transform -1 0 33120 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _515_
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _516__5
timestamp 1644511149
transform -1 0 31648 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _517_
timestamp 1644511149
transform -1 0 43792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _518__6
timestamp 1644511149
transform -1 0 23552 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _519_
timestamp 1644511149
transform -1 0 26312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _520_
timestamp 1644511149
transform 1 0 27324 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _521_
timestamp 1644511149
transform -1 0 38180 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _522_
timestamp 1644511149
transform -1 0 39928 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _523_
timestamp 1644511149
transform 1 0 26864 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _524_
timestamp 1644511149
transform -1 0 36432 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _525_
timestamp 1644511149
transform -1 0 27048 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _526_
timestamp 1644511149
transform -1 0 44160 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _527_
timestamp 1644511149
transform 1 0 15180 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _528_
timestamp 1644511149
transform -1 0 45080 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _529_
timestamp 1644511149
transform -1 0 41860 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _530_
timestamp 1644511149
transform -1 0 45172 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _531_
timestamp 1644511149
transform -1 0 46000 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _532_
timestamp 1644511149
transform 1 0 30728 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _533_
timestamp 1644511149
transform -1 0 31648 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _534_
timestamp 1644511149
transform -1 0 33304 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _535_
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _536_
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _537_
timestamp 1644511149
transform 1 0 40664 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _538_
timestamp 1644511149
transform -1 0 37352 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _539_
timestamp 1644511149
transform -1 0 29900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _540_
timestamp 1644511149
transform -1 0 36340 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _541_
timestamp 1644511149
transform -1 0 26496 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _542_
timestamp 1644511149
transform -1 0 46000 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _543_
timestamp 1644511149
transform -1 0 25484 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _544_
timestamp 1644511149
transform -1 0 31188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _545_
timestamp 1644511149
transform -1 0 46644 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _546_
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _547_
timestamp 1644511149
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _548_
timestamp 1644511149
transform 1 0 42780 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _549_
timestamp 1644511149
transform 1 0 32844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _550_
timestamp 1644511149
transform 1 0 33764 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _551_
timestamp 1644511149
transform -1 0 35328 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _552_
timestamp 1644511149
transform -1 0 35604 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _553_
timestamp 1644511149
transform -1 0 36248 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _554_
timestamp 1644511149
transform -1 0 35512 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _555_
timestamp 1644511149
transform -1 0 46644 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _556_
timestamp 1644511149
transform 1 0 18124 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _557_
timestamp 1644511149
transform 1 0 16836 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _558_
timestamp 1644511149
transform -1 0 38180 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _559__7
timestamp 1644511149
transform -1 0 43240 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _560_
timestamp 1644511149
transform 1 0 36800 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _561__8
timestamp 1644511149
transform 1 0 37444 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _562_
timestamp 1644511149
transform -1 0 42228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _563__9
timestamp 1644511149
transform -1 0 33764 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _564_
timestamp 1644511149
transform -1 0 43332 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _565__10
timestamp 1644511149
transform 1 0 43792 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _566_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 31280 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _567_
timestamp 1644511149
transform -1 0 31924 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _568_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _569_
timestamp 1644511149
transform 1 0 27232 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _570_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23920 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _571_
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _572_
timestamp 1644511149
transform -1 0 33948 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _573_
timestamp 1644511149
transform 1 0 29808 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _574_
timestamp 1644511149
transform -1 0 24932 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _575_
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _576_
timestamp 1644511149
transform -1 0 36248 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _577_
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _578_
timestamp 1644511149
transform 1 0 31004 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _579_
timestamp 1644511149
transform -1 0 31464 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _580_
timestamp 1644511149
transform 1 0 29808 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _581_
timestamp 1644511149
transform 1 0 27232 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _582_
timestamp 1644511149
transform -1 0 29348 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _583_
timestamp 1644511149
transform 1 0 27508 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _584_
timestamp 1644511149
transform 1 0 24932 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _585_
timestamp 1644511149
transform 1 0 24656 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _586_
timestamp 1644511149
transform -1 0 26772 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _587_
timestamp 1644511149
transform 1 0 29532 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _588_
timestamp 1644511149
transform -1 0 29072 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _589_
timestamp 1644511149
transform 1 0 24656 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _590_
timestamp 1644511149
transform 1 0 27232 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _591_
timestamp 1644511149
transform 1 0 25024 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _592_
timestamp 1644511149
transform 1 0 36984 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _593_
timestamp 1644511149
transform 1 0 29716 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _594_
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _595_
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _596_
timestamp 1644511149
transform -1 0 29072 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _597_
timestamp 1644511149
transform -1 0 26496 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _598_
timestamp 1644511149
transform 1 0 24656 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _599_
timestamp 1644511149
transform -1 0 26864 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29900 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _601_
timestamp 1644511149
transform -1 0 31372 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _602_
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _603_
timestamp 1644511149
transform -1 0 36524 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _604_
timestamp 1644511149
transform 1 0 25024 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _605_
timestamp 1644511149
transform 1 0 22448 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _606_
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _607_
timestamp 1644511149
transform 1 0 29716 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _608_
timestamp 1644511149
transform -1 0 36156 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _609_
timestamp 1644511149
transform 1 0 36984 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _610_
timestamp 1644511149
transform 1 0 34408 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _611_
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _612_
timestamp 1644511149
transform 1 0 29716 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _613_
timestamp 1644511149
transform 1 0 29716 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _614_
timestamp 1644511149
transform 1 0 27416 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _615_
timestamp 1644511149
transform 1 0 32016 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _616_
timestamp 1644511149
transform 1 0 29808 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _617_
timestamp 1644511149
transform -1 0 29072 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _618_
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _619_
timestamp 1644511149
transform 1 0 22080 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _620_
timestamp 1644511149
transform -1 0 39100 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _621_
timestamp 1644511149
transform 1 0 22080 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _622_
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _623_
timestamp 1644511149
transform 1 0 24656 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _624_
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _625_
timestamp 1644511149
transform 1 0 22448 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _626_
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _627_
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _628_
timestamp 1644511149
transform -1 0 33764 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _629_
timestamp 1644511149
transform -1 0 31832 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _630_
timestamp 1644511149
transform 1 0 27600 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _631_
timestamp 1644511149
transform 1 0 22448 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _632_
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _633_
timestamp 1644511149
transform 1 0 27324 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _634_
timestamp 1644511149
transform 1 0 27232 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _635_
timestamp 1644511149
transform 1 0 25024 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _636_
timestamp 1644511149
transform 1 0 29900 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _637_
timestamp 1644511149
transform 1 0 39560 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _638_
timestamp 1644511149
transform 1 0 31924 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _639_
timestamp 1644511149
transform -1 0 41676 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _640_
timestamp 1644511149
transform 1 0 29716 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _641_
timestamp 1644511149
transform 1 0 29716 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _642_
timestamp 1644511149
transform -1 0 41676 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _643_
timestamp 1644511149
transform 1 0 32016 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _644_
timestamp 1644511149
transform 1 0 27232 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _645_
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _646_
timestamp 1644511149
transform -1 0 33948 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _647_
timestamp 1644511149
transform 1 0 32200 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _648_
timestamp 1644511149
transform 1 0 24656 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _649_
timestamp 1644511149
transform 1 0 27048 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _650_
timestamp 1644511149
transform -1 0 26496 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _651_
timestamp 1644511149
transform -1 0 36524 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _652_
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _653_
timestamp 1644511149
transform -1 0 41308 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _654_
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _655_
timestamp 1644511149
transform 1 0 22080 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _656_
timestamp 1644511149
transform -1 0 34040 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _657_
timestamp 1644511149
transform -1 0 32384 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _658_
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _659_
timestamp 1644511149
transform -1 0 34960 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _660_
timestamp 1644511149
transform -1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _661_
timestamp 1644511149
transform -1 0 20240 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _662_
timestamp 1644511149
transform 1 0 20792 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _663_
timestamp 1644511149
transform -1 0 40112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _664_
timestamp 1644511149
transform 1 0 10396 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _665_
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _666_
timestamp 1644511149
transform 1 0 12144 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _667_
timestamp 1644511149
transform 1 0 11316 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _668_
timestamp 1644511149
transform 1 0 10580 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _669_
timestamp 1644511149
transform 1 0 11224 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _670_
timestamp 1644511149
transform 1 0 13064 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _671_
timestamp 1644511149
transform 1 0 13156 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _672_
timestamp 1644511149
transform 1 0 12052 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _673_
timestamp 1644511149
transform -1 0 12604 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _674_
timestamp 1644511149
transform -1 0 29900 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _675_
timestamp 1644511149
transform -1 0 16928 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _676_
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _677_
timestamp 1644511149
transform -1 0 44436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _678_
timestamp 1644511149
transform -1 0 14812 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _679_
timestamp 1644511149
transform -1 0 47840 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _680_
timestamp 1644511149
transform -1 0 14812 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _681_
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _682_
timestamp 1644511149
transform 1 0 37628 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _683_
timestamp 1644511149
transform -1 0 14812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__075_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__219_
timestamp 1644511149
transform -1 0 36984 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_master
timestamp 1644511149
transform -1 0 30268 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__075_
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__219_
timestamp 1644511149
transform -1 0 34960 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_clk_master
timestamp 1644511149
transform -1 0 25760 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__075_
timestamp 1644511149
transform -1 0 41124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__219_
timestamp 1644511149
transform 1 0 40572 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_clk_master
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 34132 0 1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn
timestamp 1644511149
transform 1 0 27876 0 -1 22848
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
timestamp 1644511149
transform -1 0 34040 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn
timestamp 1644511149
transform 1 0 25576 0 1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
timestamp 1644511149
transform 1 0 32200 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn
timestamp 1644511149
transform 1 0 23000 0 -1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
timestamp 1644511149
transform 1 0 34408 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn
timestamp 1644511149
transform 1 0 20424 0 1 17408
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
timestamp 1644511149
transform 1 0 32292 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn
timestamp 1644511149
transform 1 0 25208 0 -1 21760
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
timestamp 1644511149
transform 1 0 30820 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn
timestamp 1644511149
transform 1 0 22632 0 1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
timestamp 1644511149
transform -1 0 32660 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn
timestamp 1644511149
transform -1 0 21344 0 -1 17408
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
timestamp 1644511149
transform -1 0 34040 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn
timestamp 1644511149
transform 1 0 20056 0 -1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
timestamp 1644511149
transform -1 0 31648 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn
timestamp 1644511149
transform 1 0 29716 0 -1 25024
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
timestamp 1644511149
transform -1 0 29072 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
timestamp 1644511149
transform -1 0 29072 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
timestamp 1644511149
transform -1 0 36616 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn
timestamp 1644511149
transform 1 0 36340 0 1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
timestamp 1644511149
transform 1 0 34408 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
timestamp 1644511149
transform -1 0 36340 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn
timestamp 1644511149
transform 1 0 38916 0 -1 15232
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
timestamp 1644511149
transform 1 0 29716 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn
timestamp 1644511149
transform -1 0 41124 0 1 15232
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
timestamp 1644511149
transform -1 0 29348 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn
timestamp 1644511149
transform 1 0 31924 0 1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
timestamp 1644511149
transform -1 0 29164 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_6  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 58236 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform -1 0 14352 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform -1 0 30268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 58236 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input5
timestamp 1644511149
transform -1 0 58236 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  input6
timestamp 1644511149
transform -1 0 58236 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input7
timestamp 1644511149
transform -1 0 58236 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input8
timestamp 1644511149
transform -1 0 58236 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input9
timestamp 1644511149
transform -1 0 58236 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input10
timestamp 1644511149
transform -1 0 58236 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input11
timestamp 1644511149
transform -1 0 58236 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input12
timestamp 1644511149
transform -1 0 58236 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input13
timestamp 1644511149
transform -1 0 58236 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1644511149
transform -1 0 58236 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1644511149
transform -1 0 58236 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 57408 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1644511149
transform 1 0 40848 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1644511149
transform 1 0 46368 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  input19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 57408 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  input20
timestamp 1644511149
transform -1 0 58236 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1644511149
transform -1 0 30360 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1644511149
transform 1 0 35420 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output23
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1644511149
transform -1 0 3128 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1644511149
transform 1 0 24564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1644511149
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1644511149
transform -1 0 9292 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1644511149
transform -1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1644511149
transform -1 0 19596 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1644511149
transform -1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1644511149
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1644511149
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1644511149
transform -1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1644511149
transform -1 0 1748 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1644511149
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1644511149
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1644511149
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1644511149
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1644511149
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1644511149
transform -1 0 1748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1644511149
transform -1 0 1748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1644511149
transform -1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1644511149
transform 1 0 51796 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1644511149
transform -1 0 1748 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1644511149
transform 1 0 57868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1644511149
transform -1 0 1748 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1644511149
transform -1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1644511149
transform -1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1644511149
transform 1 0 54004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1644511149
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  ro_block_I.ro_pol.tribuf.t_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35880 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  ro_block_I.ro_pol_eve.tribuf.t_buf
timestamp 1644511149
transform -1 0 24288 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  ro_block_Q.ro_pol.tribuf.t_buf
timestamp 1644511149
transform 1 0 38824 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  ro_block_Q.ro_pol_eve.tribuf.t_buf
timestamp 1644511149
transform -1 0 26404 0 -1 22848
box -38 -48 866 592
<< labels >>
rlabel metal2 s 29918 29200 29974 30000 6 cclk_I
port 0 nsew signal tristate
rlabel metal2 s 35346 29200 35402 30000 6 cclk_Q
port 1 nsew signal tristate
rlabel metal3 s 59200 2592 60000 2712 6 clk_master
port 2 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 clk_master_out
port 3 nsew signal tristate
rlabel metal3 s 59200 4360 60000 4480 6 clkdiv2
port 4 nsew signal input
rlabel metal2 s 13542 29200 13598 30000 6 comp_high_I
port 5 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 comp_high_Q
port 6 nsew signal input
rlabel metal2 s 2686 29200 2742 30000 6 cos_out
port 7 nsew signal tristate
rlabel metal2 s 24490 29200 24546 30000 6 cos_outb
port 8 nsew signal tristate
rlabel metal3 s 0 3816 800 3936 6 div2out
port 9 nsew signal tristate
rlabel metal2 s 8114 29200 8170 30000 6 fb1_I
port 10 nsew signal tristate
rlabel metal2 s 17958 0 18014 800 6 fb1_Q
port 11 nsew signal tristate
rlabel metal2 s 18970 29200 19026 30000 6 fb2_I
port 12 nsew signal tristate
rlabel metal2 s 41970 0 42026 800 6 fb2_Q
port 13 nsew signal tristate
rlabel metal3 s 59200 7896 60000 8016 6 gray_clk_in[0]
port 14 nsew signal input
rlabel metal3 s 59200 9664 60000 9784 6 gray_clk_in[1]
port 15 nsew signal input
rlabel metal3 s 59200 11432 60000 11552 6 gray_clk_in[2]
port 16 nsew signal input
rlabel metal3 s 59200 13200 60000 13320 6 gray_clk_in[3]
port 17 nsew signal input
rlabel metal3 s 59200 14968 60000 15088 6 gray_clk_in[4]
port 18 nsew signal input
rlabel metal3 s 59200 16736 60000 16856 6 gray_clk_in[5]
port 19 nsew signal input
rlabel metal3 s 59200 18504 60000 18624 6 gray_clk_in[6]
port 20 nsew signal input
rlabel metal3 s 59200 20272 60000 20392 6 gray_clk_in[7]
port 21 nsew signal input
rlabel metal3 s 59200 22040 60000 22160 6 gray_clk_in[8]
port 22 nsew signal input
rlabel metal3 s 59200 23808 60000 23928 6 gray_clk_in[9]
port 23 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 gray_clk_out[10]
port 24 nsew signal tristate
rlabel metal3 s 0 6944 800 7064 6 gray_clk_out[1]
port 25 nsew signal tristate
rlabel metal3 s 0 8576 800 8696 6 gray_clk_out[2]
port 26 nsew signal tristate
rlabel metal3 s 0 10072 800 10192 6 gray_clk_out[3]
port 27 nsew signal tristate
rlabel metal3 s 0 11704 800 11824 6 gray_clk_out[4]
port 28 nsew signal tristate
rlabel metal3 s 0 13336 800 13456 6 gray_clk_out[5]
port 29 nsew signal tristate
rlabel metal3 s 0 14832 800 14952 6 gray_clk_out[6]
port 30 nsew signal tristate
rlabel metal3 s 0 16464 800 16584 6 gray_clk_out[7]
port 31 nsew signal tristate
rlabel metal3 s 0 17960 800 18080 6 gray_clk_out[8]
port 32 nsew signal tristate
rlabel metal3 s 0 19592 800 19712 6 gray_clk_out[9]
port 33 nsew signal tristate
rlabel metal3 s 59200 25576 60000 25696 6 no_ones_below_in[0]
port 34 nsew signal input
rlabel metal3 s 59200 27344 60000 27464 6 no_ones_below_in[1]
port 35 nsew signal input
rlabel metal3 s 59200 29112 60000 29232 6 no_ones_below_in[2]
port 36 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 no_ones_below_out[0]
port 37 nsew signal tristate
rlabel metal3 s 0 24352 800 24472 6 no_ones_below_out[1]
port 38 nsew signal tristate
rlabel metal3 s 0 25984 800 26104 6 no_ones_below_out[2]
port 39 nsew signal tristate
rlabel metal2 s 40774 29200 40830 30000 6 phi1b_dig_I
port 40 nsew signal input
rlabel metal2 s 46294 29200 46350 30000 6 phi1b_dig_Q
port 41 nsew signal input
rlabel metal2 s 51722 29200 51778 30000 6 read_out_I[0]
port 42 nsew signal tristate
rlabel metal3 s 0 27480 800 27600 6 read_out_I[1]
port 43 nsew signal tristate
rlabel metal2 s 57150 29200 57206 30000 6 read_out_Q[0]
port 44 nsew signal tristate
rlabel metal3 s 0 29112 800 29232 6 read_out_Q[1]
port 45 nsew signal tristate
rlabel metal3 s 59200 824 60000 944 6 rstb
port 46 nsew signal input
rlabel metal3 s 0 688 800 808 6 rstb_out
port 47 nsew signal tristate
rlabel metal2 s 5998 0 6054 800 6 sin_out
port 48 nsew signal tristate
rlabel metal2 s 53930 0 53986 800 6 sin_outb
port 49 nsew signal tristate
rlabel metal3 s 59200 6128 60000 6248 6 ud_en
port 50 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 ud_en_out
port 51 nsew signal tristate
rlabel metal4 s 10576 2128 10896 27792 6 vccd1
port 52 nsew power input
rlabel metal4 s 29840 2128 30160 27792 6 vccd1
port 52 nsew power input
rlabel metal4 s 49104 2128 49424 27792 6 vccd1
port 52 nsew power input
rlabel metal4 s 20208 2128 20528 27792 6 vssd1
port 53 nsew ground input
rlabel metal4 s 39472 2128 39792 27792 6 vssd1
port 53 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 60000 30000
<< end >>
