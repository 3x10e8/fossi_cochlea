magic
tech sky130A
magscale 1 2
timestamp 1654387106
<< nwell >>
rect 1715 1373 2125 1605
<< nmos >>
rect 711 1130 741 1250
rect 797 1130 827 1250
rect 884 1130 914 1250
rect 970 1130 1000 1250
rect 1057 1130 1087 1250
rect 1143 1130 1173 1250
rect 1230 1130 1260 1250
rect 1316 1130 1346 1250
rect 1403 1130 1433 1250
rect 1489 1130 1519 1250
rect 1576 1130 1606 1250
rect 1662 1130 1692 1250
rect 1749 1130 1779 1250
rect 1835 1130 1865 1250
rect 1922 1130 1952 1250
rect 2008 1130 2038 1250
rect 2095 1130 2125 1250
rect 2181 1130 2211 1250
rect 2268 1130 2298 1250
rect 2354 1130 2384 1250
rect 2441 1130 2471 1250
rect 2527 1130 2557 1250
rect 2614 1130 2644 1250
rect 2700 1130 2730 1250
rect 2787 1130 2817 1250
rect 2873 1130 2903 1250
rect 2960 1130 2990 1250
rect 3046 1130 3076 1250
rect 711 690 741 810
rect 797 690 827 810
rect 884 690 914 810
rect 970 690 1000 810
rect 1057 690 1087 810
rect 1143 690 1173 810
rect 1230 690 1260 810
rect 1316 690 1346 810
rect 1403 690 1433 810
rect 1489 690 1519 810
rect 1576 690 1606 810
rect 1662 690 1692 810
rect 1749 690 1779 810
rect 1835 690 1865 810
rect 1922 690 1952 810
rect 2008 690 2038 810
rect 2095 690 2125 810
rect 2181 690 2211 810
rect 2268 690 2298 810
rect 2354 690 2384 810
rect 2441 690 2471 810
rect 2527 690 2557 810
rect 2614 690 2644 810
rect 2700 690 2730 810
rect 2787 690 2817 810
rect 2873 690 2903 810
rect 2960 690 2990 810
rect 3046 690 3076 810
<< pmos >>
rect 1829 1445 1859 1529
rect 1930 1445 1960 1529
<< ndiff >>
rect 654 1238 711 1250
rect 654 1204 666 1238
rect 700 1204 711 1238
rect 654 1130 711 1204
rect 741 1176 797 1250
rect 741 1142 752 1176
rect 786 1142 797 1176
rect 741 1130 797 1142
rect 827 1238 884 1250
rect 827 1204 839 1238
rect 873 1204 884 1238
rect 827 1130 884 1204
rect 914 1176 970 1250
rect 914 1142 925 1176
rect 959 1142 970 1176
rect 914 1130 970 1142
rect 1000 1238 1057 1250
rect 1000 1204 1012 1238
rect 1046 1204 1057 1238
rect 1000 1130 1057 1204
rect 1087 1176 1143 1250
rect 1087 1142 1098 1176
rect 1132 1142 1143 1176
rect 1087 1130 1143 1142
rect 1173 1238 1230 1250
rect 1173 1204 1185 1238
rect 1219 1204 1230 1238
rect 1173 1130 1230 1204
rect 1260 1176 1316 1250
rect 1260 1142 1271 1176
rect 1305 1142 1316 1176
rect 1260 1130 1316 1142
rect 1346 1238 1403 1250
rect 1346 1204 1358 1238
rect 1392 1204 1403 1238
rect 1346 1130 1403 1204
rect 1433 1176 1489 1250
rect 1433 1142 1444 1176
rect 1478 1142 1489 1176
rect 1433 1130 1489 1142
rect 1519 1238 1576 1250
rect 1519 1204 1531 1238
rect 1565 1204 1576 1238
rect 1519 1130 1576 1204
rect 1606 1176 1662 1250
rect 1606 1142 1617 1176
rect 1651 1142 1662 1176
rect 1606 1130 1662 1142
rect 1692 1238 1749 1250
rect 1692 1204 1704 1238
rect 1738 1204 1749 1238
rect 1692 1130 1749 1204
rect 1779 1176 1835 1250
rect 1779 1142 1790 1176
rect 1824 1142 1835 1176
rect 1779 1130 1835 1142
rect 1865 1238 1922 1250
rect 1865 1204 1877 1238
rect 1911 1204 1922 1238
rect 1865 1130 1922 1204
rect 1952 1176 2008 1250
rect 1952 1142 1963 1176
rect 1997 1142 2008 1176
rect 1952 1130 2008 1142
rect 2038 1238 2095 1250
rect 2038 1204 2050 1238
rect 2084 1204 2095 1238
rect 2038 1130 2095 1204
rect 2125 1176 2181 1250
rect 2125 1142 2136 1176
rect 2170 1142 2181 1176
rect 2125 1130 2181 1142
rect 2211 1238 2268 1250
rect 2211 1204 2223 1238
rect 2257 1204 2268 1238
rect 2211 1130 2268 1204
rect 2298 1176 2354 1250
rect 2298 1142 2309 1176
rect 2343 1142 2354 1176
rect 2298 1130 2354 1142
rect 2384 1238 2441 1250
rect 2384 1204 2396 1238
rect 2430 1204 2441 1238
rect 2384 1130 2441 1204
rect 2471 1176 2527 1250
rect 2471 1142 2482 1176
rect 2516 1142 2527 1176
rect 2471 1130 2527 1142
rect 2557 1238 2614 1250
rect 2557 1204 2569 1238
rect 2603 1204 2614 1238
rect 2557 1130 2614 1204
rect 2644 1176 2700 1250
rect 2644 1142 2655 1176
rect 2689 1142 2700 1176
rect 2644 1130 2700 1142
rect 2730 1238 2787 1250
rect 2730 1204 2742 1238
rect 2776 1204 2787 1238
rect 2730 1130 2787 1204
rect 2817 1176 2873 1250
rect 2817 1142 2828 1176
rect 2862 1142 2873 1176
rect 2817 1130 2873 1142
rect 2903 1238 2960 1250
rect 2903 1204 2915 1238
rect 2949 1204 2960 1238
rect 2903 1130 2960 1204
rect 2990 1176 3046 1250
rect 2990 1142 3001 1176
rect 3035 1142 3046 1176
rect 2990 1130 3046 1142
rect 3076 1238 3133 1250
rect 3076 1204 3088 1238
rect 3122 1204 3133 1238
rect 3076 1130 3133 1204
rect 651 798 711 810
rect 651 764 666 798
rect 700 764 711 798
rect 651 690 711 764
rect 741 736 797 810
rect 741 702 752 736
rect 786 702 797 736
rect 741 690 797 702
rect 827 798 884 810
rect 827 764 839 798
rect 873 764 884 798
rect 827 690 884 764
rect 914 736 970 810
rect 914 702 925 736
rect 959 702 970 736
rect 914 690 970 702
rect 1000 798 1057 810
rect 1000 764 1012 798
rect 1046 764 1057 798
rect 1000 690 1057 764
rect 1087 736 1143 810
rect 1087 702 1098 736
rect 1132 702 1143 736
rect 1087 690 1143 702
rect 1173 798 1230 810
rect 1173 764 1185 798
rect 1219 764 1230 798
rect 1173 690 1230 764
rect 1260 736 1316 810
rect 1260 702 1271 736
rect 1305 702 1316 736
rect 1260 690 1316 702
rect 1346 798 1403 810
rect 1346 764 1358 798
rect 1392 764 1403 798
rect 1346 690 1403 764
rect 1433 736 1489 810
rect 1433 702 1444 736
rect 1478 702 1489 736
rect 1433 690 1489 702
rect 1519 798 1576 810
rect 1519 764 1531 798
rect 1565 764 1576 798
rect 1519 690 1576 764
rect 1606 736 1662 810
rect 1606 702 1617 736
rect 1651 702 1662 736
rect 1606 690 1662 702
rect 1692 798 1749 810
rect 1692 764 1704 798
rect 1738 764 1749 798
rect 1692 690 1749 764
rect 1779 736 1835 810
rect 1779 702 1790 736
rect 1824 702 1835 736
rect 1779 690 1835 702
rect 1865 798 1922 810
rect 1865 764 1877 798
rect 1911 764 1922 798
rect 1865 690 1922 764
rect 1952 736 2008 810
rect 1952 702 1963 736
rect 1997 702 2008 736
rect 1952 690 2008 702
rect 2038 798 2095 810
rect 2038 764 2050 798
rect 2084 764 2095 798
rect 2038 690 2095 764
rect 2125 736 2181 810
rect 2125 702 2136 736
rect 2170 702 2181 736
rect 2125 690 2181 702
rect 2211 798 2268 810
rect 2211 764 2223 798
rect 2257 764 2268 798
rect 2211 690 2268 764
rect 2298 736 2354 810
rect 2298 702 2309 736
rect 2343 702 2354 736
rect 2298 690 2354 702
rect 2384 798 2441 810
rect 2384 764 2396 798
rect 2430 764 2441 798
rect 2384 690 2441 764
rect 2471 736 2527 810
rect 2471 702 2482 736
rect 2516 702 2527 736
rect 2471 690 2527 702
rect 2557 798 2614 810
rect 2557 764 2569 798
rect 2603 764 2614 798
rect 2557 690 2614 764
rect 2644 736 2700 810
rect 2644 702 2655 736
rect 2689 702 2700 736
rect 2644 690 2700 702
rect 2730 798 2787 810
rect 2730 764 2742 798
rect 2776 764 2787 798
rect 2730 690 2787 764
rect 2817 736 2873 810
rect 2817 702 2828 736
rect 2862 702 2873 736
rect 2817 690 2873 702
rect 2903 798 2960 810
rect 2903 764 2915 798
rect 2949 764 2960 798
rect 2903 690 2960 764
rect 2990 736 3046 810
rect 2990 702 3001 736
rect 3035 702 3046 736
rect 2990 690 3046 702
rect 3076 798 3137 810
rect 3076 764 3088 798
rect 3122 764 3137 798
rect 3076 690 3137 764
<< pdiff >>
rect 1763 1505 1829 1529
rect 1763 1471 1783 1505
rect 1817 1471 1829 1505
rect 1763 1445 1829 1471
rect 1859 1505 1930 1529
rect 1859 1471 1877 1505
rect 1911 1471 1930 1505
rect 1859 1445 1930 1471
rect 1960 1505 2020 1529
rect 1960 1471 1975 1505
rect 2009 1471 2020 1505
rect 1960 1445 2020 1471
<< ndiffc >>
rect 666 1204 700 1238
rect 752 1142 786 1176
rect 839 1204 873 1238
rect 925 1142 959 1176
rect 1012 1204 1046 1238
rect 1098 1142 1132 1176
rect 1185 1204 1219 1238
rect 1271 1142 1305 1176
rect 1358 1204 1392 1238
rect 1444 1142 1478 1176
rect 1531 1204 1565 1238
rect 1617 1142 1651 1176
rect 1704 1204 1738 1238
rect 1790 1142 1824 1176
rect 1877 1204 1911 1238
rect 1963 1142 1997 1176
rect 2050 1204 2084 1238
rect 2136 1142 2170 1176
rect 2223 1204 2257 1238
rect 2309 1142 2343 1176
rect 2396 1204 2430 1238
rect 2482 1142 2516 1176
rect 2569 1204 2603 1238
rect 2655 1142 2689 1176
rect 2742 1204 2776 1238
rect 2828 1142 2862 1176
rect 2915 1204 2949 1238
rect 3001 1142 3035 1176
rect 3088 1204 3122 1238
rect 666 764 700 798
rect 752 702 786 736
rect 839 764 873 798
rect 925 702 959 736
rect 1012 764 1046 798
rect 1098 702 1132 736
rect 1185 764 1219 798
rect 1271 702 1305 736
rect 1358 764 1392 798
rect 1444 702 1478 736
rect 1531 764 1565 798
rect 1617 702 1651 736
rect 1704 764 1738 798
rect 1790 702 1824 736
rect 1877 764 1911 798
rect 1963 702 1997 736
rect 2050 764 2084 798
rect 2136 702 2170 736
rect 2223 764 2257 798
rect 2309 702 2343 736
rect 2396 764 2430 798
rect 2482 702 2516 736
rect 2569 764 2603 798
rect 2655 702 2689 736
rect 2742 764 2776 798
rect 2828 702 2862 736
rect 2915 764 2949 798
rect 3001 702 3035 736
rect 3088 764 3122 798
<< pdiffc >>
rect 1783 1471 1817 1505
rect 1877 1471 1911 1505
rect 1975 1471 2009 1505
<< psubdiff >>
rect 593 777 651 810
rect 593 743 594 777
rect 628 743 651 777
rect 593 690 651 743
rect 3137 783 3210 810
rect 3137 749 3166 783
rect 3200 749 3210 783
rect 3137 690 3210 749
<< nsubdiff >>
rect 2020 1505 2089 1529
rect 2020 1471 2043 1505
rect 2077 1471 2089 1505
rect 2020 1445 2089 1471
<< psubdiffcont >>
rect 594 743 628 777
rect 3166 749 3200 783
<< nsubdiffcont >>
rect 2043 1471 2077 1505
<< poly >>
rect 1817 1610 1871 1620
rect 1811 1576 1827 1610
rect 1861 1576 1877 1610
rect 1817 1566 1871 1576
rect 1829 1529 1859 1566
rect 1930 1529 1960 1555
rect 1829 1419 1859 1445
rect 1930 1408 1960 1445
rect 1918 1398 1972 1408
rect 1912 1364 1928 1398
rect 1962 1364 1978 1398
rect 1918 1354 1972 1364
rect 711 1276 1865 1306
rect 711 1250 741 1276
rect 797 1250 827 1276
rect 884 1250 914 1276
rect 970 1250 1000 1276
rect 1057 1250 1087 1276
rect 1143 1250 1173 1276
rect 1230 1250 1260 1276
rect 1316 1250 1346 1276
rect 1403 1250 1433 1276
rect 1489 1250 1519 1276
rect 1576 1250 1606 1276
rect 1662 1250 1692 1276
rect 1749 1250 1779 1276
rect 1835 1250 1865 1276
rect 1922 1276 3076 1306
rect 1922 1250 1952 1276
rect 2008 1250 2038 1276
rect 2095 1250 2125 1276
rect 2181 1250 2211 1276
rect 2268 1250 2298 1276
rect 2354 1250 2384 1276
rect 2441 1250 2471 1276
rect 2527 1250 2557 1276
rect 2614 1250 2644 1276
rect 2700 1250 2730 1276
rect 2787 1250 2817 1276
rect 2873 1250 2903 1276
rect 2960 1250 2990 1276
rect 3046 1250 3076 1276
rect 711 1104 741 1130
rect 797 1104 827 1130
rect 884 1104 914 1130
rect 970 1104 1000 1130
rect 1057 1104 1087 1130
rect 1143 1104 1173 1130
rect 1230 1104 1260 1130
rect 1316 1104 1346 1130
rect 1403 1104 1433 1130
rect 1489 1104 1519 1130
rect 1576 1104 1606 1130
rect 1662 1104 1692 1130
rect 1749 1104 1779 1130
rect 1835 1104 1865 1130
rect 711 1084 1865 1104
rect 711 1074 726 1084
rect 716 1050 726 1074
rect 761 1074 1865 1084
rect 1922 1104 1952 1130
rect 2008 1104 2038 1130
rect 2095 1104 2125 1130
rect 2181 1104 2211 1130
rect 2268 1104 2298 1130
rect 2354 1104 2384 1130
rect 2441 1104 2471 1130
rect 2527 1104 2557 1130
rect 2614 1104 2644 1130
rect 2700 1104 2730 1130
rect 2787 1104 2817 1130
rect 2873 1104 2903 1130
rect 2960 1104 2990 1130
rect 3046 1104 3076 1130
rect 1922 1074 3076 1104
rect 761 1050 771 1074
rect 716 1034 771 1050
rect 1778 1040 1788 1074
rect 1823 1040 1833 1074
rect 1778 1024 1833 1040
rect 1922 982 1952 1074
rect 1785 952 1952 982
rect 716 890 771 906
rect 716 866 726 890
rect 711 856 726 866
rect 761 866 771 890
rect 1785 866 1815 952
rect 1977 900 2032 916
rect 1977 866 1987 900
rect 2022 866 2032 900
rect 761 856 1865 866
rect 711 836 1865 856
rect 711 810 741 836
rect 797 810 827 836
rect 884 810 914 836
rect 970 810 1000 836
rect 1057 810 1087 836
rect 1143 810 1173 836
rect 1230 810 1260 836
rect 1316 810 1346 836
rect 1403 810 1433 836
rect 1489 810 1519 836
rect 1576 810 1606 836
rect 1662 810 1692 836
rect 1749 810 1779 836
rect 1835 810 1865 836
rect 1922 836 3076 866
rect 1922 810 1952 836
rect 2008 810 2038 836
rect 2095 810 2125 836
rect 2181 810 2211 836
rect 2268 810 2298 836
rect 2354 810 2384 836
rect 2441 810 2471 836
rect 2527 810 2557 836
rect 2614 810 2644 836
rect 2700 810 2730 836
rect 2787 810 2817 836
rect 2873 810 2903 836
rect 2960 810 2990 836
rect 3046 810 3076 836
rect 711 664 741 690
rect 797 664 827 690
rect 884 664 914 690
rect 970 664 1000 690
rect 1057 664 1087 690
rect 1143 664 1173 690
rect 1230 664 1260 690
rect 1316 664 1346 690
rect 1403 664 1433 690
rect 1489 664 1519 690
rect 1576 664 1606 690
rect 1662 664 1692 690
rect 1749 664 1779 690
rect 1835 664 1865 690
rect 711 634 1865 664
rect 1922 664 1952 690
rect 2008 664 2038 690
rect 2095 664 2125 690
rect 2181 664 2211 690
rect 2268 664 2298 690
rect 2354 664 2384 690
rect 2441 664 2471 690
rect 2527 664 2557 690
rect 2614 664 2644 690
rect 2700 664 2730 690
rect 2787 664 2817 690
rect 2873 664 2903 690
rect 2960 664 2990 690
rect 3046 664 3076 690
rect 1922 634 3076 664
<< polycont >>
rect 1827 1576 1861 1610
rect 1928 1364 1962 1398
rect 726 1050 761 1084
rect 1788 1040 1823 1074
rect 726 856 761 890
rect 1987 866 2022 900
<< locali >>
rect 1811 1576 1827 1610
rect 1861 1576 2170 1610
rect 1783 1505 1817 1521
rect 1783 1398 1817 1471
rect 1877 1505 1911 1521
rect 1877 1455 1911 1471
rect 1975 1505 2009 1576
rect 1975 1455 2009 1471
rect 2043 1505 2077 1521
rect 2043 1455 2077 1471
rect 1783 1364 1928 1398
rect 1962 1364 1978 1398
rect 666 1238 700 1254
rect 666 1188 700 1204
rect 839 1238 873 1254
rect 752 1176 786 1192
rect 839 1188 873 1204
rect 1012 1238 1046 1254
rect 752 1126 786 1142
rect 925 1176 959 1192
rect 1012 1188 1046 1204
rect 1185 1238 1219 1254
rect 925 1126 959 1142
rect 1098 1176 1132 1192
rect 1185 1188 1219 1204
rect 1358 1238 1392 1254
rect 1098 1126 1132 1142
rect 1271 1176 1305 1192
rect 1358 1188 1392 1204
rect 1531 1238 1565 1254
rect 1271 1126 1305 1142
rect 1444 1176 1478 1192
rect 1531 1188 1565 1204
rect 1704 1238 1738 1254
rect 1444 1126 1478 1142
rect 1617 1176 1651 1192
rect 1704 1188 1738 1204
rect 1617 1126 1651 1142
rect 1790 1176 1824 1364
rect 1877 1238 1911 1254
rect 1877 1188 1911 1204
rect 2050 1238 2084 1254
rect 1790 1126 1824 1142
rect 1963 1176 1997 1192
rect 2050 1188 2084 1204
rect 1963 1126 1997 1142
rect 2136 1176 2170 1576
rect 2223 1238 2257 1254
rect 2223 1188 2257 1204
rect 2396 1238 2430 1254
rect 2136 1126 2170 1142
rect 2309 1176 2343 1192
rect 2396 1188 2430 1204
rect 2569 1238 2603 1254
rect 2309 1126 2343 1142
rect 2482 1176 2516 1192
rect 2569 1188 2603 1204
rect 2742 1238 2776 1254
rect 2482 1126 2516 1142
rect 2655 1176 2689 1192
rect 2742 1188 2776 1204
rect 2915 1238 2949 1254
rect 2655 1126 2689 1142
rect 2828 1176 2862 1192
rect 2915 1188 2949 1204
rect 3088 1238 3122 1254
rect 2828 1126 2862 1142
rect 3001 1176 3035 1192
rect 3088 1188 3122 1204
rect 3001 1126 3035 1142
rect 710 1050 726 1084
rect 761 1050 777 1084
rect 1772 1040 1788 1074
rect 1823 1040 1839 1074
rect 1788 900 1823 1040
rect 710 856 726 890
rect 761 856 777 890
rect 1788 866 1987 900
rect 2022 866 2038 900
rect 666 798 700 814
rect 594 777 628 793
rect 666 748 700 764
rect 839 798 873 814
rect 594 727 628 743
rect 752 736 786 752
rect 839 748 873 764
rect 1012 798 1046 814
rect 752 686 786 702
rect 925 736 959 752
rect 1012 748 1046 764
rect 1185 798 1219 814
rect 925 686 959 702
rect 1098 736 1132 752
rect 1185 748 1219 764
rect 1358 798 1392 814
rect 1098 686 1132 702
rect 1271 736 1305 752
rect 1358 748 1392 764
rect 1531 798 1565 814
rect 1271 686 1305 702
rect 1444 736 1478 752
rect 1531 748 1565 764
rect 1704 798 1738 814
rect 1444 686 1478 702
rect 1617 736 1651 752
rect 1704 748 1738 764
rect 1877 798 1911 814
rect 1617 686 1651 702
rect 1790 736 1824 752
rect 1877 748 1911 764
rect 2050 798 2084 814
rect 1790 686 1824 702
rect 1963 736 1997 752
rect 2050 748 2084 764
rect 2223 798 2257 814
rect 1963 686 1997 702
rect 2136 736 2170 752
rect 2223 748 2257 764
rect 2396 798 2430 814
rect 2136 686 2170 702
rect 2309 736 2343 752
rect 2396 748 2430 764
rect 2569 798 2603 814
rect 2309 686 2343 702
rect 2482 736 2516 752
rect 2569 748 2603 764
rect 2742 798 2776 814
rect 2482 686 2516 702
rect 2655 736 2689 752
rect 2742 748 2776 764
rect 2915 798 2949 814
rect 2655 686 2689 702
rect 2828 736 2862 752
rect 2915 748 2949 764
rect 3088 798 3122 814
rect 2828 686 2862 702
rect 3001 736 3035 752
rect 3088 748 3122 764
rect 3166 783 3200 799
rect 3166 733 3200 749
rect 3001 686 3035 702
<< viali >>
rect 1877 1471 1911 1505
rect 2043 1471 2077 1505
rect 666 1204 700 1238
rect 839 1204 873 1238
rect 1012 1204 1046 1238
rect 752 1142 786 1176
rect 1185 1204 1219 1238
rect 925 1142 959 1176
rect 1358 1204 1392 1238
rect 1098 1142 1132 1176
rect 1531 1204 1565 1238
rect 1271 1142 1305 1176
rect 1704 1204 1738 1238
rect 1444 1142 1478 1176
rect 1617 1142 1651 1176
rect 1877 1204 1911 1238
rect 2050 1204 2084 1238
rect 1790 1142 1824 1176
rect 1963 1142 1997 1176
rect 2223 1204 2257 1238
rect 2396 1204 2430 1238
rect 2136 1142 2170 1176
rect 2569 1204 2603 1238
rect 2309 1142 2343 1176
rect 2742 1204 2776 1238
rect 2482 1142 2516 1176
rect 2915 1204 2949 1238
rect 2655 1142 2689 1176
rect 3088 1204 3122 1238
rect 2828 1142 2862 1176
rect 3001 1142 3035 1176
rect 726 1050 761 1084
rect 726 856 761 890
rect 594 743 628 777
rect 666 764 700 798
rect 839 764 873 798
rect 1012 764 1046 798
rect 752 702 786 736
rect 1185 764 1219 798
rect 925 702 959 736
rect 1358 764 1392 798
rect 1098 702 1132 736
rect 1531 764 1565 798
rect 1271 702 1305 736
rect 1704 764 1738 798
rect 1444 702 1478 736
rect 1877 764 1911 798
rect 1617 702 1651 736
rect 2050 764 2084 798
rect 1790 702 1824 736
rect 2223 764 2257 798
rect 1963 702 1997 736
rect 2396 764 2430 798
rect 2136 702 2170 736
rect 2569 764 2603 798
rect 2309 702 2343 736
rect 2742 764 2776 798
rect 2482 702 2516 736
rect 2915 764 2949 798
rect 2655 702 2689 736
rect 3088 764 3122 798
rect 2828 702 2862 736
rect 3166 749 3200 783
rect 3001 702 3035 736
<< metal1 >>
rect 429 1690 3342 1760
rect 1910 1517 1998 1690
rect 1871 1505 1998 1517
rect 2037 1505 2083 1511
rect 1871 1471 1877 1505
rect 1911 1471 2043 1505
rect 2077 1471 2089 1505
rect 1871 1465 1917 1471
rect 2037 1465 2083 1471
rect 1877 1244 1911 1465
rect 654 1238 3134 1244
rect 654 1204 666 1238
rect 700 1212 839 1238
rect 700 1204 712 1212
rect 654 1198 712 1204
rect 827 1204 839 1212
rect 873 1212 1012 1238
rect 873 1204 885 1212
rect 827 1198 885 1204
rect 1000 1204 1012 1212
rect 1046 1212 1185 1238
rect 1046 1204 1058 1212
rect 1000 1198 1058 1204
rect 1173 1204 1185 1212
rect 1219 1212 1358 1238
rect 1219 1204 1231 1212
rect 1173 1198 1231 1204
rect 1346 1204 1358 1212
rect 1392 1212 1531 1238
rect 1392 1204 1404 1212
rect 1346 1198 1404 1204
rect 1519 1204 1531 1212
rect 1565 1212 1704 1238
rect 1565 1204 1577 1212
rect 1519 1198 1577 1204
rect 1692 1204 1704 1212
rect 1738 1212 1877 1238
rect 1738 1204 1750 1212
rect 1692 1198 1750 1204
rect 1865 1204 1877 1212
rect 1911 1212 2050 1238
rect 1911 1204 1923 1212
rect 1865 1198 1923 1204
rect 2038 1204 2050 1212
rect 2084 1212 2223 1238
rect 2084 1204 2096 1212
rect 2038 1198 2096 1204
rect 2211 1204 2223 1212
rect 2257 1212 2396 1238
rect 2257 1204 2269 1212
rect 2211 1198 2269 1204
rect 2384 1204 2396 1212
rect 2430 1212 2569 1238
rect 2430 1204 2442 1212
rect 2384 1198 2442 1204
rect 2557 1204 2569 1212
rect 2603 1212 2742 1238
rect 2603 1204 2615 1212
rect 2557 1198 2615 1204
rect 2730 1204 2742 1212
rect 2776 1212 2915 1238
rect 2776 1204 2788 1212
rect 2730 1198 2788 1204
rect 2903 1204 2915 1212
rect 2949 1212 3088 1238
rect 2949 1204 2961 1212
rect 2903 1198 2961 1204
rect 3076 1204 3088 1212
rect 3122 1204 3134 1238
rect 3076 1198 3134 1204
rect 740 1176 801 1184
rect 740 1142 752 1176
rect 786 1167 801 1176
rect 913 1176 974 1184
rect 913 1167 925 1176
rect 786 1142 925 1167
rect 959 1167 974 1176
rect 1086 1176 1147 1184
rect 1086 1167 1098 1176
rect 959 1142 1098 1167
rect 1132 1167 1147 1176
rect 1259 1176 1320 1184
rect 1259 1167 1271 1176
rect 1132 1142 1271 1167
rect 1305 1167 1320 1176
rect 1432 1176 1493 1184
rect 1432 1167 1444 1176
rect 1305 1142 1444 1167
rect 1478 1167 1493 1176
rect 1603 1167 1609 1184
rect 1478 1142 1609 1167
rect 1661 1167 1667 1184
rect 1778 1176 1839 1184
rect 1778 1167 1790 1176
rect 1661 1142 1790 1167
rect 1824 1142 1839 1176
rect 1951 1176 2012 1184
rect 1951 1167 1963 1176
rect 740 1136 1609 1142
rect 1603 1132 1609 1136
rect 1661 1136 1839 1142
rect 1950 1142 1963 1167
rect 1997 1167 2012 1176
rect 2121 1167 2127 1184
rect 1997 1142 2127 1167
rect 2179 1167 2185 1184
rect 2297 1176 2358 1184
rect 2297 1167 2309 1176
rect 2179 1142 2309 1167
rect 2343 1167 2358 1176
rect 2470 1176 2531 1184
rect 2470 1167 2482 1176
rect 2343 1142 2482 1167
rect 2516 1167 2531 1176
rect 2643 1176 2704 1184
rect 2643 1167 2655 1176
rect 2516 1142 2655 1167
rect 2689 1167 2704 1176
rect 2816 1176 2877 1184
rect 2816 1167 2828 1176
rect 2689 1142 2828 1167
rect 2862 1167 2877 1176
rect 2989 1176 3050 1184
rect 2989 1167 3001 1176
rect 2862 1142 3001 1167
rect 3035 1167 3050 1176
rect 3035 1142 3133 1167
rect 1950 1136 2127 1142
rect 1661 1132 1667 1136
rect 2121 1132 2127 1136
rect 2179 1136 3133 1142
rect 2179 1132 2185 1136
rect 1603 1131 1667 1132
rect 720 1084 773 1090
rect 429 1050 726 1084
rect 761 1050 773 1084
rect 720 1044 773 1050
rect 2120 1016 2126 1068
rect 2178 1059 2184 1068
rect 2178 1025 3342 1059
rect 2178 1016 2184 1025
rect 720 890 767 896
rect 1604 894 1610 946
rect 1662 937 1668 946
rect 1662 903 3342 937
rect 1662 894 1668 903
rect 429 856 726 890
rect 761 856 773 890
rect 720 850 767 856
rect 588 798 3206 804
rect 588 777 666 798
rect 588 743 594 777
rect 628 764 666 777
rect 700 772 839 798
rect 700 764 712 772
rect 628 758 712 764
rect 827 764 839 772
rect 873 772 1012 798
rect 873 764 885 772
rect 827 758 885 764
rect 1000 764 1012 772
rect 1046 772 1185 798
rect 1046 764 1058 772
rect 1000 758 1058 764
rect 1173 764 1185 772
rect 1219 772 1358 798
rect 1219 764 1231 772
rect 1173 758 1231 764
rect 1346 764 1358 772
rect 1392 772 1531 798
rect 1392 764 1404 772
rect 1346 758 1404 764
rect 1519 764 1531 772
rect 1565 772 1704 798
rect 1565 764 1577 772
rect 1519 758 1577 764
rect 1692 764 1704 772
rect 1738 772 1877 798
rect 1738 764 1750 772
rect 1692 758 1750 764
rect 1865 764 1877 772
rect 1911 772 2050 798
rect 1911 764 1923 772
rect 1865 758 1923 764
rect 2038 764 2050 772
rect 2084 772 2223 798
rect 2084 764 2096 772
rect 2038 758 2096 764
rect 2211 764 2223 772
rect 2257 772 2396 798
rect 2257 764 2269 772
rect 2211 758 2269 764
rect 2384 764 2396 772
rect 2430 772 2569 798
rect 2430 764 2442 772
rect 2384 758 2442 764
rect 2557 764 2569 772
rect 2603 772 2742 798
rect 2603 764 2615 772
rect 2557 758 2615 764
rect 2730 764 2742 772
rect 2776 772 2915 798
rect 2776 764 2788 772
rect 2730 758 2788 764
rect 2903 764 2915 772
rect 2949 772 3088 798
rect 2949 764 2961 772
rect 2903 758 2961 764
rect 3076 764 3088 772
rect 3122 783 3206 798
rect 3122 764 3166 783
rect 3076 758 3166 764
rect 628 743 638 758
rect 588 731 638 743
rect 740 736 801 744
rect 740 702 752 736
rect 786 727 801 736
rect 913 736 974 744
rect 913 727 925 736
rect 786 702 925 727
rect 959 727 974 736
rect 1086 736 1147 744
rect 1086 727 1098 736
rect 959 702 1098 727
rect 1132 727 1147 736
rect 1259 736 1320 744
rect 1259 727 1271 736
rect 1132 702 1271 727
rect 1305 727 1320 736
rect 1432 736 1493 744
rect 1432 727 1444 736
rect 1305 702 1444 727
rect 1478 727 1493 736
rect 1603 743 1667 744
rect 1603 727 1609 743
rect 1478 702 1609 727
rect 1661 727 1667 743
rect 1778 736 1839 744
rect 1778 727 1790 736
rect 1661 702 1790 727
rect 1824 702 1839 736
rect 740 696 1609 702
rect 1603 691 1609 696
rect 1661 696 1839 702
rect 1661 691 1667 696
rect 1877 572 1911 758
rect 3158 749 3166 758
rect 3200 749 3206 783
rect 1951 736 2012 744
rect 2124 742 2185 744
rect 1951 727 1963 736
rect 1950 702 1963 727
rect 1997 727 2012 736
rect 2123 727 2129 742
rect 1997 702 2129 727
rect 2181 727 2187 742
rect 2297 736 2358 744
rect 2297 727 2309 736
rect 2181 702 2309 727
rect 2343 727 2358 736
rect 2470 736 2531 744
rect 2470 727 2482 736
rect 2343 702 2482 727
rect 2516 727 2531 736
rect 2643 736 2704 744
rect 2643 727 2655 736
rect 2516 702 2655 727
rect 2689 727 2704 736
rect 2816 736 2877 744
rect 2816 727 2828 736
rect 2689 702 2828 727
rect 2862 727 2877 736
rect 2989 736 3050 744
rect 3158 737 3206 749
rect 2989 727 3001 736
rect 2862 702 3001 727
rect 3035 702 3050 736
rect 1950 696 2129 702
rect 2123 690 2129 696
rect 2181 696 3050 702
rect 2181 690 2187 696
rect 429 502 3342 572
<< via1 >>
rect 1609 1176 1661 1184
rect 1609 1142 1617 1176
rect 1617 1142 1651 1176
rect 1651 1142 1661 1176
rect 1609 1132 1661 1142
rect 2127 1176 2179 1184
rect 2127 1142 2136 1176
rect 2136 1142 2170 1176
rect 2170 1142 2179 1176
rect 2127 1132 2179 1142
rect 2126 1016 2178 1068
rect 1610 894 1662 946
rect 1609 736 1661 743
rect 1609 702 1617 736
rect 1617 702 1651 736
rect 1651 702 1661 736
rect 1609 691 1661 702
rect 2129 736 2181 742
rect 2129 702 2136 736
rect 2136 702 2170 736
rect 2170 702 2181 736
rect 2129 690 2181 702
<< metal2 >>
rect 1603 1132 1609 1184
rect 1661 1132 1667 1184
rect 2121 1132 2127 1184
rect 2179 1132 2185 1184
rect 1617 946 1651 1132
rect 2136 1068 2170 1132
rect 2120 1016 2126 1068
rect 2178 1016 2184 1068
rect 1604 894 1610 946
rect 1662 894 1668 946
rect 1617 743 1651 894
rect 1603 691 1609 743
rect 1661 691 1667 743
rect 2136 742 2170 1016
rect 2123 690 2129 742
rect 2181 690 2187 742
<< labels >>
flabel space 1910 1690 2001 1761 0 FreeSans 480 0 0 0 VDDA
flabel space 1850 502 1941 573 0 FreeSans 480 0 0 0 GND
flabel metal1 726 856 761 890 0 FreeSans 160 0 0 0 inb
flabel metal1 726 1050 761 1084 0 FreeSans 160 0 0 0 in
flabel via1 2126 1016 2178 1068 0 FreeSans 160 0 0 0 out
flabel via1 1610 894 1662 946 0 FreeSans 160 0 0 0 outb
<< end >>
