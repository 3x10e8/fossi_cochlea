magic
tech sky130A
magscale 1 2
timestamp 1654690121
<< obsli1 >>
rect 1104 2159 98808 47345
<< obsm1 >>
rect 14 280 98808 49496
<< metal2 >>
rect 5170 49200 5226 50000
rect 12898 49200 12954 50000
rect 20626 49200 20682 50000
rect 27710 49200 27766 50000
rect 35438 49200 35494 50000
rect 43166 49200 43222 50000
rect 50894 49200 50950 50000
rect 58622 49200 58678 50000
rect 65706 49200 65762 50000
rect 73434 49200 73490 50000
rect 81162 49200 81218 50000
rect 88890 49200 88946 50000
rect 96618 49200 96674 50000
rect 18 0 74 800
rect 7102 0 7158 800
rect 14830 0 14886 800
rect 22558 0 22614 800
rect 30286 0 30342 800
rect 37370 0 37426 800
rect 45098 0 45154 800
rect 52826 0 52882 800
rect 60554 0 60610 800
rect 68282 0 68338 800
rect 75366 0 75422 800
rect 83094 0 83150 800
rect 90822 0 90878 800
rect 98550 0 98606 800
<< obsm2 >>
rect 20 49144 5114 49881
rect 5282 49144 12842 49881
rect 13010 49144 20570 49881
rect 20738 49144 27654 49881
rect 27822 49144 35382 49881
rect 35550 49144 43110 49881
rect 43278 49144 50838 49881
rect 51006 49144 58566 49881
rect 58734 49144 65650 49881
rect 65818 49144 73378 49881
rect 73546 49144 81106 49881
rect 81274 49144 88834 49881
rect 89002 49144 96562 49881
rect 96730 49144 98604 49881
rect 20 856 98604 49144
rect 130 274 7046 856
rect 7214 274 14774 856
rect 14942 274 22502 856
rect 22670 274 30230 856
rect 30398 274 37314 856
rect 37482 274 45042 856
rect 45210 274 52770 856
rect 52938 274 60498 856
rect 60666 274 68226 856
rect 68394 274 75310 856
rect 75478 274 83038 856
rect 83206 274 90766 856
rect 90934 274 98494 856
<< metal3 >>
rect 0 47608 800 47728
rect 99200 46248 100000 46368
rect 0 39448 800 39568
rect 99200 38088 100000 38208
rect 0 31968 800 32088
rect 99200 29928 100000 30048
rect 0 23808 800 23928
rect 99200 21768 100000 21888
rect 0 15648 800 15768
rect 99200 13608 100000 13728
rect 0 7488 800 7608
rect 99200 6128 100000 6248
<< obsm3 >>
rect 26190 50000 67466 50010
rect 800 47808 99200 50000
rect 880 47528 99200 47808
rect 800 46448 99200 47528
rect 800 46168 99120 46448
rect 800 39648 99200 46168
rect 880 39368 99200 39648
rect 800 38288 99200 39368
rect 800 38008 99120 38288
rect 800 32168 99200 38008
rect 880 31888 99200 32168
rect 800 30128 99200 31888
rect 800 29848 99120 30128
rect 800 24008 99200 29848
rect 880 23728 99200 24008
rect 800 21968 99200 23728
rect 800 21688 99120 21968
rect 800 15848 99200 21688
rect 880 15568 99200 15848
rect 800 13808 99200 15568
rect 800 13528 99120 13808
rect 800 7688 99200 13528
rect 880 7408 99200 7688
rect 800 6328 99200 7408
rect 800 6048 99120 6328
rect 800 308 99200 6048
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
rect 50288 2128 50608 47376
rect 65648 2128 65968 47376
rect 81008 2128 81328 47376
rect 96368 2128 96688 47376
<< obsm4 >>
rect 16435 47456 88445 49877
rect 16435 2048 19488 47456
rect 19968 2048 34848 47456
rect 35328 2048 50208 47456
rect 50688 2048 65568 47456
rect 66048 2048 80928 47456
rect 81408 2048 88445 47456
rect 16435 307 88445 2048
<< labels >>
rlabel metal2 s 52826 0 52882 800 6 cclk_I[0]
port 1 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 cclk_I[1]
port 2 nsew signal output
rlabel metal2 s 73434 49200 73490 50000 6 cclk_Q[0]
port 3 nsew signal output
rlabel metal3 s 99200 13608 100000 13728 6 cclk_Q[1]
port 4 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 clk_master
port 5 nsew signal input
rlabel metal2 s 65706 49200 65762 50000 6 clkdiv2_I[0]
port 6 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 clkdiv2_I[1]
port 7 nsew signal output
rlabel metal2 s 35438 49200 35494 50000 6 clkdiv2_Q[0]
port 8 nsew signal output
rlabel metal3 s 99200 29928 100000 30048 6 clkdiv2_Q[1]
port 9 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 comp_high_I[0]
port 10 nsew signal input
rlabel metal2 s 96618 49200 96674 50000 6 comp_high_I[1]
port 11 nsew signal input
rlabel metal3 s 99200 38088 100000 38208 6 comp_high_Q[0]
port 12 nsew signal input
rlabel metal2 s 43166 49200 43222 50000 6 comp_high_Q[1]
port 13 nsew signal input
rlabel metal2 s 12898 49200 12954 50000 6 cos_out[0]
port 14 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 cos_out[1]
port 15 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 cos_outb[0]
port 16 nsew signal output
rlabel metal3 s 99200 21768 100000 21888 6 cos_outb[1]
port 17 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 fb1_I[0]
port 18 nsew signal output
rlabel metal2 s 18 0 74 800 6 fb1_I[1]
port 19 nsew signal output
rlabel metal2 s 81162 49200 81218 50000 6 fb1_Q[0]
port 20 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 fb1_Q[1]
port 21 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 fb2_I[0]
port 22 nsew signal output
rlabel metal2 s 27710 49200 27766 50000 6 fb2_I[1]
port 23 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 fb2_Q[0]
port 24 nsew signal output
rlabel metal2 s 88890 49200 88946 50000 6 fb2_Q[1]
port 25 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 phi1b_dig_I[0]
port 26 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 phi1b_dig_I[1]
port 27 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 phi1b_dig_Q[0]
port 28 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 phi1b_dig_Q[1]
port 29 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 read_out_I[0]
port 30 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 read_out_I[1]
port 31 nsew signal output
rlabel metal2 s 5170 49200 5226 50000 6 read_out_Q[0]
port 32 nsew signal output
rlabel metal3 s 99200 46248 100000 46368 6 read_out_Q[1]
port 33 nsew signal output
rlabel metal2 s 50894 49200 50950 50000 6 rstb
port 34 nsew signal input
rlabel metal2 s 58622 49200 58678 50000 6 sin_out[0]
port 35 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 sin_out[1]
port 36 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 sin_outb[0]
port 37 nsew signal output
rlabel metal2 s 20626 49200 20682 50000 6 sin_outb[1]
port 38 nsew signal output
rlabel metal3 s 99200 6128 100000 6248 6 ud_en
port 39 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 40 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 40 nsew power input
rlabel metal4 s 65648 2128 65968 47376 6 vccd1
port 40 nsew power input
rlabel metal4 s 96368 2128 96688 47376 6 vccd1
port 40 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 41 nsew ground input
rlabel metal4 s 50288 2128 50608 47376 6 vssd1
port 41 nsew ground input
rlabel metal4 s 81008 2128 81328 47376 6 vssd1
port 41 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 100000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7886034
string GDS_FILE /Volumes/export/isn/abhinav/fossi_cochlea/openlane/digital_unison/runs/digital_unison/results/finishing/digital_unison.magic.gds
string GDS_START 459984
<< end >>

