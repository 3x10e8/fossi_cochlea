magic
tech sky130A
magscale 1 2
timestamp 1654738073
<< obsli1 >>
rect 1104 2159 78844 53329
<< obsm1 >>
rect 1104 1232 79014 55684
<< metal2 >>
rect 2042 55200 2098 56000
rect 6182 55200 6238 56000
rect 10414 55200 10470 56000
rect 14646 55200 14702 56000
rect 18878 55200 18934 56000
rect 23018 55200 23074 56000
rect 27250 55200 27306 56000
rect 31482 55200 31538 56000
rect 35714 55200 35770 56000
rect 39946 55200 40002 56000
rect 44086 55200 44142 56000
rect 48318 55200 48374 56000
rect 52550 55200 52606 56000
rect 56782 55200 56838 56000
rect 61014 55200 61070 56000
rect 65154 55200 65210 56000
rect 69386 55200 69442 56000
rect 73618 55200 73674 56000
rect 77850 55200 77906 56000
rect 4986 0 5042 800
rect 14922 0 14978 800
rect 24950 0 25006 800
rect 34978 0 35034 800
rect 45006 0 45062 800
rect 54942 0 54998 800
rect 64970 0 65026 800
rect 74998 0 75054 800
<< obsm2 >>
rect 1398 55144 1986 55865
rect 2154 55144 6126 55865
rect 6294 55144 10358 55865
rect 10526 55144 14590 55865
rect 14758 55144 18822 55865
rect 18990 55144 22962 55865
rect 23130 55144 27194 55865
rect 27362 55144 31426 55865
rect 31594 55144 35658 55865
rect 35826 55144 39890 55865
rect 40058 55144 44030 55865
rect 44198 55144 48262 55865
rect 48430 55144 52494 55865
rect 52662 55144 56726 55865
rect 56894 55144 60958 55865
rect 61126 55144 65098 55865
rect 65266 55144 69330 55865
rect 69498 55144 73562 55865
rect 73730 55144 77794 55865
rect 77962 55144 79102 55865
rect 1398 856 79102 55144
rect 1398 734 4930 856
rect 5098 734 14866 856
rect 15034 734 24894 856
rect 25062 734 34922 856
rect 35090 734 44950 856
rect 45118 734 54886 856
rect 55054 734 64914 856
rect 65082 734 74942 856
rect 75110 734 79102 856
<< metal3 >>
rect 0 54272 800 54392
rect 79200 54136 80000 54256
rect 0 51008 800 51128
rect 79200 50600 80000 50720
rect 0 47744 800 47864
rect 79200 47064 80000 47184
rect 0 44480 800 44600
rect 79200 43664 80000 43784
rect 0 41080 800 41200
rect 79200 40128 80000 40248
rect 0 37816 800 37936
rect 79200 36592 80000 36712
rect 0 34552 800 34672
rect 79200 33056 80000 33176
rect 0 31288 800 31408
rect 79200 29656 80000 29776
rect 0 27888 800 28008
rect 79200 26120 80000 26240
rect 0 24624 800 24744
rect 79200 22584 80000 22704
rect 0 21360 800 21480
rect 79200 19048 80000 19168
rect 0 18096 800 18216
rect 79200 15648 80000 15768
rect 0 14696 800 14816
rect 79200 12112 80000 12232
rect 0 11432 800 11552
rect 79200 8576 80000 8696
rect 0 8168 800 8288
rect 0 4904 800 5024
rect 79200 5040 80000 5160
rect 0 1640 800 1760
rect 79200 1640 80000 1760
<< obsm3 >>
rect 800 54472 79200 55996
rect 880 54336 79200 54472
rect 880 54192 79120 54336
rect 800 54056 79120 54192
rect 800 51208 79200 54056
rect 880 50928 79200 51208
rect 800 50800 79200 50928
rect 800 50520 79120 50800
rect 800 47944 79200 50520
rect 880 47664 79200 47944
rect 800 47264 79200 47664
rect 800 46984 79120 47264
rect 800 44680 79200 46984
rect 880 44400 79200 44680
rect 800 43864 79200 44400
rect 800 43584 79120 43864
rect 800 41280 79200 43584
rect 880 41000 79200 41280
rect 800 40328 79200 41000
rect 800 40048 79120 40328
rect 800 38016 79200 40048
rect 880 37736 79200 38016
rect 800 36792 79200 37736
rect 800 36512 79120 36792
rect 800 34752 79200 36512
rect 880 34472 79200 34752
rect 800 33256 79200 34472
rect 800 32976 79120 33256
rect 800 31488 79200 32976
rect 880 31208 79200 31488
rect 800 29856 79200 31208
rect 800 29576 79120 29856
rect 800 28088 79200 29576
rect 880 27808 79200 28088
rect 800 26320 79200 27808
rect 800 26040 79120 26320
rect 800 24824 79200 26040
rect 880 24544 79200 24824
rect 800 22784 79200 24544
rect 800 22504 79120 22784
rect 800 21560 79200 22504
rect 880 21280 79200 21560
rect 800 19248 79200 21280
rect 800 18968 79120 19248
rect 800 18296 79200 18968
rect 880 18016 79200 18296
rect 800 15848 79200 18016
rect 800 15568 79120 15848
rect 800 14896 79200 15568
rect 880 14616 79200 14896
rect 800 12312 79200 14616
rect 800 12032 79120 12312
rect 800 11632 79200 12032
rect 880 11352 79200 11632
rect 800 8776 79200 11352
rect 800 8496 79120 8776
rect 800 8368 79200 8496
rect 880 8088 79200 8368
rect 800 5240 79200 8088
rect 800 5104 79120 5240
rect 880 4960 79120 5104
rect 880 4824 79200 4960
rect 800 1840 79200 4824
rect 880 1560 79120 1840
rect 800 1532 79200 1560
<< metal4 >>
rect 4208 2128 4528 53360
rect 19568 2128 19888 53360
rect 34928 2128 35248 53360
rect 50288 2128 50608 53360
rect 65648 2128 65968 53360
<< obsm4 >>
rect 8155 53440 76485 55997
rect 8155 2048 19488 53440
rect 19968 2048 34848 53440
rect 35328 2048 50208 53440
rect 50688 2048 65568 53440
rect 66048 2048 76485 53440
rect 8155 1531 76485 2048
<< labels >>
rlabel metal3 s 0 18096 800 18216 6 cclk_I[0]
port 1 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 cclk_I[1]
port 2 nsew signal output
rlabel metal3 s 79200 5040 80000 5160 6 cclk_Q[0]
port 3 nsew signal output
rlabel metal3 s 79200 29656 80000 29776 6 cclk_Q[1]
port 4 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 clk_master
port 5 nsew signal input
rlabel metal2 s 6182 55200 6238 56000 6 clk_master_out
port 6 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 clkdiv2_I[0]
port 7 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 clkdiv2_I[1]
port 8 nsew signal output
rlabel metal3 s 79200 8576 80000 8696 6 clkdiv2_Q[0]
port 9 nsew signal output
rlabel metal3 s 79200 33056 80000 33176 6 clkdiv2_Q[1]
port 10 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 comp_high_I[0]
port 11 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 comp_high_I[1]
port 12 nsew signal input
rlabel metal3 s 79200 12112 80000 12232 6 comp_high_Q[0]
port 13 nsew signal input
rlabel metal3 s 79200 36592 80000 36712 6 comp_high_Q[1]
port 14 nsew signal input
rlabel metal3 s 0 21360 800 21480 6 cos_out[0]
port 15 nsew signal output
rlabel metal3 s 0 44480 800 44600 6 cos_out[1]
port 16 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 cos_outb[0]
port 17 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 cos_outb[1]
port 18 nsew signal output
rlabel metal2 s 14646 55200 14702 56000 6 div2out
port 19 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 fb1_I[0]
port 20 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 fb1_I[1]
port 21 nsew signal output
rlabel metal3 s 79200 19048 80000 19168 6 fb1_Q[0]
port 22 nsew signal output
rlabel metal3 s 79200 43664 80000 43784 6 fb1_Q[1]
port 23 nsew signal output
rlabel metal2 s 73618 55200 73674 56000 6 fb2_I[0]
port 24 nsew signal output
rlabel metal2 s 77850 55200 77906 56000 6 fb2_I[1]
port 25 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 fb2_Q[0]
port 26 nsew signal output
rlabel metal3 s 0 54272 800 54392 6 fb2_Q[1]
port 27 nsew signal output
rlabel metal2 s 56782 55200 56838 56000 6 gray_clk_out[10]
port 28 nsew signal output
rlabel metal2 s 18878 55200 18934 56000 6 gray_clk_out[1]
port 29 nsew signal output
rlabel metal2 s 23018 55200 23074 56000 6 gray_clk_out[2]
port 30 nsew signal output
rlabel metal2 s 27250 55200 27306 56000 6 gray_clk_out[3]
port 31 nsew signal output
rlabel metal2 s 31482 55200 31538 56000 6 gray_clk_out[4]
port 32 nsew signal output
rlabel metal2 s 35714 55200 35770 56000 6 gray_clk_out[5]
port 33 nsew signal output
rlabel metal2 s 39946 55200 40002 56000 6 gray_clk_out[6]
port 34 nsew signal output
rlabel metal2 s 44086 55200 44142 56000 6 gray_clk_out[7]
port 35 nsew signal output
rlabel metal2 s 48318 55200 48374 56000 6 gray_clk_out[8]
port 36 nsew signal output
rlabel metal2 s 52550 55200 52606 56000 6 gray_clk_out[9]
port 37 nsew signal output
rlabel metal2 s 61014 55200 61070 56000 6 no_ones_below_out[0]
port 38 nsew signal output
rlabel metal2 s 65154 55200 65210 56000 6 no_ones_below_out[1]
port 39 nsew signal output
rlabel metal2 s 69386 55200 69442 56000 6 no_ones_below_out[2]
port 40 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 phi1b_dig_I[0]
port 41 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 phi1b_dig_I[1]
port 42 nsew signal input
rlabel metal3 s 79200 15648 80000 15768 6 phi1b_dig_Q[0]
port 43 nsew signal input
rlabel metal3 s 79200 40128 80000 40248 6 phi1b_dig_Q[1]
port 44 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 read_out_I[0]
port 45 nsew signal output
rlabel metal2 s 14922 0 14978 800 6 read_out_I[1]
port 46 nsew signal output
rlabel metal3 s 0 47744 800 47864 6 read_out_I_top[0]
port 47 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 read_out_I_top[1]
port 48 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 read_out_Q[0]
port 49 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 read_out_Q[1]
port 50 nsew signal output
rlabel metal3 s 79200 50600 80000 50720 6 read_out_Q_top[0]
port 51 nsew signal output
rlabel metal3 s 79200 54136 80000 54256 6 read_out_Q_top[1]
port 52 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 rstb
port 53 nsew signal input
rlabel metal2 s 2042 55200 2098 56000 6 rstb_out
port 54 nsew signal output
rlabel metal3 s 79200 1640 80000 1760 6 sin_out[0]
port 55 nsew signal output
rlabel metal3 s 79200 26120 80000 26240 6 sin_out[1]
port 56 nsew signal output
rlabel metal3 s 79200 22584 80000 22704 6 sin_outb[0]
port 57 nsew signal output
rlabel metal3 s 79200 47064 80000 47184 6 sin_outb[1]
port 58 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 ud_en
port 59 nsew signal input
rlabel metal2 s 10414 55200 10470 56000 6 ud_en_out
port 60 nsew signal output
rlabel metal4 s 4208 2128 4528 53360 6 vccd1
port 61 nsew power input
rlabel metal4 s 34928 2128 35248 53360 6 vccd1
port 61 nsew power input
rlabel metal4 s 65648 2128 65968 53360 6 vccd1
port 61 nsew power input
rlabel metal4 s 19568 2128 19888 53360 6 vssd1
port 62 nsew ground input
rlabel metal4 s 50288 2128 50608 53360 6 vssd1
port 62 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 80000 56000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7790494
string GDS_FILE /Volumes/export/isn/abhinav/fossi_cochlea/openlane/first_dual_core/runs/first_dual_core/results/finishing/first_dual_core.magic.gds
string GDS_START 432676
<< end >>

