magic
tech sky130A
timestamp 1647868321
<< viali >>
rect 5719 -5081 5736 -5064
rect 5772 -5081 5789 -5064
<< metal1 >>
rect 5783 -1259 5809 -1256
rect 5596 -1285 5783 -1273
rect 5809 -1285 5862 -1273
rect 5596 -1287 5862 -1285
rect 5783 -1288 5809 -1287
rect 5747 -1304 5773 -1302
rect 5597 -1305 5872 -1304
rect 5597 -1318 5747 -1305
rect 5773 -1318 5872 -1305
rect 5747 -1334 5773 -1331
rect 5600 -1347 5626 -1344
rect 5158 -1367 5600 -1350
rect 5626 -1367 5872 -1350
rect 5600 -1376 5626 -1373
rect 5713 -1581 5739 -1578
rect 5597 -1599 5713 -1585
rect 5713 -1610 5739 -1607
rect 5817 -1581 5843 -1578
rect 5843 -1599 5861 -1585
rect 5817 -1610 5843 -1607
rect 5637 -1718 5663 -1715
rect 5596 -1744 5637 -1734
rect 5663 -1744 5859 -1734
rect 5596 -1748 5859 -1744
rect 5683 -1765 5709 -1762
rect 5597 -1780 5683 -1766
rect 5709 -1780 5861 -1766
rect 5683 -1794 5709 -1791
rect 5712 -5055 5742 -5052
rect 5712 -5057 5744 -5055
rect 5742 -5087 5744 -5057
rect 5712 -5089 5744 -5087
rect 5765 -5058 5796 -5055
rect 5765 -5064 5790 -5058
rect 5765 -5081 5772 -5064
rect 5789 -5081 5790 -5064
rect 5765 -5084 5790 -5081
rect 5816 -5084 5819 -5058
rect 5712 -5092 5742 -5089
rect 5765 -5090 5796 -5084
<< via1 >>
rect 5783 -1285 5809 -1259
rect 5747 -1331 5773 -1305
rect 5600 -1373 5626 -1347
rect 5713 -1607 5739 -1581
rect 5817 -1607 5843 -1581
rect 5637 -1744 5663 -1718
rect 5683 -1791 5709 -1765
rect 5712 -5064 5742 -5057
rect 5712 -5081 5719 -5064
rect 5719 -5081 5736 -5064
rect 5736 -5081 5742 -5064
rect 5712 -5087 5742 -5081
rect 5790 -5084 5816 -5058
<< metal2 >>
rect 5613 -1344 5628 3199
rect 5600 -1347 5628 -1344
rect 5626 -1373 5628 -1347
rect 5600 -1376 5628 -1373
rect 5648 -1715 5663 3199
rect 5637 -1718 5663 -1715
rect 5637 -1747 5663 -1744
rect 5642 -1748 5663 -1747
rect 5648 -4841 5663 -1748
rect 5683 -1762 5698 3199
rect 5718 -1578 5733 3199
rect 5753 -1302 5768 3199
rect 5788 -1256 5803 3199
rect 5783 -1259 5809 -1256
rect 5783 -1288 5809 -1285
rect 5747 -1305 5773 -1302
rect 5747 -1334 5773 -1331
rect 5713 -1581 5739 -1578
rect 5713 -1610 5739 -1607
rect 5683 -1765 5709 -1762
rect 5683 -1794 5709 -1791
rect 5753 -4840 5768 -1334
rect 5823 -1578 5838 3199
rect 5817 -1581 5843 -1578
rect 5817 -1610 5843 -1607
rect 5712 -5055 5742 -5052
rect 5712 -5057 5744 -5055
rect 5742 -5087 5744 -5057
rect 5712 -5089 5744 -5087
rect 5765 -5056 5796 -5055
rect 5765 -5084 5790 -5056
rect 5819 -5084 5824 -5056
rect 5712 -5092 5742 -5089
rect 5765 -5090 5796 -5084
<< via2 >>
rect 5712 -5087 5742 -5057
rect 5790 -5058 5819 -5056
rect 5790 -5084 5816 -5058
rect 5816 -5084 5819 -5058
<< metal3 >>
rect 5705 -5055 5745 -5050
rect 5705 -5056 5712 -5055
rect 5680 -5086 5712 -5056
rect 5705 -5087 5712 -5086
rect 5744 -5087 5745 -5055
rect 5705 -5092 5745 -5087
rect 5784 -5052 5839 -5045
rect 5784 -5084 5790 -5052
rect 5822 -5084 5839 -5052
rect 5784 -5097 5839 -5084
<< via3 >>
rect 5712 -5057 5744 -5055
rect 5712 -5087 5742 -5057
rect 5742 -5087 5744 -5057
rect 5790 -5056 5822 -5052
rect 5790 -5084 5819 -5056
rect 5819 -5084 5822 -5056
<< metal4 >>
rect 5563 -4815 5592 -4814
rect 5563 -5056 5593 -4815
rect 5807 -4825 5860 -4776
rect 5807 -5024 5837 -4825
rect 5798 -5051 5837 -5024
rect 5787 -5052 5837 -5051
rect 5709 -5055 5745 -5054
rect 5709 -5056 5712 -5055
rect 5563 -5086 5712 -5056
rect 5709 -5087 5712 -5086
rect 5744 -5087 5745 -5055
rect 5787 -5084 5790 -5052
rect 5822 -5054 5837 -5052
rect 5822 -5084 5829 -5054
rect 5787 -5085 5829 -5084
rect 5709 -5088 5745 -5087
rect 5712 -5089 5744 -5088
use comparator_final  comparator_final_0
timestamp 1647868321
transform 1 0 5935 0 1 -5019
box -286 -215 609 167
use fitler_cell  fitler_cell_1
timestamp 1647840975
transform -1 0 11449 0 1 0
box -2644 -4825 5604 3103
use fitler_cell  fitler_cell_0
timestamp 1647840975
transform 1 0 2 0 1 0
box -2644 -4825 5604 3103
<< end >>
