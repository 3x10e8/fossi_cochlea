** sch_path: /local_disk/fossi_cochlea/xschem/Switched_Caps/mim_cap_stacked_12pF.sch
.subckt mim_cap_stacked_12pF sig vss
*.PININFO sig:B vss:B
XC1 sig vss sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=32 m=32
XC2 sig vss sky130_fd_pr__cap_mim_m3_2 W=10 L=10 MF=32 m=32
**** begin user architecture code
 .lib /local_disk/fossi_cochlea/dependencies/pdks/sky130B/libs.tech/ngspice/sky130.lib.spice tt
.include /local_disk/fossi_cochlea/dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
.ends
.end
