* NGSPICE file created from /local_disk/fossi_cochlea/mag/final_designs/filter/filter_p_m.ext - technology: sky130B

.subckt inv_weak_pulldown_corrected a_30_590# a_n177_50# vnb w_n204_554# in li_n276_n97#
X0 a_30_590# in w_n204_554# w_n204_554# sky130_fd_pr__pfet_01v8 ad=5.04e+11p pd=3.32e+06u as=4.914e+11p ps=3.3e+06u w=1.26e+06u l=180000u
X1 a_30_50# in a_n177_50# a_n177_50# sky130_fd_pr__nfet_01v8 ad=1.323e+11p pd=1.47e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=180000u
X2 a_30_590# vnb a_30_50# a_n177_50# sky130_fd_pr__nfet_01v8 ad=1.323e+11p pd=1.47e+06u as=0p ps=0u w=420000u l=540000u
.ends

.subckt tg inp out clk_ clk
X0 out clk_ inp clk sky130_fd_pr__pfet_01v8 ad=5.859e+11p pd=4.38e+06u as=2.52e+11p ps=2.06e+06u w=630000u l=180000u
X1 inp clk_ out clk sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=180000u
X2 out clk inp clk_ sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=2.415e+11p ps=1.99e+06u w=420000u l=180000u
.ends

.subckt inverter w_n204_204# a_n177_0# out in
X0 out in a_n177_0# a_n177_0# sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=180000u
X1 w_n204_204# in out w_n204_204# sky130_fd_pr__pfet_01v8 ad=5.859e+11p pd=4.38e+06u as=2.52e+11p ps=2.06e+06u w=630000u l=180000u
X2 out in w_n204_204# w_n204_204# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=180000u
.ends

.subckt comp_clks inverter_1/out tg_0/inp inverter_2/out w_577_332# tg_0/clk VSUBS
Xtg_0 tg_0/inp tg_0/out VSUBS tg_0/clk tg
Xinverter_0 w_577_332# VSUBS inverter_1/in tg_0/inp inverter
Xinverter_1 w_577_332# VSUBS inverter_1/out inverter_1/in inverter
Xinverter_2 tg_0/clk VSUBS inverter_2/out tg_0/out inverter
.ends

.subckt cclkgen inv_weak_pulldown_corrected_1/vnb comp_clks_0/inverter_2/out comp_clks_0/tg_0/clk
+ inv_weak_pulldown_corrected_0/vnb inv_weak_pulldown_corrected_0/in comp_clks_0/w_577_332#
+ comp_clks_0/inverter_1/out VSUBS
Xinv_weak_pulldown_corrected_0 inv_weak_pulldown_corrected_1/in VSUBS inv_weak_pulldown_corrected_0/vnb
+ comp_clks_0/w_577_332# inv_weak_pulldown_corrected_0/in comp_clks_0/tg_0/clk inv_weak_pulldown_corrected
Xinv_weak_pulldown_corrected_1 comp_clks_0/tg_0/inp VSUBS inv_weak_pulldown_corrected_1/vnb
+ comp_clks_0/w_577_332# inv_weak_pulldown_corrected_1/in comp_clks_0/tg_0/clk inv_weak_pulldown_corrected
Xcomp_clks_0 comp_clks_0/inverter_1/out comp_clks_0/tg_0/inp comp_clks_0/inverter_2/out
+ comp_clks_0/w_577_332# comp_clks_0/tg_0/clk VSUBS comp_clks
.ends

.subckt inv_weak_pullup_corrected inp w_1_458# li_n53_n248# out vpb a_40_n75#
X0 out vpb a_234_496# w_1_458# sky130_fd_pr__pfet_01v8 ad=4.536e+11p pd=3.24e+06u as=3.654e+11p ps=3.1e+06u w=1.26e+06u l=540000u
X1 a_234_496# inp w_1_458# w_1_458# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.78e+11p ps=3.12e+06u w=1.26e+06u l=180000u
X2 out inp a_40_n75# a_40_n75# sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.554e+11p ps=1.58e+06u w=420000u l=180000u
.ends

.subckt phigen comp_clks_0/inverter_2/out inv_weak_pullup_corrected_0/vpb comp_clks_0/tg_0/clk
+ inv_weak_pulldown_corrected_0/vnb w_1197_875# inv_weak_pulldown_corrected_0/in comp_clks_0/inverter_1/out
+ VSUBS
Xinv_weak_pulldown_corrected_0 inv_weak_pullup_corrected_0/inp VSUBS inv_weak_pulldown_corrected_0/vnb
+ w_1197_875# inv_weak_pulldown_corrected_0/in comp_clks_0/tg_0/clk inv_weak_pulldown_corrected
Xinv_weak_pullup_corrected_0 inv_weak_pullup_corrected_0/inp w_1197_875# comp_clks_0/tg_0/clk
+ inv_weak_pullup_corrected_0/out inv_weak_pullup_corrected_0/vpb VSUBS inv_weak_pullup_corrected
Xcomp_clks_0 comp_clks_0/inverter_1/out inv_weak_pullup_corrected_0/out comp_clks_0/inverter_2/out
+ w_1197_875# comp_clks_0/tg_0/clk VSUBS comp_clks
.ends

.subckt comp_clks_stg1 tg_0/inp tg_0/out inverter_0/out inverter_0/w_n204_204# tg_0/clk
+ VSUBS
Xtg_0 tg_0/inp tg_0/out VSUBS tg_0/clk tg
Xinverter_0 inverter_0/w_n204_204# VSUBS inverter_0/out tg_0/inp inverter
.ends

.subckt level_up_shifter_d_a comp_clks_stg1_0/tg_0/inp comp_clks_stg1_0/VSUBS w_1715_1303#
+ comp_clks_stg1_0/inverter_0/w_n204_204# a_1260_620# a_1811_1506# comp_clks_stg1_0/tg_0/clk
Xcomp_clks_stg1_0 comp_clks_stg1_0/tg_0/inp comp_clks_stg1_0/tg_0/out comp_clks_stg1_0/inverter_0/out
+ comp_clks_stg1_0/inverter_0/w_n204_204# comp_clks_stg1_0/tg_0/clk comp_clks_stg1_0/VSUBS
+ comp_clks_stg1
X0 a_1811_1506# comp_clks_stg1_0/inverter_0/out w_1715_1303# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=1.344e+12p pd=1.408e+07u as=1.6839e+12p ps=1.746e+07u w=600000u l=150000u
X1 a_1260_620# comp_clks_stg1_0/inverter_0/out comp_clks_stg1_0/VSUBS comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=1.344e+12p pd=1.408e+07u as=1.6965e+12p ps=1.749e+07u w=600000u l=150000u
X2 a_1260_620# comp_clks_stg1_0/tg_0/out w_1715_1303# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X3 comp_clks_stg1_0/VSUBS comp_clks_stg1_0/tg_0/out a_1811_1506# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X4 w_1715_1303# comp_clks_stg1_0/inverter_0/out a_1811_1506# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X5 a_1260_620# comp_clks_stg1_0/inverter_0/out comp_clks_stg1_0/VSUBS comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X6 w_1715_1303# comp_clks_stg1_0/tg_0/out a_1260_620# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X7 a_1811_1506# comp_clks_stg1_0/tg_0/out comp_clks_stg1_0/VSUBS comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X8 a_1811_1506# comp_clks_stg1_0/inverter_0/out w_1715_1303# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X9 comp_clks_stg1_0/VSUBS comp_clks_stg1_0/inverter_0/out a_1260_620# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X10 w_1715_1303# comp_clks_stg1_0/inverter_0/out a_1811_1506# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X11 a_1260_620# comp_clks_stg1_0/inverter_0/out comp_clks_stg1_0/VSUBS comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X12 comp_clks_stg1_0/VSUBS comp_clks_stg1_0/inverter_0/out a_1260_620# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X13 a_1260_620# comp_clks_stg1_0/tg_0/out w_1715_1303# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X14 a_1811_1506# a_1260_620# w_1715_1303# w_1715_1303# sky130_fd_pr__pfet_01v8 ad=1.26e+11p pd=1.44e+06u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X15 w_1715_1303# comp_clks_stg1_0/tg_0/out a_1260_620# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X16 comp_clks_stg1_0/VSUBS comp_clks_stg1_0/inverter_0/out a_1260_620# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X17 comp_clks_stg1_0/VSUBS comp_clks_stg1_0/tg_0/out a_1811_1506# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X18 a_1260_620# comp_clks_stg1_0/tg_0/out w_1715_1303# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X19 a_1811_1506# comp_clks_stg1_0/tg_0/out comp_clks_stg1_0/VSUBS comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X20 w_1715_1303# comp_clks_stg1_0/inverter_0/out a_1811_1506# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X21 w_1715_1303# comp_clks_stg1_0/tg_0/out a_1260_620# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X22 a_1811_1506# comp_clks_stg1_0/tg_0/out comp_clks_stg1_0/VSUBS comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X23 comp_clks_stg1_0/VSUBS comp_clks_stg1_0/tg_0/out a_1811_1506# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X24 w_1715_1303# a_1811_1506# a_1260_620# w_1715_1303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X25 w_1715_1303# comp_clks_stg1_0/tg_0/out a_1260_620# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X26 a_1811_1506# comp_clks_stg1_0/inverter_0/out w_1715_1303# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X27 comp_clks_stg1_0/VSUBS comp_clks_stg1_0/tg_0/out a_1811_1506# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X28 a_1260_620# comp_clks_stg1_0/inverter_0/out comp_clks_stg1_0/VSUBS comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X29 a_1811_1506# comp_clks_stg1_0/inverter_0/out w_1715_1303# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X30 comp_clks_stg1_0/VSUBS comp_clks_stg1_0/inverter_0/out a_1260_620# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X31 a_1811_1506# comp_clks_stg1_0/tg_0/out comp_clks_stg1_0/VSUBS comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X32 a_1260_620# comp_clks_stg1_0/tg_0/out w_1715_1303# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X33 w_1715_1303# comp_clks_stg1_0/inverter_0/out a_1811_1506# comp_clks_stg1_0/VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
.ends

.subckt filter_clkgen cclk div2 phi2b phi2 phi1b phi1 cclkb_ana cclk_ana vnb vpb vdda
+ vccd GND
Xcclkgen_0 vnb cclkb_ana vdda vnb cclkgen_0/inv_weak_pulldown_corrected_0/in vdda
+ cclk_ana GND cclkgen
Xphigen_0 phi2b vpb vdda vnb vdda phigen_0/inv_weak_pulldown_corrected_0/in phi2 GND
+ phigen
Xphigen_1 phi1b vpb vdda vnb vdda phigen_1/inv_weak_pulldown_corrected_0/in phi1 GND
+ phigen
Xlevel_up_shifter_d_a_0 div2 GND vdda vccd phigen_1/inv_weak_pulldown_corrected_0/in
+ phigen_0/inv_weak_pulldown_corrected_0/in vccd level_up_shifter_d_a
Xlevel_up_shifter_d_a_1 cclk GND vdda vccd level_up_shifter_d_a_1/a_1260_620# cclkgen_0/inv_weak_pulldown_corrected_0/in
+ vccd level_up_shifter_d_a
.ends

.subckt sky130_fd_sc_hd__inv_8 A VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=1.33e+12p pd=1.266e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=7.02e+11p pd=7.36e+06u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt level_shifter_low sky130_fd_sc_hd__inv_8_0/VPB sky130_fd_sc_hd__inv_8_1/VPB
+ sky130_fd_sc_hd__inv_8_1/VNB sky130_fd_sc_hd__inv_8_1/Y sky130_fd_sc_hd__inv_8_0/A
Xsky130_fd_sc_hd__inv_8_0 sky130_fd_sc_hd__inv_8_0/A sky130_fd_sc_hd__inv_8_1/VNB
+ sky130_fd_sc_hd__inv_8_0/VPB sky130_fd_sc_hd__inv_8_1/A sky130_fd_sc_hd__inv_8_1/VNB
+ sky130_fd_sc_hd__inv_8_0/VPB sky130_fd_sc_hd__inv_8
Xsky130_fd_sc_hd__inv_8_1 sky130_fd_sc_hd__inv_8_1/A sky130_fd_sc_hd__inv_8_1/VNB
+ sky130_fd_sc_hd__inv_8_1/VPB sky130_fd_sc_hd__inv_8_1/Y sky130_fd_sc_hd__inv_8_1/VNB
+ sky130_fd_sc_hd__inv_8_1/VPB sky130_fd_sc_hd__inv_8
.ends

.subckt cmos_switch out w_n94_162# phib a_92_10# in phi
X0 out phi in a_92_10# sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1 out phib in w_n94_162# sky130_fd_pr__pfet_01v8 ad=1.281e+11p pd=1.45e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
.ends

.subckt cap_20fF m3_n28_n28# c1_0_0#
X0 c1_0_0# m3_n28_n28# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=4e+06u
.ends

.subckt analog_mux m1_385_1800# cclk a_30_n10# w_n125_328# m1_239_1920# cclkb a_256_n8#
+ vref2 vref1
X0 vref2 cclkb a_30_n10# a_256_n8# sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1 a_30_n10# cclkb vref1 w_n125_328# sky130_fd_pr__pfet_01v8 ad=1.386e+11p pd=1.5e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2 a_30_n10# cclk vref1 a_256_n8# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3 vref2 cclk a_30_n10# w_n125_328# sky130_fd_pr__pfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
.ends

.subckt cap_10_10_edge_x2 m3_n712_n702# c1_n16_n6#
X0 m3_n712_n702# c1_n16_n6# sky130_fd_pr__cap_mim_m3_2 l=1e+07u w=1e+07u
X1 c1_n16_n6# m3_n712_n702# sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
.ends

.subckt cap_10_10_x2 c2_n16_n6# m3_n376_n34# c1_n16_n6#
X0 c2_n16_n6# c1_n16_n6# sky130_fd_pr__cap_mim_m3_2 l=1e+07u w=1e+07u
X1 c1_n16_n6# m3_n376_n34# sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
.ends

.subckt cap_10_10__side_x2 m3_n712_n366# c1_n16_n6#
X0 m3_n712_n366# c1_n16_n6# sky130_fd_pr__cap_mim_m3_2 l=1e+07u w=1e+07u
X1 c1_n16_n6# m3_n712_n366# sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
.ends

.subckt cap_12pF sig vss
Xcap_10_10_edge_x2_1 vss sig cap_10_10_edge_x2
Xcap_10_10_edge_x2_0 vss sig cap_10_10_edge_x2
Xcap_10_10_edge_x2_2 vss sig cap_10_10_edge_x2
Xcap_10_10_x2_0[0|0] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[1|0] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[0|1] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[1|1] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[0|2] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[1|2] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[0|3] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[1|3] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[0|4] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[1|4] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[0|5] vss vss sig cap_10_10_x2
Xcap_10_10_x2_0[1|5] vss vss sig cap_10_10_x2
Xcap_10_10_edge_x2_3 vss sig cap_10_10_edge_x2
Xcap_10_10__side_x2_0[0] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_0[1] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_0[2] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_0[3] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_0[4] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_0[5] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[0] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[1] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[2] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[3] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[4] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[5] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_2 vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_3 vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_5 vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_4 vss sig cap_10_10__side_x2
.ends

.subckt cap_10fF m3_n28_n28# c1_0_0#
X0 c1_0_0# m3_n28_n28# sky130_fd_pr__cap_mim_m3_1 l=3e+06u w=3.4e+06u
.ends

.subckt cap_40fF m3_n28_n28# c1_0_0#
X0 c1_0_0# m3_n28_n28# sky130_fd_pr__cap_mim_m3_1 l=6e+06u w=6.7e+06u
.ends

.subckt cap_10_10_center_x2 m3_n710_n366# c1_n16_n6#
X0 m3_n710_n366# c1_n16_n6# sky130_fd_pr__cap_mim_m3_2 l=1e+07u w=1e+07u
X1 c1_n16_n6# m3_n710_n366# sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
.ends

.subckt cap_10_10_side2_x2 m3_n710_n366# c1_n16_n6#
X0 m3_n710_n366# c1_n16_n6# sky130_fd_pr__cap_mim_m3_2 l=1e+07u w=1e+07u
X1 c1_n16_n6# m3_n710_n366# sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
.ends

.subckt cap_3pF sig ref
Xcap_10_10_center_x2_0[0] ref sig cap_10_10_center_x2
Xcap_10_10_center_x2_0[1] ref sig cap_10_10_center_x2
Xcap_10_10_center_x2_0[2] ref sig cap_10_10_center_x2
Xcap_10_10_center_x2_0[3] ref sig cap_10_10_center_x2
Xcap_10_10_center_x2_0[4] ref sig cap_10_10_center_x2
Xcap_10_10_center_x2_0[5] ref sig cap_10_10_center_x2
Xcap_10_10_side2_x2_0 ref sig cap_10_10_side2_x2
Xcap_10_10_side2_x2_1 ref sig cap_10_10_side2_x2
.ends

.subckt mux a_n45_373# a_n131_79# out2 VDD out1 a_n45_193# GND a_150_79#
X0 a_150_79# a_n45_193# out1 VDD sky130_fd_pr__pfet_01v8 ad=1.827e+11p pd=1.71e+06u as=2.52e+11p ps=2.04e+06u w=420000u l=150000u
X1 a_n131_79# a_n45_193# out2 VDD sky130_fd_pr__pfet_01v8 ad=4.242e+11p pd=3.7e+06u as=2.52e+11p ps=2.04e+06u w=420000u l=150000u
X2 out2 a_n45_193# a_150_79# GND sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.04e+06u as=1.827e+11p ps=1.71e+06u w=420000u l=150000u
X3 out1 a_n45_193# a_n131_79# GND sky130_fd_pr__nfet_01v8 ad=2.52e+11p pd=2.04e+06u as=4.242e+11p ps=3.7e+06u w=420000u l=150000u
X4 a_150_79# a_n45_373# out1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 out2 a_n45_373# a_150_79# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_n131_79# a_n45_373# out2 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 out1 a_n45_373# a_n131_79# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt cap_6pF sig vss
Xcap_10_10_edge_x2_0 vss sig cap_10_10_edge_x2
Xcap_10_10_edge_x2_1 vss sig cap_10_10_edge_x2
Xcap_10_10_edge_x2_2 vss sig cap_10_10_edge_x2
Xcap_10_10_edge_x2_3 vss sig cap_10_10_edge_x2
Xcap_10_10__side_x2_0[0] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_0[1] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_0[2] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_0[3] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_0[4] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_0[5] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[0] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[1] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[2] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[3] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[4] vss sig cap_10_10__side_x2
Xcap_10_10__side_x2_1[5] vss sig cap_10_10__side_x2
.ends

.subckt filter m2_n261_28387# phi2 phi1 m3_n1255_33008# analog_mux_0/cclkb ctrlb analog_mux_0/vref2
+ analog_mux_0/vref1 m3_n1255_33208# mux_0/out2 m2_n649_28654# analog_mux_0/cclk mux_0/out1
+ ctrl m1_21058_32712# cmos_switch_0/in m3_n1255_33408# mux_0/VDD phi1b phi2b m1_20912_32832#
+ cap_3pF_0/sig VSUBS
Xcmos_switch_0 cmos_switch_1/out mux_0/VDD phi1b VSUBS cmos_switch_0/in phi1 cmos_switch
Xcmos_switch_1 cmos_switch_1/out mux_0/VDD phi2b VSUBS cap_12pF_0/sig phi2 cmos_switch
Xcmos_switch_2 cmos_switch_3/out mux_0/VDD phi1b VSUBS cap_12pF_0/sig phi1 cmos_switch
Xcap_20fF_0 VSUBS cmos_switch_3/out cap_20fF
Xcmos_switch_3 cmos_switch_3/out mux_0/VDD phi2b VSUBS cap_6pF_0/sig phi2 cmos_switch
Xcmos_switch_4 cmos_switch_5/out mux_0/VDD phi1b VSUBS cap_6pF_0/sig phi1 cmos_switch
Xanalog_mux_0 m1_21058_32712# analog_mux_0/cclk cap_3pF_0/ref mux_0/VDD m1_20912_32832#
+ analog_mux_0/cclkb VSUBS analog_mux_0/vref2 analog_mux_0/vref1 analog_mux
Xcmos_switch_5 cmos_switch_5/out mux_0/VDD phi2b VSUBS cap_3pF_0/sig phi2 cmos_switch
Xcap_12pF_0 cap_12pF_0/sig VSUBS cap_12pF
Xcmos_switch_6 cmos_switch_7/out mux_0/VDD phi1b VSUBS cmos_switch_6/in phi1 cmos_switch
Xcmos_switch_7 cmos_switch_7/out mux_0/VDD phi2b VSUBS cap_12pF_0/sig phi2 cmos_switch
Xcap_10fF_0 VSUBS cmos_switch_5/out cap_10fF
Xcap_10fF_1 VSUBS cmos_switch_7/out cap_10fF
Xcap_40fF_0 VSUBS cmos_switch_1/out cap_40fF
Xcap_3pF_0 cap_3pF_0/sig cap_3pF_0/ref cap_3pF
Xmux_0 ctrlb m2_n261_28387# mux_0/out2 mux_0/VDD mux_0/out1 ctrl VSUBS m2_n649_28654#
+ mux
Xcap_6pF_0 cap_6pF_0/sig VSUBS cap_6pF
.ends

.subckt inv_LV A w_987_322# a_1138_96# a_1032_466# a_1136_466# VSUBS
X0 a_1136_466# A a_1032_466# w_987_322# sky130_fd_pr__pfet_01v8 ad=1.554e+11p pd=1.58e+06u as=1.554e+11p ps=1.58e+06u w=420000u l=150000u
X1 a_1138_96# A a_1032_466# VSUBS sky130_fd_pr__nfet_01v8 ad=1.554e+11p pd=1.58e+06u as=1.554e+11p ps=1.58e+06u w=420000u l=150000u
.ends

.subckt comparator a_10_n824# inp inv_LV_7/VSUBS a_n618_473# a_n524_n144# a_280_n337#
+ w_n359_n11#
Xinv_LV_2 inv_LV_2/A w_n359_n11# inv_LV_7/VSUBS inv_LV_3/A w_n359_n11# inv_LV_7/VSUBS
+ inv_LV
Xinv_LV_3 inv_LV_3/A w_n359_n11# inv_LV_7/VSUBS li_1873_504# w_n359_n11# inv_LV_7/VSUBS
+ inv_LV
Xinv_LV_4 inv_LV_4/A w_n359_n11# inv_LV_7/VSUBS inv_LV_4/a_1032_466# w_n359_n11# inv_LV_7/VSUBS
+ inv_LV
Xinv_LV_5 inv_LV_5/A w_n359_n11# inv_LV_7/VSUBS inv_LV_4/A w_n359_n11# inv_LV_7/VSUBS
+ inv_LV
Xinv_LV_6 inv_LV_6/A w_n359_n11# inv_LV_7/VSUBS inv_LV_5/A w_n359_n11# inv_LV_7/VSUBS
+ inv_LV
Xinv_LV_7 low w_n359_n11# inv_LV_7/VSUBS inv_LV_6/A w_n359_n11# inv_LV_7/VSUBS inv_LV
Xinv_LV_0 low w_n359_n11# inv_LV_7/VSUBS inv_LV_1/A w_n359_n11# inv_LV_7/VSUBS inv_LV
Xinv_LV_1 inv_LV_1/A w_n359_n11# inv_LV_7/VSUBS inv_LV_2/A w_n359_n11# inv_LV_7/VSUBS
+ inv_LV
X0 tail a_10_n824# inv_LV_7/VSUBS inv_LV_7/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.197e+11p pd=1.41e+06u as=1.9131e+12p ps=2.003e+07u w=420000u l=2e+06u
X1 inv_LV_7/VSUBS a_n618_473# low inv_LV_7/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.394e+11p ps=2.82e+06u w=420000u l=2e+06u
X2 low FP pfetw w_n359_n11# sky130_fd_pr__pfet_01v8 ad=5.9e+11p pd=5.18e+06u as=2.815e+11p ps=2.65e+06u w=1e+06u l=150000u
X3 inv_LV_7/VSUBS a_n618_473# low inv_LV_7/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=2e+06u
X4 pfetw low w_n359_n11# w_n359_n11# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.5981e+12p ps=1.685e+07u w=420000u l=150000u
X5 FN a_10_n824# w_n359_n11# w_n359_n11# sky130_fd_pr__pfet_01v8 ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X6 FP inp tail inv_LV_7/VSUBS sky130_fd_pr__nfet_03v3_nvt ad=2.85e+11p pd=2.57e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=500000u
X7 pfete FN low w_n359_n11# sky130_fd_pr__pfet_01v8 ad=2.815e+11p pd=2.65e+06u as=0p ps=0u w=1e+06u l=150000u
X8 w_n359_n11# low pfete w_n359_n11# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 low low inv_LV_7/VSUBS inv_LV_7/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=2e+06u
X10 FN a_280_n337# tail inv_LV_7/VSUBS sky130_fd_pr__nfet_03v3_nvt ad=2.85e+11p pd=2.57e+06u as=0p ps=0u w=1e+06u l=500000u
X11 low low inv_LV_7/VSUBS inv_LV_7/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=2e+06u
X12 w_n359_n11# a_10_n824# FP w_n359_n11# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
.ends

.subckt filter_p_m
Xfilter_clkgen_0 filter_clkgen_0/cclk filter_clkgen_0/div2 filter_1/phi2b filter_1/phi2
+ filter_1/phi1b filter_1/phi1 filter_clkgen_0/cclkb_ana filter_clkgen_0/cclk_ana
+ filter_clkgen_0/vnb filter_clkgen_0/vpb filter_clkgen_0/vdda filter_clkgen_0/vccd
+ filter_1/VSUBS filter_clkgen
Xlevel_shifter_low_0 filter_clkgen_0/vdda filter_clkgen_0/vccd filter_1/VSUBS level_shifter_low_0/sky130_fd_sc_hd__inv_8_1/Y
+ filter_1/phi1 level_shifter_low
Xlevel_shifter_low_1 filter_clkgen_0/vdda filter_clkgen_0/vccd filter_1/VSUBS level_shifter_low_1/sky130_fd_sc_hd__inv_8_1/Y
+ filter_1/phi1b level_shifter_low
Xfilter_0 filter_1/m2_n261_28387# filter_1/phi2 filter_1/phi1 filter_1/analog_mux_0/vref1
+ filter_clkgen_0/cclkb_ana filter_1/ctrlb filter_1/analog_mux_0/vref1 filter_1/analog_mux_0/vref2
+ filter_1/analog_mux_0/vref2 filter_0/mux_0/out2 filter_1/m2_n649_28654# filter_clkgen_0/cclk_ana
+ filter_0/mux_0/out1 filter_1/ctrl filter_1/ctrl filter_0/mux_0/out1 filter_clkgen_0/vccd
+ filter_clkgen_0/vdda filter_1/phi1b filter_1/phi2b filter_1/ctrlb comparator_0/inp
+ filter_1/VSUBS filter
Xfilter_1 filter_1/m2_n261_28387# filter_1/phi2 filter_1/phi1 filter_1/analog_mux_0/vref1
+ filter_clkgen_0/cclkb_ana filter_1/ctrlb filter_1/analog_mux_0/vref2 filter_1/analog_mux_0/vref1
+ filter_1/analog_mux_0/vref2 filter_1/mux_0/out2 filter_1/m2_n649_28654# filter_clkgen_0/cclk_ana
+ filter_1/mux_0/out1 filter_1/ctrl filter_1/ctrl filter_1/mux_0/out2 filter_clkgen_0/vccd
+ filter_clkgen_0/vdda filter_1/phi1b filter_1/phi2b filter_1/ctrlb filter_1/cap_3pF_0/sig
+ filter_1/VSUBS filter
Xcomparator_0 level_shifter_low_0/sky130_fd_sc_hd__inv_8_1/Y comparator_0/inp filter_1/VSUBS
+ level_shifter_low_1/sky130_fd_sc_hd__inv_8_1/Y filter_1/VSUBS filter_1/cap_3pF_0/sig
+ filter_clkgen_0/vccd comparator
Xlevel_up_shifter_d_a_0 fb1 filter_1/VSUBS filter_clkgen_0/vdda filter_clkgen_0/vccd
+ fb fb_inv filter_clkgen_0/vccd level_up_shifter_d_a
.ends

