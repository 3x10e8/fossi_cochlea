VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital_unison
  CLASS BLOCK ;
  FOREIGN digital_unison ;
  ORIGIN 0.000 0.000 ;
  SIZE 960.000 BY 100.000 ;
  PIN cclk_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 96.000 143.890 100.000 ;
    END
  END cclk_I[0]
  PIN cclk_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 96.000 381.250 100.000 ;
    END
  END cclk_I[1]
  PIN cclk_I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 96.000 618.610 100.000 ;
    END
  END cclk_I[2]
  PIN cclk_I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 96.000 855.970 100.000 ;
    END
  END cclk_I[3]
  PIN cclk_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END cclk_Q[0]
  PIN cclk_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END cclk_Q[1]
  PIN cclk_Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END cclk_Q[2]
  PIN cclk_Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 0.000 855.970 4.000 ;
    END
  END cclk_Q[3]
  PIN clk_master
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END clk_master
  PIN clkdiv2_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 96.000 104.330 100.000 ;
    END
  END clkdiv2_I[0]
  PIN clkdiv2_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 96.000 341.690 100.000 ;
    END
  END clkdiv2_I[1]
  PIN clkdiv2_I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.770 96.000 579.050 100.000 ;
    END
  END clkdiv2_I[2]
  PIN clkdiv2_I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.130 96.000 816.410 100.000 ;
    END
  END clkdiv2_I[3]
  PIN clkdiv2_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END clkdiv2_Q[0]
  PIN clkdiv2_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END clkdiv2_Q[1]
  PIN clkdiv2_Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.770 0.000 579.050 4.000 ;
    END
  END clkdiv2_Q[2]
  PIN clkdiv2_Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.130 0.000 816.410 4.000 ;
    END
  END clkdiv2_Q[3]
  PIN comp_high_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 96.000 223.010 100.000 ;
    END
  END comp_high_I[0]
  PIN comp_high_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 96.000 460.370 100.000 ;
    END
  END comp_high_I[1]
  PIN comp_high_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 96.000 697.730 100.000 ;
    END
  END comp_high_I[2]
  PIN comp_high_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.810 96.000 935.090 100.000 ;
    END
  END comp_high_I[3]
  PIN comp_high_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END comp_high_Q[0]
  PIN comp_high_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 0.000 460.370 4.000 ;
    END
  END comp_high_Q[1]
  PIN comp_high_Q[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END comp_high_Q[2]
  PIN comp_high_Q[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.810 0.000 935.090 4.000 ;
    END
  END comp_high_Q[3]
  PIN cos_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 96.000 25.210 100.000 ;
    END
  END cos_out[0]
  PIN cos_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 96.000 262.570 100.000 ;
    END
  END cos_out[1]
  PIN cos_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 96.000 499.930 100.000 ;
    END
  END cos_out[2]
  PIN cos_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 96.000 737.290 100.000 ;
    END
  END cos_out[3]
  PIN fb1_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 96.000 64.770 100.000 ;
    END
  END fb1_I[0]
  PIN fb1_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 96.000 302.130 100.000 ;
    END
  END fb1_I[1]
  PIN fb1_I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 96.000 539.490 100.000 ;
    END
  END fb1_I[2]
  PIN fb1_I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 96.000 776.850 100.000 ;
    END
  END fb1_I[3]
  PIN fb1_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END fb1_Q[0]
  PIN fb1_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END fb1_Q[1]
  PIN fb1_Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 0.000 539.490 4.000 ;
    END
  END fb1_Q[2]
  PIN fb1_Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 0.000 776.850 4.000 ;
    END
  END fb1_Q[3]
  PIN phi1b_dig_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 96.000 183.450 100.000 ;
    END
  END phi1b_dig_I[0]
  PIN phi1b_dig_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 96.000 420.810 100.000 ;
    END
  END phi1b_dig_I[1]
  PIN phi1b_dig_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 96.000 658.170 100.000 ;
    END
  END phi1b_dig_I[2]
  PIN phi1b_dig_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 96.000 895.530 100.000 ;
    END
  END phi1b_dig_I[3]
  PIN phi1b_dig_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END phi1b_dig_Q[0]
  PIN phi1b_dig_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END phi1b_dig_Q[1]
  PIN phi1b_dig_Q[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END phi1b_dig_Q[2]
  PIN phi1b_dig_Q[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 0.000 895.530 4.000 ;
    END
  END phi1b_dig_Q[3]
  PIN read_out_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 956.000 86.400 960.000 87.000 ;
    END
  END read_out_I[0]
  PIN read_out_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 956.000 61.920 960.000 62.520 ;
    END
  END read_out_I[1]
  PIN read_out_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 956.000 37.440 960.000 38.040 ;
    END
  END read_out_Q[0]
  PIN read_out_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 956.000 12.960 960.000 13.560 ;
    END
  END read_out_Q[1]
  PIN rstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END rstb
  PIN sin_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END sin_out[0]
  PIN sin_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END sin_out[1]
  PIN sin_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END sin_out[2]
  PIN sin_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 4.000 ;
    END
  END sin_out[3]
  PIN ud_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END ud_en
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 123.285 10.640 124.885 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 360.415 10.640 362.015 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 597.545 10.640 599.145 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 834.675 10.640 836.275 87.280 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 241.850 10.640 243.450 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 478.980 10.640 480.580 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 716.110 10.640 717.710 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 953.240 10.640 954.840 87.280 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 954.040 87.125 ;
      LAYER met1 ;
        RECT 5.520 7.860 954.840 88.360 ;
      LAYER met2 ;
        RECT 7.910 95.720 24.650 96.290 ;
        RECT 25.490 95.720 64.210 96.290 ;
        RECT 65.050 95.720 103.770 96.290 ;
        RECT 104.610 95.720 143.330 96.290 ;
        RECT 144.170 95.720 182.890 96.290 ;
        RECT 183.730 95.720 222.450 96.290 ;
        RECT 223.290 95.720 262.010 96.290 ;
        RECT 262.850 95.720 301.570 96.290 ;
        RECT 302.410 95.720 341.130 96.290 ;
        RECT 341.970 95.720 380.690 96.290 ;
        RECT 381.530 95.720 420.250 96.290 ;
        RECT 421.090 95.720 459.810 96.290 ;
        RECT 460.650 95.720 499.370 96.290 ;
        RECT 500.210 95.720 538.930 96.290 ;
        RECT 539.770 95.720 578.490 96.290 ;
        RECT 579.330 95.720 618.050 96.290 ;
        RECT 618.890 95.720 657.610 96.290 ;
        RECT 658.450 95.720 697.170 96.290 ;
        RECT 698.010 95.720 736.730 96.290 ;
        RECT 737.570 95.720 776.290 96.290 ;
        RECT 777.130 95.720 815.850 96.290 ;
        RECT 816.690 95.720 855.410 96.290 ;
        RECT 856.250 95.720 894.970 96.290 ;
        RECT 895.810 95.720 934.530 96.290 ;
        RECT 935.370 95.720 954.810 96.290 ;
        RECT 7.910 4.280 954.810 95.720 ;
        RECT 7.910 4.000 24.650 4.280 ;
        RECT 25.490 4.000 64.210 4.280 ;
        RECT 65.050 4.000 103.770 4.280 ;
        RECT 104.610 4.000 143.330 4.280 ;
        RECT 144.170 4.000 182.890 4.280 ;
        RECT 183.730 4.000 222.450 4.280 ;
        RECT 223.290 4.000 262.010 4.280 ;
        RECT 262.850 4.000 301.570 4.280 ;
        RECT 302.410 4.000 341.130 4.280 ;
        RECT 341.970 4.000 380.690 4.280 ;
        RECT 381.530 4.000 420.250 4.280 ;
        RECT 421.090 4.000 459.810 4.280 ;
        RECT 460.650 4.000 499.370 4.280 ;
        RECT 500.210 4.000 538.930 4.280 ;
        RECT 539.770 4.000 578.490 4.280 ;
        RECT 579.330 4.000 618.050 4.280 ;
        RECT 618.890 4.000 657.610 4.280 ;
        RECT 658.450 4.000 697.170 4.280 ;
        RECT 698.010 4.000 736.730 4.280 ;
        RECT 737.570 4.000 776.290 4.280 ;
        RECT 777.130 4.000 815.850 4.280 ;
        RECT 816.690 4.000 855.410 4.280 ;
        RECT 856.250 4.000 894.970 4.280 ;
        RECT 895.810 4.000 934.530 4.280 ;
        RECT 935.370 4.000 954.810 4.280 ;
      LAYER met3 ;
        RECT 4.000 86.000 955.600 87.205 ;
        RECT 4.000 84.000 956.000 86.000 ;
        RECT 4.400 82.600 956.000 84.000 ;
        RECT 4.000 62.920 956.000 82.600 ;
        RECT 4.000 61.520 955.600 62.920 ;
        RECT 4.000 50.680 956.000 61.520 ;
        RECT 4.400 49.280 956.000 50.680 ;
        RECT 4.000 38.440 956.000 49.280 ;
        RECT 4.000 37.040 955.600 38.440 ;
        RECT 4.000 17.360 956.000 37.040 ;
        RECT 4.400 15.960 956.000 17.360 ;
        RECT 4.000 13.960 956.000 15.960 ;
        RECT 4.000 12.560 955.600 13.960 ;
        RECT 4.000 9.695 956.000 12.560 ;
      LAYER met4 ;
        RECT 257.895 11.055 360.015 66.465 ;
        RECT 362.415 11.055 413.705 66.465 ;
  END
END digital_unison
END LIBRARY

