VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital_unison
  CLASS BLOCK ;
  FOREIGN digital_unison ;
  ORIGIN 0.000 0.000 ;
  SIZE 2040.000 BY 120.000 ;
  PIN cclk_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 116.000 67.990 120.000 ;
    END
  END cclk_I[0]
  PIN cclk_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 116.000 321.910 120.000 ;
    END
  END cclk_I[1]
  PIN cclk_I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 116.000 575.830 120.000 ;
    END
  END cclk_I[2]
  PIN cclk_I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 116.000 829.750 120.000 ;
    END
  END cclk_I[3]
  PIN cclk_I[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.390 116.000 1083.670 120.000 ;
    END
  END cclk_I[4]
  PIN cclk_I[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.310 116.000 1337.590 120.000 ;
    END
  END cclk_I[5]
  PIN cclk_I[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1591.230 116.000 1591.510 120.000 ;
    END
  END cclk_I[6]
  PIN cclk_I[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.150 116.000 1845.430 120.000 ;
    END
  END cclk_I[7]
  PIN cclk_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END cclk_Q[0]
  PIN cclk_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END cclk_Q[1]
  PIN cclk_Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 0.000 575.830 4.000 ;
    END
  END cclk_Q[2]
  PIN cclk_Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 0.000 829.750 4.000 ;
    END
  END cclk_Q[3]
  PIN cclk_Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.390 0.000 1083.670 4.000 ;
    END
  END cclk_Q[4]
  PIN cclk_Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.310 0.000 1337.590 4.000 ;
    END
  END cclk_Q[5]
  PIN cclk_Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1591.230 0.000 1591.510 4.000 ;
    END
  END cclk_Q[6]
  PIN cclk_Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.150 0.000 1845.430 4.000 ;
    END
  END cclk_Q[7]
  PIN clk_master
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END clk_master
  PIN clkdiv2_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 116.000 110.310 120.000 ;
    END
  END clkdiv2_I[0]
  PIN clkdiv2_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 116.000 364.230 120.000 ;
    END
  END clkdiv2_I[1]
  PIN clkdiv2_I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 116.000 618.150 120.000 ;
    END
  END clkdiv2_I[2]
  PIN clkdiv2_I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 116.000 872.070 120.000 ;
    END
  END clkdiv2_I[3]
  PIN clkdiv2_I[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.710 116.000 1125.990 120.000 ;
    END
  END clkdiv2_I[4]
  PIN clkdiv2_I[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.630 116.000 1379.910 120.000 ;
    END
  END clkdiv2_I[5]
  PIN clkdiv2_I[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.550 116.000 1633.830 120.000 ;
    END
  END clkdiv2_I[6]
  PIN clkdiv2_I[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.470 116.000 1887.750 120.000 ;
    END
  END clkdiv2_I[7]
  PIN clkdiv2_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END clkdiv2_Q[0]
  PIN clkdiv2_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END clkdiv2_Q[1]
  PIN clkdiv2_Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 0.000 618.150 4.000 ;
    END
  END clkdiv2_Q[2]
  PIN clkdiv2_Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 0.000 872.070 4.000 ;
    END
  END clkdiv2_Q[3]
  PIN clkdiv2_Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.710 0.000 1125.990 4.000 ;
    END
  END clkdiv2_Q[4]
  PIN clkdiv2_Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.630 0.000 1379.910 4.000 ;
    END
  END clkdiv2_Q[5]
  PIN clkdiv2_Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.550 0.000 1633.830 4.000 ;
    END
  END clkdiv2_Q[6]
  PIN clkdiv2_Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.470 0.000 1887.750 4.000 ;
    END
  END clkdiv2_Q[7]
  PIN comp_high_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 116.000 152.630 120.000 ;
    END
  END comp_high_I[0]
  PIN comp_high_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 116.000 406.550 120.000 ;
    END
  END comp_high_I[1]
  PIN comp_high_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 116.000 660.470 120.000 ;
    END
  END comp_high_I[2]
  PIN comp_high_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.110 116.000 914.390 120.000 ;
    END
  END comp_high_I[3]
  PIN comp_high_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.030 116.000 1168.310 120.000 ;
    END
  END comp_high_I[4]
  PIN comp_high_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.950 116.000 1422.230 120.000 ;
    END
  END comp_high_I[5]
  PIN comp_high_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.870 116.000 1676.150 120.000 ;
    END
  END comp_high_I[6]
  PIN comp_high_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.790 116.000 1930.070 120.000 ;
    END
  END comp_high_I[7]
  PIN comp_high_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END comp_high_Q[0]
  PIN comp_high_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END comp_high_Q[1]
  PIN comp_high_Q[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END comp_high_Q[2]
  PIN comp_high_Q[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.110 0.000 914.390 4.000 ;
    END
  END comp_high_Q[3]
  PIN comp_high_Q[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.030 0.000 1168.310 4.000 ;
    END
  END comp_high_Q[4]
  PIN comp_high_Q[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.950 0.000 1422.230 4.000 ;
    END
  END comp_high_Q[5]
  PIN comp_high_Q[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.870 0.000 1676.150 4.000 ;
    END
  END comp_high_Q[6]
  PIN comp_high_Q[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.790 0.000 1930.070 4.000 ;
    END
  END comp_high_Q[7]
  PIN cos_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 116.000 237.270 120.000 ;
    END
  END cos_out[0]
  PIN cos_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 116.000 491.190 120.000 ;
    END
  END cos_out[1]
  PIN cos_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830 116.000 745.110 120.000 ;
    END
  END cos_out[2]
  PIN cos_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 116.000 999.030 120.000 ;
    END
  END cos_out[3]
  PIN cos_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 116.000 1252.950 120.000 ;
    END
  END cos_out[4]
  PIN cos_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.590 116.000 1506.870 120.000 ;
    END
  END cos_out[5]
  PIN cos_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.510 116.000 1760.790 120.000 ;
    END
  END cos_out[6]
  PIN cos_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2014.430 116.000 2014.710 120.000 ;
    END
  END cos_out[7]
  PIN fb1_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 116.000 25.670 120.000 ;
    END
  END fb1_I[0]
  PIN fb1_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 116.000 279.590 120.000 ;
    END
  END fb1_I[1]
  PIN fb1_I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 116.000 533.510 120.000 ;
    END
  END fb1_I[2]
  PIN fb1_I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 116.000 787.430 120.000 ;
    END
  END fb1_I[3]
  PIN fb1_I[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.070 116.000 1041.350 120.000 ;
    END
  END fb1_I[4]
  PIN fb1_I[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.990 116.000 1295.270 120.000 ;
    END
  END fb1_I[5]
  PIN fb1_I[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.910 116.000 1549.190 120.000 ;
    END
  END fb1_I[6]
  PIN fb1_I[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1802.830 116.000 1803.110 120.000 ;
    END
  END fb1_I[7]
  PIN fb1_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END fb1_Q[0]
  PIN fb1_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END fb1_Q[1]
  PIN fb1_Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 0.000 533.510 4.000 ;
    END
  END fb1_Q[2]
  PIN fb1_Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 0.000 787.430 4.000 ;
    END
  END fb1_Q[3]
  PIN fb1_Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.070 0.000 1041.350 4.000 ;
    END
  END fb1_Q[4]
  PIN fb1_Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.990 0.000 1295.270 4.000 ;
    END
  END fb1_Q[5]
  PIN fb1_Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.910 0.000 1549.190 4.000 ;
    END
  END fb1_Q[6]
  PIN fb1_Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1802.830 0.000 1803.110 4.000 ;
    END
  END fb1_Q[7]
  PIN phi1b_dig_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 116.000 194.950 120.000 ;
    END
  END phi1b_dig_I[0]
  PIN phi1b_dig_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 116.000 448.870 120.000 ;
    END
  END phi1b_dig_I[1]
  PIN phi1b_dig_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 116.000 702.790 120.000 ;
    END
  END phi1b_dig_I[2]
  PIN phi1b_dig_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 116.000 956.710 120.000 ;
    END
  END phi1b_dig_I[3]
  PIN phi1b_dig_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.350 116.000 1210.630 120.000 ;
    END
  END phi1b_dig_I[4]
  PIN phi1b_dig_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1464.270 116.000 1464.550 120.000 ;
    END
  END phi1b_dig_I[5]
  PIN phi1b_dig_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.190 116.000 1718.470 120.000 ;
    END
  END phi1b_dig_I[6]
  PIN phi1b_dig_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.110 116.000 1972.390 120.000 ;
    END
  END phi1b_dig_I[7]
  PIN phi1b_dig_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END phi1b_dig_Q[0]
  PIN phi1b_dig_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 4.000 ;
    END
  END phi1b_dig_Q[1]
  PIN phi1b_dig_Q[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END phi1b_dig_Q[2]
  PIN phi1b_dig_Q[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 0.000 956.710 4.000 ;
    END
  END phi1b_dig_Q[3]
  PIN phi1b_dig_Q[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.350 0.000 1210.630 4.000 ;
    END
  END phi1b_dig_Q[4]
  PIN phi1b_dig_Q[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1464.270 0.000 1464.550 4.000 ;
    END
  END phi1b_dig_Q[5]
  PIN phi1b_dig_Q[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.190 0.000 1718.470 4.000 ;
    END
  END phi1b_dig_Q[6]
  PIN phi1b_dig_Q[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.110 0.000 1972.390 4.000 ;
    END
  END phi1b_dig_Q[7]
  PIN read_out_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END read_out_I[0]
  PIN read_out_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END read_out_I[1]
  PIN read_out_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END read_out_Q[0]
  PIN read_out_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END read_out_Q[1]
  PIN rstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END rstb
  PIN sin_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END sin_out[0]
  PIN sin_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END sin_out[1]
  PIN sin_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830 0.000 745.110 4.000 ;
    END
  END sin_out[2]
  PIN sin_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 0.000 999.030 4.000 ;
    END
  END sin_out[3]
  PIN sin_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 0.000 1252.950 4.000 ;
    END
  END sin_out[4]
  PIN sin_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.590 0.000 1506.870 4.000 ;
    END
  END sin_out[5]
  PIN sin_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.510 0.000 1760.790 4.000 ;
    END
  END sin_out[6]
  PIN sin_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2014.430 0.000 2014.710 4.000 ;
    END
  END sin_out[7]
  PIN ud_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END ud_en
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 258.295 10.640 259.895 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.445 10.640 767.045 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1272.595 10.640 1274.195 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1779.745 10.640 1781.345 109.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 511.870 10.640 513.470 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.020 10.640 1020.620 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1526.170 10.640 1527.770 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2033.320 10.640 2034.920 109.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2034.120 108.885 ;
      LAYER met1 ;
        RECT 5.520 7.180 2034.920 111.480 ;
      LAYER met2 ;
        RECT 7.910 115.720 25.110 116.690 ;
        RECT 25.950 115.720 67.430 116.690 ;
        RECT 68.270 115.720 109.750 116.690 ;
        RECT 110.590 115.720 152.070 116.690 ;
        RECT 152.910 115.720 194.390 116.690 ;
        RECT 195.230 115.720 236.710 116.690 ;
        RECT 237.550 115.720 279.030 116.690 ;
        RECT 279.870 115.720 321.350 116.690 ;
        RECT 322.190 115.720 363.670 116.690 ;
        RECT 364.510 115.720 405.990 116.690 ;
        RECT 406.830 115.720 448.310 116.690 ;
        RECT 449.150 115.720 490.630 116.690 ;
        RECT 491.470 115.720 532.950 116.690 ;
        RECT 533.790 115.720 575.270 116.690 ;
        RECT 576.110 115.720 617.590 116.690 ;
        RECT 618.430 115.720 659.910 116.690 ;
        RECT 660.750 115.720 702.230 116.690 ;
        RECT 703.070 115.720 744.550 116.690 ;
        RECT 745.390 115.720 786.870 116.690 ;
        RECT 787.710 115.720 829.190 116.690 ;
        RECT 830.030 115.720 871.510 116.690 ;
        RECT 872.350 115.720 913.830 116.690 ;
        RECT 914.670 115.720 956.150 116.690 ;
        RECT 956.990 115.720 998.470 116.690 ;
        RECT 999.310 115.720 1040.790 116.690 ;
        RECT 1041.630 115.720 1083.110 116.690 ;
        RECT 1083.950 115.720 1125.430 116.690 ;
        RECT 1126.270 115.720 1167.750 116.690 ;
        RECT 1168.590 115.720 1210.070 116.690 ;
        RECT 1210.910 115.720 1252.390 116.690 ;
        RECT 1253.230 115.720 1294.710 116.690 ;
        RECT 1295.550 115.720 1337.030 116.690 ;
        RECT 1337.870 115.720 1379.350 116.690 ;
        RECT 1380.190 115.720 1421.670 116.690 ;
        RECT 1422.510 115.720 1463.990 116.690 ;
        RECT 1464.830 115.720 1506.310 116.690 ;
        RECT 1507.150 115.720 1548.630 116.690 ;
        RECT 1549.470 115.720 1590.950 116.690 ;
        RECT 1591.790 115.720 1633.270 116.690 ;
        RECT 1634.110 115.720 1675.590 116.690 ;
        RECT 1676.430 115.720 1717.910 116.690 ;
        RECT 1718.750 115.720 1760.230 116.690 ;
        RECT 1761.070 115.720 1802.550 116.690 ;
        RECT 1803.390 115.720 1844.870 116.690 ;
        RECT 1845.710 115.720 1887.190 116.690 ;
        RECT 1888.030 115.720 1929.510 116.690 ;
        RECT 1930.350 115.720 1971.830 116.690 ;
        RECT 1972.670 115.720 2014.150 116.690 ;
        RECT 2014.990 115.720 2034.890 116.690 ;
        RECT 7.910 4.280 2034.890 115.720 ;
        RECT 7.910 3.670 25.110 4.280 ;
        RECT 25.950 3.670 67.430 4.280 ;
        RECT 68.270 3.670 109.750 4.280 ;
        RECT 110.590 3.670 152.070 4.280 ;
        RECT 152.910 3.670 194.390 4.280 ;
        RECT 195.230 3.670 236.710 4.280 ;
        RECT 237.550 3.670 279.030 4.280 ;
        RECT 279.870 3.670 321.350 4.280 ;
        RECT 322.190 3.670 363.670 4.280 ;
        RECT 364.510 3.670 405.990 4.280 ;
        RECT 406.830 3.670 448.310 4.280 ;
        RECT 449.150 3.670 490.630 4.280 ;
        RECT 491.470 3.670 532.950 4.280 ;
        RECT 533.790 3.670 575.270 4.280 ;
        RECT 576.110 3.670 617.590 4.280 ;
        RECT 618.430 3.670 659.910 4.280 ;
        RECT 660.750 3.670 702.230 4.280 ;
        RECT 703.070 3.670 744.550 4.280 ;
        RECT 745.390 3.670 786.870 4.280 ;
        RECT 787.710 3.670 829.190 4.280 ;
        RECT 830.030 3.670 871.510 4.280 ;
        RECT 872.350 3.670 913.830 4.280 ;
        RECT 914.670 3.670 956.150 4.280 ;
        RECT 956.990 3.670 998.470 4.280 ;
        RECT 999.310 3.670 1040.790 4.280 ;
        RECT 1041.630 3.670 1083.110 4.280 ;
        RECT 1083.950 3.670 1125.430 4.280 ;
        RECT 1126.270 3.670 1167.750 4.280 ;
        RECT 1168.590 3.670 1210.070 4.280 ;
        RECT 1210.910 3.670 1252.390 4.280 ;
        RECT 1253.230 3.670 1294.710 4.280 ;
        RECT 1295.550 3.670 1337.030 4.280 ;
        RECT 1337.870 3.670 1379.350 4.280 ;
        RECT 1380.190 3.670 1421.670 4.280 ;
        RECT 1422.510 3.670 1463.990 4.280 ;
        RECT 1464.830 3.670 1506.310 4.280 ;
        RECT 1507.150 3.670 1548.630 4.280 ;
        RECT 1549.470 3.670 1590.950 4.280 ;
        RECT 1591.790 3.670 1633.270 4.280 ;
        RECT 1634.110 3.670 1675.590 4.280 ;
        RECT 1676.430 3.670 1717.910 4.280 ;
        RECT 1718.750 3.670 1760.230 4.280 ;
        RECT 1761.070 3.670 1802.550 4.280 ;
        RECT 1803.390 3.670 1844.870 4.280 ;
        RECT 1845.710 3.670 1887.190 4.280 ;
        RECT 1888.030 3.670 1929.510 4.280 ;
        RECT 1930.350 3.670 1971.830 4.280 ;
        RECT 1972.670 3.670 2014.150 4.280 ;
        RECT 2014.990 3.670 2034.890 4.280 ;
      LAYER met3 ;
        RECT 4.000 111.200 2034.910 111.345 ;
        RECT 4.400 109.800 2034.910 111.200 ;
        RECT 4.000 94.200 2034.910 109.800 ;
        RECT 4.400 92.800 2034.910 94.200 ;
        RECT 4.000 77.200 2034.910 92.800 ;
        RECT 4.400 75.800 2034.910 77.200 ;
        RECT 4.000 60.200 2034.910 75.800 ;
        RECT 4.400 58.800 2034.910 60.200 ;
        RECT 4.000 43.200 2034.910 58.800 ;
        RECT 4.400 41.800 2034.910 43.200 ;
        RECT 4.000 26.200 2034.910 41.800 ;
        RECT 4.400 24.800 2034.910 26.200 ;
        RECT 4.000 9.200 2034.910 24.800 ;
        RECT 4.400 8.335 2034.910 9.200 ;
      LAYER met4 ;
        RECT 45.375 109.440 2015.425 111.345 ;
        RECT 45.375 12.415 257.895 109.440 ;
        RECT 260.295 12.415 511.470 109.440 ;
        RECT 513.870 12.415 765.045 109.440 ;
        RECT 767.445 12.415 1018.620 109.440 ;
        RECT 1021.020 12.415 1272.195 109.440 ;
        RECT 1274.595 12.415 1525.770 109.440 ;
        RECT 1528.170 12.415 1779.345 109.440 ;
        RECT 1781.745 12.415 2015.425 109.440 ;
  END
END digital_unison
END LIBRARY

