magic
tech sky130A
timestamp 1647792644
<< nwell >>
rect 841 9215 987 9299
rect 1652 9215 1874 9299
rect 2522 9215 2744 9299
rect 3117 9215 3263 9299
rect 8015 9215 8161 9299
rect 8534 9215 8756 9299
rect 9404 9215 9626 9299
rect 10291 9215 10437 9299
rect 841 -1505 987 -1421
rect 1652 -1505 1874 -1421
rect 2522 -1505 2744 -1421
rect 3117 -1505 3263 -1421
rect 8015 -1505 8161 -1421
rect 8534 -1505 8756 -1421
rect 9404 -1505 9626 -1421
rect 10291 -1505 10437 -1421
<< nmos >>
rect 894 9355 909 9397
rect 1705 9355 1720 9397
rect 1781 9355 1796 9397
rect 2575 9355 2590 9397
rect 2651 9355 2666 9397
rect 3170 9355 3185 9397
rect 8093 9355 8108 9397
rect 8612 9355 8627 9397
rect 8688 9355 8703 9397
rect 9482 9355 9497 9397
rect 9558 9355 9573 9397
rect 10369 9355 10384 9397
rect 894 -1603 909 -1561
rect 1705 -1603 1720 -1561
rect 1781 -1603 1796 -1561
rect 2575 -1603 2590 -1561
rect 2651 -1603 2666 -1561
rect 3170 -1603 3185 -1561
rect 8093 -1603 8108 -1561
rect 8612 -1603 8627 -1561
rect 8688 -1603 8703 -1561
rect 9482 -1603 9497 -1561
rect 9558 -1603 9573 -1561
rect 10369 -1603 10384 -1561
<< pmos >>
rect 894 9238 909 9280
rect 1705 9238 1720 9280
rect 1781 9238 1796 9280
rect 2575 9238 2590 9280
rect 2651 9238 2666 9280
rect 3170 9238 3185 9280
rect 8093 9238 8108 9280
rect 8612 9238 8627 9280
rect 8688 9238 8703 9280
rect 9482 9238 9497 9280
rect 9558 9238 9573 9280
rect 10369 9238 10384 9280
rect 894 -1486 909 -1444
rect 1705 -1486 1720 -1444
rect 1781 -1486 1796 -1444
rect 2575 -1486 2590 -1444
rect 2651 -1486 2666 -1444
rect 3170 -1486 3185 -1444
rect 8093 -1486 8108 -1444
rect 8612 -1486 8627 -1444
rect 8688 -1486 8703 -1444
rect 9482 -1486 9497 -1444
rect 9558 -1486 9573 -1444
rect 10369 -1486 10384 -1444
<< ndiff >>
rect 863 9385 894 9397
rect 863 9368 869 9385
rect 886 9368 894 9385
rect 863 9355 894 9368
rect 909 9385 940 9397
rect 909 9368 916 9385
rect 933 9368 940 9385
rect 909 9355 940 9368
rect 1674 9385 1705 9397
rect 1674 9368 1680 9385
rect 1697 9368 1705 9385
rect 1674 9355 1705 9368
rect 1720 9384 1781 9397
rect 1720 9367 1745 9384
rect 1762 9367 1781 9384
rect 1720 9355 1781 9367
rect 1796 9385 1827 9397
rect 1796 9368 1803 9385
rect 1820 9368 1827 9385
rect 1796 9355 1827 9368
rect 2544 9385 2575 9397
rect 2544 9368 2550 9385
rect 2567 9368 2575 9385
rect 2544 9355 2575 9368
rect 2590 9384 2651 9397
rect 2590 9367 2615 9384
rect 2632 9367 2651 9384
rect 2590 9355 2651 9367
rect 2666 9385 2697 9397
rect 2666 9368 2673 9385
rect 2690 9368 2697 9385
rect 2666 9355 2697 9368
rect 3139 9385 3170 9397
rect 3139 9368 3145 9385
rect 3162 9368 3170 9385
rect 3139 9355 3170 9368
rect 3185 9385 3216 9397
rect 3185 9368 3192 9385
rect 3209 9368 3216 9385
rect 3185 9355 3216 9368
rect 8062 9385 8093 9397
rect 8062 9368 8069 9385
rect 8086 9368 8093 9385
rect 8062 9355 8093 9368
rect 8108 9385 8139 9397
rect 8108 9368 8116 9385
rect 8133 9368 8139 9385
rect 8108 9355 8139 9368
rect 8581 9385 8612 9397
rect 8581 9368 8588 9385
rect 8605 9368 8612 9385
rect 8581 9355 8612 9368
rect 8627 9384 8688 9397
rect 8627 9367 8646 9384
rect 8663 9367 8688 9384
rect 8627 9355 8688 9367
rect 8703 9385 8734 9397
rect 8703 9368 8711 9385
rect 8728 9368 8734 9385
rect 8703 9355 8734 9368
rect 9451 9385 9482 9397
rect 9451 9368 9458 9385
rect 9475 9368 9482 9385
rect 9451 9355 9482 9368
rect 9497 9384 9558 9397
rect 9497 9367 9516 9384
rect 9533 9367 9558 9384
rect 9497 9355 9558 9367
rect 9573 9385 9604 9397
rect 9573 9368 9581 9385
rect 9598 9368 9604 9385
rect 9573 9355 9604 9368
rect 10338 9385 10369 9397
rect 10338 9368 10345 9385
rect 10362 9368 10369 9385
rect 10338 9355 10369 9368
rect 10384 9385 10415 9397
rect 10384 9368 10392 9385
rect 10409 9368 10415 9385
rect 10384 9355 10415 9368
rect 863 -1574 894 -1561
rect 863 -1591 869 -1574
rect 886 -1591 894 -1574
rect 863 -1603 894 -1591
rect 909 -1574 940 -1561
rect 909 -1591 916 -1574
rect 933 -1591 940 -1574
rect 909 -1603 940 -1591
rect 1674 -1574 1705 -1561
rect 1674 -1591 1680 -1574
rect 1697 -1591 1705 -1574
rect 1674 -1603 1705 -1591
rect 1720 -1573 1781 -1561
rect 1720 -1590 1745 -1573
rect 1762 -1590 1781 -1573
rect 1720 -1603 1781 -1590
rect 1796 -1574 1827 -1561
rect 1796 -1591 1803 -1574
rect 1820 -1591 1827 -1574
rect 1796 -1603 1827 -1591
rect 2544 -1574 2575 -1561
rect 2544 -1591 2550 -1574
rect 2567 -1591 2575 -1574
rect 2544 -1603 2575 -1591
rect 2590 -1573 2651 -1561
rect 2590 -1590 2615 -1573
rect 2632 -1590 2651 -1573
rect 2590 -1603 2651 -1590
rect 2666 -1574 2697 -1561
rect 2666 -1591 2673 -1574
rect 2690 -1591 2697 -1574
rect 2666 -1603 2697 -1591
rect 3139 -1574 3170 -1561
rect 3139 -1591 3145 -1574
rect 3162 -1591 3170 -1574
rect 3139 -1603 3170 -1591
rect 3185 -1574 3216 -1561
rect 3185 -1591 3192 -1574
rect 3209 -1591 3216 -1574
rect 3185 -1603 3216 -1591
rect 8062 -1574 8093 -1561
rect 8062 -1591 8069 -1574
rect 8086 -1591 8093 -1574
rect 8062 -1603 8093 -1591
rect 8108 -1574 8139 -1561
rect 8108 -1591 8116 -1574
rect 8133 -1591 8139 -1574
rect 8108 -1603 8139 -1591
rect 8581 -1574 8612 -1561
rect 8581 -1591 8588 -1574
rect 8605 -1591 8612 -1574
rect 8581 -1603 8612 -1591
rect 8627 -1573 8688 -1561
rect 8627 -1590 8646 -1573
rect 8663 -1590 8688 -1573
rect 8627 -1603 8688 -1590
rect 8703 -1574 8734 -1561
rect 8703 -1591 8711 -1574
rect 8728 -1591 8734 -1574
rect 8703 -1603 8734 -1591
rect 9451 -1574 9482 -1561
rect 9451 -1591 9458 -1574
rect 9475 -1591 9482 -1574
rect 9451 -1603 9482 -1591
rect 9497 -1573 9558 -1561
rect 9497 -1590 9516 -1573
rect 9533 -1590 9558 -1573
rect 9497 -1603 9558 -1590
rect 9573 -1574 9604 -1561
rect 9573 -1591 9581 -1574
rect 9598 -1591 9604 -1574
rect 9573 -1603 9604 -1591
rect 10338 -1574 10369 -1561
rect 10338 -1591 10345 -1574
rect 10362 -1591 10369 -1574
rect 10338 -1603 10369 -1591
rect 10384 -1574 10415 -1561
rect 10384 -1591 10392 -1574
rect 10409 -1591 10415 -1574
rect 10384 -1603 10415 -1591
<< pdiff >>
rect 863 9267 894 9280
rect 863 9250 869 9267
rect 886 9250 894 9267
rect 863 9238 894 9250
rect 909 9267 940 9280
rect 909 9250 916 9267
rect 933 9250 940 9267
rect 909 9238 940 9250
rect 1674 9267 1705 9280
rect 1674 9250 1680 9267
rect 1697 9250 1705 9267
rect 1674 9238 1705 9250
rect 1720 9270 1781 9280
rect 1720 9253 1741 9270
rect 1758 9253 1781 9270
rect 1720 9238 1781 9253
rect 1796 9267 1827 9280
rect 1796 9250 1803 9267
rect 1820 9250 1827 9267
rect 1796 9238 1827 9250
rect 2544 9267 2575 9280
rect 2544 9250 2550 9267
rect 2567 9250 2575 9267
rect 2544 9238 2575 9250
rect 2590 9270 2651 9280
rect 2590 9253 2611 9270
rect 2628 9253 2651 9270
rect 2590 9238 2651 9253
rect 2666 9267 2697 9280
rect 2666 9250 2673 9267
rect 2690 9250 2697 9267
rect 2666 9238 2697 9250
rect 3139 9267 3170 9280
rect 3139 9250 3145 9267
rect 3162 9250 3170 9267
rect 3139 9238 3170 9250
rect 3185 9267 3216 9280
rect 3185 9250 3192 9267
rect 3209 9250 3216 9267
rect 3185 9238 3216 9250
rect 8062 9267 8093 9280
rect 8062 9250 8069 9267
rect 8086 9250 8093 9267
rect 8062 9238 8093 9250
rect 8108 9267 8139 9280
rect 8108 9250 8116 9267
rect 8133 9250 8139 9267
rect 8108 9238 8139 9250
rect 8581 9267 8612 9280
rect 8581 9250 8588 9267
rect 8605 9250 8612 9267
rect 8581 9238 8612 9250
rect 8627 9270 8688 9280
rect 8627 9253 8650 9270
rect 8667 9253 8688 9270
rect 8627 9238 8688 9253
rect 8703 9267 8734 9280
rect 8703 9250 8711 9267
rect 8728 9250 8734 9267
rect 8703 9238 8734 9250
rect 9451 9267 9482 9280
rect 9451 9250 9458 9267
rect 9475 9250 9482 9267
rect 9451 9238 9482 9250
rect 9497 9270 9558 9280
rect 9497 9253 9520 9270
rect 9537 9253 9558 9270
rect 9497 9238 9558 9253
rect 9573 9267 9604 9280
rect 9573 9250 9581 9267
rect 9598 9250 9604 9267
rect 9573 9238 9604 9250
rect 10338 9267 10369 9280
rect 10338 9250 10345 9267
rect 10362 9250 10369 9267
rect 10338 9238 10369 9250
rect 10384 9267 10415 9280
rect 10384 9250 10392 9267
rect 10409 9250 10415 9267
rect 10384 9238 10415 9250
rect 863 -1456 894 -1444
rect 863 -1473 869 -1456
rect 886 -1473 894 -1456
rect 863 -1486 894 -1473
rect 909 -1456 940 -1444
rect 909 -1473 916 -1456
rect 933 -1473 940 -1456
rect 909 -1486 940 -1473
rect 1674 -1456 1705 -1444
rect 1674 -1473 1680 -1456
rect 1697 -1473 1705 -1456
rect 1674 -1486 1705 -1473
rect 1720 -1459 1781 -1444
rect 1720 -1476 1741 -1459
rect 1758 -1476 1781 -1459
rect 1720 -1486 1781 -1476
rect 1796 -1456 1827 -1444
rect 1796 -1473 1803 -1456
rect 1820 -1473 1827 -1456
rect 1796 -1486 1827 -1473
rect 2544 -1456 2575 -1444
rect 2544 -1473 2550 -1456
rect 2567 -1473 2575 -1456
rect 2544 -1486 2575 -1473
rect 2590 -1459 2651 -1444
rect 2590 -1476 2611 -1459
rect 2628 -1476 2651 -1459
rect 2590 -1486 2651 -1476
rect 2666 -1456 2697 -1444
rect 2666 -1473 2673 -1456
rect 2690 -1473 2697 -1456
rect 2666 -1486 2697 -1473
rect 3139 -1456 3170 -1444
rect 3139 -1473 3145 -1456
rect 3162 -1473 3170 -1456
rect 3139 -1486 3170 -1473
rect 3185 -1456 3216 -1444
rect 3185 -1473 3192 -1456
rect 3209 -1473 3216 -1456
rect 3185 -1486 3216 -1473
rect 8062 -1456 8093 -1444
rect 8062 -1473 8069 -1456
rect 8086 -1473 8093 -1456
rect 8062 -1486 8093 -1473
rect 8108 -1456 8139 -1444
rect 8108 -1473 8116 -1456
rect 8133 -1473 8139 -1456
rect 8108 -1486 8139 -1473
rect 8581 -1456 8612 -1444
rect 8581 -1473 8588 -1456
rect 8605 -1473 8612 -1456
rect 8581 -1486 8612 -1473
rect 8627 -1459 8688 -1444
rect 8627 -1476 8650 -1459
rect 8667 -1476 8688 -1459
rect 8627 -1486 8688 -1476
rect 8703 -1456 8734 -1444
rect 8703 -1473 8711 -1456
rect 8728 -1473 8734 -1456
rect 8703 -1486 8734 -1473
rect 9451 -1456 9482 -1444
rect 9451 -1473 9458 -1456
rect 9475 -1473 9482 -1456
rect 9451 -1486 9482 -1473
rect 9497 -1459 9558 -1444
rect 9497 -1476 9520 -1459
rect 9537 -1476 9558 -1459
rect 9497 -1486 9558 -1476
rect 9573 -1456 9604 -1444
rect 9573 -1473 9581 -1456
rect 9598 -1473 9604 -1456
rect 9573 -1486 9604 -1473
rect 10338 -1456 10369 -1444
rect 10338 -1473 10345 -1456
rect 10362 -1473 10369 -1456
rect 10338 -1486 10369 -1473
rect 10384 -1456 10415 -1444
rect 10384 -1473 10392 -1456
rect 10409 -1473 10415 -1456
rect 10384 -1486 10415 -1473
<< ndiffc >>
rect 869 9368 886 9385
rect 916 9368 933 9385
rect 1680 9368 1697 9385
rect 1745 9367 1762 9384
rect 1803 9368 1820 9385
rect 2550 9368 2567 9385
rect 2615 9367 2632 9384
rect 2673 9368 2690 9385
rect 3145 9368 3162 9385
rect 3192 9368 3209 9385
rect 8069 9368 8086 9385
rect 8116 9368 8133 9385
rect 8588 9368 8605 9385
rect 8646 9367 8663 9384
rect 8711 9368 8728 9385
rect 9458 9368 9475 9385
rect 9516 9367 9533 9384
rect 9581 9368 9598 9385
rect 10345 9368 10362 9385
rect 10392 9368 10409 9385
rect 869 -1591 886 -1574
rect 916 -1591 933 -1574
rect 1680 -1591 1697 -1574
rect 1745 -1590 1762 -1573
rect 1803 -1591 1820 -1574
rect 2550 -1591 2567 -1574
rect 2615 -1590 2632 -1573
rect 2673 -1591 2690 -1574
rect 3145 -1591 3162 -1574
rect 3192 -1591 3209 -1574
rect 8069 -1591 8086 -1574
rect 8116 -1591 8133 -1574
rect 8588 -1591 8605 -1574
rect 8646 -1590 8663 -1573
rect 8711 -1591 8728 -1574
rect 9458 -1591 9475 -1574
rect 9516 -1590 9533 -1573
rect 9581 -1591 9598 -1574
rect 10345 -1591 10362 -1574
rect 10392 -1591 10409 -1574
<< pdiffc >>
rect 869 9250 886 9267
rect 916 9250 933 9267
rect 1680 9250 1697 9267
rect 1741 9253 1758 9270
rect 1803 9250 1820 9267
rect 2550 9250 2567 9267
rect 2611 9253 2628 9270
rect 2673 9250 2690 9267
rect 3145 9250 3162 9267
rect 3192 9250 3209 9267
rect 8069 9250 8086 9267
rect 8116 9250 8133 9267
rect 8588 9250 8605 9267
rect 8650 9253 8667 9270
rect 8711 9250 8728 9267
rect 9458 9250 9475 9267
rect 9520 9253 9537 9270
rect 9581 9250 9598 9267
rect 10345 9250 10362 9267
rect 10392 9250 10409 9267
rect 869 -1473 886 -1456
rect 916 -1473 933 -1456
rect 1680 -1473 1697 -1456
rect 1741 -1476 1758 -1459
rect 1803 -1473 1820 -1456
rect 2550 -1473 2567 -1456
rect 2611 -1476 2628 -1459
rect 2673 -1473 2690 -1456
rect 3145 -1473 3162 -1456
rect 3192 -1473 3209 -1456
rect 8069 -1473 8086 -1456
rect 8116 -1473 8133 -1456
rect 8588 -1473 8605 -1456
rect 8650 -1476 8667 -1459
rect 8711 -1473 8728 -1456
rect 9458 -1473 9475 -1456
rect 9520 -1476 9537 -1459
rect 9581 -1473 9598 -1456
rect 10345 -1473 10362 -1456
rect 10392 -1473 10409 -1456
<< psubdiff >>
rect 940 9385 969 9397
rect 940 9368 950 9385
rect 967 9368 969 9385
rect 940 9355 969 9368
rect 1827 9385 1856 9397
rect 1827 9368 1837 9385
rect 1854 9368 1856 9385
rect 1827 9355 1856 9368
rect 2697 9385 2726 9397
rect 2697 9368 2707 9385
rect 2724 9368 2726 9385
rect 2697 9355 2726 9368
rect 3216 9385 3245 9397
rect 3216 9368 3226 9385
rect 3243 9368 3245 9385
rect 3216 9355 3245 9368
rect 8033 9385 8062 9397
rect 8033 9368 8035 9385
rect 8052 9368 8062 9385
rect 8033 9355 8062 9368
rect 8552 9385 8581 9397
rect 8552 9368 8554 9385
rect 8571 9368 8581 9385
rect 8552 9355 8581 9368
rect 9422 9385 9451 9397
rect 9422 9368 9424 9385
rect 9441 9368 9451 9385
rect 9422 9355 9451 9368
rect 10309 9385 10338 9397
rect 10309 9368 10311 9385
rect 10328 9368 10338 9385
rect 10309 9355 10338 9368
rect 940 -1574 969 -1561
rect 940 -1591 950 -1574
rect 967 -1591 969 -1574
rect 940 -1603 969 -1591
rect 1827 -1574 1856 -1561
rect 1827 -1591 1837 -1574
rect 1854 -1591 1856 -1574
rect 1827 -1603 1856 -1591
rect 2697 -1574 2726 -1561
rect 2697 -1591 2707 -1574
rect 2724 -1591 2726 -1574
rect 2697 -1603 2726 -1591
rect 3216 -1574 3245 -1561
rect 3216 -1591 3226 -1574
rect 3243 -1591 3245 -1574
rect 3216 -1603 3245 -1591
rect 8033 -1574 8062 -1561
rect 8033 -1591 8035 -1574
rect 8052 -1591 8062 -1574
rect 8033 -1603 8062 -1591
rect 8552 -1574 8581 -1561
rect 8552 -1591 8554 -1574
rect 8571 -1591 8581 -1574
rect 8552 -1603 8581 -1591
rect 9422 -1574 9451 -1561
rect 9422 -1591 9424 -1574
rect 9441 -1591 9451 -1574
rect 9422 -1603 9451 -1591
rect 10309 -1574 10338 -1561
rect 10309 -1591 10311 -1574
rect 10328 -1591 10338 -1574
rect 10309 -1603 10338 -1591
<< nsubdiff >>
rect 940 9267 969 9280
rect 940 9250 950 9267
rect 967 9250 969 9267
rect 940 9238 969 9250
rect 1827 9267 1856 9280
rect 1827 9250 1837 9267
rect 1854 9250 1856 9267
rect 1827 9238 1856 9250
rect 2697 9267 2726 9280
rect 2697 9250 2707 9267
rect 2724 9250 2726 9267
rect 2697 9238 2726 9250
rect 3216 9267 3245 9280
rect 3216 9250 3226 9267
rect 3243 9250 3245 9267
rect 3216 9238 3245 9250
rect 8033 9267 8062 9280
rect 8033 9250 8035 9267
rect 8052 9250 8062 9267
rect 8033 9238 8062 9250
rect 8552 9267 8581 9280
rect 8552 9250 8554 9267
rect 8571 9250 8581 9267
rect 8552 9238 8581 9250
rect 9422 9267 9451 9280
rect 9422 9250 9424 9267
rect 9441 9250 9451 9267
rect 9422 9238 9451 9250
rect 10309 9267 10338 9280
rect 10309 9250 10311 9267
rect 10328 9250 10338 9267
rect 10309 9238 10338 9250
rect 940 -1456 969 -1444
rect 940 -1473 950 -1456
rect 967 -1473 969 -1456
rect 940 -1486 969 -1473
rect 1827 -1456 1856 -1444
rect 1827 -1473 1837 -1456
rect 1854 -1473 1856 -1456
rect 1827 -1486 1856 -1473
rect 2697 -1456 2726 -1444
rect 2697 -1473 2707 -1456
rect 2724 -1473 2726 -1456
rect 2697 -1486 2726 -1473
rect 3216 -1456 3245 -1444
rect 3216 -1473 3226 -1456
rect 3243 -1473 3245 -1456
rect 3216 -1486 3245 -1473
rect 8033 -1456 8062 -1444
rect 8033 -1473 8035 -1456
rect 8052 -1473 8062 -1456
rect 8033 -1486 8062 -1473
rect 8552 -1456 8581 -1444
rect 8552 -1473 8554 -1456
rect 8571 -1473 8581 -1456
rect 8552 -1486 8581 -1473
rect 9422 -1456 9451 -1444
rect 9422 -1473 9424 -1456
rect 9441 -1473 9451 -1456
rect 9422 -1486 9451 -1473
rect 10309 -1456 10338 -1444
rect 10309 -1473 10311 -1456
rect 10328 -1473 10338 -1456
rect 10309 -1486 10338 -1473
<< psubdiffcont >>
rect 950 9368 967 9385
rect 1837 9368 1854 9385
rect 2707 9368 2724 9385
rect 3226 9368 3243 9385
rect 8035 9368 8052 9385
rect 8554 9368 8571 9385
rect 9424 9368 9441 9385
rect 10311 9368 10328 9385
rect 950 -1591 967 -1574
rect 1837 -1591 1854 -1574
rect 2707 -1591 2724 -1574
rect 3226 -1591 3243 -1574
rect 8035 -1591 8052 -1574
rect 8554 -1591 8571 -1574
rect 9424 -1591 9441 -1574
rect 10311 -1591 10328 -1574
<< nsubdiffcont >>
rect 950 9250 967 9267
rect 1837 9250 1854 9267
rect 2707 9250 2724 9267
rect 3226 9250 3243 9267
rect 8035 9250 8052 9267
rect 8554 9250 8571 9267
rect 9424 9250 9441 9267
rect 10311 9250 10328 9267
rect 950 -1473 967 -1456
rect 1837 -1473 1854 -1456
rect 2707 -1473 2724 -1456
rect 3226 -1473 3243 -1456
rect 8035 -1473 8052 -1456
rect 8554 -1473 8571 -1456
rect 9424 -1473 9441 -1456
rect 10311 -1473 10328 -1456
<< poly >>
rect 888 9435 915 9443
rect 1699 9435 1726 9443
rect 1775 9435 1802 9443
rect 2569 9435 2596 9443
rect 2645 9435 2672 9443
rect 3164 9435 3191 9443
rect 8087 9435 8114 9443
rect 8606 9435 8633 9443
rect 8682 9435 8709 9443
rect 9476 9435 9503 9443
rect 9552 9435 9579 9443
rect 10363 9435 10390 9443
rect 885 9418 893 9435
rect 910 9418 918 9435
rect 1696 9418 1704 9435
rect 1721 9418 1729 9435
rect 1772 9418 1780 9435
rect 1797 9418 1805 9435
rect 2566 9418 2574 9435
rect 2591 9418 2599 9435
rect 2642 9418 2650 9435
rect 2667 9418 2675 9435
rect 3161 9418 3169 9435
rect 3186 9418 3194 9435
rect 8084 9418 8092 9435
rect 8109 9418 8117 9435
rect 8603 9418 8611 9435
rect 8628 9418 8636 9435
rect 8679 9418 8687 9435
rect 8704 9418 8712 9435
rect 9473 9418 9481 9435
rect 9498 9418 9506 9435
rect 9549 9418 9557 9435
rect 9574 9418 9582 9435
rect 10360 9418 10368 9435
rect 10385 9418 10393 9435
rect 888 9413 915 9418
rect 1699 9413 1726 9418
rect 1775 9413 1802 9418
rect 2569 9413 2596 9418
rect 2645 9413 2672 9418
rect 3164 9413 3191 9418
rect 8087 9413 8114 9418
rect 8606 9413 8633 9418
rect 8682 9413 8709 9418
rect 9476 9413 9503 9418
rect 9552 9413 9579 9418
rect 10363 9413 10390 9418
rect 894 9397 909 9413
rect 1705 9397 1720 9413
rect 1781 9397 1796 9413
rect 2575 9397 2590 9413
rect 2651 9397 2666 9413
rect 3170 9397 3185 9413
rect 8093 9397 8108 9413
rect 8612 9397 8627 9413
rect 8688 9397 8703 9413
rect 9482 9397 9497 9413
rect 9558 9397 9573 9413
rect 10369 9397 10384 9413
rect 894 9342 909 9355
rect 1705 9342 1720 9355
rect 1781 9342 1796 9355
rect 2575 9342 2590 9355
rect 2651 9342 2666 9355
rect 3170 9342 3185 9355
rect 8093 9342 8108 9355
rect 8612 9342 8627 9355
rect 8688 9342 8703 9355
rect 9482 9342 9497 9355
rect 9558 9342 9573 9355
rect 10369 9342 10384 9355
rect 894 9280 909 9293
rect 1705 9280 1720 9293
rect 1781 9280 1796 9293
rect 2575 9280 2590 9293
rect 2651 9280 2666 9293
rect 3170 9280 3185 9293
rect 8093 9280 8108 9293
rect 8612 9280 8627 9293
rect 8688 9280 8703 9293
rect 9482 9280 9497 9293
rect 9558 9280 9573 9293
rect 10369 9280 10384 9293
rect 894 9219 909 9238
rect 1705 9219 1720 9238
rect 1781 9219 1796 9238
rect 2575 9219 2590 9238
rect 2651 9219 2666 9238
rect 3170 9219 3185 9238
rect 8093 9219 8108 9238
rect 8612 9219 8627 9238
rect 8688 9219 8703 9238
rect 9482 9219 9497 9238
rect 9558 9219 9573 9238
rect 10369 9219 10384 9238
rect 888 9214 915 9219
rect 1699 9214 1726 9219
rect 1775 9214 1802 9219
rect 2569 9214 2596 9219
rect 2645 9214 2672 9219
rect 3164 9214 3191 9219
rect 8087 9214 8114 9219
rect 8606 9214 8633 9219
rect 8682 9214 8709 9219
rect 9476 9214 9503 9219
rect 9552 9214 9579 9219
rect 10363 9214 10390 9219
rect 885 9197 893 9214
rect 910 9197 918 9214
rect 1696 9197 1704 9214
rect 1721 9197 1729 9214
rect 1772 9197 1780 9214
rect 1797 9197 1805 9214
rect 2566 9197 2574 9214
rect 2591 9197 2599 9214
rect 2642 9197 2650 9214
rect 2667 9197 2675 9214
rect 3161 9197 3169 9214
rect 3186 9197 3194 9214
rect 8084 9197 8092 9214
rect 8109 9197 8117 9214
rect 8603 9197 8611 9214
rect 8628 9197 8636 9214
rect 8679 9197 8687 9214
rect 8704 9197 8712 9214
rect 9473 9197 9481 9214
rect 9498 9197 9506 9214
rect 9549 9197 9557 9214
rect 9574 9197 9582 9214
rect 10360 9197 10368 9214
rect 10385 9197 10393 9214
rect 888 9189 915 9197
rect 1699 9189 1726 9197
rect 1775 9189 1802 9197
rect 2569 9189 2596 9197
rect 2645 9189 2672 9197
rect 3164 9189 3191 9197
rect 8087 9189 8114 9197
rect 8606 9189 8633 9197
rect 8682 9189 8709 9197
rect 9476 9189 9503 9197
rect 9552 9189 9579 9197
rect 10363 9189 10390 9197
rect 888 -1403 915 -1395
rect 1699 -1403 1726 -1395
rect 1775 -1403 1802 -1395
rect 2569 -1403 2596 -1395
rect 2645 -1403 2672 -1395
rect 3164 -1403 3191 -1395
rect 8087 -1403 8114 -1395
rect 8606 -1403 8633 -1395
rect 8682 -1403 8709 -1395
rect 9476 -1403 9503 -1395
rect 9552 -1403 9579 -1395
rect 10363 -1403 10390 -1395
rect 885 -1420 893 -1403
rect 910 -1420 918 -1403
rect 1696 -1420 1704 -1403
rect 1721 -1420 1729 -1403
rect 1772 -1420 1780 -1403
rect 1797 -1420 1805 -1403
rect 2566 -1420 2574 -1403
rect 2591 -1420 2599 -1403
rect 2642 -1420 2650 -1403
rect 2667 -1420 2675 -1403
rect 3161 -1420 3169 -1403
rect 3186 -1420 3194 -1403
rect 8084 -1420 8092 -1403
rect 8109 -1420 8117 -1403
rect 8603 -1420 8611 -1403
rect 8628 -1420 8636 -1403
rect 8679 -1420 8687 -1403
rect 8704 -1420 8712 -1403
rect 9473 -1420 9481 -1403
rect 9498 -1420 9506 -1403
rect 9549 -1420 9557 -1403
rect 9574 -1420 9582 -1403
rect 10360 -1420 10368 -1403
rect 10385 -1420 10393 -1403
rect 888 -1425 915 -1420
rect 1699 -1425 1726 -1420
rect 1775 -1425 1802 -1420
rect 2569 -1425 2596 -1420
rect 2645 -1425 2672 -1420
rect 3164 -1425 3191 -1420
rect 8087 -1425 8114 -1420
rect 8606 -1425 8633 -1420
rect 8682 -1425 8709 -1420
rect 9476 -1425 9503 -1420
rect 9552 -1425 9579 -1420
rect 10363 -1425 10390 -1420
rect 894 -1444 909 -1425
rect 1705 -1444 1720 -1425
rect 1781 -1444 1796 -1425
rect 2575 -1444 2590 -1425
rect 2651 -1444 2666 -1425
rect 3170 -1444 3185 -1425
rect 8093 -1444 8108 -1425
rect 8612 -1444 8627 -1425
rect 8688 -1444 8703 -1425
rect 9482 -1444 9497 -1425
rect 9558 -1444 9573 -1425
rect 10369 -1444 10384 -1425
rect 894 -1499 909 -1486
rect 1705 -1499 1720 -1486
rect 1781 -1499 1796 -1486
rect 2575 -1499 2590 -1486
rect 2651 -1499 2666 -1486
rect 3170 -1499 3185 -1486
rect 8093 -1499 8108 -1486
rect 8612 -1499 8627 -1486
rect 8688 -1499 8703 -1486
rect 9482 -1499 9497 -1486
rect 9558 -1499 9573 -1486
rect 10369 -1499 10384 -1486
rect 894 -1561 909 -1548
rect 1705 -1561 1720 -1548
rect 1781 -1561 1796 -1548
rect 2575 -1561 2590 -1548
rect 2651 -1561 2666 -1548
rect 3170 -1561 3185 -1548
rect 8093 -1561 8108 -1548
rect 8612 -1561 8627 -1548
rect 8688 -1561 8703 -1548
rect 9482 -1561 9497 -1548
rect 9558 -1561 9573 -1548
rect 10369 -1561 10384 -1548
rect 894 -1619 909 -1603
rect 1705 -1619 1720 -1603
rect 1781 -1619 1796 -1603
rect 2575 -1619 2590 -1603
rect 2651 -1619 2666 -1603
rect 3170 -1619 3185 -1603
rect 8093 -1619 8108 -1603
rect 8612 -1619 8627 -1603
rect 8688 -1619 8703 -1603
rect 9482 -1619 9497 -1603
rect 9558 -1619 9573 -1603
rect 10369 -1619 10384 -1603
rect 888 -1624 915 -1619
rect 1699 -1624 1726 -1619
rect 1775 -1624 1802 -1619
rect 2569 -1624 2596 -1619
rect 2645 -1624 2672 -1619
rect 3164 -1624 3191 -1619
rect 8087 -1624 8114 -1619
rect 8606 -1624 8633 -1619
rect 8682 -1624 8709 -1619
rect 9476 -1624 9503 -1619
rect 9552 -1624 9579 -1619
rect 10363 -1624 10390 -1619
rect 885 -1641 893 -1624
rect 910 -1641 918 -1624
rect 1696 -1641 1704 -1624
rect 1721 -1641 1729 -1624
rect 1772 -1641 1780 -1624
rect 1797 -1641 1805 -1624
rect 2566 -1641 2574 -1624
rect 2591 -1641 2599 -1624
rect 2642 -1641 2650 -1624
rect 2667 -1641 2675 -1624
rect 3161 -1641 3169 -1624
rect 3186 -1641 3194 -1624
rect 8084 -1641 8092 -1624
rect 8109 -1641 8117 -1624
rect 8603 -1641 8611 -1624
rect 8628 -1641 8636 -1624
rect 8679 -1641 8687 -1624
rect 8704 -1641 8712 -1624
rect 9473 -1641 9481 -1624
rect 9498 -1641 9506 -1624
rect 9549 -1641 9557 -1624
rect 9574 -1641 9582 -1624
rect 10360 -1641 10368 -1624
rect 10385 -1641 10393 -1624
rect 888 -1649 915 -1641
rect 1699 -1649 1726 -1641
rect 1775 -1649 1802 -1641
rect 2569 -1649 2596 -1641
rect 2645 -1649 2672 -1641
rect 3164 -1649 3191 -1641
rect 8087 -1649 8114 -1641
rect 8606 -1649 8633 -1641
rect 8682 -1649 8709 -1641
rect 9476 -1649 9503 -1641
rect 9552 -1649 9579 -1641
rect 10363 -1649 10390 -1641
<< polycont >>
rect 893 9418 910 9435
rect 1704 9418 1721 9435
rect 1780 9418 1797 9435
rect 2574 9418 2591 9435
rect 2650 9418 2667 9435
rect 3169 9418 3186 9435
rect 8092 9418 8109 9435
rect 8611 9418 8628 9435
rect 8687 9418 8704 9435
rect 9481 9418 9498 9435
rect 9557 9418 9574 9435
rect 10368 9418 10385 9435
rect 893 9197 910 9214
rect 1704 9197 1721 9214
rect 1780 9197 1797 9214
rect 2574 9197 2591 9214
rect 2650 9197 2667 9214
rect 3169 9197 3186 9214
rect 8092 9197 8109 9214
rect 8611 9197 8628 9214
rect 8687 9197 8704 9214
rect 9481 9197 9498 9214
rect 9557 9197 9574 9214
rect 10368 9197 10385 9214
rect 893 -1420 910 -1403
rect 1704 -1420 1721 -1403
rect 1780 -1420 1797 -1403
rect 2574 -1420 2591 -1403
rect 2650 -1420 2667 -1403
rect 3169 -1420 3186 -1403
rect 8092 -1420 8109 -1403
rect 8611 -1420 8628 -1403
rect 8687 -1420 8704 -1403
rect 9481 -1420 9498 -1403
rect 9557 -1420 9574 -1403
rect 10368 -1420 10385 -1403
rect 893 -1641 910 -1624
rect 1704 -1641 1721 -1624
rect 1780 -1641 1797 -1624
rect 2574 -1641 2591 -1624
rect 2650 -1641 2667 -1624
rect 3169 -1641 3186 -1624
rect 8092 -1641 8109 -1624
rect 8611 -1641 8628 -1624
rect 8687 -1641 8704 -1624
rect 9481 -1641 9498 -1624
rect 9557 -1641 9574 -1624
rect 10368 -1641 10385 -1624
<< locali >>
rect 3620 9534 3637 9545
rect 798 9477 829 9494
rect 846 9477 877 9494
rect 894 9477 925 9494
rect 942 9477 973 9494
rect 990 9477 1021 9494
rect 1038 9477 1051 9494
rect 1609 9477 1640 9494
rect 1657 9477 1688 9494
rect 1733 9477 1764 9494
rect 1781 9477 1812 9494
rect 1829 9477 1860 9494
rect 1877 9477 1908 9494
rect 1925 9477 1938 9494
rect 2479 9477 2510 9494
rect 2527 9477 2558 9494
rect 2603 9477 2634 9494
rect 2651 9477 2682 9494
rect 2699 9477 2730 9494
rect 2747 9477 2778 9494
rect 2795 9477 2808 9494
rect 3074 9477 3105 9494
rect 3122 9477 3153 9494
rect 3170 9477 3201 9494
rect 3218 9477 3249 9494
rect 3266 9477 3297 9494
rect 3314 9477 3327 9494
rect 885 9418 893 9435
rect 910 9418 918 9435
rect 869 9385 886 9393
rect 869 9267 886 9368
rect 869 9242 886 9250
rect 916 9385 933 9393
rect 916 9331 933 9368
rect 950 9385 967 9477
rect 1696 9418 1704 9435
rect 1721 9418 1729 9435
rect 1772 9418 1780 9435
rect 1797 9418 1805 9435
rect 950 9360 967 9368
rect 1680 9385 1697 9393
rect 916 9314 924 9331
rect 1680 9328 1697 9368
rect 916 9267 933 9314
rect 916 9242 933 9250
rect 950 9267 967 9275
rect 885 9197 893 9214
rect 910 9197 918 9214
rect 950 9161 967 9250
rect 1680 9267 1697 9311
rect 1680 9242 1697 9250
rect 1727 9384 1773 9393
rect 1727 9367 1745 9384
rect 1762 9367 1773 9384
rect 1727 9332 1773 9367
rect 1744 9315 1773 9332
rect 1727 9270 1773 9315
rect 1727 9253 1741 9270
rect 1758 9253 1773 9270
rect 1727 9242 1773 9253
rect 1803 9385 1820 9393
rect 1803 9331 1820 9368
rect 1837 9385 1854 9477
rect 2566 9418 2574 9435
rect 2591 9418 2599 9435
rect 2642 9418 2650 9435
rect 2667 9418 2675 9435
rect 1837 9360 1854 9368
rect 2550 9385 2567 9393
rect 1803 9314 1811 9331
rect 2550 9328 2567 9368
rect 1803 9267 1820 9314
rect 1803 9242 1820 9250
rect 1837 9267 1854 9275
rect 1696 9197 1704 9214
rect 1721 9197 1729 9214
rect 1772 9197 1780 9214
rect 1797 9197 1805 9214
rect 1837 9161 1854 9250
rect 2550 9267 2567 9311
rect 2550 9242 2567 9250
rect 2597 9384 2643 9393
rect 2597 9367 2615 9384
rect 2632 9367 2643 9384
rect 2597 9332 2643 9367
rect 2614 9315 2643 9332
rect 2597 9270 2643 9315
rect 2597 9253 2611 9270
rect 2628 9253 2643 9270
rect 2597 9242 2643 9253
rect 2673 9385 2690 9393
rect 2673 9331 2690 9368
rect 2707 9385 2724 9477
rect 3161 9418 3169 9435
rect 3186 9418 3194 9435
rect 2707 9360 2724 9368
rect 3145 9385 3162 9393
rect 2673 9314 2681 9331
rect 3145 9330 3162 9368
rect 2673 9267 2690 9314
rect 3153 9313 3162 9330
rect 2673 9242 2690 9250
rect 2707 9267 2724 9275
rect 2566 9197 2574 9214
rect 2591 9197 2599 9214
rect 2642 9197 2650 9214
rect 2667 9197 2675 9214
rect 2707 9161 2724 9250
rect 3145 9267 3162 9313
rect 3145 9242 3162 9250
rect 3192 9385 3209 9393
rect 3192 9331 3209 9368
rect 3226 9385 3243 9477
rect 3620 9419 3637 9517
rect 7641 9534 7658 9545
rect 7641 9419 7658 9517
rect 7951 9477 7964 9494
rect 7981 9477 8012 9494
rect 8029 9477 8060 9494
rect 8077 9477 8108 9494
rect 8125 9477 8156 9494
rect 8173 9477 8204 9494
rect 8470 9477 8483 9494
rect 8500 9477 8531 9494
rect 8548 9477 8579 9494
rect 8596 9477 8627 9494
rect 8644 9477 8675 9494
rect 8720 9477 8751 9494
rect 8768 9477 8799 9494
rect 9340 9477 9353 9494
rect 9370 9477 9401 9494
rect 9418 9477 9449 9494
rect 9466 9477 9497 9494
rect 9514 9477 9545 9494
rect 9590 9477 9621 9494
rect 9638 9477 9669 9494
rect 10227 9477 10240 9494
rect 10257 9477 10288 9494
rect 10305 9477 10336 9494
rect 10353 9477 10384 9494
rect 10401 9477 10432 9494
rect 10449 9477 10480 9494
rect 3226 9360 3243 9368
rect 8035 9385 8052 9477
rect 8084 9418 8092 9435
rect 8109 9418 8117 9435
rect 8035 9360 8052 9368
rect 8069 9385 8086 9393
rect 8069 9331 8086 9368
rect 3192 9314 3200 9331
rect 8078 9314 8086 9331
rect 3192 9267 3209 9314
rect 3192 9242 3209 9250
rect 3226 9267 3243 9275
rect 3161 9197 3169 9214
rect 3186 9197 3194 9214
rect 3226 9161 3243 9250
rect 8035 9267 8052 9275
rect 8035 9161 8052 9250
rect 8069 9267 8086 9314
rect 8069 9242 8086 9250
rect 8116 9385 8133 9393
rect 8116 9330 8133 9368
rect 8554 9385 8571 9477
rect 8603 9418 8611 9435
rect 8628 9418 8636 9435
rect 8679 9418 8687 9435
rect 8704 9418 8712 9435
rect 8554 9360 8571 9368
rect 8588 9385 8605 9393
rect 8588 9331 8605 9368
rect 8116 9313 8125 9330
rect 8597 9314 8605 9331
rect 8116 9267 8133 9313
rect 8116 9242 8133 9250
rect 8554 9267 8571 9275
rect 8084 9197 8092 9214
rect 8109 9197 8117 9214
rect 8554 9161 8571 9250
rect 8588 9267 8605 9314
rect 8588 9242 8605 9250
rect 8635 9384 8681 9393
rect 8635 9367 8646 9384
rect 8663 9367 8681 9384
rect 8635 9332 8681 9367
rect 8635 9315 8664 9332
rect 8635 9270 8681 9315
rect 8635 9253 8650 9270
rect 8667 9253 8681 9270
rect 8635 9242 8681 9253
rect 8711 9385 8728 9393
rect 8711 9328 8728 9368
rect 9424 9385 9441 9477
rect 9473 9418 9481 9435
rect 9498 9418 9506 9435
rect 9549 9418 9557 9435
rect 9574 9418 9582 9435
rect 9424 9360 9441 9368
rect 9458 9385 9475 9393
rect 9458 9331 9475 9368
rect 9467 9314 9475 9331
rect 8711 9267 8728 9311
rect 8711 9242 8728 9250
rect 9424 9267 9441 9275
rect 8603 9197 8611 9214
rect 8628 9197 8636 9214
rect 8679 9197 8687 9214
rect 8704 9197 8712 9214
rect 9424 9161 9441 9250
rect 9458 9267 9475 9314
rect 9458 9242 9475 9250
rect 9505 9384 9551 9393
rect 9505 9367 9516 9384
rect 9533 9367 9551 9384
rect 9505 9332 9551 9367
rect 9505 9315 9534 9332
rect 9505 9270 9551 9315
rect 9505 9253 9520 9270
rect 9537 9253 9551 9270
rect 9505 9242 9551 9253
rect 9581 9385 9598 9393
rect 9581 9328 9598 9368
rect 10311 9385 10328 9477
rect 10360 9418 10368 9435
rect 10385 9418 10393 9435
rect 10311 9360 10328 9368
rect 10345 9385 10362 9393
rect 10345 9331 10362 9368
rect 10354 9314 10362 9331
rect 9581 9267 9598 9311
rect 9581 9242 9598 9250
rect 10311 9267 10328 9275
rect 9473 9197 9481 9214
rect 9498 9197 9506 9214
rect 9549 9197 9557 9214
rect 9574 9197 9582 9214
rect 10311 9161 10328 9250
rect 10345 9267 10362 9314
rect 10345 9242 10362 9250
rect 10392 9385 10409 9393
rect 10392 9267 10409 9368
rect 10392 9242 10409 9250
rect 10360 9197 10368 9214
rect 10385 9197 10393 9214
rect 798 9144 829 9161
rect 846 9144 877 9161
rect 894 9144 925 9161
rect 942 9144 973 9161
rect 990 9144 1021 9161
rect 1038 9144 1051 9161
rect 1609 9144 1640 9161
rect 1657 9144 1688 9161
rect 1733 9144 1764 9161
rect 1781 9144 1812 9161
rect 1829 9144 1860 9161
rect 1877 9144 1908 9161
rect 1925 9144 1938 9161
rect 2479 9144 2510 9161
rect 2527 9144 2558 9161
rect 2603 9144 2634 9161
rect 2651 9144 2682 9161
rect 2699 9144 2730 9161
rect 2747 9144 2778 9161
rect 2795 9144 2808 9161
rect 3074 9144 3105 9161
rect 3122 9144 3153 9161
rect 3170 9144 3201 9161
rect 3218 9144 3249 9161
rect 3266 9144 3297 9161
rect 3314 9144 3327 9161
rect 7951 9144 7964 9161
rect 7981 9144 8012 9161
rect 8029 9144 8060 9161
rect 8077 9144 8108 9161
rect 8125 9144 8156 9161
rect 8173 9144 8204 9161
rect 8470 9144 8483 9161
rect 8500 9144 8531 9161
rect 8548 9144 8579 9161
rect 8596 9144 8627 9161
rect 8644 9144 8675 9161
rect 8720 9144 8751 9161
rect 8768 9144 8799 9161
rect 9340 9144 9353 9161
rect 9370 9144 9401 9161
rect 9418 9144 9449 9161
rect 9466 9144 9497 9161
rect 9514 9144 9545 9161
rect 9590 9144 9621 9161
rect 9638 9144 9669 9161
rect 10227 9144 10240 9161
rect 10257 9144 10288 9161
rect 10305 9144 10336 9161
rect 10353 9144 10384 9161
rect 10401 9144 10432 9161
rect 10449 9144 10480 9161
rect 798 -1367 829 -1350
rect 846 -1367 877 -1350
rect 894 -1367 925 -1350
rect 942 -1367 973 -1350
rect 990 -1367 1021 -1350
rect 1038 -1367 1051 -1350
rect 1609 -1367 1640 -1350
rect 1657 -1367 1688 -1350
rect 1733 -1367 1764 -1350
rect 1781 -1367 1812 -1350
rect 1829 -1367 1860 -1350
rect 1877 -1367 1908 -1350
rect 1925 -1367 1938 -1350
rect 2479 -1367 2510 -1350
rect 2527 -1367 2558 -1350
rect 2603 -1367 2634 -1350
rect 2651 -1367 2682 -1350
rect 2699 -1367 2730 -1350
rect 2747 -1367 2778 -1350
rect 2795 -1367 2808 -1350
rect 3074 -1367 3105 -1350
rect 3122 -1367 3153 -1350
rect 3170 -1367 3201 -1350
rect 3218 -1367 3249 -1350
rect 3266 -1367 3297 -1350
rect 3314 -1367 3327 -1350
rect 7951 -1367 7964 -1350
rect 7981 -1367 8012 -1350
rect 8029 -1367 8060 -1350
rect 8077 -1367 8108 -1350
rect 8125 -1367 8156 -1350
rect 8173 -1367 8204 -1350
rect 8470 -1367 8483 -1350
rect 8500 -1367 8531 -1350
rect 8548 -1367 8579 -1350
rect 8596 -1367 8627 -1350
rect 8644 -1367 8675 -1350
rect 8720 -1367 8751 -1350
rect 8768 -1367 8799 -1350
rect 9340 -1367 9353 -1350
rect 9370 -1367 9401 -1350
rect 9418 -1367 9449 -1350
rect 9466 -1367 9497 -1350
rect 9514 -1367 9545 -1350
rect 9590 -1367 9621 -1350
rect 9638 -1367 9669 -1350
rect 10227 -1367 10240 -1350
rect 10257 -1367 10288 -1350
rect 10305 -1367 10336 -1350
rect 10353 -1367 10384 -1350
rect 10401 -1367 10432 -1350
rect 10449 -1367 10480 -1350
rect 885 -1420 893 -1403
rect 910 -1420 918 -1403
rect 869 -1456 886 -1448
rect 869 -1574 886 -1473
rect 869 -1599 886 -1591
rect 916 -1456 933 -1448
rect 916 -1520 933 -1473
rect 950 -1456 967 -1367
rect 1696 -1420 1704 -1403
rect 1721 -1420 1729 -1403
rect 1772 -1420 1780 -1403
rect 1797 -1420 1805 -1403
rect 950 -1481 967 -1473
rect 1680 -1456 1697 -1448
rect 1680 -1517 1697 -1473
rect 916 -1537 924 -1520
rect 916 -1574 933 -1537
rect 916 -1599 933 -1591
rect 950 -1574 967 -1566
rect 885 -1641 893 -1624
rect 910 -1641 918 -1624
rect 950 -1683 967 -1591
rect 1680 -1574 1697 -1534
rect 1680 -1599 1697 -1591
rect 1727 -1459 1773 -1448
rect 1727 -1476 1741 -1459
rect 1758 -1476 1773 -1459
rect 1727 -1521 1773 -1476
rect 1744 -1538 1773 -1521
rect 1727 -1573 1773 -1538
rect 1727 -1590 1745 -1573
rect 1762 -1590 1773 -1573
rect 1727 -1599 1773 -1590
rect 1803 -1456 1820 -1448
rect 1803 -1520 1820 -1473
rect 1837 -1456 1854 -1367
rect 2566 -1420 2574 -1403
rect 2591 -1420 2599 -1403
rect 2642 -1420 2650 -1403
rect 2667 -1420 2675 -1403
rect 1837 -1481 1854 -1473
rect 2550 -1456 2567 -1448
rect 2550 -1517 2567 -1473
rect 1803 -1537 1811 -1520
rect 1803 -1574 1820 -1537
rect 1803 -1599 1820 -1591
rect 1837 -1574 1854 -1566
rect 1696 -1641 1704 -1624
rect 1721 -1641 1729 -1624
rect 1772 -1641 1780 -1624
rect 1797 -1641 1805 -1624
rect 1837 -1683 1854 -1591
rect 2550 -1574 2567 -1534
rect 2550 -1599 2567 -1591
rect 2597 -1459 2643 -1448
rect 2597 -1476 2611 -1459
rect 2628 -1476 2643 -1459
rect 2597 -1521 2643 -1476
rect 2614 -1538 2643 -1521
rect 2597 -1573 2643 -1538
rect 2597 -1590 2615 -1573
rect 2632 -1590 2643 -1573
rect 2597 -1599 2643 -1590
rect 2673 -1456 2690 -1448
rect 2673 -1520 2690 -1473
rect 2707 -1456 2724 -1367
rect 3161 -1420 3169 -1403
rect 3186 -1420 3194 -1403
rect 2707 -1481 2724 -1473
rect 3145 -1456 3162 -1448
rect 3145 -1519 3162 -1473
rect 2673 -1537 2681 -1520
rect 3153 -1536 3162 -1519
rect 2673 -1574 2690 -1537
rect 2673 -1599 2690 -1591
rect 2707 -1574 2724 -1566
rect 2566 -1641 2574 -1624
rect 2591 -1641 2599 -1624
rect 2642 -1641 2650 -1624
rect 2667 -1641 2675 -1624
rect 2707 -1683 2724 -1591
rect 3145 -1574 3162 -1536
rect 3145 -1599 3162 -1591
rect 3192 -1456 3209 -1448
rect 3192 -1520 3209 -1473
rect 3226 -1456 3243 -1367
rect 3226 -1481 3243 -1473
rect 8035 -1456 8052 -1367
rect 8084 -1420 8092 -1403
rect 8109 -1420 8117 -1403
rect 8035 -1481 8052 -1473
rect 8069 -1456 8086 -1448
rect 8069 -1520 8086 -1473
rect 3192 -1537 3200 -1520
rect 8078 -1537 8086 -1520
rect 3192 -1574 3209 -1537
rect 3192 -1599 3209 -1591
rect 3226 -1574 3243 -1566
rect 3161 -1641 3169 -1624
rect 3186 -1641 3194 -1624
rect 3226 -1683 3243 -1591
rect 8035 -1574 8052 -1566
rect 798 -1700 829 -1683
rect 846 -1700 877 -1683
rect 894 -1700 925 -1683
rect 942 -1700 973 -1683
rect 990 -1700 1021 -1683
rect 1038 -1700 1051 -1683
rect 1609 -1700 1640 -1683
rect 1657 -1700 1688 -1683
rect 1733 -1700 1764 -1683
rect 1781 -1700 1812 -1683
rect 1829 -1700 1860 -1683
rect 1877 -1700 1908 -1683
rect 1925 -1700 1938 -1683
rect 2479 -1700 2510 -1683
rect 2527 -1700 2558 -1683
rect 2603 -1700 2634 -1683
rect 2651 -1700 2682 -1683
rect 2699 -1700 2730 -1683
rect 2747 -1700 2778 -1683
rect 2795 -1700 2808 -1683
rect 3074 -1700 3105 -1683
rect 3122 -1700 3153 -1683
rect 3170 -1700 3201 -1683
rect 3218 -1700 3249 -1683
rect 3266 -1700 3297 -1683
rect 3314 -1700 3327 -1683
rect 3620 -1723 3637 -1625
rect 3620 -1751 3637 -1740
rect 7641 -1723 7658 -1625
rect 8035 -1683 8052 -1591
rect 8069 -1574 8086 -1537
rect 8069 -1599 8086 -1591
rect 8116 -1456 8133 -1448
rect 8116 -1519 8133 -1473
rect 8554 -1456 8571 -1367
rect 8603 -1420 8611 -1403
rect 8628 -1420 8636 -1403
rect 8679 -1420 8687 -1403
rect 8704 -1420 8712 -1403
rect 8554 -1481 8571 -1473
rect 8588 -1456 8605 -1448
rect 8116 -1536 8125 -1519
rect 8588 -1520 8605 -1473
rect 8116 -1574 8133 -1536
rect 8597 -1537 8605 -1520
rect 8116 -1599 8133 -1591
rect 8554 -1574 8571 -1566
rect 8084 -1641 8092 -1624
rect 8109 -1641 8117 -1624
rect 8554 -1683 8571 -1591
rect 8588 -1574 8605 -1537
rect 8588 -1599 8605 -1591
rect 8635 -1459 8681 -1448
rect 8635 -1476 8650 -1459
rect 8667 -1476 8681 -1459
rect 8635 -1521 8681 -1476
rect 8635 -1538 8664 -1521
rect 8635 -1573 8681 -1538
rect 8635 -1590 8646 -1573
rect 8663 -1590 8681 -1573
rect 8635 -1599 8681 -1590
rect 8711 -1456 8728 -1448
rect 8711 -1517 8728 -1473
rect 9424 -1456 9441 -1367
rect 9473 -1420 9481 -1403
rect 9498 -1420 9506 -1403
rect 9549 -1420 9557 -1403
rect 9574 -1420 9582 -1403
rect 9424 -1481 9441 -1473
rect 9458 -1456 9475 -1448
rect 9458 -1520 9475 -1473
rect 8711 -1574 8728 -1534
rect 9467 -1537 9475 -1520
rect 8711 -1599 8728 -1591
rect 9424 -1574 9441 -1566
rect 8603 -1641 8611 -1624
rect 8628 -1641 8636 -1624
rect 8679 -1641 8687 -1624
rect 8704 -1641 8712 -1624
rect 9424 -1683 9441 -1591
rect 9458 -1574 9475 -1537
rect 9458 -1599 9475 -1591
rect 9505 -1459 9551 -1448
rect 9505 -1476 9520 -1459
rect 9537 -1476 9551 -1459
rect 9505 -1521 9551 -1476
rect 9505 -1538 9534 -1521
rect 9505 -1573 9551 -1538
rect 9505 -1590 9516 -1573
rect 9533 -1590 9551 -1573
rect 9505 -1599 9551 -1590
rect 9581 -1456 9598 -1448
rect 9581 -1517 9598 -1473
rect 10311 -1456 10328 -1367
rect 10360 -1420 10368 -1403
rect 10385 -1420 10393 -1403
rect 10311 -1481 10328 -1473
rect 10345 -1456 10362 -1448
rect 10345 -1520 10362 -1473
rect 9581 -1574 9598 -1534
rect 10354 -1537 10362 -1520
rect 9581 -1599 9598 -1591
rect 10311 -1574 10328 -1566
rect 9473 -1641 9481 -1624
rect 9498 -1641 9506 -1624
rect 9549 -1641 9557 -1624
rect 9574 -1641 9582 -1624
rect 10311 -1683 10328 -1591
rect 10345 -1574 10362 -1537
rect 10345 -1599 10362 -1591
rect 10392 -1456 10409 -1448
rect 10392 -1574 10409 -1473
rect 10392 -1599 10409 -1591
rect 10360 -1641 10368 -1624
rect 10385 -1641 10393 -1624
rect 7951 -1700 7964 -1683
rect 7981 -1700 8012 -1683
rect 8029 -1700 8060 -1683
rect 8077 -1700 8108 -1683
rect 8125 -1700 8156 -1683
rect 8173 -1700 8204 -1683
rect 8470 -1700 8483 -1683
rect 8500 -1700 8531 -1683
rect 8548 -1700 8579 -1683
rect 8596 -1700 8627 -1683
rect 8644 -1700 8675 -1683
rect 8720 -1700 8751 -1683
rect 8768 -1700 8799 -1683
rect 9340 -1700 9353 -1683
rect 9370 -1700 9401 -1683
rect 9418 -1700 9449 -1683
rect 9466 -1700 9497 -1683
rect 9514 -1700 9545 -1683
rect 9590 -1700 9621 -1683
rect 9638 -1700 9669 -1683
rect 10227 -1700 10240 -1683
rect 10257 -1700 10288 -1683
rect 10305 -1700 10336 -1683
rect 10353 -1700 10384 -1683
rect 10401 -1700 10432 -1683
rect 10449 -1700 10480 -1683
rect 7641 -1751 7658 -1740
<< viali >>
rect 3620 9517 3637 9534
rect 829 9477 846 9494
rect 877 9477 894 9494
rect 925 9477 942 9494
rect 973 9477 990 9494
rect 1021 9477 1038 9494
rect 1640 9477 1657 9494
rect 1688 9477 1733 9494
rect 1764 9477 1781 9494
rect 1812 9477 1829 9494
rect 1860 9477 1877 9494
rect 1908 9477 1925 9494
rect 2510 9477 2527 9494
rect 2558 9477 2603 9494
rect 2634 9477 2651 9494
rect 2682 9477 2699 9494
rect 2730 9477 2747 9494
rect 2778 9477 2795 9494
rect 3105 9477 3122 9494
rect 3153 9477 3170 9494
rect 3201 9477 3218 9494
rect 3249 9477 3266 9494
rect 3297 9477 3314 9494
rect 924 9314 941 9331
rect 1680 9311 1697 9328
rect 1727 9315 1744 9332
rect 1811 9314 1828 9331
rect 2550 9311 2567 9328
rect 2597 9315 2614 9332
rect 2681 9314 2698 9331
rect 3136 9313 3153 9330
rect 7641 9517 7658 9534
rect 7964 9477 7981 9494
rect 8012 9477 8029 9494
rect 8060 9477 8077 9494
rect 8108 9477 8125 9494
rect 8156 9477 8173 9494
rect 8483 9477 8500 9494
rect 8531 9477 8548 9494
rect 8579 9477 8596 9494
rect 8627 9477 8644 9494
rect 8675 9477 8720 9494
rect 8751 9477 8768 9494
rect 9353 9477 9370 9494
rect 9401 9477 9418 9494
rect 9449 9477 9466 9494
rect 9497 9477 9514 9494
rect 9545 9477 9590 9494
rect 9621 9477 9638 9494
rect 10240 9477 10257 9494
rect 10288 9477 10305 9494
rect 10336 9477 10353 9494
rect 10384 9477 10401 9494
rect 10432 9477 10449 9494
rect 3200 9314 3217 9331
rect 8061 9314 8078 9331
rect 8125 9313 8142 9330
rect 8580 9314 8597 9331
rect 8664 9315 8681 9332
rect 8711 9311 8728 9328
rect 9450 9314 9467 9331
rect 9534 9315 9551 9332
rect 9581 9311 9598 9328
rect 10337 9314 10354 9331
rect 829 9144 846 9161
rect 877 9144 894 9161
rect 925 9144 942 9161
rect 973 9144 990 9161
rect 1021 9144 1038 9161
rect 1640 9144 1657 9161
rect 1688 9144 1733 9161
rect 1764 9144 1781 9161
rect 1812 9144 1829 9161
rect 1860 9144 1877 9161
rect 1908 9144 1925 9161
rect 2510 9144 2527 9161
rect 2558 9144 2603 9161
rect 2634 9144 2651 9161
rect 2682 9144 2699 9161
rect 2730 9144 2747 9161
rect 2778 9144 2795 9161
rect 3105 9144 3122 9161
rect 3153 9144 3170 9161
rect 3201 9144 3218 9161
rect 3249 9144 3266 9161
rect 3297 9144 3314 9161
rect 7964 9144 7981 9161
rect 8012 9144 8029 9161
rect 8060 9144 8077 9161
rect 8108 9144 8125 9161
rect 8156 9144 8173 9161
rect 8483 9144 8500 9161
rect 8531 9144 8548 9161
rect 8579 9144 8596 9161
rect 8627 9144 8644 9161
rect 8675 9144 8720 9161
rect 8751 9144 8768 9161
rect 9353 9144 9370 9161
rect 9401 9144 9418 9161
rect 9449 9144 9466 9161
rect 9497 9144 9514 9161
rect 9545 9144 9590 9161
rect 9621 9144 9638 9161
rect 10240 9144 10257 9161
rect 10288 9144 10305 9161
rect 10336 9144 10353 9161
rect 10384 9144 10401 9161
rect 10432 9144 10449 9161
rect 829 -1367 846 -1350
rect 877 -1367 894 -1350
rect 925 -1367 942 -1350
rect 973 -1367 990 -1350
rect 1021 -1367 1038 -1350
rect 1640 -1367 1657 -1350
rect 1688 -1367 1733 -1350
rect 1764 -1367 1781 -1350
rect 1812 -1367 1829 -1350
rect 1860 -1367 1877 -1350
rect 1908 -1367 1925 -1350
rect 2510 -1367 2527 -1350
rect 2558 -1367 2603 -1350
rect 2634 -1367 2651 -1350
rect 2682 -1367 2699 -1350
rect 2730 -1367 2747 -1350
rect 2778 -1367 2795 -1350
rect 3105 -1367 3122 -1350
rect 3153 -1367 3170 -1350
rect 3201 -1367 3218 -1350
rect 3249 -1367 3266 -1350
rect 3297 -1367 3314 -1350
rect 7964 -1367 7981 -1350
rect 8012 -1367 8029 -1350
rect 8060 -1367 8077 -1350
rect 8108 -1367 8125 -1350
rect 8156 -1367 8173 -1350
rect 8483 -1367 8500 -1350
rect 8531 -1367 8548 -1350
rect 8579 -1367 8596 -1350
rect 8627 -1367 8644 -1350
rect 8675 -1367 8720 -1350
rect 8751 -1367 8768 -1350
rect 9353 -1367 9370 -1350
rect 9401 -1367 9418 -1350
rect 9449 -1367 9466 -1350
rect 9497 -1367 9514 -1350
rect 9545 -1367 9590 -1350
rect 9621 -1367 9638 -1350
rect 10240 -1367 10257 -1350
rect 10288 -1367 10305 -1350
rect 10336 -1367 10353 -1350
rect 10384 -1367 10401 -1350
rect 10432 -1367 10449 -1350
rect 924 -1537 941 -1520
rect 1680 -1534 1697 -1517
rect 1727 -1538 1744 -1521
rect 1811 -1537 1828 -1520
rect 2550 -1534 2567 -1517
rect 2597 -1538 2614 -1521
rect 2681 -1537 2698 -1520
rect 3136 -1536 3153 -1519
rect 3200 -1537 3217 -1520
rect 8061 -1537 8078 -1520
rect 829 -1700 846 -1683
rect 877 -1700 894 -1683
rect 925 -1700 942 -1683
rect 973 -1700 990 -1683
rect 1021 -1700 1038 -1683
rect 1640 -1700 1657 -1683
rect 1688 -1700 1733 -1683
rect 1764 -1700 1781 -1683
rect 1812 -1700 1829 -1683
rect 1860 -1700 1877 -1683
rect 1908 -1700 1925 -1683
rect 2510 -1700 2527 -1683
rect 2558 -1700 2603 -1683
rect 2634 -1700 2651 -1683
rect 2682 -1700 2699 -1683
rect 2730 -1700 2747 -1683
rect 2778 -1700 2795 -1683
rect 3105 -1700 3122 -1683
rect 3153 -1700 3170 -1683
rect 3201 -1700 3218 -1683
rect 3249 -1700 3266 -1683
rect 3297 -1700 3314 -1683
rect 3620 -1740 3637 -1723
rect 8125 -1536 8142 -1519
rect 8580 -1537 8597 -1520
rect 8664 -1538 8681 -1521
rect 8711 -1534 8728 -1517
rect 9450 -1537 9467 -1520
rect 9534 -1538 9551 -1521
rect 9581 -1534 9598 -1517
rect 10337 -1537 10354 -1520
rect 7964 -1700 7981 -1683
rect 8012 -1700 8029 -1683
rect 8060 -1700 8077 -1683
rect 8108 -1700 8125 -1683
rect 8156 -1700 8173 -1683
rect 8483 -1700 8500 -1683
rect 8531 -1700 8548 -1683
rect 8579 -1700 8596 -1683
rect 8627 -1700 8644 -1683
rect 8675 -1700 8720 -1683
rect 8751 -1700 8768 -1683
rect 9353 -1700 9370 -1683
rect 9401 -1700 9418 -1683
rect 9449 -1700 9466 -1683
rect 9497 -1700 9514 -1683
rect 9545 -1700 9590 -1683
rect 9621 -1700 9638 -1683
rect 10240 -1700 10257 -1683
rect 10288 -1700 10305 -1683
rect 10336 -1700 10353 -1683
rect 10384 -1700 10401 -1683
rect 10432 -1700 10449 -1683
rect 7641 -1740 7658 -1723
<< metal1 >>
rect 3614 9538 3642 9542
rect 3614 9512 3616 9538
rect 798 9494 1051 9510
rect 798 9477 829 9494
rect 846 9477 877 9494
rect 894 9477 925 9494
rect 942 9477 973 9494
rect 990 9477 1021 9494
rect 1038 9477 1051 9494
rect 798 9461 1051 9477
rect 1609 9494 1938 9510
rect 1609 9477 1640 9494
rect 1657 9477 1688 9494
rect 1733 9477 1764 9494
rect 1781 9477 1812 9494
rect 1829 9477 1860 9494
rect 1877 9477 1908 9494
rect 1925 9477 1938 9494
rect 1609 9461 1938 9477
rect 2479 9494 2808 9510
rect 2479 9477 2510 9494
rect 2527 9477 2558 9494
rect 2603 9477 2634 9494
rect 2651 9477 2682 9494
rect 2699 9477 2730 9494
rect 2747 9477 2778 9494
rect 2795 9477 2808 9494
rect 2479 9461 2808 9477
rect 3074 9494 3327 9510
rect 3614 9509 3642 9512
rect 7636 9538 7664 9542
rect 7662 9512 7664 9538
rect 7636 9509 7664 9512
rect 3074 9477 3105 9494
rect 3122 9477 3153 9494
rect 3170 9477 3201 9494
rect 3218 9477 3249 9494
rect 3266 9477 3297 9494
rect 3314 9477 3327 9494
rect 3074 9461 3327 9477
rect 7951 9494 8204 9510
rect 7951 9477 7964 9494
rect 7981 9477 8012 9494
rect 8029 9477 8060 9494
rect 8077 9477 8108 9494
rect 8125 9477 8156 9494
rect 8173 9477 8204 9494
rect 7951 9461 8204 9477
rect 8470 9494 8799 9510
rect 8470 9477 8483 9494
rect 8500 9477 8531 9494
rect 8548 9477 8579 9494
rect 8596 9477 8627 9494
rect 8644 9477 8675 9494
rect 8720 9477 8751 9494
rect 8768 9477 8799 9494
rect 8470 9461 8799 9477
rect 9340 9494 9669 9510
rect 9340 9477 9353 9494
rect 9370 9477 9401 9494
rect 9418 9477 9449 9494
rect 9466 9477 9497 9494
rect 9514 9477 9545 9494
rect 9590 9477 9621 9494
rect 9638 9477 9669 9494
rect 9340 9461 9669 9477
rect 10227 9494 10480 9510
rect 10227 9477 10240 9494
rect 10257 9477 10288 9494
rect 10305 9477 10336 9494
rect 10353 9477 10384 9494
rect 10401 9477 10432 9494
rect 10449 9477 10480 9494
rect 10227 9461 10480 9477
rect 968 9338 1011 9347
rect 1636 9340 1666 9341
rect 1722 9340 1756 9343
rect 968 9334 980 9338
rect 916 9331 980 9334
rect 916 9314 924 9331
rect 941 9314 980 9331
rect 916 9312 980 9314
rect 1006 9312 1011 9338
rect 916 9310 1011 9312
rect 1633 9338 1700 9340
rect 1633 9312 1638 9338
rect 1664 9328 1700 9338
rect 1664 9312 1680 9328
rect 1633 9311 1680 9312
rect 1697 9311 1700 9328
rect 978 9309 1008 9310
rect 1633 9303 1700 9311
rect 1721 9338 1756 9340
rect 1721 9312 1724 9338
rect 1750 9312 1756 9338
rect 1855 9338 1898 9347
rect 2506 9340 2536 9341
rect 2592 9340 2626 9343
rect 1855 9334 1867 9338
rect 1721 9310 1756 9312
rect 1803 9331 1867 9334
rect 1803 9314 1811 9331
rect 1828 9314 1867 9331
rect 1803 9312 1867 9314
rect 1893 9312 1898 9338
rect 1803 9310 1898 9312
rect 2503 9338 2570 9340
rect 2503 9312 2508 9338
rect 2534 9328 2570 9338
rect 2534 9312 2550 9328
rect 2503 9311 2550 9312
rect 2567 9311 2570 9328
rect 1722 9307 1756 9310
rect 1865 9309 1895 9310
rect 2503 9303 2570 9311
rect 2591 9338 2626 9340
rect 2591 9312 2594 9338
rect 2620 9312 2626 9338
rect 2725 9338 2768 9347
rect 3123 9340 3153 9341
rect 2725 9334 2737 9338
rect 2591 9310 2626 9312
rect 2673 9331 2737 9334
rect 2673 9314 2681 9331
rect 2698 9314 2737 9331
rect 2673 9312 2737 9314
rect 2763 9312 2768 9338
rect 2673 9310 2768 9312
rect 3120 9338 3163 9340
rect 3120 9312 3125 9338
rect 3151 9330 3163 9338
rect 3244 9338 3287 9347
rect 3244 9334 3256 9338
rect 3153 9313 3163 9330
rect 3151 9312 3163 9313
rect 2592 9307 2626 9310
rect 2735 9309 2765 9310
rect 3120 9303 3163 9312
rect 3192 9331 3256 9334
rect 3192 9314 3200 9331
rect 3217 9314 3256 9331
rect 3192 9312 3256 9314
rect 3282 9312 3287 9338
rect 3192 9310 3287 9312
rect 7991 9338 8034 9347
rect 8125 9340 8155 9341
rect 7991 9312 7996 9338
rect 8022 9334 8034 9338
rect 8115 9338 8158 9340
rect 8022 9331 8086 9334
rect 8022 9314 8061 9331
rect 8078 9314 8086 9331
rect 8022 9312 8086 9314
rect 7991 9310 8086 9312
rect 8115 9330 8127 9338
rect 8115 9313 8125 9330
rect 8115 9312 8127 9313
rect 8153 9312 8158 9338
rect 3254 9309 3284 9310
rect 7994 9309 8024 9310
rect 8115 9303 8158 9312
rect 8510 9338 8553 9347
rect 8510 9312 8515 9338
rect 8541 9334 8553 9338
rect 8652 9340 8686 9343
rect 8742 9340 8772 9341
rect 8652 9338 8687 9340
rect 8541 9331 8605 9334
rect 8541 9314 8580 9331
rect 8597 9314 8605 9331
rect 8541 9312 8605 9314
rect 8510 9310 8605 9312
rect 8652 9312 8658 9338
rect 8684 9312 8687 9338
rect 8652 9310 8687 9312
rect 8708 9338 8775 9340
rect 8708 9328 8744 9338
rect 8708 9311 8711 9328
rect 8728 9312 8744 9328
rect 8770 9312 8775 9338
rect 8728 9311 8775 9312
rect 8513 9309 8543 9310
rect 8652 9307 8686 9310
rect 8708 9303 8775 9311
rect 9380 9338 9423 9347
rect 9380 9312 9385 9338
rect 9411 9334 9423 9338
rect 9522 9340 9556 9343
rect 9612 9340 9642 9341
rect 9522 9338 9557 9340
rect 9411 9331 9475 9334
rect 9411 9314 9450 9331
rect 9467 9314 9475 9331
rect 9411 9312 9475 9314
rect 9380 9310 9475 9312
rect 9522 9312 9528 9338
rect 9554 9312 9557 9338
rect 9522 9310 9557 9312
rect 9578 9338 9645 9340
rect 9578 9328 9614 9338
rect 9578 9311 9581 9328
rect 9598 9312 9614 9328
rect 9640 9312 9645 9338
rect 9598 9311 9645 9312
rect 9383 9309 9413 9310
rect 9522 9307 9556 9310
rect 9578 9303 9645 9311
rect 10267 9338 10310 9347
rect 10267 9312 10272 9338
rect 10298 9334 10310 9338
rect 10298 9331 10362 9334
rect 10298 9314 10337 9331
rect 10354 9314 10362 9331
rect 10298 9312 10362 9314
rect 10267 9310 10362 9312
rect 10270 9309 10300 9310
rect 798 9161 1051 9177
rect 798 9144 829 9161
rect 846 9144 877 9161
rect 894 9144 925 9161
rect 942 9144 973 9161
rect 990 9144 1021 9161
rect 1038 9144 1051 9161
rect 798 9128 1051 9144
rect 1609 9161 1938 9177
rect 1609 9144 1640 9161
rect 1657 9144 1688 9161
rect 1733 9144 1764 9161
rect 1781 9144 1812 9161
rect 1829 9144 1860 9161
rect 1877 9144 1908 9161
rect 1925 9144 1938 9161
rect 1609 9128 1938 9144
rect 2479 9161 2808 9177
rect 2479 9144 2510 9161
rect 2527 9144 2558 9161
rect 2603 9144 2634 9161
rect 2651 9144 2682 9161
rect 2699 9144 2730 9161
rect 2747 9144 2778 9161
rect 2795 9144 2808 9161
rect 2479 9128 2808 9144
rect 3074 9161 3327 9177
rect 3074 9144 3105 9161
rect 3122 9144 3153 9161
rect 3170 9144 3201 9161
rect 3218 9144 3249 9161
rect 3266 9144 3297 9161
rect 3314 9144 3327 9161
rect 3074 9128 3327 9144
rect 7951 9161 8204 9177
rect 7951 9144 7964 9161
rect 7981 9144 8012 9161
rect 8029 9144 8060 9161
rect 8077 9144 8108 9161
rect 8125 9144 8156 9161
rect 8173 9144 8204 9161
rect 7951 9128 8204 9144
rect 8470 9161 8799 9177
rect 8470 9144 8483 9161
rect 8500 9144 8531 9161
rect 8548 9144 8579 9161
rect 8596 9144 8627 9161
rect 8644 9144 8675 9161
rect 8720 9144 8751 9161
rect 8768 9144 8799 9161
rect 8470 9128 8799 9144
rect 9340 9161 9669 9177
rect 9340 9144 9353 9161
rect 9370 9144 9401 9161
rect 9418 9144 9449 9161
rect 9466 9144 9497 9161
rect 9514 9144 9545 9161
rect 9590 9144 9621 9161
rect 9638 9144 9669 9161
rect 9340 9128 9669 9144
rect 10227 9161 10480 9177
rect 10227 9144 10240 9161
rect 10257 9144 10288 9161
rect 10305 9144 10336 9161
rect 10353 9144 10384 9161
rect 10401 9144 10432 9161
rect 10449 9144 10480 9161
rect 10227 9128 10480 9144
rect 798 -1350 1051 -1334
rect 798 -1367 829 -1350
rect 846 -1367 877 -1350
rect 894 -1367 925 -1350
rect 942 -1367 973 -1350
rect 990 -1367 1021 -1350
rect 1038 -1367 1051 -1350
rect 798 -1383 1051 -1367
rect 1609 -1350 1938 -1334
rect 1609 -1367 1640 -1350
rect 1657 -1367 1688 -1350
rect 1733 -1367 1764 -1350
rect 1781 -1367 1812 -1350
rect 1829 -1367 1860 -1350
rect 1877 -1367 1908 -1350
rect 1925 -1367 1938 -1350
rect 1609 -1383 1938 -1367
rect 2479 -1350 2808 -1334
rect 2479 -1367 2510 -1350
rect 2527 -1367 2558 -1350
rect 2603 -1367 2634 -1350
rect 2651 -1367 2682 -1350
rect 2699 -1367 2730 -1350
rect 2747 -1367 2778 -1350
rect 2795 -1367 2808 -1350
rect 2479 -1383 2808 -1367
rect 3074 -1350 3327 -1334
rect 3074 -1367 3105 -1350
rect 3122 -1367 3153 -1350
rect 3170 -1367 3201 -1350
rect 3218 -1367 3249 -1350
rect 3266 -1367 3297 -1350
rect 3314 -1367 3327 -1350
rect 3074 -1383 3327 -1367
rect 7951 -1350 8204 -1334
rect 7951 -1367 7964 -1350
rect 7981 -1367 8012 -1350
rect 8029 -1367 8060 -1350
rect 8077 -1367 8108 -1350
rect 8125 -1367 8156 -1350
rect 8173 -1367 8204 -1350
rect 7951 -1383 8204 -1367
rect 8470 -1350 8799 -1334
rect 8470 -1367 8483 -1350
rect 8500 -1367 8531 -1350
rect 8548 -1367 8579 -1350
rect 8596 -1367 8627 -1350
rect 8644 -1367 8675 -1350
rect 8720 -1367 8751 -1350
rect 8768 -1367 8799 -1350
rect 8470 -1383 8799 -1367
rect 9340 -1350 9669 -1334
rect 9340 -1367 9353 -1350
rect 9370 -1367 9401 -1350
rect 9418 -1367 9449 -1350
rect 9466 -1367 9497 -1350
rect 9514 -1367 9545 -1350
rect 9590 -1367 9621 -1350
rect 9638 -1367 9669 -1350
rect 9340 -1383 9669 -1367
rect 10227 -1350 10480 -1334
rect 10227 -1367 10240 -1350
rect 10257 -1367 10288 -1350
rect 10305 -1367 10336 -1350
rect 10353 -1367 10384 -1350
rect 10401 -1367 10432 -1350
rect 10449 -1367 10480 -1350
rect 10227 -1383 10480 -1367
rect 978 -1516 1008 -1515
rect 916 -1518 1011 -1516
rect 916 -1520 980 -1518
rect 916 -1537 924 -1520
rect 941 -1537 980 -1520
rect 916 -1540 980 -1537
rect 968 -1544 980 -1540
rect 1006 -1544 1011 -1518
rect 968 -1553 1011 -1544
rect 1633 -1517 1700 -1509
rect 1722 -1516 1756 -1513
rect 1865 -1516 1895 -1515
rect 1633 -1518 1680 -1517
rect 1633 -1544 1638 -1518
rect 1664 -1534 1680 -1518
rect 1697 -1534 1700 -1517
rect 1664 -1544 1700 -1534
rect 1633 -1546 1700 -1544
rect 1721 -1518 1756 -1516
rect 1721 -1544 1724 -1518
rect 1750 -1544 1756 -1518
rect 1803 -1518 1898 -1516
rect 1803 -1520 1867 -1518
rect 1803 -1537 1811 -1520
rect 1828 -1537 1867 -1520
rect 1803 -1540 1867 -1537
rect 1721 -1546 1756 -1544
rect 1636 -1547 1666 -1546
rect 1722 -1549 1756 -1546
rect 1855 -1544 1867 -1540
rect 1893 -1544 1898 -1518
rect 1855 -1553 1898 -1544
rect 2503 -1517 2570 -1509
rect 2592 -1516 2626 -1513
rect 2735 -1516 2765 -1515
rect 2503 -1518 2550 -1517
rect 2503 -1544 2508 -1518
rect 2534 -1534 2550 -1518
rect 2567 -1534 2570 -1517
rect 2534 -1544 2570 -1534
rect 2503 -1546 2570 -1544
rect 2591 -1518 2626 -1516
rect 2591 -1544 2594 -1518
rect 2620 -1544 2626 -1518
rect 2673 -1518 2768 -1516
rect 2673 -1520 2737 -1518
rect 2673 -1537 2681 -1520
rect 2698 -1537 2737 -1520
rect 2673 -1540 2737 -1537
rect 2591 -1546 2626 -1544
rect 2506 -1547 2536 -1546
rect 2592 -1549 2626 -1546
rect 2725 -1544 2737 -1540
rect 2763 -1544 2768 -1518
rect 2725 -1553 2768 -1544
rect 3120 -1518 3163 -1509
rect 3254 -1516 3284 -1515
rect 7994 -1516 8024 -1515
rect 3120 -1544 3125 -1518
rect 3151 -1519 3163 -1518
rect 3153 -1536 3163 -1519
rect 3151 -1544 3163 -1536
rect 3192 -1518 3287 -1516
rect 3192 -1520 3256 -1518
rect 3192 -1537 3200 -1520
rect 3217 -1537 3256 -1520
rect 3192 -1540 3256 -1537
rect 3120 -1546 3163 -1544
rect 3244 -1544 3256 -1540
rect 3282 -1544 3287 -1518
rect 3123 -1547 3153 -1546
rect 3244 -1553 3287 -1544
rect 7991 -1518 8086 -1516
rect 7991 -1544 7996 -1518
rect 8022 -1520 8086 -1518
rect 8022 -1537 8061 -1520
rect 8078 -1537 8086 -1520
rect 8022 -1540 8086 -1537
rect 8115 -1518 8158 -1509
rect 8513 -1516 8543 -1515
rect 8652 -1516 8686 -1513
rect 8115 -1519 8127 -1518
rect 8115 -1536 8125 -1519
rect 8022 -1544 8034 -1540
rect 7991 -1553 8034 -1544
rect 8115 -1544 8127 -1536
rect 8153 -1544 8158 -1518
rect 8115 -1546 8158 -1544
rect 8510 -1518 8605 -1516
rect 8510 -1544 8515 -1518
rect 8541 -1520 8605 -1518
rect 8541 -1537 8580 -1520
rect 8597 -1537 8605 -1520
rect 8541 -1540 8605 -1537
rect 8652 -1518 8687 -1516
rect 8541 -1544 8553 -1540
rect 8125 -1547 8155 -1546
rect 8510 -1553 8553 -1544
rect 8652 -1544 8658 -1518
rect 8684 -1544 8687 -1518
rect 8652 -1546 8687 -1544
rect 8708 -1517 8775 -1509
rect 9383 -1516 9413 -1515
rect 9522 -1516 9556 -1513
rect 8708 -1534 8711 -1517
rect 8728 -1518 8775 -1517
rect 8728 -1534 8744 -1518
rect 8708 -1544 8744 -1534
rect 8770 -1544 8775 -1518
rect 8708 -1546 8775 -1544
rect 9380 -1518 9475 -1516
rect 9380 -1544 9385 -1518
rect 9411 -1520 9475 -1518
rect 9411 -1537 9450 -1520
rect 9467 -1537 9475 -1520
rect 9411 -1540 9475 -1537
rect 9522 -1518 9557 -1516
rect 9411 -1544 9423 -1540
rect 8652 -1549 8686 -1546
rect 8742 -1547 8772 -1546
rect 9380 -1553 9423 -1544
rect 9522 -1544 9528 -1518
rect 9554 -1544 9557 -1518
rect 9522 -1546 9557 -1544
rect 9578 -1517 9645 -1509
rect 10270 -1516 10300 -1515
rect 9578 -1534 9581 -1517
rect 9598 -1518 9645 -1517
rect 9598 -1534 9614 -1518
rect 9578 -1544 9614 -1534
rect 9640 -1544 9645 -1518
rect 9578 -1546 9645 -1544
rect 10267 -1518 10362 -1516
rect 10267 -1544 10272 -1518
rect 10298 -1520 10362 -1518
rect 10298 -1537 10337 -1520
rect 10354 -1537 10362 -1520
rect 10298 -1540 10362 -1537
rect 10298 -1544 10310 -1540
rect 9522 -1549 9556 -1546
rect 9612 -1547 9642 -1546
rect 10267 -1553 10310 -1544
rect 798 -1683 1051 -1667
rect 798 -1700 829 -1683
rect 846 -1700 877 -1683
rect 894 -1700 925 -1683
rect 942 -1700 973 -1683
rect 990 -1700 1021 -1683
rect 1038 -1700 1051 -1683
rect 798 -1716 1051 -1700
rect 1609 -1683 1938 -1667
rect 1609 -1700 1640 -1683
rect 1657 -1700 1688 -1683
rect 1733 -1700 1764 -1683
rect 1781 -1700 1812 -1683
rect 1829 -1700 1860 -1683
rect 1877 -1700 1908 -1683
rect 1925 -1700 1938 -1683
rect 1609 -1716 1938 -1700
rect 2479 -1683 2808 -1667
rect 2479 -1700 2510 -1683
rect 2527 -1700 2558 -1683
rect 2603 -1700 2634 -1683
rect 2651 -1700 2682 -1683
rect 2699 -1700 2730 -1683
rect 2747 -1700 2778 -1683
rect 2795 -1700 2808 -1683
rect 2479 -1716 2808 -1700
rect 3074 -1683 3327 -1667
rect 3074 -1700 3105 -1683
rect 3122 -1700 3153 -1683
rect 3170 -1700 3201 -1683
rect 3218 -1700 3249 -1683
rect 3266 -1700 3297 -1683
rect 3314 -1700 3327 -1683
rect 3074 -1716 3327 -1700
rect 7951 -1683 8204 -1667
rect 7951 -1700 7964 -1683
rect 7981 -1700 8012 -1683
rect 8029 -1700 8060 -1683
rect 8077 -1700 8108 -1683
rect 8125 -1700 8156 -1683
rect 8173 -1700 8204 -1683
rect 3614 -1718 3642 -1715
rect 3614 -1744 3616 -1718
rect 3614 -1748 3642 -1744
rect 7636 -1718 7664 -1715
rect 7951 -1716 8204 -1700
rect 8470 -1683 8799 -1667
rect 8470 -1700 8483 -1683
rect 8500 -1700 8531 -1683
rect 8548 -1700 8579 -1683
rect 8596 -1700 8627 -1683
rect 8644 -1700 8675 -1683
rect 8720 -1700 8751 -1683
rect 8768 -1700 8799 -1683
rect 8470 -1716 8799 -1700
rect 9340 -1683 9669 -1667
rect 9340 -1700 9353 -1683
rect 9370 -1700 9401 -1683
rect 9418 -1700 9449 -1683
rect 9466 -1700 9497 -1683
rect 9514 -1700 9545 -1683
rect 9590 -1700 9621 -1683
rect 9638 -1700 9669 -1683
rect 9340 -1716 9669 -1700
rect 10227 -1683 10480 -1667
rect 10227 -1700 10240 -1683
rect 10257 -1700 10288 -1683
rect 10305 -1700 10336 -1683
rect 10353 -1700 10384 -1683
rect 10401 -1700 10432 -1683
rect 10449 -1700 10480 -1683
rect 10227 -1716 10480 -1700
rect 7662 -1744 7664 -1718
rect 7636 -1748 7664 -1744
<< via1 >>
rect 3616 9534 3642 9538
rect 3616 9517 3620 9534
rect 3620 9517 3637 9534
rect 3637 9517 3642 9534
rect 3616 9512 3642 9517
rect 7636 9534 7662 9538
rect 7636 9517 7641 9534
rect 7641 9517 7658 9534
rect 7658 9517 7662 9534
rect 7636 9512 7662 9517
rect 980 9312 1006 9338
rect 1638 9312 1664 9338
rect 1724 9332 1750 9338
rect 1724 9315 1727 9332
rect 1727 9315 1744 9332
rect 1744 9315 1750 9332
rect 1724 9312 1750 9315
rect 1867 9312 1893 9338
rect 2508 9312 2534 9338
rect 2594 9332 2620 9338
rect 2594 9315 2597 9332
rect 2597 9315 2614 9332
rect 2614 9315 2620 9332
rect 2594 9312 2620 9315
rect 2737 9312 2763 9338
rect 3125 9330 3151 9338
rect 3125 9313 3136 9330
rect 3136 9313 3151 9330
rect 3125 9312 3151 9313
rect 3256 9312 3282 9338
rect 7996 9312 8022 9338
rect 8127 9330 8153 9338
rect 8127 9313 8142 9330
rect 8142 9313 8153 9330
rect 8127 9312 8153 9313
rect 8515 9312 8541 9338
rect 8658 9332 8684 9338
rect 8658 9315 8664 9332
rect 8664 9315 8681 9332
rect 8681 9315 8684 9332
rect 8658 9312 8684 9315
rect 8744 9312 8770 9338
rect 9385 9312 9411 9338
rect 9528 9332 9554 9338
rect 9528 9315 9534 9332
rect 9534 9315 9551 9332
rect 9551 9315 9554 9332
rect 9528 9312 9554 9315
rect 9614 9312 9640 9338
rect 10272 9312 10298 9338
rect 980 -1544 1006 -1518
rect 1638 -1544 1664 -1518
rect 1724 -1521 1750 -1518
rect 1724 -1538 1727 -1521
rect 1727 -1538 1744 -1521
rect 1744 -1538 1750 -1521
rect 1724 -1544 1750 -1538
rect 1867 -1544 1893 -1518
rect 2508 -1544 2534 -1518
rect 2594 -1521 2620 -1518
rect 2594 -1538 2597 -1521
rect 2597 -1538 2614 -1521
rect 2614 -1538 2620 -1521
rect 2594 -1544 2620 -1538
rect 2737 -1544 2763 -1518
rect 3125 -1519 3151 -1518
rect 3125 -1536 3136 -1519
rect 3136 -1536 3151 -1519
rect 3125 -1544 3151 -1536
rect 3256 -1544 3282 -1518
rect 7996 -1544 8022 -1518
rect 8127 -1519 8153 -1518
rect 8127 -1536 8142 -1519
rect 8142 -1536 8153 -1519
rect 8127 -1544 8153 -1536
rect 8515 -1544 8541 -1518
rect 8658 -1521 8684 -1518
rect 8658 -1538 8664 -1521
rect 8664 -1538 8681 -1521
rect 8681 -1538 8684 -1521
rect 8658 -1544 8684 -1538
rect 8744 -1544 8770 -1518
rect 9385 -1544 9411 -1518
rect 9528 -1521 9554 -1518
rect 9528 -1538 9534 -1521
rect 9534 -1538 9551 -1521
rect 9551 -1538 9554 -1521
rect 9528 -1544 9554 -1538
rect 9614 -1544 9640 -1518
rect 10272 -1544 10298 -1518
rect 3616 -1723 3642 -1718
rect 3616 -1740 3620 -1723
rect 3620 -1740 3637 -1723
rect 3637 -1740 3642 -1723
rect 3616 -1744 3642 -1740
rect 7636 -1723 7662 -1718
rect 7636 -1740 7641 -1723
rect 7641 -1740 7658 -1723
rect 7658 -1740 7662 -1723
rect 7636 -1744 7662 -1740
<< metal2 >>
rect 3613 9539 3645 9544
rect 3613 9511 3615 9539
rect 3643 9511 3645 9539
rect 3613 9506 3645 9511
rect 7633 9539 7665 9544
rect 7633 9511 7635 9539
rect 7663 9511 7665 9539
rect 7633 9506 7665 9511
rect 975 9339 1011 9344
rect 975 9311 979 9339
rect 1007 9311 1011 9339
rect 975 9306 1011 9311
rect 1633 9339 1669 9344
rect 1633 9311 1637 9339
rect 1665 9311 1669 9339
rect 1633 9306 1669 9311
rect 1718 9339 1756 9343
rect 1718 9311 1723 9339
rect 1751 9311 1756 9339
rect 1718 9307 1756 9311
rect 1862 9339 1898 9344
rect 1862 9311 1866 9339
rect 1894 9311 1898 9339
rect 1862 9306 1898 9311
rect 2503 9339 2539 9344
rect 2503 9311 2507 9339
rect 2535 9311 2539 9339
rect 2503 9306 2539 9311
rect 2588 9339 2626 9343
rect 2588 9311 2593 9339
rect 2621 9311 2626 9339
rect 2588 9307 2626 9311
rect 2732 9339 2768 9344
rect 2732 9311 2736 9339
rect 2764 9311 2768 9339
rect 2732 9306 2768 9311
rect 3120 9339 3156 9344
rect 3120 9311 3124 9339
rect 3152 9311 3156 9339
rect 3120 9306 3156 9311
rect 3251 9339 3287 9344
rect 3251 9311 3255 9339
rect 3283 9311 3287 9339
rect 3251 9306 3287 9311
rect 7991 9339 8027 9344
rect 7991 9311 7995 9339
rect 8023 9311 8027 9339
rect 7991 9306 8027 9311
rect 8122 9339 8158 9344
rect 8122 9311 8126 9339
rect 8154 9311 8158 9339
rect 8122 9306 8158 9311
rect 8510 9339 8546 9344
rect 8510 9311 8514 9339
rect 8542 9311 8546 9339
rect 8510 9306 8546 9311
rect 8652 9339 8690 9343
rect 8652 9311 8657 9339
rect 8685 9311 8690 9339
rect 8652 9307 8690 9311
rect 8739 9339 8775 9344
rect 8739 9311 8743 9339
rect 8771 9311 8775 9339
rect 8739 9306 8775 9311
rect 9380 9339 9416 9344
rect 9380 9311 9384 9339
rect 9412 9311 9416 9339
rect 9380 9306 9416 9311
rect 9522 9339 9560 9343
rect 9522 9311 9527 9339
rect 9555 9311 9560 9339
rect 9522 9307 9560 9311
rect 9609 9339 9645 9344
rect 9609 9311 9613 9339
rect 9641 9311 9645 9339
rect 9609 9306 9645 9311
rect 10267 9339 10303 9344
rect 10267 9311 10271 9339
rect 10299 9311 10303 9339
rect 10267 9306 10303 9311
rect 975 -1517 1011 -1512
rect 975 -1545 979 -1517
rect 1007 -1545 1011 -1517
rect 975 -1550 1011 -1545
rect 1633 -1517 1669 -1512
rect 1633 -1545 1637 -1517
rect 1665 -1545 1669 -1517
rect 1633 -1550 1669 -1545
rect 1718 -1517 1756 -1513
rect 1718 -1545 1723 -1517
rect 1751 -1545 1756 -1517
rect 1718 -1549 1756 -1545
rect 1862 -1517 1898 -1512
rect 1862 -1545 1866 -1517
rect 1894 -1545 1898 -1517
rect 1862 -1550 1898 -1545
rect 2503 -1517 2539 -1512
rect 2503 -1545 2507 -1517
rect 2535 -1545 2539 -1517
rect 2503 -1550 2539 -1545
rect 2588 -1517 2626 -1513
rect 2588 -1545 2593 -1517
rect 2621 -1545 2626 -1517
rect 2588 -1549 2626 -1545
rect 2732 -1517 2768 -1512
rect 2732 -1545 2736 -1517
rect 2764 -1545 2768 -1517
rect 2732 -1550 2768 -1545
rect 3120 -1517 3156 -1512
rect 3120 -1545 3124 -1517
rect 3152 -1545 3156 -1517
rect 3120 -1550 3156 -1545
rect 3251 -1517 3287 -1512
rect 3251 -1545 3255 -1517
rect 3283 -1545 3287 -1517
rect 3251 -1550 3287 -1545
rect 7991 -1517 8027 -1512
rect 7991 -1545 7995 -1517
rect 8023 -1545 8027 -1517
rect 7991 -1550 8027 -1545
rect 8122 -1517 8158 -1512
rect 8122 -1545 8126 -1517
rect 8154 -1545 8158 -1517
rect 8122 -1550 8158 -1545
rect 8510 -1517 8546 -1512
rect 8510 -1545 8514 -1517
rect 8542 -1545 8546 -1517
rect 8510 -1550 8546 -1545
rect 8652 -1517 8690 -1513
rect 8652 -1545 8657 -1517
rect 8685 -1545 8690 -1517
rect 8652 -1549 8690 -1545
rect 8739 -1517 8775 -1512
rect 8739 -1545 8743 -1517
rect 8771 -1545 8775 -1517
rect 8739 -1550 8775 -1545
rect 9380 -1517 9416 -1512
rect 9380 -1545 9384 -1517
rect 9412 -1545 9416 -1517
rect 9380 -1550 9416 -1545
rect 9522 -1517 9560 -1513
rect 9522 -1545 9527 -1517
rect 9555 -1545 9560 -1517
rect 9522 -1549 9560 -1545
rect 9609 -1517 9645 -1512
rect 9609 -1545 9613 -1517
rect 9641 -1545 9645 -1517
rect 9609 -1550 9645 -1545
rect 10267 -1517 10303 -1512
rect 10267 -1545 10271 -1517
rect 10299 -1545 10303 -1517
rect 10267 -1550 10303 -1545
rect 3613 -1717 3645 -1712
rect 3613 -1745 3615 -1717
rect 3643 -1745 3645 -1717
rect 3613 -1750 3645 -1745
rect 7633 -1717 7665 -1712
rect 7633 -1745 7635 -1717
rect 7663 -1745 7665 -1717
rect 7633 -1750 7665 -1745
<< via2 >>
rect 3615 9538 3643 9539
rect 3615 9512 3616 9538
rect 3616 9512 3642 9538
rect 3642 9512 3643 9538
rect 3615 9511 3643 9512
rect 7635 9538 7663 9539
rect 7635 9512 7636 9538
rect 7636 9512 7662 9538
rect 7662 9512 7663 9538
rect 7635 9511 7663 9512
rect 979 9338 1007 9339
rect 979 9312 980 9338
rect 980 9312 1006 9338
rect 1006 9312 1007 9338
rect 979 9311 1007 9312
rect 1637 9338 1665 9339
rect 1637 9312 1638 9338
rect 1638 9312 1664 9338
rect 1664 9312 1665 9338
rect 1637 9311 1665 9312
rect 1723 9338 1751 9339
rect 1723 9312 1724 9338
rect 1724 9312 1750 9338
rect 1750 9312 1751 9338
rect 1723 9311 1751 9312
rect 1866 9338 1894 9339
rect 1866 9312 1867 9338
rect 1867 9312 1893 9338
rect 1893 9312 1894 9338
rect 1866 9311 1894 9312
rect 2507 9338 2535 9339
rect 2507 9312 2508 9338
rect 2508 9312 2534 9338
rect 2534 9312 2535 9338
rect 2507 9311 2535 9312
rect 2593 9338 2621 9339
rect 2593 9312 2594 9338
rect 2594 9312 2620 9338
rect 2620 9312 2621 9338
rect 2593 9311 2621 9312
rect 2736 9338 2764 9339
rect 2736 9312 2737 9338
rect 2737 9312 2763 9338
rect 2763 9312 2764 9338
rect 2736 9311 2764 9312
rect 3124 9338 3152 9339
rect 3124 9312 3125 9338
rect 3125 9312 3151 9338
rect 3151 9312 3152 9338
rect 3124 9311 3152 9312
rect 3255 9338 3283 9339
rect 3255 9312 3256 9338
rect 3256 9312 3282 9338
rect 3282 9312 3283 9338
rect 3255 9311 3283 9312
rect 7995 9338 8023 9339
rect 7995 9312 7996 9338
rect 7996 9312 8022 9338
rect 8022 9312 8023 9338
rect 7995 9311 8023 9312
rect 8126 9338 8154 9339
rect 8126 9312 8127 9338
rect 8127 9312 8153 9338
rect 8153 9312 8154 9338
rect 8126 9311 8154 9312
rect 8514 9338 8542 9339
rect 8514 9312 8515 9338
rect 8515 9312 8541 9338
rect 8541 9312 8542 9338
rect 8514 9311 8542 9312
rect 8657 9338 8685 9339
rect 8657 9312 8658 9338
rect 8658 9312 8684 9338
rect 8684 9312 8685 9338
rect 8657 9311 8685 9312
rect 8743 9338 8771 9339
rect 8743 9312 8744 9338
rect 8744 9312 8770 9338
rect 8770 9312 8771 9338
rect 8743 9311 8771 9312
rect 9384 9338 9412 9339
rect 9384 9312 9385 9338
rect 9385 9312 9411 9338
rect 9411 9312 9412 9338
rect 9384 9311 9412 9312
rect 9527 9338 9555 9339
rect 9527 9312 9528 9338
rect 9528 9312 9554 9338
rect 9554 9312 9555 9338
rect 9527 9311 9555 9312
rect 9613 9338 9641 9339
rect 9613 9312 9614 9338
rect 9614 9312 9640 9338
rect 9640 9312 9641 9338
rect 9613 9311 9641 9312
rect 10271 9338 10299 9339
rect 10271 9312 10272 9338
rect 10272 9312 10298 9338
rect 10298 9312 10299 9338
rect 10271 9311 10299 9312
rect 979 -1518 1007 -1517
rect 979 -1544 980 -1518
rect 980 -1544 1006 -1518
rect 1006 -1544 1007 -1518
rect 979 -1545 1007 -1544
rect 1637 -1518 1665 -1517
rect 1637 -1544 1638 -1518
rect 1638 -1544 1664 -1518
rect 1664 -1544 1665 -1518
rect 1637 -1545 1665 -1544
rect 1723 -1518 1751 -1517
rect 1723 -1544 1724 -1518
rect 1724 -1544 1750 -1518
rect 1750 -1544 1751 -1518
rect 1723 -1545 1751 -1544
rect 1866 -1518 1894 -1517
rect 1866 -1544 1867 -1518
rect 1867 -1544 1893 -1518
rect 1893 -1544 1894 -1518
rect 1866 -1545 1894 -1544
rect 2507 -1518 2535 -1517
rect 2507 -1544 2508 -1518
rect 2508 -1544 2534 -1518
rect 2534 -1544 2535 -1518
rect 2507 -1545 2535 -1544
rect 2593 -1518 2621 -1517
rect 2593 -1544 2594 -1518
rect 2594 -1544 2620 -1518
rect 2620 -1544 2621 -1518
rect 2593 -1545 2621 -1544
rect 2736 -1518 2764 -1517
rect 2736 -1544 2737 -1518
rect 2737 -1544 2763 -1518
rect 2763 -1544 2764 -1518
rect 2736 -1545 2764 -1544
rect 3124 -1518 3152 -1517
rect 3124 -1544 3125 -1518
rect 3125 -1544 3151 -1518
rect 3151 -1544 3152 -1518
rect 3124 -1545 3152 -1544
rect 3255 -1518 3283 -1517
rect 3255 -1544 3256 -1518
rect 3256 -1544 3282 -1518
rect 3282 -1544 3283 -1518
rect 3255 -1545 3283 -1544
rect 7995 -1518 8023 -1517
rect 7995 -1544 7996 -1518
rect 7996 -1544 8022 -1518
rect 8022 -1544 8023 -1518
rect 7995 -1545 8023 -1544
rect 8126 -1518 8154 -1517
rect 8126 -1544 8127 -1518
rect 8127 -1544 8153 -1518
rect 8153 -1544 8154 -1518
rect 8126 -1545 8154 -1544
rect 8514 -1518 8542 -1517
rect 8514 -1544 8515 -1518
rect 8515 -1544 8541 -1518
rect 8541 -1544 8542 -1518
rect 8514 -1545 8542 -1544
rect 8657 -1518 8685 -1517
rect 8657 -1544 8658 -1518
rect 8658 -1544 8684 -1518
rect 8684 -1544 8685 -1518
rect 8657 -1545 8685 -1544
rect 8743 -1518 8771 -1517
rect 8743 -1544 8744 -1518
rect 8744 -1544 8770 -1518
rect 8770 -1544 8771 -1518
rect 8743 -1545 8771 -1544
rect 9384 -1518 9412 -1517
rect 9384 -1544 9385 -1518
rect 9385 -1544 9411 -1518
rect 9411 -1544 9412 -1518
rect 9384 -1545 9412 -1544
rect 9527 -1518 9555 -1517
rect 9527 -1544 9528 -1518
rect 9528 -1544 9554 -1518
rect 9554 -1544 9555 -1518
rect 9527 -1545 9555 -1544
rect 9613 -1518 9641 -1517
rect 9613 -1544 9614 -1518
rect 9614 -1544 9640 -1518
rect 9640 -1544 9641 -1518
rect 9613 -1545 9641 -1544
rect 10271 -1518 10299 -1517
rect 10271 -1544 10272 -1518
rect 10272 -1544 10298 -1518
rect 10298 -1544 10299 -1518
rect 10271 -1545 10299 -1544
rect 3615 -1718 3643 -1717
rect 3615 -1744 3616 -1718
rect 3616 -1744 3642 -1718
rect 3642 -1744 3643 -1718
rect 3615 -1745 3643 -1744
rect 7635 -1718 7663 -1717
rect 7635 -1744 7636 -1718
rect 7636 -1744 7662 -1718
rect 7662 -1744 7663 -1718
rect 7635 -1745 7663 -1744
<< metal3 >>
rect -2093 9591 3019 12619
rect 3075 9591 5604 12619
rect 5674 9591 8203 12619
rect 8259 9591 13371 12619
rect 3602 9541 3651 9591
rect 968 9341 1017 9351
rect 968 9309 977 9341
rect 1009 9309 1017 9341
rect 968 9299 1017 9309
rect 1057 9100 1585 9528
rect 3602 9509 3614 9541
rect 3646 9509 3651 9541
rect 3602 9503 3651 9509
rect 7627 9541 7676 9591
rect 7627 9509 7632 9541
rect 7664 9509 7676 9541
rect 7627 9503 7676 9509
rect 1627 9341 1676 9351
rect 1627 9309 1635 9341
rect 1667 9309 1676 9341
rect 1627 9299 1676 9309
rect 1711 9341 1763 9350
rect 1711 9309 1721 9341
rect 1753 9309 1763 9341
rect 1711 9301 1763 9309
rect 1855 9341 1904 9351
rect 1855 9309 1864 9341
rect 1896 9309 1904 9341
rect 1855 9299 1904 9309
rect 1936 9224 2464 9452
rect 2497 9341 2546 9351
rect 2497 9309 2505 9341
rect 2537 9309 2546 9341
rect 2497 9299 2546 9309
rect 2581 9341 2633 9350
rect 2581 9309 2591 9341
rect 2623 9309 2633 9341
rect 2581 9301 2633 9309
rect 2725 9341 2774 9351
rect 2725 9309 2734 9341
rect 2766 9309 2774 9341
rect 2725 9299 2774 9309
rect 2806 9217 3084 9445
rect 3114 9341 3163 9351
rect 3114 9309 3122 9341
rect 3154 9309 3163 9341
rect 3114 9299 3163 9309
rect 3244 9345 3286 9351
rect 7992 9345 8034 9351
rect 3244 9341 3293 9345
rect 3244 9309 3253 9341
rect 3285 9309 3293 9341
rect 3244 9299 3293 9309
rect 7985 9341 8034 9345
rect 7985 9309 7993 9341
rect 8025 9309 8034 9341
rect 7985 9299 8034 9309
rect 8115 9341 8164 9351
rect 8115 9309 8124 9341
rect 8156 9309 8164 9341
rect 8115 9299 8164 9309
rect 8194 9217 8472 9445
rect 8504 9341 8553 9351
rect 8504 9309 8512 9341
rect 8544 9309 8553 9341
rect 8504 9299 8553 9309
rect 8645 9341 8697 9350
rect 8645 9309 8655 9341
rect 8687 9309 8697 9341
rect 8645 9301 8697 9309
rect 8732 9341 8781 9351
rect 8732 9309 8741 9341
rect 8773 9309 8781 9341
rect 8732 9299 8781 9309
rect 8814 9224 9342 9452
rect 9374 9341 9423 9351
rect 9374 9309 9382 9341
rect 9414 9309 9423 9341
rect 9374 9299 9423 9309
rect 9515 9341 9567 9350
rect 9515 9309 9525 9341
rect 9557 9309 9567 9341
rect 9515 9301 9567 9309
rect 9602 9341 9651 9351
rect 9602 9309 9611 9341
rect 9643 9309 9651 9341
rect 9602 9299 9651 9309
rect 9693 9100 10221 9528
rect 10261 9341 10310 9351
rect 10261 9309 10269 9341
rect 10301 9309 10310 9341
rect 10261 9299 10310 9309
rect -2092 4932 5604 9044
rect 5674 4932 13370 9044
rect -2092 -1250 5604 2862
rect 5674 -1250 13370 2862
rect 968 -1515 1017 -1505
rect 968 -1547 977 -1515
rect 1009 -1547 1017 -1515
rect 968 -1557 1017 -1547
rect 1057 -1734 1585 -1306
rect 1627 -1515 1676 -1505
rect 1627 -1547 1635 -1515
rect 1667 -1547 1676 -1515
rect 1627 -1557 1676 -1547
rect 1711 -1515 1763 -1507
rect 1711 -1547 1721 -1515
rect 1753 -1547 1763 -1515
rect 1711 -1556 1763 -1547
rect 1855 -1515 1904 -1505
rect 1855 -1547 1864 -1515
rect 1896 -1547 1904 -1515
rect 1855 -1557 1904 -1547
rect 1936 -1658 2464 -1430
rect 2497 -1515 2546 -1505
rect 2497 -1547 2505 -1515
rect 2537 -1547 2546 -1515
rect 2497 -1557 2546 -1547
rect 2581 -1515 2633 -1507
rect 2581 -1547 2591 -1515
rect 2623 -1547 2633 -1515
rect 2581 -1556 2633 -1547
rect 2725 -1515 2774 -1505
rect 2725 -1547 2734 -1515
rect 2766 -1547 2774 -1515
rect 2725 -1557 2774 -1547
rect 2806 -1651 3084 -1423
rect 3114 -1515 3163 -1505
rect 3114 -1547 3122 -1515
rect 3154 -1547 3163 -1515
rect 3114 -1557 3163 -1547
rect 3244 -1515 3293 -1505
rect 3244 -1547 3253 -1515
rect 3285 -1547 3293 -1515
rect 3244 -1551 3293 -1547
rect 7985 -1515 8034 -1505
rect 7985 -1547 7993 -1515
rect 8025 -1547 8034 -1515
rect 7985 -1551 8034 -1547
rect 3244 -1557 3286 -1551
rect 7992 -1557 8034 -1551
rect 8115 -1515 8164 -1505
rect 8115 -1547 8124 -1515
rect 8156 -1547 8164 -1515
rect 8115 -1557 8164 -1547
rect 8194 -1651 8472 -1423
rect 8504 -1515 8553 -1505
rect 8504 -1547 8512 -1515
rect 8544 -1547 8553 -1515
rect 8504 -1557 8553 -1547
rect 8645 -1515 8697 -1507
rect 8645 -1547 8655 -1515
rect 8687 -1547 8697 -1515
rect 8645 -1556 8697 -1547
rect 8732 -1515 8781 -1505
rect 8732 -1547 8741 -1515
rect 8773 -1547 8781 -1515
rect 8732 -1557 8781 -1547
rect 8814 -1658 9342 -1430
rect 9374 -1515 9423 -1505
rect 9374 -1547 9382 -1515
rect 9414 -1547 9423 -1515
rect 9374 -1557 9423 -1547
rect 9515 -1515 9567 -1507
rect 9515 -1547 9525 -1515
rect 9557 -1547 9567 -1515
rect 9515 -1556 9567 -1547
rect 9602 -1515 9651 -1505
rect 9602 -1547 9611 -1515
rect 9643 -1547 9651 -1515
rect 9602 -1557 9651 -1547
rect 3602 -1715 3651 -1709
rect 3602 -1747 3614 -1715
rect 3646 -1747 3651 -1715
rect 3602 -1797 3651 -1747
rect 7627 -1715 7676 -1709
rect 7627 -1747 7632 -1715
rect 7664 -1747 7676 -1715
rect 9693 -1734 10221 -1306
rect 10261 -1515 10310 -1505
rect 10261 -1547 10269 -1515
rect 10301 -1547 10310 -1515
rect 10261 -1557 10310 -1547
rect 7627 -1797 7676 -1747
rect -2093 -4825 3019 -1797
rect 3075 -4825 5604 -1797
rect 5674 -4825 8203 -1797
rect 8259 -4825 13371 -1797
<< via3 >>
rect 977 9339 1009 9341
rect 977 9311 979 9339
rect 979 9311 1007 9339
rect 1007 9311 1009 9339
rect 977 9309 1009 9311
rect 3614 9539 3646 9541
rect 3614 9511 3615 9539
rect 3615 9511 3643 9539
rect 3643 9511 3646 9539
rect 3614 9509 3646 9511
rect 7632 9539 7664 9541
rect 7632 9511 7635 9539
rect 7635 9511 7663 9539
rect 7663 9511 7664 9539
rect 7632 9509 7664 9511
rect 1635 9339 1667 9341
rect 1635 9311 1637 9339
rect 1637 9311 1665 9339
rect 1665 9311 1667 9339
rect 1635 9309 1667 9311
rect 1721 9339 1753 9341
rect 1721 9311 1723 9339
rect 1723 9311 1751 9339
rect 1751 9311 1753 9339
rect 1721 9309 1753 9311
rect 1864 9339 1896 9341
rect 1864 9311 1866 9339
rect 1866 9311 1894 9339
rect 1894 9311 1896 9339
rect 1864 9309 1896 9311
rect 2505 9339 2537 9341
rect 2505 9311 2507 9339
rect 2507 9311 2535 9339
rect 2535 9311 2537 9339
rect 2505 9309 2537 9311
rect 2591 9339 2623 9341
rect 2591 9311 2593 9339
rect 2593 9311 2621 9339
rect 2621 9311 2623 9339
rect 2591 9309 2623 9311
rect 2734 9339 2766 9341
rect 2734 9311 2736 9339
rect 2736 9311 2764 9339
rect 2764 9311 2766 9339
rect 2734 9309 2766 9311
rect 3122 9339 3154 9341
rect 3122 9311 3124 9339
rect 3124 9311 3152 9339
rect 3152 9311 3154 9339
rect 3122 9309 3154 9311
rect 3253 9339 3285 9341
rect 3253 9311 3255 9339
rect 3255 9311 3283 9339
rect 3283 9311 3285 9339
rect 3253 9309 3285 9311
rect 7993 9339 8025 9341
rect 7993 9311 7995 9339
rect 7995 9311 8023 9339
rect 8023 9311 8025 9339
rect 7993 9309 8025 9311
rect 8124 9339 8156 9341
rect 8124 9311 8126 9339
rect 8126 9311 8154 9339
rect 8154 9311 8156 9339
rect 8124 9309 8156 9311
rect 8512 9339 8544 9341
rect 8512 9311 8514 9339
rect 8514 9311 8542 9339
rect 8542 9311 8544 9339
rect 8512 9309 8544 9311
rect 8655 9339 8687 9341
rect 8655 9311 8657 9339
rect 8657 9311 8685 9339
rect 8685 9311 8687 9339
rect 8655 9309 8687 9311
rect 8741 9339 8773 9341
rect 8741 9311 8743 9339
rect 8743 9311 8771 9339
rect 8771 9311 8773 9339
rect 8741 9309 8773 9311
rect 9382 9339 9414 9341
rect 9382 9311 9384 9339
rect 9384 9311 9412 9339
rect 9412 9311 9414 9339
rect 9382 9309 9414 9311
rect 9525 9339 9557 9341
rect 9525 9311 9527 9339
rect 9527 9311 9555 9339
rect 9555 9311 9557 9339
rect 9525 9309 9557 9311
rect 9611 9339 9643 9341
rect 9611 9311 9613 9339
rect 9613 9311 9641 9339
rect 9641 9311 9643 9339
rect 9611 9309 9643 9311
rect 10269 9339 10301 9341
rect 10269 9311 10271 9339
rect 10271 9311 10299 9339
rect 10299 9311 10301 9339
rect 10269 9309 10301 9311
rect 977 -1517 1009 -1515
rect 977 -1545 979 -1517
rect 979 -1545 1007 -1517
rect 1007 -1545 1009 -1517
rect 977 -1547 1009 -1545
rect 1635 -1517 1667 -1515
rect 1635 -1545 1637 -1517
rect 1637 -1545 1665 -1517
rect 1665 -1545 1667 -1517
rect 1635 -1547 1667 -1545
rect 1721 -1517 1753 -1515
rect 1721 -1545 1723 -1517
rect 1723 -1545 1751 -1517
rect 1751 -1545 1753 -1517
rect 1721 -1547 1753 -1545
rect 1864 -1517 1896 -1515
rect 1864 -1545 1866 -1517
rect 1866 -1545 1894 -1517
rect 1894 -1545 1896 -1517
rect 1864 -1547 1896 -1545
rect 2505 -1517 2537 -1515
rect 2505 -1545 2507 -1517
rect 2507 -1545 2535 -1517
rect 2535 -1545 2537 -1517
rect 2505 -1547 2537 -1545
rect 2591 -1517 2623 -1515
rect 2591 -1545 2593 -1517
rect 2593 -1545 2621 -1517
rect 2621 -1545 2623 -1517
rect 2591 -1547 2623 -1545
rect 2734 -1517 2766 -1515
rect 2734 -1545 2736 -1517
rect 2736 -1545 2764 -1517
rect 2764 -1545 2766 -1517
rect 2734 -1547 2766 -1545
rect 3122 -1517 3154 -1515
rect 3122 -1545 3124 -1517
rect 3124 -1545 3152 -1517
rect 3152 -1545 3154 -1517
rect 3122 -1547 3154 -1545
rect 3253 -1517 3285 -1515
rect 3253 -1545 3255 -1517
rect 3255 -1545 3283 -1517
rect 3283 -1545 3285 -1517
rect 3253 -1547 3285 -1545
rect 7993 -1517 8025 -1515
rect 7993 -1545 7995 -1517
rect 7995 -1545 8023 -1517
rect 8023 -1545 8025 -1517
rect 7993 -1547 8025 -1545
rect 8124 -1517 8156 -1515
rect 8124 -1545 8126 -1517
rect 8126 -1545 8154 -1517
rect 8154 -1545 8156 -1517
rect 8124 -1547 8156 -1545
rect 8512 -1517 8544 -1515
rect 8512 -1545 8514 -1517
rect 8514 -1545 8542 -1517
rect 8542 -1545 8544 -1517
rect 8512 -1547 8544 -1545
rect 8655 -1517 8687 -1515
rect 8655 -1545 8657 -1517
rect 8657 -1545 8685 -1517
rect 8685 -1545 8687 -1517
rect 8655 -1547 8687 -1545
rect 8741 -1517 8773 -1515
rect 8741 -1545 8743 -1517
rect 8743 -1545 8771 -1517
rect 8771 -1545 8773 -1517
rect 8741 -1547 8773 -1545
rect 9382 -1517 9414 -1515
rect 9382 -1545 9384 -1517
rect 9384 -1545 9412 -1517
rect 9412 -1545 9414 -1517
rect 9382 -1547 9414 -1545
rect 9525 -1517 9557 -1515
rect 9525 -1545 9527 -1517
rect 9527 -1545 9555 -1517
rect 9555 -1545 9557 -1517
rect 9525 -1547 9557 -1545
rect 9611 -1517 9643 -1515
rect 9611 -1545 9613 -1517
rect 9613 -1545 9641 -1517
rect 9641 -1545 9643 -1517
rect 9611 -1547 9643 -1545
rect 3614 -1717 3646 -1715
rect 3614 -1745 3615 -1717
rect 3615 -1745 3643 -1717
rect 3643 -1745 3646 -1717
rect 3614 -1747 3646 -1745
rect 7632 -1717 7664 -1715
rect 7632 -1745 7635 -1717
rect 7635 -1745 7663 -1717
rect 7663 -1745 7664 -1717
rect 7632 -1747 7664 -1745
rect 10269 -1517 10301 -1515
rect 10269 -1545 10271 -1517
rect 10271 -1545 10299 -1517
rect 10299 -1545 10301 -1517
rect 10269 -1547 10301 -1545
<< mimcap >>
rect -2079 9776 421 12605
rect -2079 9658 -1843 9776
rect -1725 9658 421 9776
rect -2079 9605 421 9658
rect 505 9759 3005 12605
rect 505 9641 725 9759
rect 843 9641 3005 9759
rect 505 9605 3005 9641
rect 3089 9776 5590 12605
rect 3089 9658 3327 9776
rect 3445 9658 5590 9776
rect 3089 9605 5590 9658
rect 5688 9776 8189 12605
rect 5688 9658 7833 9776
rect 7951 9658 8189 9776
rect 5688 9605 8189 9658
rect 8273 9759 10773 12605
rect 8273 9641 10435 9759
rect 10553 9641 10773 9759
rect 8273 9605 10773 9641
rect 10857 9776 13357 12605
rect 10857 9658 13003 9776
rect 13121 9658 13357 9776
rect 10857 9605 13357 9658
rect 1071 9344 1571 9514
rect 1071 9343 1519 9344
rect 1071 9308 1091 9343
rect 1127 9308 1519 9343
rect 1553 9308 1571 9344
rect 1071 9114 1571 9308
rect 1950 9343 2450 9438
rect 1950 9342 2405 9343
rect 1950 9306 1965 9342
rect 2000 9309 2405 9342
rect 2440 9309 2450 9343
rect 2000 9306 2450 9309
rect 1950 9238 2450 9306
rect 2820 9344 3070 9431
rect 2820 9341 3026 9344
rect 2820 9307 2830 9341
rect 2864 9309 3026 9341
rect 3060 9309 3070 9344
rect 2864 9307 3070 9309
rect 2820 9231 3070 9307
rect 8208 9344 8458 9431
rect 8208 9309 8218 9344
rect 8252 9341 8458 9344
rect 8252 9309 8414 9341
rect 8208 9307 8414 9309
rect 8448 9307 8458 9341
rect 8208 9231 8458 9307
rect 8828 9343 9328 9438
rect 8828 9309 8838 9343
rect 8873 9342 9328 9343
rect 8873 9309 9278 9342
rect 8828 9306 9278 9309
rect 9313 9306 9328 9342
rect 8828 9238 9328 9306
rect 9707 9344 10207 9514
rect 9707 9308 9725 9344
rect 9759 9343 10207 9344
rect 9759 9308 10151 9343
rect 10187 9308 10207 9343
rect 9707 9114 10207 9308
rect -2078 8983 922 9030
rect -2078 8865 -1858 8983
rect -1740 8865 922 8983
rect -2078 7372 922 8865
rect -2078 7254 767 7372
rect 885 7254 922 7372
rect -2078 7030 922 7254
rect 1006 7407 4006 9030
rect 1006 7365 3825 7407
rect 1006 7247 1040 7365
rect 1158 7289 3825 7365
rect 3943 7289 4006 7407
rect 1158 7247 4006 7289
rect 1006 7030 4006 7247
rect 4090 7424 5590 9030
rect 4090 7306 4133 7424
rect 4251 7306 5590 7424
rect 4090 7030 5590 7306
rect 5688 7424 7188 9030
rect 5688 7306 7027 7424
rect 7145 7306 7188 7424
rect 5688 7030 7188 7306
rect 7272 7407 10272 9030
rect 7272 7289 7335 7407
rect 7453 7365 10272 7407
rect 7453 7289 10120 7365
rect 7272 7247 10120 7289
rect 10238 7247 10272 7365
rect 7272 7030 10272 7247
rect 10356 8983 13356 9030
rect 10356 8865 13018 8983
rect 13136 8865 13356 8983
rect 10356 7372 13356 8865
rect 10356 7254 10393 7372
rect 10511 7254 13356 7372
rect 10356 7030 13356 7254
rect -2078 6725 922 6946
rect -2078 6607 757 6725
rect 875 6607 922 6725
rect -2078 4946 922 6607
rect 1006 6751 4006 6946
rect 1006 6728 3847 6751
rect 1006 6610 1059 6728
rect 1177 6633 3847 6728
rect 3965 6633 4006 6751
rect 1177 6610 4006 6633
rect 1006 4946 4006 6610
rect 4090 6718 5590 6946
rect 4090 6600 4143 6718
rect 4261 6600 5590 6718
rect 4090 4946 5590 6600
rect 5688 6718 7188 6946
rect 5688 6600 7017 6718
rect 7135 6600 7188 6718
rect 5688 4946 7188 6600
rect 7272 6751 10272 6946
rect 7272 6633 7313 6751
rect 7431 6728 10272 6751
rect 7431 6633 10101 6728
rect 7272 6610 10101 6633
rect 10219 6610 10272 6728
rect 7272 4946 10272 6610
rect 10356 6725 13356 6946
rect 10356 6607 10403 6725
rect 10521 6607 13356 6725
rect 10356 4946 13356 6607
rect -2078 1187 922 2848
rect -2078 1069 757 1187
rect 875 1069 922 1187
rect -2078 848 922 1069
rect 1006 1184 4006 2848
rect 1006 1066 1059 1184
rect 1177 1161 4006 1184
rect 1177 1066 3847 1161
rect 1006 1043 3847 1066
rect 3965 1043 4006 1161
rect 1006 848 4006 1043
rect 4090 1194 5590 2848
rect 4090 1076 4143 1194
rect 4261 1076 5590 1194
rect 4090 848 5590 1076
rect 5688 1194 7188 2848
rect 5688 1076 7017 1194
rect 7135 1076 7188 1194
rect 5688 848 7188 1076
rect 7272 1184 10272 2848
rect 7272 1161 10101 1184
rect 7272 1043 7313 1161
rect 7431 1066 10101 1161
rect 10219 1066 10272 1184
rect 7431 1043 10272 1066
rect 7272 848 10272 1043
rect 10356 1187 13356 2848
rect 10356 1069 10403 1187
rect 10521 1069 13356 1187
rect 10356 848 13356 1069
rect -2078 540 922 764
rect -2078 422 767 540
rect 885 422 922 540
rect -2078 -1071 922 422
rect -2078 -1189 -1858 -1071
rect -1740 -1189 922 -1071
rect -2078 -1236 922 -1189
rect 1006 547 4006 764
rect 1006 429 1040 547
rect 1158 505 4006 547
rect 1158 429 3825 505
rect 1006 387 3825 429
rect 3943 387 4006 505
rect 1006 -1236 4006 387
rect 4090 488 5590 764
rect 4090 370 4133 488
rect 4251 370 5590 488
rect 4090 -1236 5590 370
rect 5688 488 7188 764
rect 5688 370 7027 488
rect 7145 370 7188 488
rect 5688 -1236 7188 370
rect 7272 547 10272 764
rect 7272 505 10120 547
rect 7272 387 7335 505
rect 7453 429 10120 505
rect 10238 429 10272 547
rect 7453 387 10272 429
rect 7272 -1236 10272 387
rect 10356 540 13356 764
rect 10356 422 10393 540
rect 10511 422 13356 540
rect 10356 -1071 13356 422
rect 10356 -1189 13018 -1071
rect 13136 -1189 13356 -1071
rect 10356 -1236 13356 -1189
rect 1071 -1514 1571 -1320
rect 1071 -1549 1091 -1514
rect 1127 -1549 1519 -1514
rect 1071 -1550 1519 -1549
rect 1553 -1550 1571 -1514
rect 1071 -1720 1571 -1550
rect 1950 -1512 2450 -1444
rect 1950 -1548 1965 -1512
rect 2000 -1515 2450 -1512
rect 2000 -1548 2405 -1515
rect 1950 -1549 2405 -1548
rect 2440 -1549 2450 -1515
rect 1950 -1644 2450 -1549
rect 2820 -1513 3070 -1437
rect 2820 -1547 2830 -1513
rect 2864 -1515 3070 -1513
rect 2864 -1547 3026 -1515
rect 2820 -1550 3026 -1547
rect 3060 -1550 3070 -1515
rect 2820 -1637 3070 -1550
rect 8208 -1513 8458 -1437
rect 8208 -1515 8414 -1513
rect 8208 -1550 8218 -1515
rect 8252 -1547 8414 -1515
rect 8448 -1547 8458 -1513
rect 8252 -1550 8458 -1547
rect 8208 -1637 8458 -1550
rect 8828 -1512 9328 -1444
rect 8828 -1515 9278 -1512
rect 8828 -1549 8838 -1515
rect 8873 -1548 9278 -1515
rect 9313 -1548 9328 -1512
rect 8873 -1549 9328 -1548
rect 8828 -1644 9328 -1549
rect 9707 -1514 10207 -1320
rect 9707 -1550 9725 -1514
rect 9759 -1549 10151 -1514
rect 10187 -1549 10207 -1514
rect 9759 -1550 10207 -1549
rect 9707 -1720 10207 -1550
rect -2079 -1864 421 -1811
rect -2079 -1982 -1843 -1864
rect -1725 -1982 421 -1864
rect -2079 -4811 421 -1982
rect 505 -1847 3005 -1811
rect 505 -1965 725 -1847
rect 843 -1965 3005 -1847
rect 505 -4811 3005 -1965
rect 3089 -1864 5590 -1811
rect 3089 -1982 3327 -1864
rect 3445 -1982 5590 -1864
rect 3089 -4811 5590 -1982
rect 5688 -1864 8189 -1811
rect 5688 -1982 7833 -1864
rect 7951 -1982 8189 -1864
rect 5688 -4811 8189 -1982
rect 8273 -1847 10773 -1811
rect 8273 -1965 10435 -1847
rect 10553 -1965 10773 -1847
rect 8273 -4811 10773 -1965
rect 10857 -1864 13357 -1811
rect 10857 -1982 13003 -1864
rect 13121 -1982 13357 -1864
rect 10857 -4811 13357 -1982
<< mimcapcontact >>
rect -1843 9658 -1725 9776
rect 725 9641 843 9759
rect 3327 9658 3445 9776
rect 7833 9658 7951 9776
rect 10435 9641 10553 9759
rect 13003 9658 13121 9776
rect 1091 9308 1127 9343
rect 1519 9308 1553 9344
rect 1965 9306 2000 9342
rect 2405 9309 2440 9343
rect 2830 9307 2864 9341
rect 3026 9309 3060 9344
rect 8218 9309 8252 9344
rect 8414 9307 8448 9341
rect 8838 9309 8873 9343
rect 9278 9306 9313 9342
rect 9725 9308 9759 9344
rect 10151 9308 10187 9343
rect -1858 8865 -1740 8983
rect 767 7254 885 7372
rect 1040 7247 1158 7365
rect 3825 7289 3943 7407
rect 4133 7306 4251 7424
rect 7027 7306 7145 7424
rect 7335 7289 7453 7407
rect 10120 7247 10238 7365
rect 13018 8865 13136 8983
rect 10393 7254 10511 7372
rect 757 6607 875 6725
rect 1059 6610 1177 6728
rect 3847 6633 3965 6751
rect 4143 6600 4261 6718
rect 7017 6600 7135 6718
rect 7313 6633 7431 6751
rect 10101 6610 10219 6728
rect 10403 6607 10521 6725
rect 757 1069 875 1187
rect 1059 1066 1177 1184
rect 3847 1043 3965 1161
rect 4143 1076 4261 1194
rect 7017 1076 7135 1194
rect 7313 1043 7431 1161
rect 10101 1066 10219 1184
rect 10403 1069 10521 1187
rect 767 422 885 540
rect -1858 -1189 -1740 -1071
rect 1040 429 1158 547
rect 3825 387 3943 505
rect 4133 370 4251 488
rect 7027 370 7145 488
rect 7335 387 7453 505
rect 10120 429 10238 547
rect 10393 422 10511 540
rect 13018 -1189 13136 -1071
rect 1091 -1549 1127 -1514
rect 1519 -1550 1553 -1514
rect 1965 -1548 2000 -1512
rect 2405 -1549 2440 -1515
rect 2830 -1547 2864 -1513
rect 3026 -1550 3060 -1515
rect 8218 -1550 8252 -1515
rect 8414 -1547 8448 -1513
rect 8838 -1549 8873 -1515
rect 9278 -1548 9313 -1512
rect 9725 -1550 9759 -1514
rect 10151 -1549 10187 -1514
rect -1843 -1982 -1725 -1864
rect 725 -1965 843 -1847
rect 3327 -1982 3445 -1864
rect 7833 -1982 7951 -1864
rect 10435 -1965 10553 -1847
rect 13003 -1982 13121 -1864
<< metal4 >>
rect -2093 9776 3019 12619
rect -2093 9658 -1843 9776
rect -1725 9759 3019 9776
rect -1725 9658 725 9759
rect -2093 9641 725 9658
rect 843 9641 3019 9759
rect -2093 9591 3019 9641
rect 3075 9776 5604 12619
rect 3075 9658 3327 9776
rect 3445 9658 5604 9776
rect 3075 9591 5604 9658
rect 5674 9776 8203 12619
rect 5674 9658 7833 9776
rect 7951 9658 8203 9776
rect 5674 9591 8203 9658
rect 8259 9776 13371 12619
rect 8259 9759 13003 9776
rect 8259 9641 10435 9759
rect 10553 9658 13003 9759
rect 13121 9658 13371 9776
rect 10553 9641 13371 9658
rect 8259 9591 13371 9641
rect 1518 9344 1556 9345
rect 1090 9343 1128 9344
rect 1090 9342 1091 9343
rect 976 9341 1091 9342
rect 976 9309 977 9341
rect 1009 9309 1091 9341
rect 976 9308 1091 9309
rect 1127 9308 1128 9343
rect 976 9306 1128 9308
rect 1518 9308 1519 9344
rect 1553 9341 1668 9344
rect 2404 9343 2538 9344
rect 1553 9309 1635 9341
rect 1667 9309 1668 9341
rect 1553 9308 1668 9309
rect 1718 9341 1754 9342
rect 1718 9309 1721 9341
rect 1753 9309 1754 9341
rect 1518 9307 1556 9308
rect 1718 9044 1754 9309
rect 1863 9341 1965 9342
rect 1863 9309 1864 9341
rect 1896 9309 1965 9341
rect 1863 9306 1965 9309
rect 2000 9306 2010 9342
rect 2404 9309 2405 9343
rect 2440 9341 2538 9343
rect 2591 9342 2623 9591
rect 2440 9309 2505 9341
rect 2537 9309 2538 9341
rect 2404 9308 2538 9309
rect 2588 9341 2624 9342
rect 2588 9309 2591 9341
rect 2623 9309 2624 9341
rect 2588 9307 2624 9309
rect 2733 9341 2876 9342
rect 2733 9309 2734 9341
rect 2766 9309 2830 9341
rect 2733 9307 2830 9309
rect 2864 9307 2876 9341
rect 3024 9309 3026 9344
rect 3060 9341 3155 9344
rect 3060 9309 3122 9341
rect 3154 9309 3155 9341
rect 3024 9308 3155 9309
rect 3248 9341 3298 9591
rect 3248 9309 3253 9341
rect 3285 9309 3298 9341
rect 2733 9306 2876 9307
rect 3248 9303 3298 9309
rect 7980 9341 8030 9591
rect 7980 9309 7993 9341
rect 8025 9309 8030 9341
rect 7980 9303 8030 9309
rect 8123 9341 8218 9344
rect 8123 9309 8124 9341
rect 8156 9309 8218 9341
rect 8252 9309 8254 9344
rect 8655 9342 8687 9591
rect 9722 9344 9760 9345
rect 8740 9343 8874 9344
rect 8123 9308 8254 9309
rect 8402 9341 8545 9342
rect 8402 9307 8414 9341
rect 8448 9309 8512 9341
rect 8544 9309 8545 9341
rect 8448 9307 8545 9309
rect 8654 9341 8690 9342
rect 8654 9309 8655 9341
rect 8687 9309 8690 9341
rect 8654 9307 8690 9309
rect 8740 9341 8838 9343
rect 8740 9309 8741 9341
rect 8773 9309 8838 9341
rect 8873 9309 8874 9343
rect 8740 9308 8874 9309
rect 8402 9306 8545 9307
rect 9268 9306 9278 9342
rect 9313 9341 9415 9342
rect 9313 9309 9382 9341
rect 9414 9309 9415 9341
rect 9313 9306 9415 9309
rect 9524 9341 9560 9342
rect 9524 9309 9525 9341
rect 9557 9309 9560 9341
rect 9524 9044 9560 9309
rect 9610 9341 9725 9344
rect 9610 9309 9611 9341
rect 9643 9309 9725 9341
rect 9610 9308 9725 9309
rect 9759 9308 9760 9344
rect 9722 9307 9760 9308
rect 10150 9343 10188 9344
rect 10150 9308 10151 9343
rect 10187 9342 10188 9343
rect 10187 9341 10302 9342
rect 10187 9309 10269 9341
rect 10301 9309 10302 9341
rect 10187 9308 10302 9309
rect 10150 9306 10302 9308
rect -2092 8983 5604 9044
rect -2092 8865 -1858 8983
rect -1740 8865 5604 8983
rect -2092 7424 5604 8865
rect -2092 7407 4133 7424
rect -2092 7372 3825 7407
rect -2092 7254 767 7372
rect 885 7365 3825 7372
rect 885 7254 1040 7365
rect -2092 7247 1040 7254
rect 1158 7289 3825 7365
rect 3943 7306 4133 7407
rect 4251 7306 5604 7424
rect 3943 7289 5604 7306
rect 1158 7247 5604 7289
rect -2092 6751 5604 7247
rect -2092 6728 3847 6751
rect -2092 6725 1059 6728
rect -2092 6607 757 6725
rect 875 6610 1059 6725
rect 1177 6633 3847 6728
rect 3965 6718 5604 6751
rect 3965 6633 4143 6718
rect 1177 6610 4143 6633
rect 875 6607 4143 6610
rect -2092 6600 4143 6607
rect 4261 6600 5604 6718
rect -2092 4932 5604 6600
rect 5674 8983 13370 9044
rect 5674 8865 13018 8983
rect 13136 8865 13370 8983
rect 5674 7424 13370 8865
rect 5674 7306 7027 7424
rect 7145 7407 13370 7424
rect 7145 7306 7335 7407
rect 5674 7289 7335 7306
rect 7453 7372 13370 7407
rect 7453 7365 10393 7372
rect 7453 7289 10120 7365
rect 5674 7247 10120 7289
rect 10238 7254 10393 7365
rect 10511 7254 13370 7372
rect 10238 7247 13370 7254
rect 5674 6751 13370 7247
rect 5674 6718 7313 6751
rect 5674 6600 7017 6718
rect 7135 6633 7313 6718
rect 7431 6728 13370 6751
rect 7431 6633 10101 6728
rect 7135 6610 10101 6633
rect 10219 6725 13370 6728
rect 10219 6610 10403 6725
rect 7135 6607 10403 6610
rect 10521 6607 13370 6725
rect 7135 6600 13370 6607
rect 5674 4932 13370 6600
rect -2092 1194 5604 2862
rect -2092 1187 4143 1194
rect -2092 1069 757 1187
rect 875 1184 4143 1187
rect 875 1069 1059 1184
rect -2092 1066 1059 1069
rect 1177 1161 4143 1184
rect 1177 1066 3847 1161
rect -2092 1043 3847 1066
rect 3965 1076 4143 1161
rect 4261 1076 5604 1194
rect 3965 1043 5604 1076
rect -2092 547 5604 1043
rect -2092 540 1040 547
rect -2092 422 767 540
rect 885 429 1040 540
rect 1158 505 5604 547
rect 1158 429 3825 505
rect 885 422 3825 429
rect -2092 387 3825 422
rect 3943 488 5604 505
rect 3943 387 4133 488
rect -2092 370 4133 387
rect 4251 370 5604 488
rect -2092 -1071 5604 370
rect -2092 -1189 -1858 -1071
rect -1740 -1189 5604 -1071
rect -2092 -1250 5604 -1189
rect 5674 1194 13370 2862
rect 5674 1076 7017 1194
rect 7135 1187 13370 1194
rect 7135 1184 10403 1187
rect 7135 1161 10101 1184
rect 7135 1076 7313 1161
rect 5674 1043 7313 1076
rect 7431 1066 10101 1161
rect 10219 1069 10403 1184
rect 10521 1069 13370 1187
rect 10219 1066 13370 1069
rect 7431 1043 13370 1066
rect 5674 547 13370 1043
rect 5674 505 10120 547
rect 5674 488 7335 505
rect 5674 370 7027 488
rect 7145 387 7335 488
rect 7453 429 10120 505
rect 10238 540 13370 547
rect 10238 429 10393 540
rect 7453 422 10393 429
rect 10511 422 13370 540
rect 7453 387 13370 422
rect 7145 370 13370 387
rect 5674 -1071 13370 370
rect 5674 -1189 13018 -1071
rect 13136 -1189 13370 -1071
rect 5674 -1250 13370 -1189
rect 976 -1514 1128 -1512
rect 976 -1515 1091 -1514
rect 976 -1547 977 -1515
rect 1009 -1547 1091 -1515
rect 976 -1548 1091 -1547
rect 1090 -1549 1091 -1548
rect 1127 -1549 1128 -1514
rect 1090 -1550 1128 -1549
rect 1518 -1514 1556 -1513
rect 1518 -1550 1519 -1514
rect 1553 -1515 1668 -1514
rect 1553 -1547 1635 -1515
rect 1667 -1547 1668 -1515
rect 1553 -1550 1668 -1547
rect 1718 -1515 1754 -1250
rect 1718 -1547 1721 -1515
rect 1753 -1547 1754 -1515
rect 1718 -1548 1754 -1547
rect 1863 -1515 1965 -1512
rect 1863 -1547 1864 -1515
rect 1896 -1547 1965 -1515
rect 1863 -1548 1965 -1547
rect 2000 -1548 2010 -1512
rect 2733 -1513 2876 -1512
rect 2404 -1515 2538 -1514
rect 2404 -1549 2405 -1515
rect 2440 -1547 2505 -1515
rect 2537 -1547 2538 -1515
rect 2440 -1549 2538 -1547
rect 2588 -1515 2624 -1513
rect 2588 -1547 2591 -1515
rect 2623 -1547 2624 -1515
rect 2588 -1548 2624 -1547
rect 2733 -1515 2830 -1513
rect 2733 -1547 2734 -1515
rect 2766 -1547 2830 -1515
rect 2864 -1547 2876 -1513
rect 2733 -1548 2876 -1547
rect 3024 -1515 3155 -1514
rect 2404 -1550 2538 -1549
rect 1518 -1551 1556 -1550
rect 2591 -1797 2623 -1548
rect 3024 -1550 3026 -1515
rect 3060 -1547 3122 -1515
rect 3154 -1547 3155 -1515
rect 3060 -1550 3155 -1547
rect 3248 -1515 3298 -1509
rect 3248 -1547 3253 -1515
rect 3285 -1547 3298 -1515
rect 3248 -1797 3298 -1547
rect 7980 -1515 8030 -1509
rect 8402 -1513 8545 -1512
rect 7980 -1547 7993 -1515
rect 8025 -1547 8030 -1515
rect 7980 -1797 8030 -1547
rect 8123 -1515 8254 -1514
rect 8123 -1547 8124 -1515
rect 8156 -1547 8218 -1515
rect 8123 -1550 8218 -1547
rect 8252 -1550 8254 -1515
rect 8402 -1547 8414 -1513
rect 8448 -1515 8545 -1513
rect 8448 -1547 8512 -1515
rect 8544 -1547 8545 -1515
rect 8402 -1548 8545 -1547
rect 8654 -1515 8690 -1513
rect 8654 -1547 8655 -1515
rect 8687 -1547 8690 -1515
rect 8654 -1548 8690 -1547
rect 8740 -1515 8874 -1514
rect 8740 -1547 8741 -1515
rect 8773 -1547 8838 -1515
rect 8655 -1797 8687 -1548
rect 8740 -1549 8838 -1547
rect 8873 -1549 8874 -1515
rect 9268 -1548 9278 -1512
rect 9313 -1515 9415 -1512
rect 9313 -1547 9382 -1515
rect 9414 -1547 9415 -1515
rect 9313 -1548 9415 -1547
rect 9524 -1515 9560 -1250
rect 9722 -1514 9760 -1513
rect 9524 -1547 9525 -1515
rect 9557 -1547 9560 -1515
rect 9524 -1548 9560 -1547
rect 9610 -1515 9725 -1514
rect 9610 -1547 9611 -1515
rect 9643 -1547 9725 -1515
rect 8740 -1550 8874 -1549
rect 9610 -1550 9725 -1547
rect 9759 -1550 9760 -1514
rect 10150 -1514 10302 -1512
rect 10150 -1549 10151 -1514
rect 10187 -1515 10302 -1514
rect 10187 -1547 10269 -1515
rect 10301 -1547 10302 -1515
rect 10187 -1548 10302 -1547
rect 10187 -1549 10188 -1548
rect 10150 -1550 10188 -1549
rect 9722 -1551 9760 -1550
rect -2093 -1847 3019 -1797
rect -2093 -1864 725 -1847
rect -2093 -1982 -1843 -1864
rect -1725 -1965 725 -1864
rect 843 -1965 3019 -1847
rect -1725 -1982 3019 -1965
rect -2093 -4825 3019 -1982
rect 3075 -1864 5604 -1797
rect 3075 -1982 3327 -1864
rect 3445 -1982 5604 -1864
rect 3075 -4825 5604 -1982
rect 5674 -1864 8203 -1797
rect 5674 -1982 7833 -1864
rect 7951 -1982 8203 -1864
rect 5674 -4825 8203 -1982
rect 8259 -1847 13371 -1797
rect 8259 -1965 10435 -1847
rect 10553 -1864 13371 -1847
rect 10553 -1965 13003 -1864
rect 8259 -1982 13003 -1965
rect 13121 -1982 13371 -1864
rect 8259 -4825 13371 -1982
<< via4 >>
rect 3570 9541 3689 9551
rect 3570 9509 3614 9541
rect 3614 9509 3646 9541
rect 3646 9509 3689 9541
rect 3570 9433 3689 9509
rect 7589 9541 7708 9551
rect 7589 9509 7632 9541
rect 7632 9509 7664 9541
rect 7664 9509 7708 9541
rect 7589 9433 7708 9509
rect 3570 -1715 3689 -1639
rect 3570 -1747 3614 -1715
rect 3614 -1747 3646 -1715
rect 3646 -1747 3689 -1715
rect 3570 -1757 3689 -1747
rect 7589 -1715 7708 -1639
rect 7589 -1747 7632 -1715
rect 7632 -1747 7664 -1715
rect 7664 -1747 7708 -1715
rect 7589 -1757 7708 -1747
<< mimcap2 >>
rect -2079 9777 421 12605
rect -2079 9659 241 9777
rect 359 9659 421 9777
rect -2079 9605 421 9659
rect 505 9777 3005 12605
rect 505 9659 554 9777
rect 672 9659 3005 9777
rect 505 9605 3005 9659
rect 3089 9770 5590 12605
rect 3089 9652 3571 9770
rect 3689 9652 5590 9770
rect 3089 9605 5590 9652
rect 5688 9770 8189 12605
rect 5688 9652 7589 9770
rect 7707 9652 8189 9770
rect 5688 9605 8189 9652
rect 8273 9777 10773 12605
rect 8273 9659 10606 9777
rect 10724 9659 10773 9777
rect 8273 9605 10773 9659
rect 10857 9777 13357 12605
rect 10857 9659 10919 9777
rect 11037 9659 13357 9777
rect 10857 9605 13357 9659
rect -2078 7186 922 9030
rect -2078 7068 762 7186
rect 880 7068 922 7186
rect -2078 7030 922 7068
rect 1006 7204 4006 9030
rect 1006 7183 3830 7204
rect 1006 7065 1044 7183
rect 1162 7086 3830 7183
rect 3948 7086 4006 7204
rect 1162 7065 4006 7086
rect 1006 7030 4006 7065
rect 4090 7206 5590 9030
rect 4090 7088 4122 7206
rect 4240 7088 5590 7206
rect 4090 7030 5590 7088
rect 5688 7206 7188 9030
rect 5688 7088 7038 7206
rect 7156 7088 7188 7206
rect 5688 7030 7188 7088
rect 7272 7204 10272 9030
rect 7272 7086 7330 7204
rect 7448 7183 10272 7204
rect 7448 7086 10116 7183
rect 7272 7065 10116 7086
rect 10234 7065 10272 7183
rect 7272 7030 10272 7065
rect 10356 7186 13356 9030
rect 10356 7068 10398 7186
rect 10516 7068 13356 7186
rect 10356 7030 13356 7068
rect -2078 6909 922 6946
rect -2078 6791 763 6909
rect 881 6791 922 6909
rect -2078 4946 922 6791
rect 1006 6925 4006 6946
rect 1006 6907 3833 6925
rect 1006 6789 1047 6907
rect 1165 6807 3833 6907
rect 3951 6807 4006 6925
rect 1165 6789 4006 6807
rect 1006 4946 4006 6789
rect 4090 6920 5590 6946
rect 4090 6802 4124 6920
rect 4242 6802 5590 6920
rect 4090 4946 5590 6802
rect 5688 6920 7188 6946
rect 5688 6802 7036 6920
rect 7154 6802 7188 6920
rect 5688 4946 7188 6802
rect 7272 6925 10272 6946
rect 7272 6807 7327 6925
rect 7445 6907 10272 6925
rect 7445 6807 10113 6907
rect 7272 6789 10113 6807
rect 10231 6789 10272 6907
rect 7272 4946 10272 6789
rect 10356 6909 13356 6946
rect 10356 6791 10397 6909
rect 10515 6791 13356 6909
rect 10356 4946 13356 6791
rect -2078 1003 922 2848
rect -2078 885 763 1003
rect 881 885 922 1003
rect -2078 848 922 885
rect 1006 1005 4006 2848
rect 1006 887 1047 1005
rect 1165 987 4006 1005
rect 1165 887 3833 987
rect 1006 869 3833 887
rect 3951 869 4006 987
rect 1006 848 4006 869
rect 4090 992 5590 2848
rect 4090 874 4124 992
rect 4242 874 5590 992
rect 4090 848 5590 874
rect 5688 992 7188 2848
rect 5688 874 7036 992
rect 7154 874 7188 992
rect 5688 848 7188 874
rect 7272 1005 10272 2848
rect 7272 987 10113 1005
rect 7272 869 7327 987
rect 7445 887 10113 987
rect 10231 887 10272 1005
rect 7445 869 10272 887
rect 7272 848 10272 869
rect 10356 1003 13356 2848
rect 10356 885 10397 1003
rect 10515 885 13356 1003
rect 10356 848 13356 885
rect -2078 726 922 764
rect -2078 608 762 726
rect 880 608 922 726
rect -2078 -1236 922 608
rect 1006 729 4006 764
rect 1006 611 1044 729
rect 1162 708 4006 729
rect 1162 611 3830 708
rect 1006 590 3830 611
rect 3948 590 4006 708
rect 1006 -1236 4006 590
rect 4090 706 5590 764
rect 4090 588 4122 706
rect 4240 588 5590 706
rect 4090 -1236 5590 588
rect 5688 706 7188 764
rect 5688 588 7038 706
rect 7156 588 7188 706
rect 5688 -1236 7188 588
rect 7272 729 10272 764
rect 7272 708 10116 729
rect 7272 590 7330 708
rect 7448 611 10116 708
rect 10234 611 10272 729
rect 7448 590 10272 611
rect 7272 -1236 10272 590
rect 10356 726 13356 764
rect 10356 608 10398 726
rect 10516 608 13356 726
rect 10356 -1236 13356 608
rect -2079 -1865 421 -1811
rect -2079 -1983 241 -1865
rect 359 -1983 421 -1865
rect -2079 -4811 421 -1983
rect 505 -1865 3005 -1811
rect 505 -1983 554 -1865
rect 672 -1983 3005 -1865
rect 505 -4811 3005 -1983
rect 3089 -1858 5590 -1811
rect 3089 -1976 3571 -1858
rect 3689 -1976 5590 -1858
rect 3089 -4811 5590 -1976
rect 5688 -1858 8189 -1811
rect 5688 -1976 7589 -1858
rect 7707 -1976 8189 -1858
rect 5688 -4811 8189 -1976
rect 8273 -1865 10773 -1811
rect 8273 -1983 10606 -1865
rect 10724 -1983 10773 -1865
rect 8273 -4811 10773 -1983
rect 10857 -1865 13357 -1811
rect 10857 -1983 10919 -1865
rect 11037 -1983 13357 -1865
rect 10857 -4811 13357 -1983
<< mimcap2contact >>
rect 241 9659 359 9777
rect 554 9659 672 9777
rect 3571 9652 3689 9770
rect 7589 9652 7707 9770
rect 10606 9659 10724 9777
rect 10919 9659 11037 9777
rect 762 7068 880 7186
rect 1044 7065 1162 7183
rect 3830 7086 3948 7204
rect 4122 7088 4240 7206
rect 7038 7088 7156 7206
rect 7330 7086 7448 7204
rect 10116 7065 10234 7183
rect 10398 7068 10516 7186
rect 763 6791 881 6909
rect 1047 6789 1165 6907
rect 3833 6807 3951 6925
rect 4124 6802 4242 6920
rect 7036 6802 7154 6920
rect 7327 6807 7445 6925
rect 10113 6789 10231 6907
rect 10397 6791 10515 6909
rect 763 885 881 1003
rect 1047 887 1165 1005
rect 3833 869 3951 987
rect 4124 874 4242 992
rect 7036 874 7154 992
rect 7327 869 7445 987
rect 10113 887 10231 1005
rect 10397 885 10515 1003
rect 762 608 880 726
rect 1044 611 1162 729
rect 3830 590 3948 708
rect 4122 588 4240 706
rect 7038 588 7156 706
rect 7330 590 7448 708
rect 10116 611 10234 729
rect 10398 608 10516 726
rect 241 -1983 359 -1865
rect 554 -1983 672 -1865
rect 3571 -1976 3689 -1858
rect 7589 -1976 7707 -1858
rect 10606 -1983 10724 -1865
rect 10919 -1983 11037 -1865
<< metal5 >>
rect 218 9777 700 9794
rect 218 9659 241 9777
rect 359 9659 554 9777
rect 672 9659 700 9777
rect 218 9633 700 9659
rect 3555 9770 3716 9788
rect 3555 9652 3571 9770
rect 3689 9652 3716 9770
rect 3555 9630 3716 9652
rect 7562 9770 7723 9788
rect 7562 9652 7589 9770
rect 7707 9652 7723 9770
rect 7562 9630 7723 9652
rect 10578 9777 11060 9794
rect 10578 9659 10606 9777
rect 10724 9659 10919 9777
rect 11037 9659 11060 9777
rect 10578 9633 11060 9659
rect 3555 9551 3719 9630
rect 3555 9433 3570 9551
rect 3689 9433 3719 9551
rect 3555 9420 3719 9433
rect 7559 9551 7723 9630
rect 7559 9433 7589 9551
rect 7708 9433 7723 9551
rect 7559 9420 7723 9433
rect 3809 7206 4266 7225
rect 3809 7204 4122 7206
rect 730 7186 1188 7202
rect 730 7068 762 7186
rect 880 7183 1188 7186
rect 880 7068 1044 7183
rect 730 7065 1044 7068
rect 1162 7065 1188 7183
rect 730 6909 1188 7065
rect 730 6791 763 6909
rect 881 6907 1188 6909
rect 881 6791 1047 6907
rect 730 6789 1047 6791
rect 1165 6789 1188 6907
rect 730 6765 1188 6789
rect 3809 7086 3830 7204
rect 3948 7088 4122 7204
rect 4240 7088 4266 7206
rect 3948 7086 4266 7088
rect 3809 6925 4266 7086
rect 3809 6807 3833 6925
rect 3951 6920 4266 6925
rect 3951 6807 4124 6920
rect 3809 6802 4124 6807
rect 4242 6802 4266 6920
rect 3809 6781 4266 6802
rect 7012 7206 7469 7225
rect 7012 7088 7038 7206
rect 7156 7204 7469 7206
rect 7156 7088 7330 7204
rect 7012 7086 7330 7088
rect 7448 7086 7469 7204
rect 7012 6925 7469 7086
rect 7012 6920 7327 6925
rect 7012 6802 7036 6920
rect 7154 6807 7327 6920
rect 7445 6807 7469 6925
rect 7154 6802 7469 6807
rect 7012 6781 7469 6802
rect 10090 7186 10548 7202
rect 10090 7183 10398 7186
rect 10090 7065 10116 7183
rect 10234 7068 10398 7183
rect 10516 7068 10548 7186
rect 10234 7065 10548 7068
rect 10090 6909 10548 7065
rect 10090 6907 10397 6909
rect 10090 6789 10113 6907
rect 10231 6791 10397 6907
rect 10515 6791 10548 6909
rect 10231 6789 10548 6791
rect 10090 6765 10548 6789
rect 730 1005 1188 1029
rect 730 1003 1047 1005
rect 730 885 763 1003
rect 881 887 1047 1003
rect 1165 887 1188 1005
rect 881 885 1188 887
rect 730 729 1188 885
rect 730 726 1044 729
rect 730 608 762 726
rect 880 611 1044 726
rect 1162 611 1188 729
rect 880 608 1188 611
rect 730 592 1188 608
rect 3809 992 4266 1013
rect 3809 987 4124 992
rect 3809 869 3833 987
rect 3951 874 4124 987
rect 4242 874 4266 992
rect 3951 869 4266 874
rect 3809 708 4266 869
rect 3809 590 3830 708
rect 3948 706 4266 708
rect 3948 590 4122 706
rect 3809 588 4122 590
rect 4240 588 4266 706
rect 3809 569 4266 588
rect 7012 992 7469 1013
rect 7012 874 7036 992
rect 7154 987 7469 992
rect 7154 874 7327 987
rect 7012 869 7327 874
rect 7445 869 7469 987
rect 7012 708 7469 869
rect 7012 706 7330 708
rect 7012 588 7038 706
rect 7156 590 7330 706
rect 7448 590 7469 708
rect 10090 1005 10548 1029
rect 10090 887 10113 1005
rect 10231 1003 10548 1005
rect 10231 887 10397 1003
rect 10090 885 10397 887
rect 10515 885 10548 1003
rect 10090 729 10548 885
rect 10090 611 10116 729
rect 10234 726 10548 729
rect 10234 611 10398 726
rect 10090 608 10398 611
rect 10516 608 10548 726
rect 10090 592 10548 608
rect 7156 588 7469 590
rect 7012 569 7469 588
rect 3555 -1639 3719 -1626
rect 3555 -1757 3570 -1639
rect 3689 -1757 3719 -1639
rect 3555 -1836 3719 -1757
rect 7559 -1639 7723 -1626
rect 7559 -1757 7589 -1639
rect 7708 -1757 7723 -1639
rect 7559 -1836 7723 -1757
rect 218 -1865 700 -1839
rect 218 -1983 241 -1865
rect 359 -1983 554 -1865
rect 672 -1983 700 -1865
rect 218 -2000 700 -1983
rect 3555 -1858 3716 -1836
rect 3555 -1976 3571 -1858
rect 3689 -1976 3716 -1858
rect 3555 -1994 3716 -1976
rect 7562 -1858 7723 -1836
rect 7562 -1976 7589 -1858
rect 7707 -1976 7723 -1858
rect 7562 -1994 7723 -1976
rect 10578 -1865 11060 -1839
rect 10578 -1983 10606 -1865
rect 10724 -1983 10919 -1865
rect 11037 -1983 11060 -1865
rect 10578 -2000 11060 -1983
<< labels >>
flabel metal4 1885 -36 2909 887 0 FreeSans 800 0 0 0 C1
flabel mimcap 1256 -1622 1447 -1471 0 FreeSans 800 0 0 0 Cs1
rlabel metal4 1033 -1512 1033 -1512 1 cs1
flabel mimcap 2115 -1620 2306 -1469 0 FreeSans 800 0 0 0 Cs2
flabel metal4 -82 -3740 942 -2817 0 FreeSans 800 0 0 0 C2
flabel mimcap2 3912 -3489 4936 -2566 0 FreeSans 800 0 0 0 C3
flabel mimcap 2863 -1593 3054 -1442 0 FreeSans 800 0 0 0 Cs3
rlabel metal4 1754 -1270 1754 -1270 3 c1
rlabel metal4 1922 -1548 1922 -1548 5 cs2
rlabel metal4 2623 -1752 2623 -1752 3 c2
rlabel metal4 3098 -1550 3098 -1550 5 cs3
rlabel metal4 3298 -1734 3298 -1734 3 c3
flabel metal4 8369 -36 9393 887 0 FreeSans 800 180 0 0 C1
flabel mimcap 9831 -1622 10022 -1471 0 FreeSans 800 180 0 0 Cs1
rlabel metal4 10245 -1512 10245 -1512 1 cs1
flabel mimcap 8972 -1620 9163 -1469 0 FreeSans 800 180 0 0 Cs2
flabel metal4 10336 -3740 11360 -2817 0 FreeSans 800 180 0 0 C2
flabel mimcap2 6342 -3489 7366 -2566 0 FreeSans 800 180 0 0 C3
flabel mimcap 8224 -1593 8415 -1442 0 FreeSans 800 180 0 0 Cs3
rlabel metal4 9524 -1270 9524 -1270 7 c1
rlabel metal4 9356 -1548 9356 -1548 5 cs2
rlabel metal4 8655 -1752 8655 -1752 7 c2
rlabel metal4 8180 -1550 8180 -1550 5 cs3
rlabel metal4 7980 -1734 7980 -1734 7 c3
flabel metal4 1885 6907 2909 7830 0 FreeSans 800 0 0 0 C1
flabel mimcap 1256 9265 1447 9416 0 FreeSans 800 0 0 0 Cs1
rlabel metal4 1033 9306 1033 9306 5 cs1
flabel mimcap 2115 9263 2306 9414 0 FreeSans 800 0 0 0 Cs2
flabel metal4 -82 10611 942 11534 0 FreeSans 800 0 0 0 C2
flabel mimcap2 3912 10360 4936 11283 0 FreeSans 800 0 0 0 C3
flabel mimcap 2863 9236 3054 9387 0 FreeSans 800 0 0 0 Cs3
rlabel metal4 1754 9064 1754 9064 3 c1
rlabel metal4 1922 9342 1922 9342 1 cs2
rlabel metal4 2623 9546 2623 9546 3 c2
rlabel metal4 3098 9344 3098 9344 1 cs3
rlabel metal4 3298 9528 3298 9528 3 c3
flabel metal4 8369 6907 9393 7830 0 FreeSans 800 180 0 0 C1
flabel mimcap 9831 9265 10022 9416 0 FreeSans 800 180 0 0 Cs1
rlabel metal4 10245 9306 10245 9306 5 cs1
flabel mimcap 8972 9263 9163 9414 0 FreeSans 800 180 0 0 Cs2
flabel metal4 10336 10611 11360 11534 0 FreeSans 800 180 0 0 C2
flabel mimcap2 6342 10360 7366 11283 0 FreeSans 800 180 0 0 C3
flabel mimcap 8224 9236 8415 9387 0 FreeSans 800 180 0 0 Cs3
rlabel metal4 9524 9064 9524 9064 7 c1
rlabel metal4 9356 9342 9356 9342 1 cs2
rlabel metal4 8655 9546 8655 9546 7 c2
rlabel metal4 8180 9344 8180 9344 1 cs3
rlabel metal4 7980 9528 7980 9528 7 c3
<< end >>
