** sch_path: /local_disk/fossi_cochlea/xschem/Switched_Caps/mim_cap_stacked_6pF.sch
.subckt mim_cap_stacked_6pF sig vss
*.PININFO sig:B vss:B
XC1 sig vss sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=16 m=16
XC2 vss sig sky130_fd_pr__cap_mim_m3_2 W=10 L=10 VM=16 m=16
.ends
.end
