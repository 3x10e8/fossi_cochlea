magic
tech sky130A
magscale 1 2
timestamp 1647885722
<< viali >>
rect 4077 5321 4111 5355
rect 4905 5321 4939 5355
rect 8493 5321 8527 5355
rect 9413 5321 9447 5355
rect 16865 5321 16899 5355
rect 2237 5253 2271 5287
rect 15117 5253 15151 5287
rect 17509 5253 17543 5287
rect 3065 5185 3099 5219
rect 4261 5185 4295 5219
rect 5089 5185 5123 5219
rect 8677 5185 8711 5219
rect 9229 5185 9263 5219
rect 10149 5185 10183 5219
rect 10793 5185 10827 5219
rect 15393 5185 15427 5219
rect 15945 5185 15979 5219
rect 16681 5185 16715 5219
rect 17417 5185 17451 5219
rect 2513 5117 2547 5151
rect 5733 5117 5767 5151
rect 6009 5117 6043 5151
rect 11069 5117 11103 5151
rect 765 4981 799 5015
rect 3249 4981 3283 5015
rect 7481 4981 7515 5015
rect 10149 4981 10183 5015
rect 12541 4981 12575 5015
rect 13645 4981 13679 5015
rect 16129 4981 16163 5015
rect 1409 4777 1443 4811
rect 3249 4777 3283 4811
rect 6469 4777 6503 4811
rect 7389 4777 7423 4811
rect 8217 4777 8251 4811
rect 9689 4777 9723 4811
rect 11989 4777 12023 4811
rect 12725 4777 12759 4811
rect 16681 4777 16715 4811
rect 17417 4777 17451 4811
rect 9229 4709 9263 4743
rect 3985 4641 4019 4675
rect 4261 4641 4295 4675
rect 11161 4641 11195 4675
rect 14565 4641 14599 4675
rect 16037 4641 16071 4675
rect 1225 4573 1259 4607
rect 2237 4573 2271 4607
rect 3065 4573 3099 4607
rect 6653 4573 6687 4607
rect 7573 4573 7607 4607
rect 8217 4573 8251 4607
rect 8401 4573 8435 4607
rect 9045 4573 9079 4607
rect 9229 4573 9263 4607
rect 11437 4573 11471 4607
rect 12173 4573 12207 4607
rect 12817 4573 12851 4607
rect 13645 4573 13679 4607
rect 14289 4573 14323 4607
rect 16497 4573 16531 4607
rect 17233 4573 17267 4607
rect 1961 4505 1995 4539
rect 13369 4505 13403 4539
rect 5733 4437 5767 4471
rect 2973 4233 3007 4267
rect 14657 4233 14691 4267
rect 1501 4165 1535 4199
rect 3801 4165 3835 4199
rect 13185 4165 13219 4199
rect 4997 4097 5031 4131
rect 6469 4097 6503 4131
rect 7481 4097 7515 4131
rect 10241 4097 10275 4131
rect 11069 4097 11103 4131
rect 11621 4097 11655 4131
rect 12449 4097 12483 4131
rect 12909 4097 12943 4131
rect 15209 4097 15243 4131
rect 15301 4097 15335 4131
rect 15945 4097 15979 4131
rect 16037 4097 16071 4131
rect 16129 4097 16163 4131
rect 16589 4097 16623 4131
rect 16773 4097 16807 4131
rect 17325 4097 17359 4131
rect 1225 4029 1259 4063
rect 4721 4029 4755 4063
rect 7757 4029 7791 4063
rect 3617 3961 3651 3995
rect 6285 3961 6319 3995
rect 10057 3961 10091 3995
rect 12265 3961 12299 3995
rect 16589 3961 16623 3995
rect 17509 3961 17543 3995
rect 9229 3893 9263 3927
rect 8309 3689 8343 3723
rect 12633 3689 12667 3723
rect 8953 3621 8987 3655
rect 7389 3553 7423 3587
rect 13369 3553 13403 3587
rect 1317 3485 1351 3519
rect 2421 3485 2455 3519
rect 7665 3485 7699 3519
rect 8309 3485 8343 3519
rect 8953 3485 8987 3519
rect 10333 3485 10367 3519
rect 10885 3485 10919 3519
rect 11989 3485 12023 3519
rect 12173 3485 12207 3519
rect 12633 3485 12667 3519
rect 12817 3485 12851 3519
rect 15577 3485 15611 3519
rect 1869 3417 1903 3451
rect 3433 3417 3467 3451
rect 11253 3417 11287 3451
rect 13645 3417 13679 3451
rect 15853 3417 15887 3451
rect 1133 3349 1167 3383
rect 4721 3349 4755 3383
rect 5917 3349 5951 3383
rect 10241 3349 10275 3383
rect 12081 3349 12115 3383
rect 15117 3349 15151 3383
rect 17325 3349 17359 3383
rect 1409 3145 1443 3179
rect 5733 3145 5767 3179
rect 13645 3145 13679 3179
rect 14381 3145 14415 3179
rect 16037 3145 16071 3179
rect 17509 3145 17543 3179
rect 857 3077 891 3111
rect 2881 3077 2915 3111
rect 6377 3077 6411 3111
rect 11069 3077 11103 3111
rect 765 3009 799 3043
rect 949 3009 983 3043
rect 3617 3009 3651 3043
rect 3884 3009 3918 3043
rect 5641 3009 5675 3043
rect 6285 3009 6319 3043
rect 6929 3009 6963 3043
rect 9505 3009 9539 3043
rect 13645 3009 13679 3043
rect 14289 3009 14323 3043
rect 14473 3009 14507 3043
rect 14933 3009 14967 3043
rect 15117 3009 15151 3043
rect 16037 3009 16071 3043
rect 16681 3009 16715 3043
rect 16865 3009 16899 3043
rect 17325 3009 17359 3043
rect 3157 2941 3191 2975
rect 7205 2941 7239 2975
rect 8677 2941 8711 2975
rect 10793 2941 10827 2975
rect 15025 2941 15059 2975
rect 16773 2941 16807 2975
rect 4997 2873 5031 2907
rect 10149 2805 10183 2839
rect 12541 2805 12575 2839
rect 1133 2601 1167 2635
rect 1685 2601 1719 2635
rect 3065 2533 3099 2567
rect 6285 2533 6319 2567
rect 6745 2533 6779 2567
rect 7389 2533 7423 2567
rect 8309 2533 8343 2567
rect 9597 2533 9631 2567
rect 13369 2533 13403 2567
rect 15393 2533 15427 2567
rect 4445 2465 4479 2499
rect 4997 2465 5031 2499
rect 11437 2465 11471 2499
rect 12633 2465 12667 2499
rect 949 2397 983 2431
rect 1133 2397 1167 2431
rect 1777 2397 1811 2431
rect 2513 2397 2547 2431
rect 4905 2397 4939 2431
rect 5641 2397 5675 2431
rect 6745 2397 6779 2431
rect 6929 2397 6963 2431
rect 7389 2397 7423 2431
rect 7573 2397 7607 2431
rect 8401 2397 8435 2431
rect 9137 2397 9171 2431
rect 10241 2397 10275 2431
rect 10885 2397 10919 2431
rect 12081 2397 12115 2431
rect 13369 2397 13403 2431
rect 13553 2397 13587 2431
rect 14013 2397 14047 2431
rect 14197 2397 14231 2431
rect 15209 2397 15243 2431
rect 15393 2397 15427 2431
rect 16037 2397 16071 2431
rect 16221 2397 16255 2431
rect 16865 2397 16899 2431
rect 2329 2329 2363 2363
rect 4200 2329 4234 2363
rect 14105 2329 14139 2363
rect 8953 2261 8987 2295
rect 16129 2261 16163 2295
rect 16681 2261 16715 2295
<< metal1 >>
rect 10778 5584 10784 5636
rect 10836 5624 10842 5636
rect 10836 5596 16574 5624
rect 10836 5584 10842 5596
rect 14090 5516 14096 5568
rect 14148 5556 14154 5568
rect 16114 5556 16120 5568
rect 14148 5528 16120 5556
rect 14148 5516 14154 5528
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 16546 5556 16574 5596
rect 16666 5556 16672 5568
rect 16546 5528 16672 5556
rect 16666 5516 16672 5528
rect 16724 5516 16730 5568
rect 368 5466 18308 5488
rect 368 5414 6194 5466
rect 6246 5414 6258 5466
rect 6310 5414 6322 5466
rect 6374 5414 6386 5466
rect 6438 5414 6450 5466
rect 6502 5414 12174 5466
rect 12226 5414 12238 5466
rect 12290 5414 12302 5466
rect 12354 5414 12366 5466
rect 12418 5414 12430 5466
rect 12482 5414 18308 5466
rect 368 5392 18308 5414
rect 3878 5352 3884 5364
rect 2148 5324 3884 5352
rect 2148 5284 2176 5324
rect 3878 5312 3884 5324
rect 3936 5312 3942 5364
rect 4062 5352 4068 5364
rect 4023 5324 4068 5352
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4890 5352 4896 5364
rect 4851 5324 4896 5352
rect 4890 5312 4896 5324
rect 4948 5312 4954 5364
rect 8478 5352 8484 5364
rect 8439 5324 8484 5352
rect 8478 5312 8484 5324
rect 8536 5312 8542 5364
rect 9398 5352 9404 5364
rect 9359 5324 9404 5352
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 15194 5312 15200 5364
rect 15252 5352 15258 5364
rect 16853 5355 16911 5361
rect 16853 5352 16865 5355
rect 15252 5324 16865 5352
rect 15252 5312 15258 5324
rect 16853 5321 16865 5324
rect 16899 5321 16911 5355
rect 16853 5315 16911 5321
rect 1794 5256 2176 5284
rect 2225 5287 2283 5293
rect 2225 5253 2237 5287
rect 2271 5284 2283 5287
rect 5626 5284 5632 5296
rect 2271 5256 5632 5284
rect 2271 5253 2283 5256
rect 2225 5247 2283 5253
rect 5626 5244 5632 5256
rect 5684 5244 5690 5296
rect 8202 5284 8208 5296
rect 7222 5256 8208 5284
rect 8202 5244 8208 5256
rect 8260 5244 8266 5296
rect 12434 5284 12440 5296
rect 12282 5256 12440 5284
rect 12434 5244 12440 5256
rect 12492 5244 12498 5296
rect 15010 5284 15016 5296
rect 14674 5256 15016 5284
rect 15010 5244 15016 5256
rect 15068 5244 15074 5296
rect 15105 5287 15163 5293
rect 15105 5253 15117 5287
rect 15151 5284 15163 5287
rect 17497 5287 17555 5293
rect 17497 5284 17509 5287
rect 15151 5256 17509 5284
rect 15151 5253 15163 5256
rect 15105 5247 15163 5253
rect 17497 5253 17509 5256
rect 17543 5253 17555 5287
rect 17497 5247 17555 5253
rect 3050 5216 3056 5228
rect 3011 5188 3056 5216
rect 3050 5176 3056 5188
rect 3108 5176 3114 5228
rect 3970 5216 3976 5228
rect 3160 5188 3976 5216
rect 2501 5151 2559 5157
rect 2501 5117 2513 5151
rect 2547 5148 2559 5151
rect 2958 5148 2964 5160
rect 2547 5120 2964 5148
rect 2547 5117 2559 5120
rect 2501 5111 2559 5117
rect 2958 5108 2964 5120
rect 3016 5108 3022 5160
rect 753 5015 811 5021
rect 753 4981 765 5015
rect 799 5012 811 5015
rect 3160 5012 3188 5188
rect 3970 5176 3976 5188
rect 4028 5216 4034 5228
rect 4249 5219 4307 5225
rect 4249 5216 4261 5219
rect 4028 5188 4261 5216
rect 4028 5176 4034 5188
rect 4249 5185 4261 5188
rect 4295 5185 4307 5219
rect 4249 5179 4307 5185
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5216 5135 5219
rect 8662 5216 8668 5228
rect 5123 5188 5764 5216
rect 8623 5188 8668 5216
rect 5123 5185 5135 5188
rect 5077 5179 5135 5185
rect 4264 5148 4292 5179
rect 5736 5160 5764 5188
rect 8662 5176 8668 5188
rect 8720 5176 8726 5228
rect 9030 5176 9036 5228
rect 9088 5216 9094 5228
rect 9217 5219 9275 5225
rect 9217 5216 9229 5219
rect 9088 5188 9229 5216
rect 9088 5176 9094 5188
rect 9217 5185 9229 5188
rect 9263 5185 9275 5219
rect 9217 5179 9275 5185
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5216 10195 5219
rect 10778 5216 10784 5228
rect 10183 5188 10784 5216
rect 10183 5185 10195 5188
rect 10137 5179 10195 5185
rect 10778 5176 10784 5188
rect 10836 5176 10842 5228
rect 15381 5219 15439 5225
rect 15381 5185 15393 5219
rect 15427 5216 15439 5219
rect 15746 5216 15752 5228
rect 15427 5188 15752 5216
rect 15427 5185 15439 5188
rect 15381 5179 15439 5185
rect 15746 5176 15752 5188
rect 15804 5176 15810 5228
rect 15930 5216 15936 5228
rect 15891 5188 15936 5216
rect 15930 5176 15936 5188
rect 15988 5176 15994 5228
rect 16666 5216 16672 5228
rect 16627 5188 16672 5216
rect 16666 5176 16672 5188
rect 16724 5176 16730 5228
rect 17310 5176 17316 5228
rect 17368 5216 17374 5228
rect 17405 5219 17463 5225
rect 17405 5216 17417 5219
rect 17368 5188 17417 5216
rect 17368 5176 17374 5188
rect 17405 5185 17417 5188
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 5534 5148 5540 5160
rect 4264 5120 5540 5148
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 5718 5148 5724 5160
rect 5679 5120 5724 5148
rect 5718 5108 5724 5120
rect 5776 5108 5782 5160
rect 5997 5151 6055 5157
rect 5997 5117 6009 5151
rect 6043 5148 6055 5151
rect 6454 5148 6460 5160
rect 6043 5120 6460 5148
rect 6043 5117 6055 5120
rect 5997 5111 6055 5117
rect 6454 5108 6460 5120
rect 6512 5108 6518 5160
rect 11057 5151 11115 5157
rect 11057 5117 11069 5151
rect 11103 5148 11115 5151
rect 12618 5148 12624 5160
rect 11103 5120 12624 5148
rect 11103 5117 11115 5120
rect 11057 5111 11115 5117
rect 12618 5108 12624 5120
rect 12676 5108 12682 5160
rect 17310 5080 17316 5092
rect 15304 5052 17316 5080
rect 799 4984 3188 5012
rect 3237 5015 3295 5021
rect 799 4981 811 4984
rect 753 4975 811 4981
rect 3237 4981 3249 5015
rect 3283 5012 3295 5015
rect 3786 5012 3792 5024
rect 3283 4984 3792 5012
rect 3283 4981 3295 4984
rect 3237 4975 3295 4981
rect 3786 4972 3792 4984
rect 3844 4972 3850 5024
rect 3878 4972 3884 5024
rect 3936 5012 3942 5024
rect 6730 5012 6736 5024
rect 3936 4984 6736 5012
rect 3936 4972 3942 4984
rect 6730 4972 6736 4984
rect 6788 4972 6794 5024
rect 7466 5012 7472 5024
rect 7427 4984 7472 5012
rect 7466 4972 7472 4984
rect 7524 4972 7530 5024
rect 10137 5015 10195 5021
rect 10137 4981 10149 5015
rect 10183 5012 10195 5015
rect 11146 5012 11152 5024
rect 10183 4984 11152 5012
rect 10183 4981 10195 4984
rect 10137 4975 10195 4981
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 12526 5012 12532 5024
rect 12487 4984 12532 5012
rect 12526 4972 12532 4984
rect 12584 4972 12590 5024
rect 13633 5015 13691 5021
rect 13633 4981 13645 5015
rect 13679 5012 13691 5015
rect 15304 5012 15332 5052
rect 17310 5040 17316 5052
rect 17368 5040 17374 5092
rect 16114 5012 16120 5024
rect 13679 4984 15332 5012
rect 16075 4984 16120 5012
rect 13679 4981 13691 4984
rect 13633 4975 13691 4981
rect 16114 4972 16120 4984
rect 16172 4972 16178 5024
rect 368 4922 18308 4944
rect 368 4870 3204 4922
rect 3256 4870 3268 4922
rect 3320 4870 3332 4922
rect 3384 4870 3396 4922
rect 3448 4870 3460 4922
rect 3512 4870 9184 4922
rect 9236 4870 9248 4922
rect 9300 4870 9312 4922
rect 9364 4870 9376 4922
rect 9428 4870 9440 4922
rect 9492 4870 15164 4922
rect 15216 4870 15228 4922
rect 15280 4870 15292 4922
rect 15344 4870 15356 4922
rect 15408 4870 15420 4922
rect 15472 4870 18308 4922
rect 368 4848 18308 4870
rect 1394 4808 1400 4820
rect 1355 4780 1400 4808
rect 1394 4768 1400 4780
rect 1452 4768 1458 4820
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 3237 4811 3295 4817
rect 3237 4808 3249 4811
rect 2832 4780 3249 4808
rect 2832 4768 2838 4780
rect 3237 4777 3249 4780
rect 3283 4777 3295 4811
rect 6454 4808 6460 4820
rect 6415 4780 6460 4808
rect 3237 4771 3295 4777
rect 6454 4768 6460 4780
rect 6512 4768 6518 4820
rect 7190 4768 7196 4820
rect 7248 4808 7254 4820
rect 7377 4811 7435 4817
rect 7377 4808 7389 4811
rect 7248 4780 7389 4808
rect 7248 4768 7254 4780
rect 7377 4777 7389 4780
rect 7423 4777 7435 4811
rect 8202 4808 8208 4820
rect 8163 4780 8208 4808
rect 7377 4771 7435 4777
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 10778 4808 10784 4820
rect 9723 4780 10784 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 11606 4768 11612 4820
rect 11664 4808 11670 4820
rect 11977 4811 12035 4817
rect 11977 4808 11989 4811
rect 11664 4780 11989 4808
rect 11664 4768 11670 4780
rect 11977 4777 11989 4780
rect 12023 4777 12035 4811
rect 11977 4771 12035 4777
rect 12618 4768 12624 4820
rect 12676 4808 12682 4820
rect 12713 4811 12771 4817
rect 12713 4808 12725 4811
rect 12676 4780 12725 4808
rect 12676 4768 12682 4780
rect 12713 4777 12725 4780
rect 12759 4777 12771 4811
rect 12713 4771 12771 4777
rect 16022 4768 16028 4820
rect 16080 4808 16086 4820
rect 16669 4811 16727 4817
rect 16669 4808 16681 4811
rect 16080 4780 16681 4808
rect 16080 4768 16086 4780
rect 16669 4777 16681 4780
rect 16715 4777 16727 4811
rect 17402 4808 17408 4820
rect 17363 4780 17408 4808
rect 16669 4771 16727 4777
rect 17402 4768 17408 4780
rect 17460 4768 17466 4820
rect 9217 4743 9275 4749
rect 9217 4709 9229 4743
rect 9263 4740 9275 4743
rect 9263 4712 10088 4740
rect 9263 4709 9275 4712
rect 9217 4703 9275 4709
rect 3970 4672 3976 4684
rect 3931 4644 3976 4672
rect 3970 4632 3976 4644
rect 4028 4632 4034 4684
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 5994 4672 6000 4684
rect 4295 4644 6000 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 5994 4632 6000 4644
rect 6052 4632 6058 4684
rect 6914 4632 6920 4684
rect 6972 4672 6978 4684
rect 6972 4644 8248 4672
rect 6972 4632 6978 4644
rect 1210 4604 1216 4616
rect 1171 4576 1216 4604
rect 1210 4564 1216 4576
rect 1268 4564 1274 4616
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4604 2283 4607
rect 2958 4604 2964 4616
rect 2271 4576 2964 4604
rect 2271 4573 2283 4576
rect 2225 4567 2283 4573
rect 2958 4564 2964 4576
rect 3016 4604 3022 4616
rect 3053 4607 3111 4613
rect 3053 4604 3065 4607
rect 3016 4576 3065 4604
rect 3016 4564 3022 4576
rect 3053 4573 3065 4576
rect 3099 4573 3111 4607
rect 3053 4567 3111 4573
rect 5350 4564 5356 4616
rect 5408 4564 5414 4616
rect 6641 4607 6699 4613
rect 6641 4573 6653 4607
rect 6687 4604 6699 4607
rect 7466 4604 7472 4616
rect 6687 4576 7472 4604
rect 6687 4573 6699 4576
rect 6641 4567 6699 4573
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 7561 4607 7619 4613
rect 7561 4573 7573 4607
rect 7607 4604 7619 4607
rect 8110 4604 8116 4616
rect 7607 4576 8116 4604
rect 7607 4573 7619 4576
rect 7561 4567 7619 4573
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 8220 4613 8248 4644
rect 8205 4607 8263 4613
rect 8205 4573 8217 4607
rect 8251 4573 8263 4607
rect 8205 4567 8263 4573
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 9033 4607 9091 4613
rect 9033 4573 9045 4607
rect 9079 4604 9091 4607
rect 9122 4604 9128 4616
rect 9079 4576 9128 4604
rect 9079 4573 9091 4576
rect 9033 4567 9091 4573
rect 1486 4496 1492 4548
rect 1544 4536 1550 4548
rect 1949 4539 2007 4545
rect 1949 4536 1961 4539
rect 1544 4508 1961 4536
rect 1544 4496 1550 4508
rect 1949 4505 1961 4508
rect 1995 4505 2007 4539
rect 1949 4499 2007 4505
rect 7374 4496 7380 4548
rect 7432 4536 7438 4548
rect 8404 4536 8432 4567
rect 9122 4564 9128 4576
rect 9180 4564 9186 4616
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4604 9275 4607
rect 9263 4576 9812 4604
rect 10060 4590 10088 4712
rect 11146 4672 11152 4684
rect 11107 4644 11152 4672
rect 11146 4632 11152 4644
rect 11204 4632 11210 4684
rect 12526 4632 12532 4684
rect 12584 4672 12590 4684
rect 14553 4675 14611 4681
rect 12584 4644 14320 4672
rect 12584 4632 12590 4644
rect 11425 4607 11483 4613
rect 9263 4573 9275 4576
rect 9217 4567 9275 4573
rect 7432 4508 8432 4536
rect 7432 4496 7438 4508
rect 5718 4468 5724 4480
rect 5679 4440 5724 4468
rect 5718 4428 5724 4440
rect 5776 4428 5782 4480
rect 9784 4468 9812 4576
rect 11425 4573 11437 4607
rect 11471 4573 11483 4607
rect 11425 4567 11483 4573
rect 12161 4607 12219 4613
rect 12161 4573 12173 4607
rect 12207 4604 12219 4607
rect 12618 4604 12624 4616
rect 12207 4576 12624 4604
rect 12207 4573 12219 4576
rect 12161 4567 12219 4573
rect 11440 4536 11468 4567
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 12820 4613 12848 4644
rect 12805 4607 12863 4613
rect 12805 4573 12817 4607
rect 12851 4573 12863 4607
rect 13633 4607 13691 4613
rect 13633 4604 13645 4607
rect 12805 4567 12863 4573
rect 12912 4576 13645 4604
rect 12912 4536 12940 4576
rect 13633 4573 13645 4576
rect 13679 4604 13691 4607
rect 14182 4604 14188 4616
rect 13679 4576 14188 4604
rect 13679 4573 13691 4576
rect 13633 4567 13691 4573
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 14292 4613 14320 4644
rect 14553 4641 14565 4675
rect 14599 4672 14611 4675
rect 15194 4672 15200 4684
rect 14599 4644 15200 4672
rect 14599 4641 14611 4644
rect 14553 4635 14611 4641
rect 15194 4632 15200 4644
rect 15252 4632 15258 4684
rect 15746 4632 15752 4684
rect 15804 4672 15810 4684
rect 16025 4675 16083 4681
rect 16025 4672 16037 4675
rect 15804 4644 16037 4672
rect 15804 4632 15810 4644
rect 16025 4641 16037 4644
rect 16071 4672 16083 4675
rect 16071 4644 17264 4672
rect 16071 4641 16083 4644
rect 16025 4635 16083 4641
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 11440 4508 12940 4536
rect 13170 4496 13176 4548
rect 13228 4536 13234 4548
rect 13357 4539 13415 4545
rect 13357 4536 13369 4539
rect 13228 4508 13369 4536
rect 13228 4496 13234 4508
rect 13357 4505 13369 4508
rect 13403 4505 13415 4539
rect 14292 4536 14320 4567
rect 15654 4564 15660 4616
rect 15712 4564 15718 4616
rect 17236 4613 17264 4644
rect 16485 4607 16543 4613
rect 16485 4573 16497 4607
rect 16531 4573 16543 4607
rect 16485 4567 16543 4573
rect 17221 4607 17279 4613
rect 17221 4573 17233 4607
rect 17267 4573 17279 4607
rect 17221 4567 17279 4573
rect 16500 4536 16528 4567
rect 14292 4508 14412 4536
rect 13357 4499 13415 4505
rect 11054 4468 11060 4480
rect 9784 4440 11060 4468
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 14384 4468 14412 4508
rect 15856 4508 16528 4536
rect 15856 4468 15884 4508
rect 14384 4440 15884 4468
rect 368 4378 18308 4400
rect 368 4326 6194 4378
rect 6246 4326 6258 4378
rect 6310 4326 6322 4378
rect 6374 4326 6386 4378
rect 6438 4326 6450 4378
rect 6502 4326 12174 4378
rect 12226 4326 12238 4378
rect 12290 4326 12302 4378
rect 12354 4326 12366 4378
rect 12418 4326 12430 4378
rect 12482 4326 18308 4378
rect 368 4304 18308 4326
rect 1118 4224 1124 4276
rect 1176 4264 1182 4276
rect 2958 4264 2964 4276
rect 1176 4236 1624 4264
rect 2919 4236 2964 4264
rect 1176 4224 1182 4236
rect 1486 4196 1492 4208
rect 1447 4168 1492 4196
rect 1486 4156 1492 4168
rect 1544 4156 1550 4208
rect 1596 4196 1624 4236
rect 2958 4224 2964 4236
rect 3016 4224 3022 4276
rect 9122 4224 9128 4276
rect 9180 4264 9186 4276
rect 11238 4264 11244 4276
rect 9180 4236 11244 4264
rect 9180 4224 9186 4236
rect 11238 4224 11244 4236
rect 11296 4224 11302 4276
rect 14090 4264 14096 4276
rect 13004 4236 14096 4264
rect 3789 4199 3847 4205
rect 1596 4168 1978 4196
rect 3789 4165 3801 4199
rect 3835 4196 3847 4199
rect 4154 4196 4160 4208
rect 3835 4168 4160 4196
rect 3835 4165 3847 4168
rect 3789 4159 3847 4165
rect 4154 4156 4160 4168
rect 4212 4156 4218 4208
rect 13004 4196 13032 4236
rect 14090 4224 14096 4236
rect 14148 4224 14154 4276
rect 14182 4224 14188 4276
rect 14240 4264 14246 4276
rect 14645 4267 14703 4273
rect 14645 4264 14657 4267
rect 14240 4236 14657 4264
rect 14240 4224 14246 4236
rect 14645 4233 14657 4236
rect 14691 4264 14703 4267
rect 15930 4264 15936 4276
rect 14691 4236 15936 4264
rect 14691 4233 14703 4236
rect 14645 4227 14703 4233
rect 15930 4224 15936 4236
rect 15988 4224 15994 4276
rect 13170 4196 13176 4208
rect 8970 4168 13032 4196
rect 13131 4168 13176 4196
rect 13170 4156 13176 4168
rect 13228 4156 13234 4208
rect 14398 4168 16068 4196
rect 4982 4128 4988 4140
rect 4943 4100 4988 4128
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 6457 4131 6515 4137
rect 6457 4097 6469 4131
rect 6503 4128 6515 4131
rect 7466 4128 7472 4140
rect 6503 4100 7472 4128
rect 6503 4097 6515 4100
rect 6457 4091 6515 4097
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 10229 4131 10287 4137
rect 10229 4097 10241 4131
rect 10275 4128 10287 4131
rect 10318 4128 10324 4140
rect 10275 4100 10324 4128
rect 10275 4097 10287 4100
rect 10229 4091 10287 4097
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 11054 4128 11060 4140
rect 11015 4100 11060 4128
rect 11054 4088 11060 4100
rect 11112 4088 11118 4140
rect 11606 4128 11612 4140
rect 11567 4100 11612 4128
rect 11606 4088 11612 4100
rect 11664 4088 11670 4140
rect 12437 4131 12495 4137
rect 12437 4097 12449 4131
rect 12483 4128 12495 4131
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12483 4100 12909 4128
rect 12483 4097 12495 4100
rect 12437 4091 12495 4097
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 15194 4128 15200 4140
rect 15155 4100 15200 4128
rect 12897 4091 12955 4097
rect 1210 4060 1216 4072
rect 1171 4032 1216 4060
rect 1210 4020 1216 4032
rect 1268 4020 1274 4072
rect 4709 4063 4767 4069
rect 4709 4060 4721 4063
rect 1320 4032 4721 4060
rect 750 3952 756 4004
rect 808 3992 814 4004
rect 1320 3992 1348 4032
rect 4709 4029 4721 4032
rect 4755 4060 4767 4063
rect 7006 4060 7012 4072
rect 4755 4032 7012 4060
rect 4755 4029 4767 4032
rect 4709 4023 4767 4029
rect 7006 4020 7012 4032
rect 7064 4060 7070 4072
rect 7374 4060 7380 4072
rect 7064 4032 7380 4060
rect 7064 4020 7070 4032
rect 7374 4020 7380 4032
rect 7432 4020 7438 4072
rect 7745 4063 7803 4069
rect 7745 4029 7757 4063
rect 7791 4060 7803 4063
rect 8294 4060 8300 4072
rect 7791 4032 8300 4060
rect 7791 4029 7803 4032
rect 7745 4023 7803 4029
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 11238 4020 11244 4072
rect 11296 4060 11302 4072
rect 12802 4060 12808 4072
rect 11296 4032 12808 4060
rect 11296 4020 11302 4032
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 12912 4060 12940 4091
rect 15194 4088 15200 4100
rect 15252 4088 15258 4140
rect 15289 4131 15347 4137
rect 15289 4097 15301 4131
rect 15335 4128 15347 4131
rect 15746 4128 15752 4140
rect 15335 4100 15752 4128
rect 15335 4097 15347 4100
rect 15289 4091 15347 4097
rect 15746 4088 15752 4100
rect 15804 4088 15810 4140
rect 15930 4128 15936 4140
rect 15891 4100 15936 4128
rect 15930 4088 15936 4100
rect 15988 4088 15994 4140
rect 16040 4137 16068 4168
rect 16025 4131 16083 4137
rect 16025 4097 16037 4131
rect 16071 4097 16083 4131
rect 16025 4091 16083 4097
rect 16114 4088 16120 4140
rect 16172 4128 16178 4140
rect 16172 4100 16217 4128
rect 16172 4088 16178 4100
rect 16574 4088 16580 4140
rect 16632 4128 16638 4140
rect 16761 4131 16819 4137
rect 16632 4100 16677 4128
rect 16632 4088 16638 4100
rect 16761 4097 16773 4131
rect 16807 4097 16819 4131
rect 17310 4128 17316 4140
rect 17271 4100 17316 4128
rect 16761 4091 16819 4097
rect 13538 4060 13544 4072
rect 12912 4032 13544 4060
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 16132 4060 16160 4088
rect 16776 4060 16804 4091
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 16132 4032 16804 4060
rect 808 3964 1348 3992
rect 808 3952 814 3964
rect 2958 3952 2964 4004
rect 3016 3992 3022 4004
rect 3605 3995 3663 4001
rect 3605 3992 3617 3995
rect 3016 3964 3617 3992
rect 3016 3952 3022 3964
rect 3605 3961 3617 3964
rect 3651 3961 3663 3995
rect 3605 3955 3663 3961
rect 6086 3952 6092 4004
rect 6144 3992 6150 4004
rect 6273 3995 6331 4001
rect 6273 3992 6285 3995
rect 6144 3964 6285 3992
rect 6144 3952 6150 3964
rect 6273 3961 6285 3964
rect 6319 3961 6331 3995
rect 6273 3955 6331 3961
rect 10045 3995 10103 4001
rect 10045 3961 10057 3995
rect 10091 3992 10103 3995
rect 10502 3992 10508 4004
rect 10091 3964 10508 3992
rect 10091 3961 10103 3964
rect 10045 3955 10103 3961
rect 10502 3952 10508 3964
rect 10560 3952 10566 4004
rect 12253 3995 12311 4001
rect 12253 3961 12265 3995
rect 12299 3992 12311 3995
rect 12710 3992 12716 4004
rect 12299 3964 12716 3992
rect 12299 3961 12311 3964
rect 12253 3955 12311 3961
rect 12710 3952 12716 3964
rect 12768 3952 12774 4004
rect 15654 3952 15660 4004
rect 15712 3992 15718 4004
rect 16577 3995 16635 4001
rect 16577 3992 16589 3995
rect 15712 3964 16589 3992
rect 15712 3952 15718 3964
rect 16577 3961 16589 3964
rect 16623 3961 16635 3995
rect 16577 3955 16635 3961
rect 17497 3995 17555 4001
rect 17497 3961 17509 3995
rect 17543 3992 17555 3995
rect 18230 3992 18236 4004
rect 17543 3964 18236 3992
rect 17543 3961 17555 3964
rect 17497 3955 17555 3961
rect 18230 3952 18236 3964
rect 18288 3952 18294 4004
rect 8202 3884 8208 3936
rect 8260 3924 8266 3936
rect 9217 3927 9275 3933
rect 9217 3924 9229 3927
rect 8260 3896 9229 3924
rect 8260 3884 8266 3896
rect 9217 3893 9229 3896
rect 9263 3893 9275 3927
rect 9217 3887 9275 3893
rect 12342 3884 12348 3936
rect 12400 3924 12406 3936
rect 15930 3924 15936 3936
rect 12400 3896 15936 3924
rect 12400 3884 12406 3896
rect 15930 3884 15936 3896
rect 15988 3924 15994 3936
rect 16482 3924 16488 3936
rect 15988 3896 16488 3924
rect 15988 3884 15994 3896
rect 16482 3884 16488 3896
rect 16540 3884 16546 3936
rect 368 3834 18308 3856
rect 368 3782 3204 3834
rect 3256 3782 3268 3834
rect 3320 3782 3332 3834
rect 3384 3782 3396 3834
rect 3448 3782 3460 3834
rect 3512 3782 9184 3834
rect 9236 3782 9248 3834
rect 9300 3782 9312 3834
rect 9364 3782 9376 3834
rect 9428 3782 9440 3834
rect 9492 3782 15164 3834
rect 15216 3782 15228 3834
rect 15280 3782 15292 3834
rect 15344 3782 15356 3834
rect 15408 3782 15420 3834
rect 15472 3782 18308 3834
rect 368 3760 18308 3782
rect 8294 3720 8300 3732
rect 2424 3692 8156 3720
rect 8255 3692 8300 3720
rect 1302 3516 1308 3528
rect 1263 3488 1308 3516
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 2424 3525 2452 3692
rect 8128 3652 8156 3692
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 12526 3680 12532 3732
rect 12584 3720 12590 3732
rect 12621 3723 12679 3729
rect 12621 3720 12633 3723
rect 12584 3692 12633 3720
rect 12584 3680 12590 3692
rect 12621 3689 12633 3692
rect 12667 3689 12679 3723
rect 12621 3683 12679 3689
rect 12802 3680 12808 3732
rect 12860 3720 12866 3732
rect 16022 3720 16028 3732
rect 12860 3692 16028 3720
rect 12860 3680 12866 3692
rect 16022 3680 16028 3692
rect 16080 3680 16086 3732
rect 8846 3652 8852 3664
rect 8128 3624 8852 3652
rect 8846 3612 8852 3624
rect 8904 3612 8910 3664
rect 8941 3655 8999 3661
rect 8941 3621 8953 3655
rect 8987 3621 8999 3655
rect 8941 3615 8999 3621
rect 7377 3587 7435 3593
rect 7377 3553 7389 3587
rect 7423 3584 7435 3587
rect 8956 3584 8984 3615
rect 10686 3612 10692 3664
rect 10744 3652 10750 3664
rect 10744 3624 13492 3652
rect 10744 3612 10750 3624
rect 13357 3587 13415 3593
rect 13357 3584 13369 3587
rect 7423 3556 8984 3584
rect 10336 3556 13369 3584
rect 7423 3553 7435 3556
rect 7377 3547 7435 3553
rect 10336 3528 10364 3556
rect 13357 3553 13369 3556
rect 13403 3553 13415 3587
rect 13464 3584 13492 3624
rect 14182 3584 14188 3596
rect 13464 3556 14188 3584
rect 13357 3547 13415 3553
rect 14182 3544 14188 3556
rect 14240 3584 14246 3596
rect 15102 3584 15108 3596
rect 14240 3556 15108 3584
rect 14240 3544 14246 3556
rect 15102 3544 15108 3556
rect 15160 3544 15166 3596
rect 2409 3519 2467 3525
rect 2409 3485 2421 3519
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 7653 3519 7711 3525
rect 7653 3485 7665 3519
rect 7699 3516 7711 3519
rect 8202 3516 8208 3528
rect 7699 3488 8208 3516
rect 7699 3485 7711 3488
rect 7653 3479 7711 3485
rect 8202 3476 8208 3488
rect 8260 3516 8266 3528
rect 8297 3519 8355 3525
rect 8297 3516 8309 3519
rect 8260 3488 8309 3516
rect 8260 3476 8266 3488
rect 8297 3485 8309 3488
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 8662 3476 8668 3528
rect 8720 3516 8726 3528
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8720 3488 8953 3516
rect 8720 3476 8726 3488
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 10318 3516 10324 3528
rect 10279 3488 10324 3516
rect 8941 3479 8999 3485
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 10686 3476 10692 3528
rect 10744 3516 10750 3528
rect 10873 3519 10931 3525
rect 10873 3516 10885 3519
rect 10744 3488 10885 3516
rect 10744 3476 10750 3488
rect 10873 3485 10885 3488
rect 10919 3485 10931 3519
rect 10873 3479 10931 3485
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11974 3516 11980 3528
rect 11112 3488 11836 3516
rect 11935 3488 11980 3516
rect 11112 3476 11118 3488
rect 1026 3408 1032 3460
rect 1084 3448 1090 3460
rect 1857 3451 1915 3457
rect 1857 3448 1869 3451
rect 1084 3420 1869 3448
rect 1084 3408 1090 3420
rect 1857 3417 1869 3420
rect 1903 3417 1915 3451
rect 3418 3448 3424 3460
rect 3379 3420 3424 3448
rect 1857 3411 1915 3417
rect 3418 3408 3424 3420
rect 3476 3408 3482 3460
rect 11146 3448 11152 3460
rect 6946 3420 11152 3448
rect 11146 3408 11152 3420
rect 11204 3408 11210 3460
rect 11238 3408 11244 3460
rect 11296 3448 11302 3460
rect 11808 3448 11836 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 12161 3519 12219 3525
rect 12161 3485 12173 3519
rect 12207 3516 12219 3519
rect 12526 3516 12532 3528
rect 12207 3488 12532 3516
rect 12207 3485 12219 3488
rect 12161 3479 12219 3485
rect 12526 3476 12532 3488
rect 12584 3476 12590 3528
rect 12621 3519 12679 3525
rect 12621 3485 12633 3519
rect 12667 3485 12679 3519
rect 12802 3516 12808 3528
rect 12763 3488 12808 3516
rect 12621 3479 12679 3485
rect 12342 3448 12348 3460
rect 11296 3420 11341 3448
rect 11808 3420 12348 3448
rect 11296 3408 11302 3420
rect 12342 3408 12348 3420
rect 12400 3448 12406 3460
rect 12636 3448 12664 3479
rect 12802 3476 12808 3488
rect 12860 3476 12866 3528
rect 15565 3519 15623 3525
rect 15565 3516 15577 3519
rect 15120 3488 15577 3516
rect 13630 3448 13636 3460
rect 12400 3420 12664 3448
rect 13591 3420 13636 3448
rect 12400 3408 12406 3420
rect 13630 3408 13636 3420
rect 13688 3408 13694 3460
rect 14366 3408 14372 3460
rect 14424 3408 14430 3460
rect 1121 3383 1179 3389
rect 1121 3349 1133 3383
rect 1167 3380 1179 3383
rect 2866 3380 2872 3392
rect 1167 3352 2872 3380
rect 1167 3349 1179 3352
rect 1121 3343 1179 3349
rect 2866 3340 2872 3352
rect 2924 3340 2930 3392
rect 4154 3340 4160 3392
rect 4212 3380 4218 3392
rect 4709 3383 4767 3389
rect 4709 3380 4721 3383
rect 4212 3352 4721 3380
rect 4212 3340 4218 3352
rect 4709 3349 4721 3352
rect 4755 3349 4767 3383
rect 5902 3380 5908 3392
rect 5863 3352 5908 3380
rect 4709 3343 4767 3349
rect 5902 3340 5908 3352
rect 5960 3340 5966 3392
rect 10229 3383 10287 3389
rect 10229 3349 10241 3383
rect 10275 3380 10287 3383
rect 11054 3380 11060 3392
rect 10275 3352 11060 3380
rect 10275 3349 10287 3352
rect 10229 3343 10287 3349
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 12066 3380 12072 3392
rect 12027 3352 12072 3380
rect 12066 3340 12072 3352
rect 12124 3340 12130 3392
rect 13722 3340 13728 3392
rect 13780 3380 13786 3392
rect 15120 3389 15148 3488
rect 15565 3485 15577 3488
rect 15611 3485 15623 3519
rect 15565 3479 15623 3485
rect 15838 3448 15844 3460
rect 15799 3420 15844 3448
rect 15838 3408 15844 3420
rect 15896 3408 15902 3460
rect 16298 3408 16304 3460
rect 16356 3408 16362 3460
rect 15105 3383 15163 3389
rect 15105 3380 15117 3383
rect 13780 3352 15117 3380
rect 13780 3340 13786 3352
rect 15105 3349 15117 3352
rect 15151 3349 15163 3383
rect 15105 3343 15163 3349
rect 16114 3340 16120 3392
rect 16172 3380 16178 3392
rect 17313 3383 17371 3389
rect 17313 3380 17325 3383
rect 16172 3352 17325 3380
rect 16172 3340 16178 3352
rect 17313 3349 17325 3352
rect 17359 3349 17371 3383
rect 17313 3343 17371 3349
rect 368 3290 18308 3312
rect 368 3238 6194 3290
rect 6246 3238 6258 3290
rect 6310 3238 6322 3290
rect 6374 3238 6386 3290
rect 6438 3238 6450 3290
rect 6502 3238 12174 3290
rect 12226 3238 12238 3290
rect 12290 3238 12302 3290
rect 12354 3238 12366 3290
rect 12418 3238 12430 3290
rect 12482 3238 18308 3290
rect 368 3216 18308 3238
rect 1302 3136 1308 3188
rect 1360 3176 1366 3188
rect 1397 3179 1455 3185
rect 1397 3176 1409 3179
rect 1360 3148 1409 3176
rect 1360 3136 1366 3148
rect 1397 3145 1409 3148
rect 1443 3145 1455 3179
rect 1397 3139 1455 3145
rect 5534 3136 5540 3188
rect 5592 3136 5598 3188
rect 5626 3136 5632 3188
rect 5684 3176 5690 3188
rect 5721 3179 5779 3185
rect 5721 3176 5733 3179
rect 5684 3148 5733 3176
rect 5684 3136 5690 3148
rect 5721 3145 5733 3148
rect 5767 3145 5779 3179
rect 5721 3139 5779 3145
rect 5902 3136 5908 3188
rect 5960 3176 5966 3188
rect 8662 3176 8668 3188
rect 5960 3148 8668 3176
rect 5960 3136 5966 3148
rect 845 3111 903 3117
rect 845 3077 857 3111
rect 891 3108 903 3111
rect 2866 3108 2872 3120
rect 891 3080 1702 3108
rect 2827 3080 2872 3108
rect 891 3077 903 3080
rect 845 3071 903 3077
rect 2866 3068 2872 3080
rect 2924 3068 2930 3120
rect 5552 3108 5580 3136
rect 5552 3080 5672 3108
rect 750 3040 756 3052
rect 711 3012 756 3040
rect 750 3000 756 3012
rect 808 3000 814 3052
rect 937 3043 995 3049
rect 937 3009 949 3043
rect 983 3040 995 3043
rect 1026 3040 1032 3052
rect 983 3012 1032 3040
rect 983 3009 995 3012
rect 937 3003 995 3009
rect 1026 3000 1032 3012
rect 1084 3000 1090 3052
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3040 3663 3043
rect 3694 3040 3700 3052
rect 3651 3012 3700 3040
rect 3651 3009 3663 3012
rect 3605 3003 3663 3009
rect 3694 3000 3700 3012
rect 3752 3000 3758 3052
rect 3872 3043 3930 3049
rect 3872 3009 3884 3043
rect 3918 3040 3930 3043
rect 5534 3040 5540 3052
rect 3918 3012 5540 3040
rect 3918 3009 3930 3012
rect 3872 3003 3930 3009
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 5644 3049 5672 3080
rect 5994 3068 6000 3120
rect 6052 3108 6058 3120
rect 6365 3111 6423 3117
rect 6365 3108 6377 3111
rect 6052 3080 6377 3108
rect 6052 3068 6058 3080
rect 6365 3077 6377 3080
rect 6411 3077 6423 3111
rect 6365 3071 6423 3077
rect 5629 3043 5687 3049
rect 5629 3009 5641 3043
rect 5675 3009 5687 3043
rect 5629 3003 5687 3009
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 6932 3049 6960 3148
rect 8662 3136 8668 3148
rect 8720 3136 8726 3188
rect 12066 3176 12072 3188
rect 10888 3148 12072 3176
rect 10888 3108 10916 3148
rect 12066 3136 12072 3148
rect 12124 3136 12130 3188
rect 13630 3176 13636 3188
rect 13591 3148 13636 3176
rect 13630 3136 13636 3148
rect 13688 3136 13694 3188
rect 14366 3176 14372 3188
rect 14327 3148 14372 3176
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 15838 3136 15844 3188
rect 15896 3176 15902 3188
rect 16025 3179 16083 3185
rect 16025 3176 16037 3179
rect 15896 3148 16037 3176
rect 15896 3136 15902 3148
rect 16025 3145 16037 3148
rect 16071 3145 16083 3179
rect 17494 3176 17500 3188
rect 17455 3148 17500 3176
rect 16025 3139 16083 3145
rect 17494 3136 17500 3148
rect 17552 3136 17558 3188
rect 11054 3108 11060 3120
rect 8418 3080 10916 3108
rect 11015 3080 11060 3108
rect 11054 3068 11060 3080
rect 11112 3068 11118 3120
rect 13354 3108 13360 3120
rect 12282 3080 13360 3108
rect 13354 3068 13360 3080
rect 13412 3068 13418 3120
rect 13538 3068 13544 3120
rect 13596 3108 13602 3120
rect 16114 3108 16120 3120
rect 13596 3080 16120 3108
rect 13596 3068 13602 3080
rect 6273 3043 6331 3049
rect 6273 3040 6285 3043
rect 5776 3012 6285 3040
rect 5776 3000 5782 3012
rect 6273 3009 6285 3012
rect 6319 3009 6331 3043
rect 6273 3003 6331 3009
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 9493 3043 9551 3049
rect 9493 3009 9505 3043
rect 9539 3040 9551 3043
rect 9582 3040 9588 3052
rect 9539 3012 9588 3040
rect 9539 3009 9551 3012
rect 9493 3003 9551 3009
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 12618 3000 12624 3052
rect 12676 3040 12682 3052
rect 13633 3043 13691 3049
rect 13633 3040 13645 3043
rect 12676 3012 13645 3040
rect 12676 3000 12682 3012
rect 13633 3009 13645 3012
rect 13679 3040 13691 3043
rect 13722 3040 13728 3052
rect 13679 3012 13728 3040
rect 13679 3009 13691 3012
rect 13633 3003 13691 3009
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 14458 3040 14464 3052
rect 14419 3012 14464 3040
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 14826 3000 14832 3052
rect 14884 3040 14890 3052
rect 14921 3043 14979 3049
rect 14921 3040 14933 3043
rect 14884 3012 14933 3040
rect 14884 3000 14890 3012
rect 14921 3009 14933 3012
rect 14967 3009 14979 3043
rect 15102 3040 15108 3052
rect 15063 3012 15108 3040
rect 14921 3003 14979 3009
rect 15102 3000 15108 3012
rect 15160 3000 15166 3052
rect 16040 3049 16068 3080
rect 16114 3068 16120 3080
rect 16172 3068 16178 3120
rect 16390 3068 16396 3120
rect 16448 3108 16454 3120
rect 16448 3080 16896 3108
rect 16448 3068 16454 3080
rect 16025 3043 16083 3049
rect 16025 3009 16037 3043
rect 16071 3009 16083 3043
rect 16025 3003 16083 3009
rect 16482 3000 16488 3052
rect 16540 3040 16546 3052
rect 16868 3049 16896 3080
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 16540 3012 16681 3040
rect 16540 3000 16546 3012
rect 16669 3009 16681 3012
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 17313 3043 17371 3049
rect 17313 3009 17325 3043
rect 17359 3009 17371 3043
rect 17313 3003 17371 3009
rect 3145 2975 3203 2981
rect 3145 2941 3157 2975
rect 3191 2972 3203 2975
rect 7193 2975 7251 2981
rect 3191 2944 3648 2972
rect 3191 2941 3203 2944
rect 3145 2935 3203 2941
rect 3620 2916 3648 2944
rect 7193 2941 7205 2975
rect 7239 2972 7251 2975
rect 7239 2944 8248 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 3602 2864 3608 2916
rect 3660 2864 3666 2916
rect 4982 2904 4988 2916
rect 4895 2876 4988 2904
rect 4982 2864 4988 2876
rect 5040 2904 5046 2916
rect 8220 2904 8248 2944
rect 8386 2932 8392 2984
rect 8444 2972 8450 2984
rect 8665 2975 8723 2981
rect 8665 2972 8677 2975
rect 8444 2944 8677 2972
rect 8444 2932 8450 2944
rect 8665 2941 8677 2944
rect 8711 2972 8723 2975
rect 9030 2972 9036 2984
rect 8711 2944 9036 2972
rect 8711 2941 8723 2944
rect 8665 2935 8723 2941
rect 9030 2932 9036 2944
rect 9088 2972 9094 2984
rect 10781 2975 10839 2981
rect 10781 2972 10793 2975
rect 9088 2944 10793 2972
rect 9088 2932 9094 2944
rect 10781 2941 10793 2944
rect 10827 2941 10839 2975
rect 10781 2935 10839 2941
rect 11146 2932 11152 2984
rect 11204 2972 11210 2984
rect 15013 2975 15071 2981
rect 15013 2972 15025 2975
rect 11204 2944 15025 2972
rect 11204 2932 11210 2944
rect 15013 2941 15025 2944
rect 15059 2941 15071 2975
rect 15013 2935 15071 2941
rect 16761 2975 16819 2981
rect 16761 2941 16773 2975
rect 16807 2972 16819 2975
rect 17328 2972 17356 3003
rect 16807 2944 17356 2972
rect 16807 2941 16819 2944
rect 16761 2935 16819 2941
rect 8294 2904 8300 2916
rect 5040 2876 6914 2904
rect 8220 2876 8300 2904
rect 5040 2864 5046 2876
rect 6886 2836 6914 2876
rect 8294 2864 8300 2876
rect 8352 2864 8358 2916
rect 10686 2904 10692 2916
rect 9968 2876 10692 2904
rect 9968 2836 9996 2876
rect 10686 2864 10692 2876
rect 10744 2864 10750 2916
rect 12066 2864 12072 2916
rect 12124 2904 12130 2916
rect 14274 2904 14280 2916
rect 12124 2876 14280 2904
rect 12124 2864 12130 2876
rect 14274 2864 14280 2876
rect 14332 2864 14338 2916
rect 10134 2836 10140 2848
rect 6886 2808 9996 2836
rect 10095 2808 10140 2836
rect 10134 2796 10140 2808
rect 10192 2796 10198 2848
rect 10318 2796 10324 2848
rect 10376 2836 10382 2848
rect 12529 2839 12587 2845
rect 12529 2836 12541 2839
rect 10376 2808 12541 2836
rect 10376 2796 10382 2808
rect 12529 2805 12541 2808
rect 12575 2805 12587 2839
rect 12529 2799 12587 2805
rect 368 2746 18308 2768
rect 368 2694 3204 2746
rect 3256 2694 3268 2746
rect 3320 2694 3332 2746
rect 3384 2694 3396 2746
rect 3448 2694 3460 2746
rect 3512 2694 9184 2746
rect 9236 2694 9248 2746
rect 9300 2694 9312 2746
rect 9364 2694 9376 2746
rect 9428 2694 9440 2746
rect 9492 2694 15164 2746
rect 15216 2694 15228 2746
rect 15280 2694 15292 2746
rect 15344 2694 15356 2746
rect 15408 2694 15420 2746
rect 15472 2694 18308 2746
rect 368 2672 18308 2694
rect 1118 2632 1124 2644
rect 1079 2604 1124 2632
rect 1118 2592 1124 2604
rect 1176 2592 1182 2644
rect 1673 2635 1731 2641
rect 1673 2601 1685 2635
rect 1719 2632 1731 2635
rect 3694 2632 3700 2644
rect 1719 2604 3700 2632
rect 1719 2601 1731 2604
rect 1673 2595 1731 2601
rect 3694 2592 3700 2604
rect 3752 2592 3758 2644
rect 3786 2592 3792 2644
rect 3844 2632 3850 2644
rect 3844 2604 16574 2632
rect 3844 2592 3850 2604
rect 3053 2567 3111 2573
rect 3053 2533 3065 2567
rect 3099 2564 3111 2567
rect 3418 2564 3424 2576
rect 3099 2536 3424 2564
rect 3099 2533 3111 2536
rect 3053 2527 3111 2533
rect 3418 2524 3424 2536
rect 3476 2524 3482 2576
rect 5534 2524 5540 2576
rect 5592 2564 5598 2576
rect 6273 2567 6331 2573
rect 6273 2564 6285 2567
rect 5592 2536 6285 2564
rect 5592 2524 5598 2536
rect 6273 2533 6285 2536
rect 6319 2533 6331 2567
rect 6730 2564 6736 2576
rect 6691 2536 6736 2564
rect 6273 2527 6331 2533
rect 6730 2524 6736 2536
rect 6788 2524 6794 2576
rect 7190 2524 7196 2576
rect 7248 2564 7254 2576
rect 7377 2567 7435 2573
rect 7377 2564 7389 2567
rect 7248 2536 7389 2564
rect 7248 2524 7254 2536
rect 7377 2533 7389 2536
rect 7423 2533 7435 2567
rect 8294 2564 8300 2576
rect 8255 2536 8300 2564
rect 7377 2527 7435 2533
rect 8294 2524 8300 2536
rect 8352 2524 8358 2576
rect 8846 2524 8852 2576
rect 8904 2564 8910 2576
rect 9585 2567 9643 2573
rect 9585 2564 9597 2567
rect 8904 2536 9597 2564
rect 8904 2524 8910 2536
rect 9585 2533 9597 2536
rect 9631 2533 9643 2567
rect 13354 2564 13360 2576
rect 13315 2536 13360 2564
rect 9585 2527 9643 2533
rect 13354 2524 13360 2536
rect 13412 2524 13418 2576
rect 14274 2564 14280 2576
rect 13832 2536 14280 2564
rect 2958 2496 2964 2508
rect 1780 2468 2964 2496
rect 750 2388 756 2440
rect 808 2428 814 2440
rect 937 2431 995 2437
rect 937 2428 949 2431
rect 808 2400 949 2428
rect 808 2388 814 2400
rect 937 2397 949 2400
rect 983 2397 995 2431
rect 1118 2428 1124 2440
rect 1079 2400 1124 2428
rect 937 2391 995 2397
rect 1118 2388 1124 2400
rect 1176 2388 1182 2440
rect 1780 2437 1808 2468
rect 2958 2456 2964 2468
rect 3016 2456 3022 2508
rect 4433 2499 4491 2505
rect 4433 2465 4445 2499
rect 4479 2496 4491 2499
rect 4985 2499 5043 2505
rect 4985 2496 4997 2499
rect 4479 2468 4997 2496
rect 4479 2465 4491 2468
rect 4433 2459 4491 2465
rect 4985 2465 4997 2468
rect 5031 2465 5043 2499
rect 11425 2499 11483 2505
rect 4985 2459 5043 2465
rect 7024 2468 7604 2496
rect 7024 2440 7052 2468
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2428 2559 2431
rect 3602 2428 3608 2440
rect 2547 2400 3608 2428
rect 2547 2397 2559 2400
rect 2501 2391 2559 2397
rect 3602 2388 3608 2400
rect 3660 2428 3666 2440
rect 4893 2431 4951 2437
rect 4893 2428 4905 2431
rect 3660 2400 4905 2428
rect 3660 2388 3666 2400
rect 4893 2397 4905 2400
rect 4939 2397 4951 2431
rect 5626 2428 5632 2440
rect 5587 2400 5632 2428
rect 4893 2391 4951 2397
rect 5626 2388 5632 2400
rect 5684 2388 5690 2440
rect 6733 2431 6791 2437
rect 6104 2400 6500 2428
rect 566 2320 572 2372
rect 624 2360 630 2372
rect 2317 2363 2375 2369
rect 624 2332 2268 2360
rect 624 2320 630 2332
rect 2240 2292 2268 2332
rect 2317 2329 2329 2363
rect 2363 2360 2375 2363
rect 4062 2360 4068 2372
rect 2363 2332 4068 2360
rect 2363 2329 2375 2332
rect 2317 2323 2375 2329
rect 4062 2320 4068 2332
rect 4120 2320 4126 2372
rect 4188 2363 4246 2369
rect 4188 2329 4200 2363
rect 4234 2360 4246 2363
rect 6104 2360 6132 2400
rect 6472 2360 6500 2400
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 6822 2428 6828 2440
rect 6779 2400 6828 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 6822 2388 6828 2400
rect 6880 2388 6886 2440
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2428 6975 2431
rect 7006 2428 7012 2440
rect 6963 2400 7012 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 7006 2388 7012 2400
rect 7064 2388 7070 2440
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7576 2437 7604 2468
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 11974 2496 11980 2508
rect 11471 2468 11980 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 11974 2456 11980 2468
rect 12032 2456 12038 2508
rect 12526 2456 12532 2508
rect 12584 2496 12590 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12584 2468 12633 2496
rect 12584 2456 12590 2468
rect 12621 2465 12633 2468
rect 12667 2496 12679 2499
rect 12667 2468 13400 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 7156 2400 7389 2428
rect 7156 2388 7162 2400
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2397 7619 2431
rect 8386 2428 8392 2440
rect 8347 2400 8392 2428
rect 7561 2391 7619 2397
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 10134 2428 10140 2440
rect 9171 2400 10140 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 10229 2431 10287 2437
rect 10229 2397 10241 2431
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 10244 2360 10272 2391
rect 10686 2388 10692 2440
rect 10744 2428 10750 2440
rect 13372 2437 13400 2468
rect 10873 2431 10931 2437
rect 10744 2422 10824 2428
rect 10873 2422 10885 2431
rect 10744 2400 10885 2422
rect 10744 2388 10750 2400
rect 10796 2397 10885 2400
rect 10919 2397 10931 2431
rect 10796 2394 10931 2397
rect 10873 2391 10931 2394
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 13357 2431 13415 2437
rect 12115 2400 13308 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 11606 2360 11612 2372
rect 4234 2332 6132 2360
rect 6196 2332 6408 2360
rect 6472 2332 7604 2360
rect 4234 2329 4246 2332
rect 4188 2323 4246 2329
rect 6196 2292 6224 2332
rect 2240 2264 6224 2292
rect 6380 2292 6408 2332
rect 7374 2292 7380 2304
rect 6380 2264 7380 2292
rect 7374 2252 7380 2264
rect 7432 2252 7438 2304
rect 7576 2292 7604 2332
rect 9692 2332 11612 2360
rect 8941 2295 8999 2301
rect 8941 2292 8953 2295
rect 7576 2264 8953 2292
rect 8941 2261 8953 2264
rect 8987 2292 8999 2295
rect 9692 2292 9720 2332
rect 11606 2320 11612 2332
rect 11664 2360 11670 2372
rect 12084 2360 12112 2391
rect 11664 2332 12112 2360
rect 11664 2320 11670 2332
rect 8987 2264 9720 2292
rect 13280 2292 13308 2400
rect 13357 2397 13369 2431
rect 13403 2397 13415 2431
rect 13357 2391 13415 2397
rect 13541 2431 13599 2437
rect 13541 2397 13553 2431
rect 13587 2422 13599 2431
rect 13832 2428 13860 2536
rect 14274 2524 14280 2536
rect 14332 2524 14338 2576
rect 15381 2567 15439 2573
rect 15381 2533 15393 2567
rect 15427 2564 15439 2567
rect 16298 2564 16304 2576
rect 15427 2536 16304 2564
rect 15427 2533 15439 2536
rect 15381 2527 15439 2533
rect 16298 2524 16304 2536
rect 16356 2524 16362 2576
rect 14458 2496 14464 2508
rect 13648 2422 13860 2428
rect 13587 2400 13860 2422
rect 13924 2468 14464 2496
rect 13587 2397 13676 2400
rect 13541 2394 13676 2397
rect 13541 2391 13599 2394
rect 13372 2360 13400 2391
rect 13924 2360 13952 2468
rect 14458 2456 14464 2468
rect 14516 2496 14522 2508
rect 16390 2496 16396 2508
rect 14516 2468 16396 2496
rect 14516 2456 14522 2468
rect 14001 2431 14059 2437
rect 14001 2397 14013 2431
rect 14047 2397 14059 2431
rect 14001 2391 14059 2397
rect 13372 2332 13952 2360
rect 14016 2292 14044 2391
rect 14182 2388 14188 2440
rect 14240 2428 14246 2440
rect 15396 2437 15424 2468
rect 16390 2456 16396 2468
rect 16448 2456 16454 2508
rect 15197 2431 15255 2437
rect 14240 2400 14285 2428
rect 14240 2388 14246 2400
rect 15197 2397 15209 2431
rect 15243 2397 15255 2431
rect 15197 2391 15255 2397
rect 15381 2431 15439 2437
rect 15381 2397 15393 2431
rect 15427 2397 15439 2431
rect 15381 2391 15439 2397
rect 14090 2320 14096 2372
rect 14148 2360 14154 2372
rect 14148 2332 14193 2360
rect 14148 2320 14154 2332
rect 14274 2320 14280 2372
rect 14332 2360 14338 2372
rect 15212 2360 15240 2391
rect 15930 2388 15936 2440
rect 15988 2428 15994 2440
rect 16025 2431 16083 2437
rect 16025 2428 16037 2431
rect 15988 2400 16037 2428
rect 15988 2388 15994 2400
rect 16025 2397 16037 2400
rect 16071 2397 16083 2431
rect 16025 2391 16083 2397
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16209 2431 16267 2437
rect 16209 2428 16221 2431
rect 16172 2400 16221 2428
rect 16172 2388 16178 2400
rect 16209 2397 16221 2400
rect 16255 2397 16267 2431
rect 16546 2428 16574 2604
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16546 2400 16865 2428
rect 16209 2391 16267 2397
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 16482 2360 16488 2372
rect 14332 2332 16488 2360
rect 14332 2320 14338 2332
rect 16482 2320 16488 2332
rect 16540 2320 16546 2372
rect 14826 2292 14832 2304
rect 13280 2264 14832 2292
rect 8987 2261 8999 2264
rect 8941 2255 8999 2261
rect 14826 2252 14832 2264
rect 14884 2252 14890 2304
rect 15010 2252 15016 2304
rect 15068 2292 15074 2304
rect 16117 2295 16175 2301
rect 16117 2292 16129 2295
rect 15068 2264 16129 2292
rect 15068 2252 15074 2264
rect 16117 2261 16129 2264
rect 16163 2261 16175 2295
rect 16117 2255 16175 2261
rect 16206 2252 16212 2304
rect 16264 2292 16270 2304
rect 16669 2295 16727 2301
rect 16669 2292 16681 2295
rect 16264 2264 16681 2292
rect 16264 2252 16270 2264
rect 16669 2261 16681 2264
rect 16715 2261 16727 2295
rect 16669 2255 16727 2261
rect 368 2202 18308 2224
rect 368 2150 6194 2202
rect 6246 2150 6258 2202
rect 6310 2150 6322 2202
rect 6374 2150 6386 2202
rect 6438 2150 6450 2202
rect 6502 2150 12174 2202
rect 12226 2150 12238 2202
rect 12290 2150 12302 2202
rect 12354 2150 12366 2202
rect 12418 2150 12430 2202
rect 12482 2150 18308 2202
rect 368 2128 18308 2150
rect 3418 2048 3424 2100
rect 3476 2088 3482 2100
rect 5626 2088 5632 2100
rect 3476 2060 5632 2088
rect 3476 2048 3482 2060
rect 5626 2048 5632 2060
rect 5684 2048 5690 2100
rect 7374 2048 7380 2100
rect 7432 2088 7438 2100
rect 16206 2088 16212 2100
rect 7432 2060 16212 2088
rect 7432 2048 7438 2060
rect 16206 2048 16212 2060
rect 16264 2048 16270 2100
rect 5350 1980 5356 2032
rect 5408 2020 5414 2032
rect 7190 2020 7196 2032
rect 5408 1992 7196 2020
rect 5408 1980 5414 1992
rect 7190 1980 7196 1992
rect 7248 1980 7254 2032
rect 1118 1912 1124 1964
rect 1176 1952 1182 1964
rect 6914 1952 6920 1964
rect 1176 1924 6920 1952
rect 1176 1912 1182 1924
rect 6914 1912 6920 1924
rect 6972 1912 6978 1964
<< via1 >>
rect 10784 5584 10836 5636
rect 14096 5516 14148 5568
rect 16120 5516 16172 5568
rect 16672 5516 16724 5568
rect 6194 5414 6246 5466
rect 6258 5414 6310 5466
rect 6322 5414 6374 5466
rect 6386 5414 6438 5466
rect 6450 5414 6502 5466
rect 12174 5414 12226 5466
rect 12238 5414 12290 5466
rect 12302 5414 12354 5466
rect 12366 5414 12418 5466
rect 12430 5414 12482 5466
rect 3884 5312 3936 5364
rect 4068 5355 4120 5364
rect 4068 5321 4077 5355
rect 4077 5321 4111 5355
rect 4111 5321 4120 5355
rect 4068 5312 4120 5321
rect 4896 5355 4948 5364
rect 4896 5321 4905 5355
rect 4905 5321 4939 5355
rect 4939 5321 4948 5355
rect 4896 5312 4948 5321
rect 8484 5355 8536 5364
rect 8484 5321 8493 5355
rect 8493 5321 8527 5355
rect 8527 5321 8536 5355
rect 8484 5312 8536 5321
rect 9404 5355 9456 5364
rect 9404 5321 9413 5355
rect 9413 5321 9447 5355
rect 9447 5321 9456 5355
rect 9404 5312 9456 5321
rect 15200 5312 15252 5364
rect 5632 5244 5684 5296
rect 8208 5244 8260 5296
rect 12440 5244 12492 5296
rect 15016 5244 15068 5296
rect 3056 5219 3108 5228
rect 3056 5185 3065 5219
rect 3065 5185 3099 5219
rect 3099 5185 3108 5219
rect 3056 5176 3108 5185
rect 2964 5108 3016 5160
rect 3976 5176 4028 5228
rect 8668 5219 8720 5228
rect 8668 5185 8677 5219
rect 8677 5185 8711 5219
rect 8711 5185 8720 5219
rect 8668 5176 8720 5185
rect 9036 5176 9088 5228
rect 10784 5219 10836 5228
rect 10784 5185 10793 5219
rect 10793 5185 10827 5219
rect 10827 5185 10836 5219
rect 10784 5176 10836 5185
rect 15752 5176 15804 5228
rect 15936 5219 15988 5228
rect 15936 5185 15945 5219
rect 15945 5185 15979 5219
rect 15979 5185 15988 5219
rect 15936 5176 15988 5185
rect 16672 5219 16724 5228
rect 16672 5185 16681 5219
rect 16681 5185 16715 5219
rect 16715 5185 16724 5219
rect 16672 5176 16724 5185
rect 17316 5176 17368 5228
rect 5540 5108 5592 5160
rect 5724 5151 5776 5160
rect 5724 5117 5733 5151
rect 5733 5117 5767 5151
rect 5767 5117 5776 5151
rect 5724 5108 5776 5117
rect 6460 5108 6512 5160
rect 12624 5108 12676 5160
rect 3792 4972 3844 5024
rect 3884 4972 3936 5024
rect 6736 4972 6788 5024
rect 7472 5015 7524 5024
rect 7472 4981 7481 5015
rect 7481 4981 7515 5015
rect 7515 4981 7524 5015
rect 7472 4972 7524 4981
rect 11152 4972 11204 5024
rect 12532 5015 12584 5024
rect 12532 4981 12541 5015
rect 12541 4981 12575 5015
rect 12575 4981 12584 5015
rect 12532 4972 12584 4981
rect 17316 5040 17368 5092
rect 16120 5015 16172 5024
rect 16120 4981 16129 5015
rect 16129 4981 16163 5015
rect 16163 4981 16172 5015
rect 16120 4972 16172 4981
rect 3204 4870 3256 4922
rect 3268 4870 3320 4922
rect 3332 4870 3384 4922
rect 3396 4870 3448 4922
rect 3460 4870 3512 4922
rect 9184 4870 9236 4922
rect 9248 4870 9300 4922
rect 9312 4870 9364 4922
rect 9376 4870 9428 4922
rect 9440 4870 9492 4922
rect 15164 4870 15216 4922
rect 15228 4870 15280 4922
rect 15292 4870 15344 4922
rect 15356 4870 15408 4922
rect 15420 4870 15472 4922
rect 1400 4811 1452 4820
rect 1400 4777 1409 4811
rect 1409 4777 1443 4811
rect 1443 4777 1452 4811
rect 1400 4768 1452 4777
rect 2780 4768 2832 4820
rect 6460 4811 6512 4820
rect 6460 4777 6469 4811
rect 6469 4777 6503 4811
rect 6503 4777 6512 4811
rect 6460 4768 6512 4777
rect 7196 4768 7248 4820
rect 8208 4811 8260 4820
rect 8208 4777 8217 4811
rect 8217 4777 8251 4811
rect 8251 4777 8260 4811
rect 8208 4768 8260 4777
rect 10784 4768 10836 4820
rect 11612 4768 11664 4820
rect 12624 4768 12676 4820
rect 16028 4768 16080 4820
rect 17408 4811 17460 4820
rect 17408 4777 17417 4811
rect 17417 4777 17451 4811
rect 17451 4777 17460 4811
rect 17408 4768 17460 4777
rect 3976 4675 4028 4684
rect 3976 4641 3985 4675
rect 3985 4641 4019 4675
rect 4019 4641 4028 4675
rect 3976 4632 4028 4641
rect 6000 4632 6052 4684
rect 6920 4632 6972 4684
rect 1216 4607 1268 4616
rect 1216 4573 1225 4607
rect 1225 4573 1259 4607
rect 1259 4573 1268 4607
rect 1216 4564 1268 4573
rect 2964 4564 3016 4616
rect 5356 4564 5408 4616
rect 7472 4564 7524 4616
rect 8116 4564 8168 4616
rect 1492 4496 1544 4548
rect 7380 4496 7432 4548
rect 9128 4564 9180 4616
rect 11152 4675 11204 4684
rect 11152 4641 11161 4675
rect 11161 4641 11195 4675
rect 11195 4641 11204 4675
rect 11152 4632 11204 4641
rect 12532 4632 12584 4684
rect 5724 4471 5776 4480
rect 5724 4437 5733 4471
rect 5733 4437 5767 4471
rect 5767 4437 5776 4471
rect 5724 4428 5776 4437
rect 12624 4564 12676 4616
rect 14188 4564 14240 4616
rect 15200 4632 15252 4684
rect 15752 4632 15804 4684
rect 13176 4496 13228 4548
rect 15660 4564 15712 4616
rect 11060 4428 11112 4480
rect 6194 4326 6246 4378
rect 6258 4326 6310 4378
rect 6322 4326 6374 4378
rect 6386 4326 6438 4378
rect 6450 4326 6502 4378
rect 12174 4326 12226 4378
rect 12238 4326 12290 4378
rect 12302 4326 12354 4378
rect 12366 4326 12418 4378
rect 12430 4326 12482 4378
rect 1124 4224 1176 4276
rect 2964 4267 3016 4276
rect 1492 4199 1544 4208
rect 1492 4165 1501 4199
rect 1501 4165 1535 4199
rect 1535 4165 1544 4199
rect 1492 4156 1544 4165
rect 2964 4233 2973 4267
rect 2973 4233 3007 4267
rect 3007 4233 3016 4267
rect 2964 4224 3016 4233
rect 9128 4224 9180 4276
rect 11244 4224 11296 4276
rect 4160 4156 4212 4208
rect 14096 4224 14148 4276
rect 14188 4224 14240 4276
rect 15936 4224 15988 4276
rect 13176 4199 13228 4208
rect 13176 4165 13185 4199
rect 13185 4165 13219 4199
rect 13219 4165 13228 4199
rect 13176 4156 13228 4165
rect 4988 4131 5040 4140
rect 4988 4097 4997 4131
rect 4997 4097 5031 4131
rect 5031 4097 5040 4131
rect 4988 4088 5040 4097
rect 7472 4131 7524 4140
rect 7472 4097 7481 4131
rect 7481 4097 7515 4131
rect 7515 4097 7524 4131
rect 7472 4088 7524 4097
rect 10324 4088 10376 4140
rect 11060 4131 11112 4140
rect 11060 4097 11069 4131
rect 11069 4097 11103 4131
rect 11103 4097 11112 4131
rect 11060 4088 11112 4097
rect 11612 4131 11664 4140
rect 11612 4097 11621 4131
rect 11621 4097 11655 4131
rect 11655 4097 11664 4131
rect 11612 4088 11664 4097
rect 15200 4131 15252 4140
rect 1216 4063 1268 4072
rect 1216 4029 1225 4063
rect 1225 4029 1259 4063
rect 1259 4029 1268 4063
rect 1216 4020 1268 4029
rect 756 3952 808 4004
rect 7012 4020 7064 4072
rect 7380 4020 7432 4072
rect 8300 4020 8352 4072
rect 11244 4020 11296 4072
rect 12808 4020 12860 4072
rect 15200 4097 15209 4131
rect 15209 4097 15243 4131
rect 15243 4097 15252 4131
rect 15200 4088 15252 4097
rect 15752 4088 15804 4140
rect 15936 4131 15988 4140
rect 15936 4097 15945 4131
rect 15945 4097 15979 4131
rect 15979 4097 15988 4131
rect 15936 4088 15988 4097
rect 16120 4131 16172 4140
rect 16120 4097 16129 4131
rect 16129 4097 16163 4131
rect 16163 4097 16172 4131
rect 16120 4088 16172 4097
rect 16580 4131 16632 4140
rect 16580 4097 16589 4131
rect 16589 4097 16623 4131
rect 16623 4097 16632 4131
rect 16580 4088 16632 4097
rect 17316 4131 17368 4140
rect 13544 4020 13596 4072
rect 17316 4097 17325 4131
rect 17325 4097 17359 4131
rect 17359 4097 17368 4131
rect 17316 4088 17368 4097
rect 2964 3952 3016 4004
rect 6092 3952 6144 4004
rect 10508 3952 10560 4004
rect 12716 3952 12768 4004
rect 15660 3952 15712 4004
rect 18236 3952 18288 4004
rect 8208 3884 8260 3936
rect 12348 3884 12400 3936
rect 15936 3884 15988 3936
rect 16488 3884 16540 3936
rect 3204 3782 3256 3834
rect 3268 3782 3320 3834
rect 3332 3782 3384 3834
rect 3396 3782 3448 3834
rect 3460 3782 3512 3834
rect 9184 3782 9236 3834
rect 9248 3782 9300 3834
rect 9312 3782 9364 3834
rect 9376 3782 9428 3834
rect 9440 3782 9492 3834
rect 15164 3782 15216 3834
rect 15228 3782 15280 3834
rect 15292 3782 15344 3834
rect 15356 3782 15408 3834
rect 15420 3782 15472 3834
rect 8300 3723 8352 3732
rect 1308 3519 1360 3528
rect 1308 3485 1317 3519
rect 1317 3485 1351 3519
rect 1351 3485 1360 3519
rect 1308 3476 1360 3485
rect 8300 3689 8309 3723
rect 8309 3689 8343 3723
rect 8343 3689 8352 3723
rect 8300 3680 8352 3689
rect 12532 3680 12584 3732
rect 12808 3680 12860 3732
rect 16028 3680 16080 3732
rect 8852 3612 8904 3664
rect 10692 3612 10744 3664
rect 14188 3544 14240 3596
rect 15108 3544 15160 3596
rect 8208 3476 8260 3528
rect 8668 3476 8720 3528
rect 10324 3519 10376 3528
rect 10324 3485 10333 3519
rect 10333 3485 10367 3519
rect 10367 3485 10376 3519
rect 10324 3476 10376 3485
rect 10692 3476 10744 3528
rect 11060 3476 11112 3528
rect 11980 3519 12032 3528
rect 1032 3408 1084 3460
rect 3424 3451 3476 3460
rect 3424 3417 3433 3451
rect 3433 3417 3467 3451
rect 3467 3417 3476 3451
rect 3424 3408 3476 3417
rect 11152 3408 11204 3460
rect 11244 3451 11296 3460
rect 11244 3417 11253 3451
rect 11253 3417 11287 3451
rect 11287 3417 11296 3451
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 12532 3476 12584 3528
rect 12808 3519 12860 3528
rect 11244 3408 11296 3417
rect 12348 3408 12400 3460
rect 12808 3485 12817 3519
rect 12817 3485 12851 3519
rect 12851 3485 12860 3519
rect 12808 3476 12860 3485
rect 13636 3451 13688 3460
rect 13636 3417 13645 3451
rect 13645 3417 13679 3451
rect 13679 3417 13688 3451
rect 13636 3408 13688 3417
rect 14372 3408 14424 3460
rect 2872 3340 2924 3392
rect 4160 3340 4212 3392
rect 5908 3383 5960 3392
rect 5908 3349 5917 3383
rect 5917 3349 5951 3383
rect 5951 3349 5960 3383
rect 5908 3340 5960 3349
rect 11060 3340 11112 3392
rect 12072 3383 12124 3392
rect 12072 3349 12081 3383
rect 12081 3349 12115 3383
rect 12115 3349 12124 3383
rect 12072 3340 12124 3349
rect 13728 3340 13780 3392
rect 15844 3451 15896 3460
rect 15844 3417 15853 3451
rect 15853 3417 15887 3451
rect 15887 3417 15896 3451
rect 15844 3408 15896 3417
rect 16304 3408 16356 3460
rect 16120 3340 16172 3392
rect 6194 3238 6246 3290
rect 6258 3238 6310 3290
rect 6322 3238 6374 3290
rect 6386 3238 6438 3290
rect 6450 3238 6502 3290
rect 12174 3238 12226 3290
rect 12238 3238 12290 3290
rect 12302 3238 12354 3290
rect 12366 3238 12418 3290
rect 12430 3238 12482 3290
rect 1308 3136 1360 3188
rect 5540 3136 5592 3188
rect 5632 3136 5684 3188
rect 5908 3136 5960 3188
rect 2872 3111 2924 3120
rect 2872 3077 2881 3111
rect 2881 3077 2915 3111
rect 2915 3077 2924 3111
rect 2872 3068 2924 3077
rect 756 3043 808 3052
rect 756 3009 765 3043
rect 765 3009 799 3043
rect 799 3009 808 3043
rect 756 3000 808 3009
rect 1032 3000 1084 3052
rect 3700 3000 3752 3052
rect 5540 3000 5592 3052
rect 6000 3068 6052 3120
rect 5724 3000 5776 3052
rect 8668 3136 8720 3188
rect 12072 3136 12124 3188
rect 13636 3179 13688 3188
rect 13636 3145 13645 3179
rect 13645 3145 13679 3179
rect 13679 3145 13688 3179
rect 13636 3136 13688 3145
rect 14372 3179 14424 3188
rect 14372 3145 14381 3179
rect 14381 3145 14415 3179
rect 14415 3145 14424 3179
rect 14372 3136 14424 3145
rect 15844 3136 15896 3188
rect 17500 3179 17552 3188
rect 17500 3145 17509 3179
rect 17509 3145 17543 3179
rect 17543 3145 17552 3179
rect 17500 3136 17552 3145
rect 11060 3111 11112 3120
rect 11060 3077 11069 3111
rect 11069 3077 11103 3111
rect 11103 3077 11112 3111
rect 11060 3068 11112 3077
rect 13360 3068 13412 3120
rect 13544 3068 13596 3120
rect 9588 3000 9640 3052
rect 12624 3000 12676 3052
rect 13728 3000 13780 3052
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 14464 3043 14516 3052
rect 14464 3009 14473 3043
rect 14473 3009 14507 3043
rect 14507 3009 14516 3043
rect 14464 3000 14516 3009
rect 14832 3000 14884 3052
rect 15108 3043 15160 3052
rect 15108 3009 15117 3043
rect 15117 3009 15151 3043
rect 15151 3009 15160 3043
rect 15108 3000 15160 3009
rect 16120 3068 16172 3120
rect 16396 3068 16448 3120
rect 16488 3000 16540 3052
rect 3608 2864 3660 2916
rect 4988 2907 5040 2916
rect 4988 2873 4997 2907
rect 4997 2873 5031 2907
rect 5031 2873 5040 2907
rect 8392 2932 8444 2984
rect 9036 2932 9088 2984
rect 11152 2932 11204 2984
rect 4988 2864 5040 2873
rect 8300 2864 8352 2916
rect 10692 2864 10744 2916
rect 12072 2864 12124 2916
rect 14280 2864 14332 2916
rect 10140 2839 10192 2848
rect 10140 2805 10149 2839
rect 10149 2805 10183 2839
rect 10183 2805 10192 2839
rect 10140 2796 10192 2805
rect 10324 2796 10376 2848
rect 3204 2694 3256 2746
rect 3268 2694 3320 2746
rect 3332 2694 3384 2746
rect 3396 2694 3448 2746
rect 3460 2694 3512 2746
rect 9184 2694 9236 2746
rect 9248 2694 9300 2746
rect 9312 2694 9364 2746
rect 9376 2694 9428 2746
rect 9440 2694 9492 2746
rect 15164 2694 15216 2746
rect 15228 2694 15280 2746
rect 15292 2694 15344 2746
rect 15356 2694 15408 2746
rect 15420 2694 15472 2746
rect 1124 2635 1176 2644
rect 1124 2601 1133 2635
rect 1133 2601 1167 2635
rect 1167 2601 1176 2635
rect 1124 2592 1176 2601
rect 3700 2592 3752 2644
rect 3792 2592 3844 2644
rect 3424 2524 3476 2576
rect 5540 2524 5592 2576
rect 6736 2567 6788 2576
rect 6736 2533 6745 2567
rect 6745 2533 6779 2567
rect 6779 2533 6788 2567
rect 6736 2524 6788 2533
rect 7196 2524 7248 2576
rect 8300 2567 8352 2576
rect 8300 2533 8309 2567
rect 8309 2533 8343 2567
rect 8343 2533 8352 2567
rect 8300 2524 8352 2533
rect 8852 2524 8904 2576
rect 13360 2567 13412 2576
rect 13360 2533 13369 2567
rect 13369 2533 13403 2567
rect 13403 2533 13412 2567
rect 13360 2524 13412 2533
rect 756 2388 808 2440
rect 1124 2431 1176 2440
rect 1124 2397 1133 2431
rect 1133 2397 1167 2431
rect 1167 2397 1176 2431
rect 1124 2388 1176 2397
rect 2964 2456 3016 2508
rect 3608 2388 3660 2440
rect 5632 2431 5684 2440
rect 5632 2397 5641 2431
rect 5641 2397 5675 2431
rect 5675 2397 5684 2431
rect 5632 2388 5684 2397
rect 572 2320 624 2372
rect 4068 2320 4120 2372
rect 6828 2388 6880 2440
rect 7012 2388 7064 2440
rect 7104 2388 7156 2440
rect 11980 2456 12032 2508
rect 12532 2456 12584 2508
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 10140 2388 10192 2440
rect 10692 2388 10744 2440
rect 7380 2252 7432 2304
rect 11612 2320 11664 2372
rect 14280 2524 14332 2576
rect 16304 2524 16356 2576
rect 14464 2456 14516 2508
rect 14188 2431 14240 2440
rect 14188 2397 14197 2431
rect 14197 2397 14231 2431
rect 14231 2397 14240 2431
rect 16396 2456 16448 2508
rect 14188 2388 14240 2397
rect 14096 2363 14148 2372
rect 14096 2329 14105 2363
rect 14105 2329 14139 2363
rect 14139 2329 14148 2363
rect 14096 2320 14148 2329
rect 14280 2320 14332 2372
rect 15936 2388 15988 2440
rect 16120 2388 16172 2440
rect 16488 2320 16540 2372
rect 14832 2252 14884 2304
rect 15016 2252 15068 2304
rect 16212 2252 16264 2304
rect 6194 2150 6246 2202
rect 6258 2150 6310 2202
rect 6322 2150 6374 2202
rect 6386 2150 6438 2202
rect 6450 2150 6502 2202
rect 12174 2150 12226 2202
rect 12238 2150 12290 2202
rect 12302 2150 12354 2202
rect 12366 2150 12418 2202
rect 12430 2150 12482 2202
rect 3424 2048 3476 2100
rect 5632 2048 5684 2100
rect 7380 2048 7432 2100
rect 16212 2048 16264 2100
rect 5356 1980 5408 2032
rect 7196 1980 7248 2032
rect 1124 1912 1176 1964
rect 6920 1912 6972 1964
<< metal2 >>
rect 570 5922 626 6322
rect 1674 6066 1730 6322
rect 1412 6038 1730 6066
rect 584 2378 612 5922
rect 1412 4826 1440 6038
rect 1674 5922 1730 6038
rect 2778 5922 2834 6322
rect 3882 6066 3938 6322
rect 4986 6066 5042 6322
rect 3882 6038 4108 6066
rect 3882 5922 3938 6038
rect 2792 4826 2820 5922
rect 4080 5370 4108 6038
rect 4908 6038 5042 6066
rect 4908 5370 4936 6038
rect 4986 5922 5042 6038
rect 6090 5922 6146 6322
rect 7194 5922 7250 6322
rect 8298 6066 8354 6322
rect 8298 6038 8524 6066
rect 8298 5922 8354 6038
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2976 4622 3004 5102
rect 1216 4616 1268 4622
rect 1216 4558 1268 4564
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 1124 4276 1176 4282
rect 1124 4218 1176 4224
rect 756 4004 808 4010
rect 756 3946 808 3952
rect 768 3058 796 3946
rect 1032 3460 1084 3466
rect 1032 3402 1084 3408
rect 1044 3058 1072 3402
rect 756 3052 808 3058
rect 756 2994 808 3000
rect 1032 3052 1084 3058
rect 1032 2994 1084 3000
rect 768 2446 796 2994
rect 1044 2530 1072 2994
rect 1136 2650 1164 4218
rect 1228 4078 1256 4558
rect 1492 4548 1544 4554
rect 1492 4490 1544 4496
rect 1504 4214 1532 4490
rect 2976 4282 3004 4558
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 1492 4208 1544 4214
rect 1492 4150 1544 4156
rect 1216 4072 1268 4078
rect 3068 4026 3096 5170
rect 3896 5030 3924 5306
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3204 4924 3512 4944
rect 3204 4922 3210 4924
rect 3266 4922 3290 4924
rect 3346 4922 3370 4924
rect 3426 4922 3450 4924
rect 3506 4922 3512 4924
rect 3266 4870 3268 4922
rect 3448 4870 3450 4922
rect 3204 4868 3210 4870
rect 3266 4868 3290 4870
rect 3346 4868 3370 4870
rect 3426 4868 3450 4870
rect 3506 4868 3512 4870
rect 3204 4848 3512 4868
rect 1216 4014 1268 4020
rect 1228 3890 1256 4014
rect 2976 4010 3096 4026
rect 2964 4004 3096 4010
rect 3016 3998 3096 4004
rect 2964 3946 3016 3952
rect 1228 3862 1348 3890
rect 1320 3534 1348 3862
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1320 3194 1348 3470
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 1308 3188 1360 3194
rect 1308 3130 1360 3136
rect 2884 3126 2912 3334
rect 2872 3120 2924 3126
rect 2872 3062 2924 3068
rect 1124 2644 1176 2650
rect 1124 2586 1176 2592
rect 1044 2502 1164 2530
rect 2976 2514 3004 3946
rect 3204 3836 3512 3856
rect 3204 3834 3210 3836
rect 3266 3834 3290 3836
rect 3346 3834 3370 3836
rect 3426 3834 3450 3836
rect 3506 3834 3512 3836
rect 3266 3782 3268 3834
rect 3448 3782 3450 3834
rect 3204 3780 3210 3782
rect 3266 3780 3290 3782
rect 3346 3780 3370 3782
rect 3426 3780 3450 3782
rect 3506 3780 3512 3782
rect 3204 3760 3512 3780
rect 3424 3460 3476 3466
rect 3424 3402 3476 3408
rect 3436 3233 3464 3402
rect 3422 3224 3478 3233
rect 3422 3159 3478 3168
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3608 2916 3660 2922
rect 3608 2858 3660 2864
rect 3204 2748 3512 2768
rect 3204 2746 3210 2748
rect 3266 2746 3290 2748
rect 3346 2746 3370 2748
rect 3426 2746 3450 2748
rect 3506 2746 3512 2748
rect 3266 2694 3268 2746
rect 3448 2694 3450 2746
rect 3204 2692 3210 2694
rect 3266 2692 3290 2694
rect 3346 2692 3370 2694
rect 3426 2692 3450 2694
rect 3506 2692 3512 2694
rect 3204 2672 3512 2692
rect 3424 2576 3476 2582
rect 3424 2518 3476 2524
rect 1136 2446 1164 2502
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 756 2440 808 2446
rect 756 2382 808 2388
rect 1124 2440 1176 2446
rect 1124 2382 1176 2388
rect 572 2372 624 2378
rect 572 2314 624 2320
rect 1136 1970 1164 2382
rect 3436 2106 3464 2518
rect 3620 2446 3648 2858
rect 3712 2650 3740 2994
rect 3804 2650 3832 4966
rect 3988 4690 4016 5170
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 3976 4684 4028 4690
rect 3976 4626 4028 4632
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 4172 3398 4200 4150
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 3700 2644 3752 2650
rect 3700 2586 3752 2592
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3608 2440 3660 2446
rect 4172 2394 4200 3334
rect 5000 2922 5028 4082
rect 4988 2916 5040 2922
rect 4988 2858 5040 2864
rect 3608 2382 3660 2388
rect 4080 2378 4200 2394
rect 4068 2372 4200 2378
rect 4120 2366 4200 2372
rect 4068 2314 4120 2320
rect 3424 2100 3476 2106
rect 3424 2042 3476 2048
rect 5368 2038 5396 4558
rect 5552 3194 5580 5102
rect 5644 3194 5672 5238
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5736 4486 5764 5102
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5736 3058 5764 4422
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 5920 3194 5948 3334
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 6012 3126 6040 4626
rect 6104 4010 6132 5922
rect 6194 5468 6502 5488
rect 6194 5466 6200 5468
rect 6256 5466 6280 5468
rect 6336 5466 6360 5468
rect 6416 5466 6440 5468
rect 6496 5466 6502 5468
rect 6256 5414 6258 5466
rect 6438 5414 6440 5466
rect 6194 5412 6200 5414
rect 6256 5412 6280 5414
rect 6336 5412 6360 5414
rect 6416 5412 6440 5414
rect 6496 5412 6502 5414
rect 6194 5392 6502 5412
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6472 4826 6500 5102
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6194 4380 6502 4400
rect 6194 4378 6200 4380
rect 6256 4378 6280 4380
rect 6336 4378 6360 4380
rect 6416 4378 6440 4380
rect 6496 4378 6502 4380
rect 6256 4326 6258 4378
rect 6438 4326 6440 4378
rect 6194 4324 6200 4326
rect 6256 4324 6280 4326
rect 6336 4324 6360 4326
rect 6416 4324 6440 4326
rect 6496 4324 6502 4326
rect 6194 4304 6502 4324
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 6194 3292 6502 3312
rect 6194 3290 6200 3292
rect 6256 3290 6280 3292
rect 6336 3290 6360 3292
rect 6416 3290 6440 3292
rect 6496 3290 6502 3292
rect 6256 3238 6258 3290
rect 6438 3238 6440 3290
rect 6194 3236 6200 3238
rect 6256 3236 6280 3238
rect 6336 3236 6360 3238
rect 6416 3236 6440 3238
rect 6496 3236 6502 3238
rect 6194 3216 6502 3236
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5552 2582 5580 2994
rect 6748 2582 6776 4966
rect 7208 4826 7236 5922
rect 8496 5370 8524 6038
rect 9402 5922 9458 6322
rect 10506 5922 10562 6322
rect 11610 5922 11666 6322
rect 12714 5922 12770 6322
rect 13818 6066 13874 6322
rect 13818 6038 14136 6066
rect 13818 5922 13874 6038
rect 9416 5370 9444 5922
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 6736 2576 6788 2582
rect 6736 2518 6788 2524
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 6828 2440 6880 2446
rect 6932 2394 6960 4626
rect 7484 4622 7512 4966
rect 8220 4826 8248 5238
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 8116 4616 8168 4622
rect 8168 4564 8248 4570
rect 8116 4558 8248 4564
rect 7380 4548 7432 4554
rect 7380 4490 7432 4496
rect 7392 4078 7420 4490
rect 7484 4146 7512 4558
rect 8128 4542 8248 4558
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7024 2446 7052 4014
rect 8220 3942 8248 4542
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8220 3534 8248 3878
rect 8312 3738 8340 4014
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8680 3534 8708 5170
rect 8852 3664 8904 3670
rect 8852 3606 8904 3612
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8680 3194 8708 3470
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8312 2582 8340 2858
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 6880 2388 6960 2394
rect 6828 2382 6960 2388
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 5644 2106 5672 2382
rect 6840 2366 6960 2382
rect 6932 2258 6960 2366
rect 7116 2258 7144 2382
rect 6932 2230 7144 2258
rect 6194 2204 6502 2224
rect 6194 2202 6200 2204
rect 6256 2202 6280 2204
rect 6336 2202 6360 2204
rect 6416 2202 6440 2204
rect 6496 2202 6502 2204
rect 6256 2150 6258 2202
rect 6438 2150 6440 2202
rect 6194 2148 6200 2150
rect 6256 2148 6280 2150
rect 6336 2148 6360 2150
rect 6416 2148 6440 2150
rect 6496 2148 6502 2150
rect 6194 2128 6502 2148
rect 5632 2100 5684 2106
rect 5632 2042 5684 2048
rect 5356 2032 5408 2038
rect 5356 1974 5408 1980
rect 6932 1970 6960 2230
rect 7208 2038 7236 2518
rect 8404 2446 8432 2926
rect 8864 2582 8892 3606
rect 9048 2990 9076 5170
rect 9184 4924 9492 4944
rect 9184 4922 9190 4924
rect 9246 4922 9270 4924
rect 9326 4922 9350 4924
rect 9406 4922 9430 4924
rect 9486 4922 9492 4924
rect 9246 4870 9248 4922
rect 9428 4870 9430 4922
rect 9184 4868 9190 4870
rect 9246 4868 9270 4870
rect 9326 4868 9350 4870
rect 9406 4868 9430 4870
rect 9486 4868 9492 4870
rect 9184 4848 9492 4868
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9140 4282 9168 4558
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 9184 3836 9492 3856
rect 9184 3834 9190 3836
rect 9246 3834 9270 3836
rect 9326 3834 9350 3836
rect 9406 3834 9430 3836
rect 9486 3834 9492 3836
rect 9246 3782 9248 3834
rect 9428 3782 9430 3834
rect 9184 3780 9190 3782
rect 9246 3780 9270 3782
rect 9326 3780 9350 3782
rect 9406 3780 9430 3782
rect 9486 3780 9492 3782
rect 9184 3760 9492 3780
rect 10336 3534 10364 4082
rect 10520 4010 10548 5922
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 10796 5234 10824 5578
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10796 4826 10824 5170
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 11164 4690 11192 4966
rect 11624 4826 11652 5922
rect 12174 5468 12482 5488
rect 12174 5466 12180 5468
rect 12236 5466 12260 5468
rect 12316 5466 12340 5468
rect 12396 5466 12420 5468
rect 12476 5466 12482 5468
rect 12236 5414 12238 5466
rect 12418 5414 12420 5466
rect 12174 5412 12180 5414
rect 12236 5412 12260 5414
rect 12316 5412 12340 5414
rect 12396 5412 12420 5414
rect 12476 5412 12482 5414
rect 12174 5392 12482 5412
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 12452 4570 12480 5238
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12544 4690 12572 4966
rect 12636 4826 12664 5102
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12624 4616 12676 4622
rect 12452 4542 12572 4570
rect 12624 4558 12676 4564
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11072 4146 11100 4422
rect 12174 4380 12482 4400
rect 12174 4378 12180 4380
rect 12236 4378 12260 4380
rect 12316 4378 12340 4380
rect 12396 4378 12420 4380
rect 12476 4378 12482 4380
rect 12236 4326 12238 4378
rect 12418 4326 12420 4378
rect 12174 4324 12180 4326
rect 12236 4324 12260 4326
rect 12316 4324 12340 4326
rect 12396 4324 12420 4326
rect 12476 4324 12482 4326
rect 12174 4304 12482 4324
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 10508 4004 10560 4010
rect 10508 3946 10560 3952
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10704 3534 10732 3606
rect 11072 3534 11100 4082
rect 11256 4078 11284 4218
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 9184 2748 9492 2768
rect 9184 2746 9190 2748
rect 9246 2746 9270 2748
rect 9326 2746 9350 2748
rect 9406 2746 9430 2748
rect 9486 2746 9492 2748
rect 9246 2694 9248 2746
rect 9428 2694 9430 2746
rect 9184 2692 9190 2694
rect 9246 2692 9270 2694
rect 9326 2692 9350 2694
rect 9406 2692 9430 2694
rect 9486 2692 9492 2694
rect 9184 2672 9492 2692
rect 8852 2576 8904 2582
rect 8852 2518 8904 2524
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 7380 2304 7432 2310
rect 7380 2246 7432 2252
rect 7392 2106 7420 2246
rect 7380 2100 7432 2106
rect 7380 2042 7432 2048
rect 7196 2032 7248 2038
rect 7196 1974 7248 1980
rect 1124 1964 1176 1970
rect 1124 1906 1176 1912
rect 6920 1964 6972 1970
rect 6920 1906 6972 1912
rect 9600 1578 9628 2994
rect 10336 2854 10364 3470
rect 10704 2922 10732 3470
rect 11256 3466 11284 4014
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 11072 3126 11100 3334
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 11164 2990 11192 3402
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 10692 2916 10744 2922
rect 10692 2858 10744 2864
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 10152 2446 10180 2790
rect 10704 2446 10732 2858
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 11624 2378 11652 4082
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11992 2938 12020 3470
rect 12360 3466 12388 3878
rect 12544 3738 12572 4542
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 12084 3194 12112 3334
rect 12174 3292 12482 3312
rect 12174 3290 12180 3292
rect 12236 3290 12260 3292
rect 12316 3290 12340 3292
rect 12396 3290 12420 3292
rect 12476 3290 12482 3292
rect 12236 3238 12238 3290
rect 12418 3238 12420 3290
rect 12174 3236 12180 3238
rect 12236 3236 12260 3238
rect 12316 3236 12340 3238
rect 12396 3236 12420 3238
rect 12476 3236 12482 3238
rect 12174 3216 12482 3236
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 11992 2922 12112 2938
rect 11992 2916 12124 2922
rect 11992 2910 12072 2916
rect 11992 2514 12020 2910
rect 12072 2858 12124 2864
rect 12544 2514 12572 3470
rect 12636 3058 12664 4558
rect 12728 4010 12756 5922
rect 14108 5574 14136 6038
rect 14922 5930 14978 6322
rect 15028 6038 15240 6066
rect 15028 5930 15056 6038
rect 14922 5922 15056 5930
rect 14936 5902 15056 5922
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 15212 5370 15240 6038
rect 16026 5922 16082 6322
rect 17130 6066 17186 6322
rect 17130 6038 17448 6066
rect 17130 5922 17186 6038
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15016 5296 15068 5302
rect 15016 5238 15068 5244
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 13188 4214 13216 4490
rect 14200 4282 14228 4558
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 13176 4208 13228 4214
rect 13176 4150 13228 4156
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 12716 4004 12768 4010
rect 12716 3946 12768 3952
rect 12820 3738 12848 4014
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12820 3534 12848 3674
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 13556 3126 13584 4014
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13648 3194 13676 3402
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 13544 3120 13596 3126
rect 13544 3062 13596 3068
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 13372 2582 13400 3062
rect 13740 3058 13768 3334
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13360 2576 13412 2582
rect 13360 2518 13412 2524
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 14108 2378 14136 4218
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 14200 2446 14228 3538
rect 14372 3460 14424 3466
rect 14372 3402 14424 3408
rect 14384 3194 14412 3402
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 14292 2922 14320 2994
rect 14280 2916 14332 2922
rect 14280 2858 14332 2864
rect 14292 2582 14320 2858
rect 14280 2576 14332 2582
rect 14280 2518 14332 2524
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14292 2378 14320 2518
rect 14476 2514 14504 2994
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 14096 2372 14148 2378
rect 14096 2314 14148 2320
rect 14280 2372 14332 2378
rect 14280 2314 14332 2320
rect 14844 2310 14872 2994
rect 15028 2310 15056 5238
rect 15752 5228 15804 5234
rect 15752 5170 15804 5176
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 15164 4924 15472 4944
rect 15164 4922 15170 4924
rect 15226 4922 15250 4924
rect 15306 4922 15330 4924
rect 15386 4922 15410 4924
rect 15466 4922 15472 4924
rect 15226 4870 15228 4922
rect 15408 4870 15410 4922
rect 15164 4868 15170 4870
rect 15226 4868 15250 4870
rect 15306 4868 15330 4870
rect 15386 4868 15410 4870
rect 15466 4868 15472 4870
rect 15164 4848 15472 4868
rect 15764 4690 15792 5170
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15212 4146 15240 4626
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15672 4010 15700 4558
rect 15764 4146 15792 4626
rect 15948 4282 15976 5170
rect 16040 4826 16068 5922
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16132 5030 16160 5510
rect 16684 5234 16712 5510
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17328 5098 17356 5170
rect 17316 5092 17368 5098
rect 17316 5034 17368 5040
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 17328 4146 17356 5034
rect 17420 4826 17448 6038
rect 18234 5922 18290 6322
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15936 4140 15988 4146
rect 16120 4140 16172 4146
rect 15936 4082 15988 4088
rect 16040 4100 16120 4128
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 15948 3942 15976 4082
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15164 3836 15472 3856
rect 15164 3834 15170 3836
rect 15226 3834 15250 3836
rect 15306 3834 15330 3836
rect 15386 3834 15410 3836
rect 15466 3834 15472 3836
rect 15226 3782 15228 3834
rect 15408 3782 15410 3834
rect 15164 3780 15170 3782
rect 15226 3780 15250 3782
rect 15306 3780 15330 3782
rect 15386 3780 15410 3782
rect 15466 3780 15472 3782
rect 15164 3760 15472 3780
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15120 3058 15148 3538
rect 15844 3460 15896 3466
rect 15844 3402 15896 3408
rect 15856 3194 15884 3402
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 15164 2748 15472 2768
rect 15164 2746 15170 2748
rect 15226 2746 15250 2748
rect 15306 2746 15330 2748
rect 15386 2746 15410 2748
rect 15466 2746 15472 2748
rect 15226 2694 15228 2746
rect 15408 2694 15410 2746
rect 15164 2692 15170 2694
rect 15226 2692 15250 2694
rect 15306 2692 15330 2694
rect 15386 2692 15410 2694
rect 15466 2692 15472 2694
rect 15164 2672 15472 2692
rect 15948 2446 15976 3878
rect 16040 3738 16068 4100
rect 16120 4082 16172 4088
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 16592 4026 16620 4082
rect 16500 3998 16620 4026
rect 18248 4010 18276 5922
rect 18236 4004 18288 4010
rect 16500 3942 16528 3998
rect 18236 3946 18288 3952
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 15936 2440 15988 2446
rect 16040 2428 16068 3674
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 16132 3126 16160 3334
rect 16120 3120 16172 3126
rect 16120 3062 16172 3068
rect 16316 2582 16344 3402
rect 17498 3224 17554 3233
rect 17498 3159 17500 3168
rect 17552 3159 17554 3168
rect 17500 3130 17552 3136
rect 16396 3120 16448 3126
rect 16396 3062 16448 3068
rect 16304 2576 16356 2582
rect 16304 2518 16356 2524
rect 16408 2514 16436 3062
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16396 2508 16448 2514
rect 16396 2450 16448 2456
rect 16120 2440 16172 2446
rect 16040 2400 16120 2428
rect 15936 2382 15988 2388
rect 16120 2382 16172 2388
rect 16500 2378 16528 2994
rect 16488 2372 16540 2378
rect 16488 2314 16540 2320
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 15016 2304 15068 2310
rect 15016 2246 15068 2252
rect 16212 2304 16264 2310
rect 16212 2246 16264 2252
rect 12174 2204 12482 2224
rect 12174 2202 12180 2204
rect 12236 2202 12260 2204
rect 12316 2202 12340 2204
rect 12396 2202 12420 2204
rect 12476 2202 12482 2204
rect 12236 2150 12238 2202
rect 12418 2150 12420 2202
rect 12174 2148 12180 2150
rect 12236 2148 12260 2150
rect 12316 2148 12340 2150
rect 12396 2148 12420 2150
rect 12476 2148 12482 2150
rect 12174 2128 12482 2148
rect 16224 2106 16252 2246
rect 16212 2100 16264 2106
rect 16212 2042 16264 2048
rect 9416 1550 9628 1578
rect 9416 400 9444 1550
rect 9402 0 9458 400
<< via2 >>
rect 3210 4922 3266 4924
rect 3290 4922 3346 4924
rect 3370 4922 3426 4924
rect 3450 4922 3506 4924
rect 3210 4870 3256 4922
rect 3256 4870 3266 4922
rect 3290 4870 3320 4922
rect 3320 4870 3332 4922
rect 3332 4870 3346 4922
rect 3370 4870 3384 4922
rect 3384 4870 3396 4922
rect 3396 4870 3426 4922
rect 3450 4870 3460 4922
rect 3460 4870 3506 4922
rect 3210 4868 3266 4870
rect 3290 4868 3346 4870
rect 3370 4868 3426 4870
rect 3450 4868 3506 4870
rect 3210 3834 3266 3836
rect 3290 3834 3346 3836
rect 3370 3834 3426 3836
rect 3450 3834 3506 3836
rect 3210 3782 3256 3834
rect 3256 3782 3266 3834
rect 3290 3782 3320 3834
rect 3320 3782 3332 3834
rect 3332 3782 3346 3834
rect 3370 3782 3384 3834
rect 3384 3782 3396 3834
rect 3396 3782 3426 3834
rect 3450 3782 3460 3834
rect 3460 3782 3506 3834
rect 3210 3780 3266 3782
rect 3290 3780 3346 3782
rect 3370 3780 3426 3782
rect 3450 3780 3506 3782
rect 3422 3168 3478 3224
rect 3210 2746 3266 2748
rect 3290 2746 3346 2748
rect 3370 2746 3426 2748
rect 3450 2746 3506 2748
rect 3210 2694 3256 2746
rect 3256 2694 3266 2746
rect 3290 2694 3320 2746
rect 3320 2694 3332 2746
rect 3332 2694 3346 2746
rect 3370 2694 3384 2746
rect 3384 2694 3396 2746
rect 3396 2694 3426 2746
rect 3450 2694 3460 2746
rect 3460 2694 3506 2746
rect 3210 2692 3266 2694
rect 3290 2692 3346 2694
rect 3370 2692 3426 2694
rect 3450 2692 3506 2694
rect 6200 5466 6256 5468
rect 6280 5466 6336 5468
rect 6360 5466 6416 5468
rect 6440 5466 6496 5468
rect 6200 5414 6246 5466
rect 6246 5414 6256 5466
rect 6280 5414 6310 5466
rect 6310 5414 6322 5466
rect 6322 5414 6336 5466
rect 6360 5414 6374 5466
rect 6374 5414 6386 5466
rect 6386 5414 6416 5466
rect 6440 5414 6450 5466
rect 6450 5414 6496 5466
rect 6200 5412 6256 5414
rect 6280 5412 6336 5414
rect 6360 5412 6416 5414
rect 6440 5412 6496 5414
rect 6200 4378 6256 4380
rect 6280 4378 6336 4380
rect 6360 4378 6416 4380
rect 6440 4378 6496 4380
rect 6200 4326 6246 4378
rect 6246 4326 6256 4378
rect 6280 4326 6310 4378
rect 6310 4326 6322 4378
rect 6322 4326 6336 4378
rect 6360 4326 6374 4378
rect 6374 4326 6386 4378
rect 6386 4326 6416 4378
rect 6440 4326 6450 4378
rect 6450 4326 6496 4378
rect 6200 4324 6256 4326
rect 6280 4324 6336 4326
rect 6360 4324 6416 4326
rect 6440 4324 6496 4326
rect 6200 3290 6256 3292
rect 6280 3290 6336 3292
rect 6360 3290 6416 3292
rect 6440 3290 6496 3292
rect 6200 3238 6246 3290
rect 6246 3238 6256 3290
rect 6280 3238 6310 3290
rect 6310 3238 6322 3290
rect 6322 3238 6336 3290
rect 6360 3238 6374 3290
rect 6374 3238 6386 3290
rect 6386 3238 6416 3290
rect 6440 3238 6450 3290
rect 6450 3238 6496 3290
rect 6200 3236 6256 3238
rect 6280 3236 6336 3238
rect 6360 3236 6416 3238
rect 6440 3236 6496 3238
rect 6200 2202 6256 2204
rect 6280 2202 6336 2204
rect 6360 2202 6416 2204
rect 6440 2202 6496 2204
rect 6200 2150 6246 2202
rect 6246 2150 6256 2202
rect 6280 2150 6310 2202
rect 6310 2150 6322 2202
rect 6322 2150 6336 2202
rect 6360 2150 6374 2202
rect 6374 2150 6386 2202
rect 6386 2150 6416 2202
rect 6440 2150 6450 2202
rect 6450 2150 6496 2202
rect 6200 2148 6256 2150
rect 6280 2148 6336 2150
rect 6360 2148 6416 2150
rect 6440 2148 6496 2150
rect 9190 4922 9246 4924
rect 9270 4922 9326 4924
rect 9350 4922 9406 4924
rect 9430 4922 9486 4924
rect 9190 4870 9236 4922
rect 9236 4870 9246 4922
rect 9270 4870 9300 4922
rect 9300 4870 9312 4922
rect 9312 4870 9326 4922
rect 9350 4870 9364 4922
rect 9364 4870 9376 4922
rect 9376 4870 9406 4922
rect 9430 4870 9440 4922
rect 9440 4870 9486 4922
rect 9190 4868 9246 4870
rect 9270 4868 9326 4870
rect 9350 4868 9406 4870
rect 9430 4868 9486 4870
rect 9190 3834 9246 3836
rect 9270 3834 9326 3836
rect 9350 3834 9406 3836
rect 9430 3834 9486 3836
rect 9190 3782 9236 3834
rect 9236 3782 9246 3834
rect 9270 3782 9300 3834
rect 9300 3782 9312 3834
rect 9312 3782 9326 3834
rect 9350 3782 9364 3834
rect 9364 3782 9376 3834
rect 9376 3782 9406 3834
rect 9430 3782 9440 3834
rect 9440 3782 9486 3834
rect 9190 3780 9246 3782
rect 9270 3780 9326 3782
rect 9350 3780 9406 3782
rect 9430 3780 9486 3782
rect 12180 5466 12236 5468
rect 12260 5466 12316 5468
rect 12340 5466 12396 5468
rect 12420 5466 12476 5468
rect 12180 5414 12226 5466
rect 12226 5414 12236 5466
rect 12260 5414 12290 5466
rect 12290 5414 12302 5466
rect 12302 5414 12316 5466
rect 12340 5414 12354 5466
rect 12354 5414 12366 5466
rect 12366 5414 12396 5466
rect 12420 5414 12430 5466
rect 12430 5414 12476 5466
rect 12180 5412 12236 5414
rect 12260 5412 12316 5414
rect 12340 5412 12396 5414
rect 12420 5412 12476 5414
rect 12180 4378 12236 4380
rect 12260 4378 12316 4380
rect 12340 4378 12396 4380
rect 12420 4378 12476 4380
rect 12180 4326 12226 4378
rect 12226 4326 12236 4378
rect 12260 4326 12290 4378
rect 12290 4326 12302 4378
rect 12302 4326 12316 4378
rect 12340 4326 12354 4378
rect 12354 4326 12366 4378
rect 12366 4326 12396 4378
rect 12420 4326 12430 4378
rect 12430 4326 12476 4378
rect 12180 4324 12236 4326
rect 12260 4324 12316 4326
rect 12340 4324 12396 4326
rect 12420 4324 12476 4326
rect 9190 2746 9246 2748
rect 9270 2746 9326 2748
rect 9350 2746 9406 2748
rect 9430 2746 9486 2748
rect 9190 2694 9236 2746
rect 9236 2694 9246 2746
rect 9270 2694 9300 2746
rect 9300 2694 9312 2746
rect 9312 2694 9326 2746
rect 9350 2694 9364 2746
rect 9364 2694 9376 2746
rect 9376 2694 9406 2746
rect 9430 2694 9440 2746
rect 9440 2694 9486 2746
rect 9190 2692 9246 2694
rect 9270 2692 9326 2694
rect 9350 2692 9406 2694
rect 9430 2692 9486 2694
rect 12180 3290 12236 3292
rect 12260 3290 12316 3292
rect 12340 3290 12396 3292
rect 12420 3290 12476 3292
rect 12180 3238 12226 3290
rect 12226 3238 12236 3290
rect 12260 3238 12290 3290
rect 12290 3238 12302 3290
rect 12302 3238 12316 3290
rect 12340 3238 12354 3290
rect 12354 3238 12366 3290
rect 12366 3238 12396 3290
rect 12420 3238 12430 3290
rect 12430 3238 12476 3290
rect 12180 3236 12236 3238
rect 12260 3236 12316 3238
rect 12340 3236 12396 3238
rect 12420 3236 12476 3238
rect 15170 4922 15226 4924
rect 15250 4922 15306 4924
rect 15330 4922 15386 4924
rect 15410 4922 15466 4924
rect 15170 4870 15216 4922
rect 15216 4870 15226 4922
rect 15250 4870 15280 4922
rect 15280 4870 15292 4922
rect 15292 4870 15306 4922
rect 15330 4870 15344 4922
rect 15344 4870 15356 4922
rect 15356 4870 15386 4922
rect 15410 4870 15420 4922
rect 15420 4870 15466 4922
rect 15170 4868 15226 4870
rect 15250 4868 15306 4870
rect 15330 4868 15386 4870
rect 15410 4868 15466 4870
rect 15170 3834 15226 3836
rect 15250 3834 15306 3836
rect 15330 3834 15386 3836
rect 15410 3834 15466 3836
rect 15170 3782 15216 3834
rect 15216 3782 15226 3834
rect 15250 3782 15280 3834
rect 15280 3782 15292 3834
rect 15292 3782 15306 3834
rect 15330 3782 15344 3834
rect 15344 3782 15356 3834
rect 15356 3782 15386 3834
rect 15410 3782 15420 3834
rect 15420 3782 15466 3834
rect 15170 3780 15226 3782
rect 15250 3780 15306 3782
rect 15330 3780 15386 3782
rect 15410 3780 15466 3782
rect 15170 2746 15226 2748
rect 15250 2746 15306 2748
rect 15330 2746 15386 2748
rect 15410 2746 15466 2748
rect 15170 2694 15216 2746
rect 15216 2694 15226 2746
rect 15250 2694 15280 2746
rect 15280 2694 15292 2746
rect 15292 2694 15306 2746
rect 15330 2694 15344 2746
rect 15344 2694 15356 2746
rect 15356 2694 15386 2746
rect 15410 2694 15420 2746
rect 15420 2694 15466 2746
rect 15170 2692 15226 2694
rect 15250 2692 15306 2694
rect 15330 2692 15386 2694
rect 15410 2692 15466 2694
rect 17498 3188 17554 3224
rect 17498 3168 17500 3188
rect 17500 3168 17552 3188
rect 17552 3168 17554 3188
rect 12180 2202 12236 2204
rect 12260 2202 12316 2204
rect 12340 2202 12396 2204
rect 12420 2202 12476 2204
rect 12180 2150 12226 2202
rect 12226 2150 12236 2202
rect 12260 2150 12290 2202
rect 12290 2150 12302 2202
rect 12302 2150 12316 2202
rect 12340 2150 12354 2202
rect 12354 2150 12366 2202
rect 12366 2150 12396 2202
rect 12420 2150 12430 2202
rect 12430 2150 12476 2202
rect 12180 2148 12236 2150
rect 12260 2148 12316 2150
rect 12340 2148 12396 2150
rect 12420 2148 12476 2150
<< metal3 >>
rect 6188 5472 6508 5473
rect 6188 5408 6196 5472
rect 6260 5408 6276 5472
rect 6340 5408 6356 5472
rect 6420 5408 6436 5472
rect 6500 5408 6508 5472
rect 6188 5407 6508 5408
rect 12168 5472 12488 5473
rect 12168 5408 12176 5472
rect 12240 5408 12256 5472
rect 12320 5408 12336 5472
rect 12400 5408 12416 5472
rect 12480 5408 12488 5472
rect 12168 5407 12488 5408
rect 3198 4928 3518 4929
rect 3198 4864 3206 4928
rect 3270 4864 3286 4928
rect 3350 4864 3366 4928
rect 3430 4864 3446 4928
rect 3510 4864 3518 4928
rect 3198 4863 3518 4864
rect 9178 4928 9498 4929
rect 9178 4864 9186 4928
rect 9250 4864 9266 4928
rect 9330 4864 9346 4928
rect 9410 4864 9426 4928
rect 9490 4864 9498 4928
rect 9178 4863 9498 4864
rect 15158 4928 15478 4929
rect 15158 4864 15166 4928
rect 15230 4864 15246 4928
rect 15310 4864 15326 4928
rect 15390 4864 15406 4928
rect 15470 4864 15478 4928
rect 15158 4863 15478 4864
rect 6188 4384 6508 4385
rect 6188 4320 6196 4384
rect 6260 4320 6276 4384
rect 6340 4320 6356 4384
rect 6420 4320 6436 4384
rect 6500 4320 6508 4384
rect 6188 4319 6508 4320
rect 12168 4384 12488 4385
rect 12168 4320 12176 4384
rect 12240 4320 12256 4384
rect 12320 4320 12336 4384
rect 12400 4320 12416 4384
rect 12480 4320 12488 4384
rect 12168 4319 12488 4320
rect 3198 3840 3518 3841
rect 3198 3776 3206 3840
rect 3270 3776 3286 3840
rect 3350 3776 3366 3840
rect 3430 3776 3446 3840
rect 3510 3776 3518 3840
rect 3198 3775 3518 3776
rect 9178 3840 9498 3841
rect 9178 3776 9186 3840
rect 9250 3776 9266 3840
rect 9330 3776 9346 3840
rect 9410 3776 9426 3840
rect 9490 3776 9498 3840
rect 9178 3775 9498 3776
rect 15158 3840 15478 3841
rect 15158 3776 15166 3840
rect 15230 3776 15246 3840
rect 15310 3776 15326 3840
rect 15390 3776 15406 3840
rect 15470 3776 15478 3840
rect 15158 3775 15478 3776
rect 6188 3296 6508 3297
rect 0 3226 400 3256
rect 6188 3232 6196 3296
rect 6260 3232 6276 3296
rect 6340 3232 6356 3296
rect 6420 3232 6436 3296
rect 6500 3232 6508 3296
rect 6188 3231 6508 3232
rect 12168 3296 12488 3297
rect 12168 3232 12176 3296
rect 12240 3232 12256 3296
rect 12320 3232 12336 3296
rect 12400 3232 12416 3296
rect 12480 3232 12488 3296
rect 12168 3231 12488 3232
rect 3417 3226 3483 3229
rect 0 3224 3483 3226
rect 0 3168 3422 3224
rect 3478 3168 3483 3224
rect 0 3166 3483 3168
rect 0 3136 400 3166
rect 3417 3163 3483 3166
rect 17493 3226 17559 3229
rect 18345 3226 18745 3256
rect 17493 3224 18745 3226
rect 17493 3168 17498 3224
rect 17554 3168 18745 3224
rect 17493 3166 18745 3168
rect 17493 3163 17559 3166
rect 18345 3136 18745 3166
rect 3198 2752 3518 2753
rect 3198 2688 3206 2752
rect 3270 2688 3286 2752
rect 3350 2688 3366 2752
rect 3430 2688 3446 2752
rect 3510 2688 3518 2752
rect 3198 2687 3518 2688
rect 9178 2752 9498 2753
rect 9178 2688 9186 2752
rect 9250 2688 9266 2752
rect 9330 2688 9346 2752
rect 9410 2688 9426 2752
rect 9490 2688 9498 2752
rect 9178 2687 9498 2688
rect 15158 2752 15478 2753
rect 15158 2688 15166 2752
rect 15230 2688 15246 2752
rect 15310 2688 15326 2752
rect 15390 2688 15406 2752
rect 15470 2688 15478 2752
rect 15158 2687 15478 2688
rect 6188 2208 6508 2209
rect 6188 2144 6196 2208
rect 6260 2144 6276 2208
rect 6340 2144 6356 2208
rect 6420 2144 6436 2208
rect 6500 2144 6508 2208
rect 6188 2143 6508 2144
rect 12168 2208 12488 2209
rect 12168 2144 12176 2208
rect 12240 2144 12256 2208
rect 12320 2144 12336 2208
rect 12400 2144 12416 2208
rect 12480 2144 12488 2208
rect 12168 2143 12488 2144
<< via3 >>
rect 6196 5468 6260 5472
rect 6196 5412 6200 5468
rect 6200 5412 6256 5468
rect 6256 5412 6260 5468
rect 6196 5408 6260 5412
rect 6276 5468 6340 5472
rect 6276 5412 6280 5468
rect 6280 5412 6336 5468
rect 6336 5412 6340 5468
rect 6276 5408 6340 5412
rect 6356 5468 6420 5472
rect 6356 5412 6360 5468
rect 6360 5412 6416 5468
rect 6416 5412 6420 5468
rect 6356 5408 6420 5412
rect 6436 5468 6500 5472
rect 6436 5412 6440 5468
rect 6440 5412 6496 5468
rect 6496 5412 6500 5468
rect 6436 5408 6500 5412
rect 12176 5468 12240 5472
rect 12176 5412 12180 5468
rect 12180 5412 12236 5468
rect 12236 5412 12240 5468
rect 12176 5408 12240 5412
rect 12256 5468 12320 5472
rect 12256 5412 12260 5468
rect 12260 5412 12316 5468
rect 12316 5412 12320 5468
rect 12256 5408 12320 5412
rect 12336 5468 12400 5472
rect 12336 5412 12340 5468
rect 12340 5412 12396 5468
rect 12396 5412 12400 5468
rect 12336 5408 12400 5412
rect 12416 5468 12480 5472
rect 12416 5412 12420 5468
rect 12420 5412 12476 5468
rect 12476 5412 12480 5468
rect 12416 5408 12480 5412
rect 3206 4924 3270 4928
rect 3206 4868 3210 4924
rect 3210 4868 3266 4924
rect 3266 4868 3270 4924
rect 3206 4864 3270 4868
rect 3286 4924 3350 4928
rect 3286 4868 3290 4924
rect 3290 4868 3346 4924
rect 3346 4868 3350 4924
rect 3286 4864 3350 4868
rect 3366 4924 3430 4928
rect 3366 4868 3370 4924
rect 3370 4868 3426 4924
rect 3426 4868 3430 4924
rect 3366 4864 3430 4868
rect 3446 4924 3510 4928
rect 3446 4868 3450 4924
rect 3450 4868 3506 4924
rect 3506 4868 3510 4924
rect 3446 4864 3510 4868
rect 9186 4924 9250 4928
rect 9186 4868 9190 4924
rect 9190 4868 9246 4924
rect 9246 4868 9250 4924
rect 9186 4864 9250 4868
rect 9266 4924 9330 4928
rect 9266 4868 9270 4924
rect 9270 4868 9326 4924
rect 9326 4868 9330 4924
rect 9266 4864 9330 4868
rect 9346 4924 9410 4928
rect 9346 4868 9350 4924
rect 9350 4868 9406 4924
rect 9406 4868 9410 4924
rect 9346 4864 9410 4868
rect 9426 4924 9490 4928
rect 9426 4868 9430 4924
rect 9430 4868 9486 4924
rect 9486 4868 9490 4924
rect 9426 4864 9490 4868
rect 15166 4924 15230 4928
rect 15166 4868 15170 4924
rect 15170 4868 15226 4924
rect 15226 4868 15230 4924
rect 15166 4864 15230 4868
rect 15246 4924 15310 4928
rect 15246 4868 15250 4924
rect 15250 4868 15306 4924
rect 15306 4868 15310 4924
rect 15246 4864 15310 4868
rect 15326 4924 15390 4928
rect 15326 4868 15330 4924
rect 15330 4868 15386 4924
rect 15386 4868 15390 4924
rect 15326 4864 15390 4868
rect 15406 4924 15470 4928
rect 15406 4868 15410 4924
rect 15410 4868 15466 4924
rect 15466 4868 15470 4924
rect 15406 4864 15470 4868
rect 6196 4380 6260 4384
rect 6196 4324 6200 4380
rect 6200 4324 6256 4380
rect 6256 4324 6260 4380
rect 6196 4320 6260 4324
rect 6276 4380 6340 4384
rect 6276 4324 6280 4380
rect 6280 4324 6336 4380
rect 6336 4324 6340 4380
rect 6276 4320 6340 4324
rect 6356 4380 6420 4384
rect 6356 4324 6360 4380
rect 6360 4324 6416 4380
rect 6416 4324 6420 4380
rect 6356 4320 6420 4324
rect 6436 4380 6500 4384
rect 6436 4324 6440 4380
rect 6440 4324 6496 4380
rect 6496 4324 6500 4380
rect 6436 4320 6500 4324
rect 12176 4380 12240 4384
rect 12176 4324 12180 4380
rect 12180 4324 12236 4380
rect 12236 4324 12240 4380
rect 12176 4320 12240 4324
rect 12256 4380 12320 4384
rect 12256 4324 12260 4380
rect 12260 4324 12316 4380
rect 12316 4324 12320 4380
rect 12256 4320 12320 4324
rect 12336 4380 12400 4384
rect 12336 4324 12340 4380
rect 12340 4324 12396 4380
rect 12396 4324 12400 4380
rect 12336 4320 12400 4324
rect 12416 4380 12480 4384
rect 12416 4324 12420 4380
rect 12420 4324 12476 4380
rect 12476 4324 12480 4380
rect 12416 4320 12480 4324
rect 3206 3836 3270 3840
rect 3206 3780 3210 3836
rect 3210 3780 3266 3836
rect 3266 3780 3270 3836
rect 3206 3776 3270 3780
rect 3286 3836 3350 3840
rect 3286 3780 3290 3836
rect 3290 3780 3346 3836
rect 3346 3780 3350 3836
rect 3286 3776 3350 3780
rect 3366 3836 3430 3840
rect 3366 3780 3370 3836
rect 3370 3780 3426 3836
rect 3426 3780 3430 3836
rect 3366 3776 3430 3780
rect 3446 3836 3510 3840
rect 3446 3780 3450 3836
rect 3450 3780 3506 3836
rect 3506 3780 3510 3836
rect 3446 3776 3510 3780
rect 9186 3836 9250 3840
rect 9186 3780 9190 3836
rect 9190 3780 9246 3836
rect 9246 3780 9250 3836
rect 9186 3776 9250 3780
rect 9266 3836 9330 3840
rect 9266 3780 9270 3836
rect 9270 3780 9326 3836
rect 9326 3780 9330 3836
rect 9266 3776 9330 3780
rect 9346 3836 9410 3840
rect 9346 3780 9350 3836
rect 9350 3780 9406 3836
rect 9406 3780 9410 3836
rect 9346 3776 9410 3780
rect 9426 3836 9490 3840
rect 9426 3780 9430 3836
rect 9430 3780 9486 3836
rect 9486 3780 9490 3836
rect 9426 3776 9490 3780
rect 15166 3836 15230 3840
rect 15166 3780 15170 3836
rect 15170 3780 15226 3836
rect 15226 3780 15230 3836
rect 15166 3776 15230 3780
rect 15246 3836 15310 3840
rect 15246 3780 15250 3836
rect 15250 3780 15306 3836
rect 15306 3780 15310 3836
rect 15246 3776 15310 3780
rect 15326 3836 15390 3840
rect 15326 3780 15330 3836
rect 15330 3780 15386 3836
rect 15386 3780 15390 3836
rect 15326 3776 15390 3780
rect 15406 3836 15470 3840
rect 15406 3780 15410 3836
rect 15410 3780 15466 3836
rect 15466 3780 15470 3836
rect 15406 3776 15470 3780
rect 6196 3292 6260 3296
rect 6196 3236 6200 3292
rect 6200 3236 6256 3292
rect 6256 3236 6260 3292
rect 6196 3232 6260 3236
rect 6276 3292 6340 3296
rect 6276 3236 6280 3292
rect 6280 3236 6336 3292
rect 6336 3236 6340 3292
rect 6276 3232 6340 3236
rect 6356 3292 6420 3296
rect 6356 3236 6360 3292
rect 6360 3236 6416 3292
rect 6416 3236 6420 3292
rect 6356 3232 6420 3236
rect 6436 3292 6500 3296
rect 6436 3236 6440 3292
rect 6440 3236 6496 3292
rect 6496 3236 6500 3292
rect 6436 3232 6500 3236
rect 12176 3292 12240 3296
rect 12176 3236 12180 3292
rect 12180 3236 12236 3292
rect 12236 3236 12240 3292
rect 12176 3232 12240 3236
rect 12256 3292 12320 3296
rect 12256 3236 12260 3292
rect 12260 3236 12316 3292
rect 12316 3236 12320 3292
rect 12256 3232 12320 3236
rect 12336 3292 12400 3296
rect 12336 3236 12340 3292
rect 12340 3236 12396 3292
rect 12396 3236 12400 3292
rect 12336 3232 12400 3236
rect 12416 3292 12480 3296
rect 12416 3236 12420 3292
rect 12420 3236 12476 3292
rect 12476 3236 12480 3292
rect 12416 3232 12480 3236
rect 3206 2748 3270 2752
rect 3206 2692 3210 2748
rect 3210 2692 3266 2748
rect 3266 2692 3270 2748
rect 3206 2688 3270 2692
rect 3286 2748 3350 2752
rect 3286 2692 3290 2748
rect 3290 2692 3346 2748
rect 3346 2692 3350 2748
rect 3286 2688 3350 2692
rect 3366 2748 3430 2752
rect 3366 2692 3370 2748
rect 3370 2692 3426 2748
rect 3426 2692 3430 2748
rect 3366 2688 3430 2692
rect 3446 2748 3510 2752
rect 3446 2692 3450 2748
rect 3450 2692 3506 2748
rect 3506 2692 3510 2748
rect 3446 2688 3510 2692
rect 9186 2748 9250 2752
rect 9186 2692 9190 2748
rect 9190 2692 9246 2748
rect 9246 2692 9250 2748
rect 9186 2688 9250 2692
rect 9266 2748 9330 2752
rect 9266 2692 9270 2748
rect 9270 2692 9326 2748
rect 9326 2692 9330 2748
rect 9266 2688 9330 2692
rect 9346 2748 9410 2752
rect 9346 2692 9350 2748
rect 9350 2692 9406 2748
rect 9406 2692 9410 2748
rect 9346 2688 9410 2692
rect 9426 2748 9490 2752
rect 9426 2692 9430 2748
rect 9430 2692 9486 2748
rect 9486 2692 9490 2748
rect 9426 2688 9490 2692
rect 15166 2748 15230 2752
rect 15166 2692 15170 2748
rect 15170 2692 15226 2748
rect 15226 2692 15230 2748
rect 15166 2688 15230 2692
rect 15246 2748 15310 2752
rect 15246 2692 15250 2748
rect 15250 2692 15306 2748
rect 15306 2692 15310 2748
rect 15246 2688 15310 2692
rect 15326 2748 15390 2752
rect 15326 2692 15330 2748
rect 15330 2692 15386 2748
rect 15386 2692 15390 2748
rect 15326 2688 15390 2692
rect 15406 2748 15470 2752
rect 15406 2692 15410 2748
rect 15410 2692 15466 2748
rect 15466 2692 15470 2748
rect 15406 2688 15470 2692
rect 6196 2204 6260 2208
rect 6196 2148 6200 2204
rect 6200 2148 6256 2204
rect 6256 2148 6260 2204
rect 6196 2144 6260 2148
rect 6276 2204 6340 2208
rect 6276 2148 6280 2204
rect 6280 2148 6336 2204
rect 6336 2148 6340 2204
rect 6276 2144 6340 2148
rect 6356 2204 6420 2208
rect 6356 2148 6360 2204
rect 6360 2148 6416 2204
rect 6416 2148 6420 2204
rect 6356 2144 6420 2148
rect 6436 2204 6500 2208
rect 6436 2148 6440 2204
rect 6440 2148 6496 2204
rect 6496 2148 6500 2204
rect 6436 2144 6500 2148
rect 12176 2204 12240 2208
rect 12176 2148 12180 2204
rect 12180 2148 12236 2204
rect 12236 2148 12240 2204
rect 12176 2144 12240 2148
rect 12256 2204 12320 2208
rect 12256 2148 12260 2204
rect 12260 2148 12316 2204
rect 12316 2148 12320 2204
rect 12256 2144 12320 2148
rect 12336 2204 12400 2208
rect 12336 2148 12340 2204
rect 12340 2148 12396 2204
rect 12396 2148 12400 2204
rect 12336 2144 12400 2148
rect 12416 2204 12480 2208
rect 12416 2148 12420 2204
rect 12420 2148 12476 2204
rect 12476 2148 12480 2204
rect 12416 2144 12480 2148
<< metal4 >>
rect 3198 4928 3518 5488
rect 3198 4864 3206 4928
rect 3270 4864 3286 4928
rect 3350 4864 3366 4928
rect 3430 4864 3446 4928
rect 3510 4864 3518 4928
rect 3198 3840 3518 4864
rect 3198 3776 3206 3840
rect 3270 3776 3286 3840
rect 3350 3776 3366 3840
rect 3430 3776 3446 3840
rect 3510 3776 3518 3840
rect 3198 2752 3518 3776
rect 3198 2688 3206 2752
rect 3270 2688 3286 2752
rect 3350 2688 3366 2752
rect 3430 2688 3446 2752
rect 3510 2688 3518 2752
rect 3198 2128 3518 2688
rect 6188 5472 6508 5488
rect 6188 5408 6196 5472
rect 6260 5408 6276 5472
rect 6340 5408 6356 5472
rect 6420 5408 6436 5472
rect 6500 5408 6508 5472
rect 6188 4384 6508 5408
rect 6188 4320 6196 4384
rect 6260 4320 6276 4384
rect 6340 4320 6356 4384
rect 6420 4320 6436 4384
rect 6500 4320 6508 4384
rect 6188 3296 6508 4320
rect 6188 3232 6196 3296
rect 6260 3232 6276 3296
rect 6340 3232 6356 3296
rect 6420 3232 6436 3296
rect 6500 3232 6508 3296
rect 6188 2208 6508 3232
rect 6188 2144 6196 2208
rect 6260 2144 6276 2208
rect 6340 2144 6356 2208
rect 6420 2144 6436 2208
rect 6500 2144 6508 2208
rect 6188 2128 6508 2144
rect 9178 4928 9498 5488
rect 9178 4864 9186 4928
rect 9250 4864 9266 4928
rect 9330 4864 9346 4928
rect 9410 4864 9426 4928
rect 9490 4864 9498 4928
rect 9178 3840 9498 4864
rect 9178 3776 9186 3840
rect 9250 3776 9266 3840
rect 9330 3776 9346 3840
rect 9410 3776 9426 3840
rect 9490 3776 9498 3840
rect 9178 2752 9498 3776
rect 9178 2688 9186 2752
rect 9250 2688 9266 2752
rect 9330 2688 9346 2752
rect 9410 2688 9426 2752
rect 9490 2688 9498 2752
rect 9178 2128 9498 2688
rect 12168 5472 12488 5488
rect 12168 5408 12176 5472
rect 12240 5408 12256 5472
rect 12320 5408 12336 5472
rect 12400 5408 12416 5472
rect 12480 5408 12488 5472
rect 12168 4384 12488 5408
rect 12168 4320 12176 4384
rect 12240 4320 12256 4384
rect 12320 4320 12336 4384
rect 12400 4320 12416 4384
rect 12480 4320 12488 4384
rect 12168 3296 12488 4320
rect 12168 3232 12176 3296
rect 12240 3232 12256 3296
rect 12320 3232 12336 3296
rect 12400 3232 12416 3296
rect 12480 3232 12488 3296
rect 12168 2208 12488 3232
rect 12168 2144 12176 2208
rect 12240 2144 12256 2208
rect 12320 2144 12336 2208
rect 12400 2144 12416 2208
rect 12480 2144 12488 2208
rect 12168 2128 12488 2144
rect 15158 4928 15478 5488
rect 15158 4864 15166 4928
rect 15230 4864 15246 4928
rect 15310 4864 15326 4928
rect 15390 4864 15406 4928
rect 15470 4864 15478 4928
rect 15158 3840 15478 4864
rect 15158 3776 15166 3840
rect 15230 3776 15246 3840
rect 15310 3776 15326 3840
rect 15390 3776 15406 3840
rect 15470 3776 15478 3840
rect 15158 2752 15478 3776
rect 15158 2688 15166 2752
rect 15230 2688 15246 2752
rect 15310 2688 15326 2752
rect 15390 2688 15406 2752
rect 15470 2688 15478 2752
rect 15158 2128 15478 2688
use sky130_fd_sc_hd__decap_3  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1196 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16
timestamp 1644511149
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1644511149
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45
timestamp 1644511149
transform 1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1644511149
transform 1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1644511149
transform 1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79
timestamp 1644511149
transform 1 0 7636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8004 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1644511149
transform 1 0 9200 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1644511149
transform 1 0 10304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_122
timestamp 1644511149
transform 1 0 11592 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135
timestamp 1644511149
transform 1 0 12788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1644511149
transform 1 0 13156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_144
timestamp 1644511149
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_151 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_159 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1644511149
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_169
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_180 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16928 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3
timestamp 1644511149
transform 1 0 644 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7
timestamp 1644511149
transform 1 0 1012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_31
timestamp 1644511149
transform 1 0 3220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_60
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_67
timestamp 1644511149
transform 1 0 6532 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_91
timestamp 1644511149
transform 1 0 8740 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1644511149
transform 1 0 10212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 10580 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_133
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_141
timestamp 1644511149
transform 1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_147
timestamp 1644511149
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_154
timestamp 1644511149
transform 1 0 14536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15180 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 15732 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_173
timestamp 1644511149
transform 1 0 16284 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1644511149
transform 1 0 16928 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1644511149
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 644 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_11
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 2576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_53
timestamp 1644511149
transform 1 0 5244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_59
timestamp 1644511149
transform 1 0 5796 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 7728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_89
timestamp 1644511149
transform 1 0 8556 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_97
timestamp 1644511149
transform 1 0 9292 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_105
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_109
timestamp 1644511149
transform 1 0 10396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_122
timestamp 1644511149
transform 1 0 11592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_129
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 12880 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_161
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_185
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_191
timestamp 1644511149
transform 1 0 17940 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1644511149
transform 1 0 644 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_29
timestamp 1644511149
transform 1 0 3036 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_39
timestamp 1644511149
transform 1 0 3956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_57
timestamp 1644511149
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_67
timestamp 1644511149
transform 1 0 6532 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_75
timestamp 1644511149
transform 1 0 7268 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_97
timestamp 1644511149
transform 1 0 9292 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_103
timestamp 1644511149
transform 1 0 9844 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1644511149
transform 1 0 10304 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_124
timestamp 1644511149
transform 1 0 11776 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1644511149
transform 1 0 12512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_156
timestamp 1644511149
transform 1 0 14720 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp 1644511149
transform 1 0 15364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 15732 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1644511149
transform 1 0 16836 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_183
timestamp 1644511149
transform 1 0 17204 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_188
timestamp 1644511149
transform 1 0 17664 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1644511149
transform 1 0 644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_13
timestamp 1644511149
transform 1 0 1564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp 1644511149
transform 1 0 2300 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 2852 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_33
timestamp 1644511149
transform 1 0 3404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_59
timestamp 1644511149
transform 1 0 5796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_69
timestamp 1644511149
transform 1 0 6716 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_79
timestamp 1644511149
transform 1 0 7636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8004 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_88
timestamp 1644511149
transform 1 0 8464 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_97
timestamp 1644511149
transform 1 0 9292 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_121
timestamp 1644511149
transform 1 0 11500 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_129
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1644511149
transform 1 0 12880 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_145
timestamp 1644511149
transform 1 0 13708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_171
timestamp 1644511149
transform 1 0 16100 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_179
timestamp 1644511149
transform 1 0 16836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_187
timestamp 1644511149
transform 1 0 17572 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_191
timestamp 1644511149
transform 1 0 17940 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1644511149
transform 1 0 644 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_24
timestamp 1644511149
transform 1 0 2576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_33
timestamp 1644511149
transform 1 0 3404 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_43
timestamp 1644511149
transform 1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_47
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1644511149
transform 1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1644511149
transform 1 0 5612 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_78
timestamp 1644511149
transform 1 0 7544 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_85
timestamp 1644511149
transform 1 0 8188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_91
timestamp 1644511149
transform 1 0 8740 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_95
timestamp 1644511149
transform 1 0 9108 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_100
timestamp 1644511149
transform 1 0 9568 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1644511149
transform 1 0 10304 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_133
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_139
timestamp 1644511149
transform 1 0 13156 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_141
timestamp 1644511149
transform 1 0 13340 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1644511149
transform 1 0 15456 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_173
timestamp 1644511149
transform 1 0 16284 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_181
timestamp 1644511149
transform 1 0 17020 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_188
timestamp 1644511149
transform 1 0 17664 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 368 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 368 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 368 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 368 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 18308 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 368 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_13
timestamp 1644511149
transform 1 0 5520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_14
timestamp 1644511149
transform 1 0 8096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_15
timestamp 1644511149
transform 1 0 10672 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_16
timestamp 1644511149
transform 1 0 13248 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_17
timestamp 1644511149
transform 1 0 15824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_18
timestamp 1644511149
transform 1 0 5520 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_19
timestamp 1644511149
transform 1 0 10672 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20
timestamp 1644511149
transform 1 0 15824 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1644511149
transform 1 0 2944 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1644511149
transform 1 0 8096 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1644511149
transform 1 0 13248 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1644511149
transform 1 0 5520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1644511149
transform 1 0 10672 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1644511149
transform 1 0 15824 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1644511149
transform 1 0 2944 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1644511149
transform 1 0 8096 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1644511149
transform 1 0 13248 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1644511149
transform 1 0 2944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1644511149
transform 1 0 5520 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1644511149
transform 1 0 8096 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1644511149
transform 1 0 10672 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1644511149
transform 1 0 13248 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1644511149
transform 1 0 15824 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _24_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _25_
timestamp 1644511149
transform -1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _26_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _27_
timestamp 1644511149
transform -1 0 16284 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _28_
timestamp 1644511149
transform -1 0 13708 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _29_
timestamp 1644511149
transform 1 0 9936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _30_
timestamp 1644511149
transform -1 0 12880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _31_
timestamp 1644511149
transform -1 0 15364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _32_
timestamp 1644511149
transform 1 0 17388 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _33_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10764 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _34_
timestamp 1644511149
transform 1 0 11960 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _35_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _36_
timestamp 1644511149
transform -1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _37_
timestamp 1644511149
transform -1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _38_
timestamp 1644511149
transform 1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _39_
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _40_
timestamp 1644511149
transform -1 0 6716 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _41_
timestamp 1644511149
transform -1 0 8556 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _42_
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _43_
timestamp 1644511149
transform -1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _44_
timestamp 1644511149
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _45_
timestamp 1644511149
transform -1 0 14536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _46_
timestamp 1644511149
transform -1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _47_
timestamp 1644511149
transform 1 0 10764 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _48_
timestamp 1644511149
transform -1 0 11776 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _49_
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _50_
timestamp 1644511149
transform -1 0 9292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _51_
timestamp 1644511149
transform 1 0 12604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _52_
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _53_
timestamp 1644511149
transform 1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _54__1
timestamp 1644511149
transform -1 0 1840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _55__2
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _56_
timestamp 1644511149
transform -1 0 5152 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _57_
timestamp 1644511149
transform -1 0 2576 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _58_
timestamp 1644511149
transform -1 0 1012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _59_
timestamp 1644511149
transform -1 0 1196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _60_
timestamp 1644511149
transform 1 0 6716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _61_
timestamp 1644511149
transform 1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _62_
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _63_
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _64_
timestamp 1644511149
transform 1 0 14904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _65_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6900 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _66_
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _67_
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _68_
timestamp 1644511149
transform 1 0 15548 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _69_
timestamp 1644511149
transform 1 0 12880 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _70_
timestamp 1644511149
transform -1 0 11500 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _71_
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _72_
timestamp 1644511149
transform 1 0 14260 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _73_
timestamp 1644511149
transform -1 0 15456 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_2  _74_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _75_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 4508 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _76_
timestamp 1644511149
transform -1 0 3220 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _77_
timestamp 1644511149
transform 1 0 1196 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _78_
timestamp 1644511149
transform -1 0 2576 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _79_
timestamp 1644511149
transform 1 0 3956 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _80_
timestamp 1644511149
transform 1 0 5704 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _81_
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _82_
timestamp 1644511149
transform -1 0 7728 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  _83_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3036 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_ext $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3404 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_clk_ext $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_clk_ext
timestamp 1644511149
transform -1 0 3956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 10304 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9476 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1644511149
transform 1 0 5612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1644511149
transform -1 0 9200 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1644511149
transform -1 0 12236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1644511149
transform -1 0 12512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1644511149
transform 1 0 16468 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1644511149
transform 1 0 17204 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1644511149
transform 1 0 17296 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1644511149
transform 1 0 1196 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1644511149
transform 1 0 3036 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1644511149
transform -1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1644511149
transform -1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1644511149
transform -1 0 6532 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1644511149
transform -1 0 7636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1644511149
transform -1 0 8740 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1644511149
transform 1 0 9200 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1644511149
transform -1 0 10304 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1644511149
transform 1 0 17296 0 -1 3264
box -38 -48 406 592
<< labels >>
rlabel metal4 s 6188 2128 6508 5488 6 VGND
port 0 nsew ground input
rlabel metal4 s 12168 2128 12488 5488 6 VGND
port 0 nsew ground input
rlabel metal4 s 3198 2128 3518 5488 6 VPWR
port 1 nsew power input
rlabel metal4 s 9178 2128 9498 5488 6 VPWR
port 1 nsew power input
rlabel metal4 s 15158 2128 15478 5488 6 VPWR
port 1 nsew power input
rlabel metal3 s 0 3136 400 3256 6 clk_ext
port 2 nsew signal input
rlabel metal2 s 570 5922 626 6322 6 f_out[0]
port 3 nsew signal tristate
rlabel metal2 s 11610 5922 11666 6322 6 f_out[10]
port 4 nsew signal tristate
rlabel metal2 s 12714 5922 12770 6322 6 f_out[11]
port 5 nsew signal tristate
rlabel metal2 s 13818 5922 13874 6322 6 f_out[12]
port 6 nsew signal tristate
rlabel metal2 s 14922 5922 14978 6322 6 f_out[13]
port 7 nsew signal tristate
rlabel metal2 s 16026 5922 16082 6322 6 f_out[14]
port 8 nsew signal tristate
rlabel metal2 s 17130 5922 17186 6322 6 f_out[15]
port 9 nsew signal tristate
rlabel metal2 s 18234 5922 18290 6322 6 f_out[16]
port 10 nsew signal tristate
rlabel metal2 s 1674 5922 1730 6322 6 f_out[1]
port 11 nsew signal tristate
rlabel metal2 s 2778 5922 2834 6322 6 f_out[2]
port 12 nsew signal tristate
rlabel metal2 s 3882 5922 3938 6322 6 f_out[3]
port 13 nsew signal tristate
rlabel metal2 s 4986 5922 5042 6322 6 f_out[4]
port 14 nsew signal tristate
rlabel metal2 s 6090 5922 6146 6322 6 f_out[5]
port 15 nsew signal tristate
rlabel metal2 s 7194 5922 7250 6322 6 f_out[6]
port 16 nsew signal tristate
rlabel metal2 s 8298 5922 8354 6322 6 f_out[7]
port 17 nsew signal tristate
rlabel metal2 s 9402 5922 9458 6322 6 f_out[8]
port 18 nsew signal tristate
rlabel metal2 s 10506 5922 10562 6322 6 f_out[9]
port 19 nsew signal tristate
rlabel metal2 s 9402 0 9458 400 6 rst_ext
port 20 nsew signal input
rlabel metal3 s 18345 3136 18745 3256 6 rstb
port 21 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 18745 6322
<< end >>
