VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO filter_p_m
  CLASS BLOCK ;
  FOREIGN filter_p_m ;
  ORIGIN 0.130 1.640 ;
  SIZE 253.920 BY 187.340 ;
  PIN cclk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.580 165.160 67.860 185.700 ;
    END
  END cclk
  PIN fb1
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.260 175.700 25.540 185.700 ;
    END
  END fb1
  PIN div2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.900 177.350 110.180 185.700 ;
    END
  END div2
  PIN high_buf
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 152.220 177.405 152.500 185.700 ;
    END
  END high_buf
  PIN phi1b_dig
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 194.540 177.285 194.820 185.700 ;
    END
  END phi1b_dig
  PIN lo
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.860 174.915 237.140 185.700 ;
    END
  END lo
  OBS
      LAYER li1 ;
        RECT 3.100 125.140 237.280 175.850 ;
      LAYER met1 ;
        RECT 2.435 125.505 237.945 177.380 ;
      LAYER met2 ;
        RECT 2.460 175.420 24.980 177.450 ;
        RECT 25.820 175.420 67.300 177.450 ;
        RECT 2.460 164.880 67.300 175.420 ;
        RECT 68.140 177.070 109.620 177.450 ;
        RECT 110.460 177.125 151.940 177.450 ;
        RECT 152.780 177.125 194.260 177.450 ;
        RECT 110.460 177.070 194.260 177.125 ;
        RECT 68.140 177.005 194.260 177.070 ;
        RECT 195.100 177.005 236.580 177.450 ;
        RECT 68.140 174.635 236.580 177.005 ;
        RECT 237.420 174.635 237.920 177.450 ;
        RECT 68.140 164.880 237.920 174.635 ;
        RECT 2.460 126.325 237.920 164.880 ;
      LAYER met3 ;
        RECT -0.130 0.000 253.790 177.430 ;
      LAYER met4 ;
        RECT -0.130 -1.640 253.790 177.430 ;
      LAYER met5 ;
        RECT -0.130 -1.640 253.790 140.315 ;
  END
END filter_p_m
END LIBRARY

