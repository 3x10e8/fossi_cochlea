VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital_unison
  CLASS BLOCK ;
  FOREIGN digital_unison ;
  ORIGIN 0.000 0.000 ;
  SIZE 1440.000 BY 120.000 ;
  PIN cclk_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 116.000 146.190 120.000 ;
    END
  END cclk_I[0]
  PIN cclk_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 116.000 383.550 120.000 ;
    END
  END cclk_I[1]
  PIN cclk_I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 116.000 620.910 120.000 ;
    END
  END cclk_I[2]
  PIN cclk_I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.990 116.000 858.270 120.000 ;
    END
  END cclk_I[3]
  PIN cclk_I[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.350 116.000 1095.630 120.000 ;
    END
  END cclk_I[4]
  PIN cclk_I[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.710 116.000 1332.990 120.000 ;
    END
  END cclk_I[5]
  PIN cclk_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END cclk_Q[0]
  PIN cclk_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END cclk_Q[1]
  PIN cclk_Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 0.000 620.910 4.000 ;
    END
  END cclk_Q[2]
  PIN cclk_Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.990 0.000 858.270 4.000 ;
    END
  END cclk_Q[3]
  PIN cclk_Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.350 0.000 1095.630 4.000 ;
    END
  END cclk_Q[4]
  PIN cclk_Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.710 0.000 1332.990 4.000 ;
    END
  END cclk_Q[5]
  PIN clk_master
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END clk_master
  PIN clkdiv2_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 116.000 106.630 120.000 ;
    END
  END clkdiv2_I[0]
  PIN clkdiv2_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 116.000 343.990 120.000 ;
    END
  END clkdiv2_I[1]
  PIN clkdiv2_I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 116.000 581.350 120.000 ;
    END
  END clkdiv2_I[2]
  PIN clkdiv2_I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 116.000 818.710 120.000 ;
    END
  END clkdiv2_I[3]
  PIN clkdiv2_I[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.790 116.000 1056.070 120.000 ;
    END
  END clkdiv2_I[4]
  PIN clkdiv2_I[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.150 116.000 1293.430 120.000 ;
    END
  END clkdiv2_I[5]
  PIN clkdiv2_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END clkdiv2_Q[0]
  PIN clkdiv2_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END clkdiv2_Q[1]
  PIN clkdiv2_Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 4.000 ;
    END
  END clkdiv2_Q[2]
  PIN clkdiv2_Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 0.000 818.710 4.000 ;
    END
  END clkdiv2_Q[3]
  PIN clkdiv2_Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.790 0.000 1056.070 4.000 ;
    END
  END clkdiv2_Q[4]
  PIN clkdiv2_Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.150 0.000 1293.430 4.000 ;
    END
  END clkdiv2_Q[5]
  PIN comp_high_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 116.000 225.310 120.000 ;
    END
  END comp_high_I[0]
  PIN comp_high_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 116.000 462.670 120.000 ;
    END
  END comp_high_I[1]
  PIN comp_high_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 116.000 700.030 120.000 ;
    END
  END comp_high_I[2]
  PIN comp_high_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 116.000 937.390 120.000 ;
    END
  END comp_high_I[3]
  PIN comp_high_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.470 116.000 1174.750 120.000 ;
    END
  END comp_high_I[4]
  PIN comp_high_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1411.830 116.000 1412.110 120.000 ;
    END
  END comp_high_I[5]
  PIN comp_high_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END comp_high_Q[0]
  PIN comp_high_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END comp_high_Q[1]
  PIN comp_high_Q[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 0.000 700.030 4.000 ;
    END
  END comp_high_Q[2]
  PIN comp_high_Q[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 0.000 937.390 4.000 ;
    END
  END comp_high_Q[3]
  PIN comp_high_Q[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.470 0.000 1174.750 4.000 ;
    END
  END comp_high_Q[4]
  PIN comp_high_Q[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1411.830 0.000 1412.110 4.000 ;
    END
  END comp_high_Q[5]
  PIN cos_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 116.000 27.510 120.000 ;
    END
  END cos_out[0]
  PIN cos_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 116.000 264.870 120.000 ;
    END
  END cos_out[1]
  PIN cos_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 116.000 502.230 120.000 ;
    END
  END cos_out[2]
  PIN cos_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 116.000 739.590 120.000 ;
    END
  END cos_out[3]
  PIN cos_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 116.000 976.950 120.000 ;
    END
  END cos_out[4]
  PIN cos_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.030 116.000 1214.310 120.000 ;
    END
  END cos_out[5]
  PIN fb1_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 116.000 67.070 120.000 ;
    END
  END fb1_I[0]
  PIN fb1_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 116.000 304.430 120.000 ;
    END
  END fb1_I[1]
  PIN fb1_I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 116.000 541.790 120.000 ;
    END
  END fb1_I[2]
  PIN fb1_I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.870 116.000 779.150 120.000 ;
    END
  END fb1_I[3]
  PIN fb1_I[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.230 116.000 1016.510 120.000 ;
    END
  END fb1_I[4]
  PIN fb1_I[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.590 116.000 1253.870 120.000 ;
    END
  END fb1_I[5]
  PIN fb1_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END fb1_Q[0]
  PIN fb1_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END fb1_Q[1]
  PIN fb1_Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 0.000 541.790 4.000 ;
    END
  END fb1_Q[2]
  PIN fb1_Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.870 0.000 779.150 4.000 ;
    END
  END fb1_Q[3]
  PIN fb1_Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.230 0.000 1016.510 4.000 ;
    END
  END fb1_Q[4]
  PIN fb1_Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.590 0.000 1253.870 4.000 ;
    END
  END fb1_Q[5]
  PIN phi1b_dig_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 116.000 185.750 120.000 ;
    END
  END phi1b_dig_I[0]
  PIN phi1b_dig_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 116.000 423.110 120.000 ;
    END
  END phi1b_dig_I[1]
  PIN phi1b_dig_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 116.000 660.470 120.000 ;
    END
  END phi1b_dig_I[2]
  PIN phi1b_dig_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 116.000 897.830 120.000 ;
    END
  END phi1b_dig_I[3]
  PIN phi1b_dig_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.910 116.000 1135.190 120.000 ;
    END
  END phi1b_dig_I[4]
  PIN phi1b_dig_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1372.270 116.000 1372.550 120.000 ;
    END
  END phi1b_dig_I[5]
  PIN phi1b_dig_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END phi1b_dig_Q[0]
  PIN phi1b_dig_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END phi1b_dig_Q[1]
  PIN phi1b_dig_Q[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END phi1b_dig_Q[2]
  PIN phi1b_dig_Q[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 0.000 897.830 4.000 ;
    END
  END phi1b_dig_Q[3]
  PIN phi1b_dig_Q[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.910 0.000 1135.190 4.000 ;
    END
  END phi1b_dig_Q[4]
  PIN phi1b_dig_Q[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1372.270 0.000 1372.550 4.000 ;
    END
  END phi1b_dig_Q[5]
  PIN read_out_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1436.000 104.080 1440.000 104.680 ;
    END
  END read_out_I[0]
  PIN read_out_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1436.000 74.160 1440.000 74.760 ;
    END
  END read_out_I[1]
  PIN read_out_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1436.000 44.240 1440.000 44.840 ;
    END
  END read_out_Q[0]
  PIN read_out_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1436.000 14.320 1440.000 14.920 ;
    END
  END read_out_Q[1]
  PIN rstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END rstb
  PIN sin_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END sin_out[0]
  PIN sin_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END sin_out[1]
  PIN sin_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END sin_out[2]
  PIN sin_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 0.000 739.590 4.000 ;
    END
  END sin_out[3]
  PIN sin_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 0.000 976.950 4.000 ;
    END
  END sin_out[4]
  PIN sin_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.030 0.000 1214.310 4.000 ;
    END
  END sin_out[5]
  PIN ud_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END ud_en
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 183.315 10.640 184.915 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 540.505 10.640 542.105 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 897.695 10.640 899.295 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.885 10.640 1256.485 109.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 361.910 10.640 363.510 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 719.100 10.640 720.700 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1076.290 10.640 1077.890 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1433.480 10.640 1435.080 109.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1434.280 108.885 ;
      LAYER met1 ;
        RECT 5.520 10.640 1435.080 117.260 ;
      LAYER met2 ;
        RECT 7.910 115.720 26.950 117.290 ;
        RECT 27.790 115.720 66.510 117.290 ;
        RECT 67.350 115.720 106.070 117.290 ;
        RECT 106.910 115.720 145.630 117.290 ;
        RECT 146.470 115.720 185.190 117.290 ;
        RECT 186.030 115.720 224.750 117.290 ;
        RECT 225.590 115.720 264.310 117.290 ;
        RECT 265.150 115.720 303.870 117.290 ;
        RECT 304.710 115.720 343.430 117.290 ;
        RECT 344.270 115.720 382.990 117.290 ;
        RECT 383.830 115.720 422.550 117.290 ;
        RECT 423.390 115.720 462.110 117.290 ;
        RECT 462.950 115.720 501.670 117.290 ;
        RECT 502.510 115.720 541.230 117.290 ;
        RECT 542.070 115.720 580.790 117.290 ;
        RECT 581.630 115.720 620.350 117.290 ;
        RECT 621.190 115.720 659.910 117.290 ;
        RECT 660.750 115.720 699.470 117.290 ;
        RECT 700.310 115.720 739.030 117.290 ;
        RECT 739.870 115.720 778.590 117.290 ;
        RECT 779.430 115.720 818.150 117.290 ;
        RECT 818.990 115.720 857.710 117.290 ;
        RECT 858.550 115.720 897.270 117.290 ;
        RECT 898.110 115.720 936.830 117.290 ;
        RECT 937.670 115.720 976.390 117.290 ;
        RECT 977.230 115.720 1015.950 117.290 ;
        RECT 1016.790 115.720 1055.510 117.290 ;
        RECT 1056.350 115.720 1095.070 117.290 ;
        RECT 1095.910 115.720 1134.630 117.290 ;
        RECT 1135.470 115.720 1174.190 117.290 ;
        RECT 1175.030 115.720 1213.750 117.290 ;
        RECT 1214.590 115.720 1253.310 117.290 ;
        RECT 1254.150 115.720 1292.870 117.290 ;
        RECT 1293.710 115.720 1332.430 117.290 ;
        RECT 1333.270 115.720 1371.990 117.290 ;
        RECT 1372.830 115.720 1411.550 117.290 ;
        RECT 1412.390 115.720 1435.050 117.290 ;
        RECT 7.910 4.280 1435.050 115.720 ;
        RECT 7.910 4.000 26.950 4.280 ;
        RECT 27.790 4.000 66.510 4.280 ;
        RECT 67.350 4.000 106.070 4.280 ;
        RECT 106.910 4.000 145.630 4.280 ;
        RECT 146.470 4.000 185.190 4.280 ;
        RECT 186.030 4.000 224.750 4.280 ;
        RECT 225.590 4.000 264.310 4.280 ;
        RECT 265.150 4.000 303.870 4.280 ;
        RECT 304.710 4.000 343.430 4.280 ;
        RECT 344.270 4.000 382.990 4.280 ;
        RECT 383.830 4.000 422.550 4.280 ;
        RECT 423.390 4.000 462.110 4.280 ;
        RECT 462.950 4.000 501.670 4.280 ;
        RECT 502.510 4.000 541.230 4.280 ;
        RECT 542.070 4.000 580.790 4.280 ;
        RECT 581.630 4.000 620.350 4.280 ;
        RECT 621.190 4.000 659.910 4.280 ;
        RECT 660.750 4.000 699.470 4.280 ;
        RECT 700.310 4.000 739.030 4.280 ;
        RECT 739.870 4.000 778.590 4.280 ;
        RECT 779.430 4.000 818.150 4.280 ;
        RECT 818.990 4.000 857.710 4.280 ;
        RECT 858.550 4.000 897.270 4.280 ;
        RECT 898.110 4.000 936.830 4.280 ;
        RECT 937.670 4.000 976.390 4.280 ;
        RECT 977.230 4.000 1015.950 4.280 ;
        RECT 1016.790 4.000 1055.510 4.280 ;
        RECT 1056.350 4.000 1095.070 4.280 ;
        RECT 1095.910 4.000 1134.630 4.280 ;
        RECT 1135.470 4.000 1174.190 4.280 ;
        RECT 1175.030 4.000 1213.750 4.280 ;
        RECT 1214.590 4.000 1253.310 4.280 ;
        RECT 1254.150 4.000 1292.870 4.280 ;
        RECT 1293.710 4.000 1332.430 4.280 ;
        RECT 1333.270 4.000 1371.990 4.280 ;
        RECT 1372.830 4.000 1411.550 4.280 ;
        RECT 1412.390 4.000 1435.050 4.280 ;
      LAYER met3 ;
        RECT 4.000 105.080 1436.000 111.345 ;
        RECT 4.000 103.680 1435.600 105.080 ;
        RECT 4.000 99.640 1436.000 103.680 ;
        RECT 4.400 98.240 1436.000 99.640 ;
        RECT 4.000 75.160 1436.000 98.240 ;
        RECT 4.000 73.760 1435.600 75.160 ;
        RECT 4.000 60.200 1436.000 73.760 ;
        RECT 4.400 58.800 1436.000 60.200 ;
        RECT 4.000 45.240 1436.000 58.800 ;
        RECT 4.000 43.840 1435.600 45.240 ;
        RECT 4.000 20.760 1436.000 43.840 ;
        RECT 4.400 19.360 1436.000 20.760 ;
        RECT 4.000 15.320 1436.000 19.360 ;
        RECT 4.000 13.920 1435.600 15.320 ;
        RECT 4.000 10.715 1436.000 13.920 ;
      LAYER met4 ;
        RECT 39.855 109.440 1394.425 111.345 ;
        RECT 39.855 11.735 182.915 109.440 ;
        RECT 185.315 11.735 361.510 109.440 ;
        RECT 363.910 11.735 540.105 109.440 ;
        RECT 542.505 11.735 718.700 109.440 ;
        RECT 721.100 11.735 897.295 109.440 ;
        RECT 899.695 11.735 1075.890 109.440 ;
        RECT 1078.290 11.735 1254.485 109.440 ;
        RECT 1256.885 11.735 1394.425 109.440 ;
  END
END digital_unison
END LIBRARY

