magic
tech sky130A
timestamp 1647573571
<< nwell >>
rect 2694 -1643 3074 -1555
rect 8615 -1643 8995 -1555
<< nmos >>
rect 2739 -1803 2754 -1761
rect 2783 -1803 2798 -1761
rect 2827 -1803 2842 -1761
rect 2871 -1803 2886 -1761
rect 2915 -1803 2930 -1761
rect 2959 -1803 2974 -1761
rect 8715 -1803 8730 -1761
rect 8759 -1803 8774 -1761
rect 8803 -1803 8818 -1761
rect 8847 -1803 8862 -1761
rect 8891 -1803 8906 -1761
rect 8935 -1803 8950 -1761
<< pmos >>
rect 2739 -1625 2754 -1583
rect 2783 -1625 2798 -1583
rect 2827 -1625 2842 -1583
rect 2871 -1625 2886 -1583
rect 2915 -1625 2930 -1583
rect 2959 -1625 2974 -1583
rect 8715 -1625 8730 -1583
rect 8759 -1625 8774 -1583
rect 8803 -1625 8818 -1583
rect 8847 -1625 8862 -1583
rect 8891 -1625 8906 -1583
rect 8935 -1625 8950 -1583
<< ndiff >>
rect 2712 -1773 2739 -1761
rect 2712 -1790 2716 -1773
rect 2733 -1790 2739 -1773
rect 2712 -1803 2739 -1790
rect 2754 -1773 2783 -1761
rect 2754 -1790 2760 -1773
rect 2777 -1790 2783 -1773
rect 2754 -1803 2783 -1790
rect 2798 -1773 2827 -1761
rect 2798 -1790 2804 -1773
rect 2821 -1790 2827 -1773
rect 2798 -1803 2827 -1790
rect 2842 -1773 2871 -1761
rect 2842 -1790 2848 -1773
rect 2865 -1790 2871 -1773
rect 2842 -1803 2871 -1790
rect 2886 -1773 2915 -1761
rect 2886 -1790 2892 -1773
rect 2909 -1790 2915 -1773
rect 2886 -1803 2915 -1790
rect 2930 -1773 2959 -1761
rect 2930 -1790 2936 -1773
rect 2953 -1790 2959 -1773
rect 2930 -1803 2959 -1790
rect 2974 -1773 3001 -1761
rect 2974 -1790 2980 -1773
rect 2997 -1790 3001 -1773
rect 2974 -1803 3001 -1790
rect 8688 -1773 8715 -1761
rect 8688 -1790 8692 -1773
rect 8709 -1790 8715 -1773
rect 8688 -1803 8715 -1790
rect 8730 -1773 8759 -1761
rect 8730 -1790 8736 -1773
rect 8753 -1790 8759 -1773
rect 8730 -1803 8759 -1790
rect 8774 -1773 8803 -1761
rect 8774 -1790 8780 -1773
rect 8797 -1790 8803 -1773
rect 8774 -1803 8803 -1790
rect 8818 -1773 8847 -1761
rect 8818 -1790 8824 -1773
rect 8841 -1790 8847 -1773
rect 8818 -1803 8847 -1790
rect 8862 -1773 8891 -1761
rect 8862 -1790 8868 -1773
rect 8885 -1790 8891 -1773
rect 8862 -1803 8891 -1790
rect 8906 -1773 8935 -1761
rect 8906 -1790 8912 -1773
rect 8929 -1790 8935 -1773
rect 8906 -1803 8935 -1790
rect 8950 -1773 8977 -1761
rect 8950 -1790 8956 -1773
rect 8973 -1790 8977 -1773
rect 8950 -1803 8977 -1790
<< pdiff >>
rect 2712 -1595 2739 -1583
rect 2712 -1612 2716 -1595
rect 2733 -1612 2739 -1595
rect 2712 -1625 2739 -1612
rect 2754 -1595 2783 -1583
rect 2754 -1612 2760 -1595
rect 2777 -1612 2783 -1595
rect 2754 -1625 2783 -1612
rect 2798 -1595 2827 -1583
rect 2798 -1612 2804 -1595
rect 2821 -1612 2827 -1595
rect 2798 -1625 2827 -1612
rect 2842 -1595 2871 -1583
rect 2842 -1612 2848 -1595
rect 2865 -1612 2871 -1595
rect 2842 -1625 2871 -1612
rect 2886 -1595 2915 -1583
rect 2886 -1612 2892 -1595
rect 2909 -1612 2915 -1595
rect 2886 -1625 2915 -1612
rect 2930 -1595 2959 -1583
rect 2930 -1612 2936 -1595
rect 2953 -1612 2959 -1595
rect 2930 -1625 2959 -1612
rect 2974 -1595 3001 -1583
rect 2974 -1612 2980 -1595
rect 2997 -1612 3001 -1595
rect 2974 -1625 3001 -1612
rect 8688 -1595 8715 -1583
rect 8688 -1612 8692 -1595
rect 8709 -1612 8715 -1595
rect 8688 -1625 8715 -1612
rect 8730 -1595 8759 -1583
rect 8730 -1612 8736 -1595
rect 8753 -1612 8759 -1595
rect 8730 -1625 8759 -1612
rect 8774 -1595 8803 -1583
rect 8774 -1612 8780 -1595
rect 8797 -1612 8803 -1595
rect 8774 -1625 8803 -1612
rect 8818 -1595 8847 -1583
rect 8818 -1612 8824 -1595
rect 8841 -1612 8847 -1595
rect 8818 -1625 8847 -1612
rect 8862 -1595 8891 -1583
rect 8862 -1612 8868 -1595
rect 8885 -1612 8891 -1595
rect 8862 -1625 8891 -1612
rect 8906 -1595 8935 -1583
rect 8906 -1612 8912 -1595
rect 8929 -1612 8935 -1595
rect 8906 -1625 8935 -1612
rect 8950 -1595 8977 -1583
rect 8950 -1612 8956 -1595
rect 8973 -1612 8977 -1595
rect 8950 -1625 8977 -1612
<< ndiffc >>
rect 2716 -1790 2733 -1773
rect 2760 -1790 2777 -1773
rect 2804 -1790 2821 -1773
rect 2848 -1790 2865 -1773
rect 2892 -1790 2909 -1773
rect 2936 -1790 2953 -1773
rect 2980 -1790 2997 -1773
rect 8692 -1790 8709 -1773
rect 8736 -1790 8753 -1773
rect 8780 -1790 8797 -1773
rect 8824 -1790 8841 -1773
rect 8868 -1790 8885 -1773
rect 8912 -1790 8929 -1773
rect 8956 -1790 8973 -1773
<< pdiffc >>
rect 2716 -1612 2733 -1595
rect 2760 -1612 2777 -1595
rect 2804 -1612 2821 -1595
rect 2848 -1612 2865 -1595
rect 2892 -1612 2909 -1595
rect 2936 -1612 2953 -1595
rect 2980 -1612 2997 -1595
rect 8692 -1612 8709 -1595
rect 8736 -1612 8753 -1595
rect 8780 -1612 8797 -1595
rect 8824 -1612 8841 -1595
rect 8868 -1612 8885 -1595
rect 8912 -1612 8929 -1595
rect 8956 -1612 8973 -1595
<< psubdiff >>
rect 2841 -1879 2868 -1866
rect 2841 -1896 2846 -1879
rect 2863 -1896 2868 -1879
rect 2841 -1908 2868 -1896
rect 8821 -1879 8848 -1866
rect 8821 -1896 8826 -1879
rect 8843 -1896 8848 -1879
rect 8821 -1908 8848 -1896
<< nsubdiff >>
rect 3029 -1596 3056 -1583
rect 3029 -1613 3034 -1596
rect 3051 -1613 3056 -1596
rect 3029 -1625 3056 -1613
rect 8633 -1596 8660 -1583
rect 8633 -1613 8638 -1596
rect 8655 -1613 8660 -1596
rect 8633 -1625 8660 -1613
<< psubdiffcont >>
rect 2846 -1896 2863 -1879
rect 8826 -1896 8843 -1879
<< nsubdiffcont >>
rect 3034 -1613 3051 -1596
rect 8638 -1613 8655 -1596
<< poly >>
rect 2735 -1531 2762 -1523
rect 2735 -1548 2740 -1531
rect 2757 -1534 2762 -1531
rect 8927 -1531 8954 -1523
rect 8927 -1534 8932 -1531
rect 2757 -1548 2930 -1534
rect 2735 -1549 2930 -1548
rect 2735 -1557 2762 -1549
rect 2739 -1583 2754 -1557
rect 2783 -1583 2798 -1570
rect 2827 -1583 2842 -1549
rect 2871 -1583 2886 -1570
rect 2915 -1583 2930 -1549
rect 8759 -1548 8932 -1534
rect 8949 -1548 8954 -1531
rect 8759 -1549 8954 -1548
rect 2959 -1583 2974 -1570
rect 8715 -1583 8730 -1570
rect 8759 -1583 8774 -1549
rect 8803 -1583 8818 -1570
rect 8847 -1583 8862 -1549
rect 8927 -1557 8954 -1549
rect 8891 -1583 8906 -1570
rect 8935 -1583 8950 -1557
rect 2739 -1638 2754 -1625
rect 2675 -1653 2702 -1645
rect 2675 -1670 2680 -1653
rect 2697 -1659 2702 -1653
rect 2783 -1659 2798 -1625
rect 2827 -1638 2842 -1625
rect 2871 -1659 2886 -1625
rect 2915 -1638 2930 -1625
rect 2959 -1659 2974 -1625
rect 2697 -1670 2974 -1659
rect 2675 -1674 2974 -1670
rect 8715 -1659 8730 -1625
rect 8759 -1638 8774 -1625
rect 8803 -1659 8818 -1625
rect 8847 -1638 8862 -1625
rect 8891 -1659 8906 -1625
rect 8935 -1638 8950 -1625
rect 8987 -1653 9014 -1645
rect 8987 -1659 8992 -1653
rect 8715 -1670 8992 -1659
rect 9009 -1670 9014 -1653
rect 8715 -1674 9014 -1670
rect 2675 -1679 2702 -1674
rect 8987 -1679 9014 -1674
rect 2675 -1709 2702 -1701
rect 2675 -1726 2680 -1709
rect 2697 -1712 2702 -1709
rect 8987 -1709 9014 -1701
rect 8987 -1712 8992 -1709
rect 2697 -1726 2930 -1712
rect 2675 -1727 2930 -1726
rect 2675 -1735 2702 -1727
rect 2739 -1761 2754 -1727
rect 2783 -1761 2798 -1748
rect 2827 -1761 2842 -1727
rect 2871 -1761 2886 -1748
rect 2915 -1761 2930 -1727
rect 8759 -1726 8992 -1712
rect 9009 -1726 9014 -1709
rect 8759 -1727 9014 -1726
rect 2959 -1761 2974 -1748
rect 8715 -1761 8730 -1748
rect 8759 -1761 8774 -1727
rect 8803 -1761 8818 -1748
rect 8847 -1761 8862 -1727
rect 8891 -1761 8906 -1748
rect 8935 -1761 8950 -1727
rect 8987 -1735 9014 -1727
rect 2739 -1816 2754 -1803
rect 2783 -1823 2798 -1803
rect 2827 -1816 2842 -1803
rect 2779 -1831 2806 -1823
rect 2779 -1848 2784 -1831
rect 2801 -1837 2806 -1831
rect 2871 -1837 2886 -1803
rect 2915 -1816 2930 -1803
rect 2959 -1837 2974 -1803
rect 2801 -1848 2974 -1837
rect 2779 -1852 2974 -1848
rect 8715 -1837 8730 -1803
rect 8759 -1816 8774 -1803
rect 8803 -1837 8818 -1803
rect 8847 -1816 8862 -1803
rect 8891 -1823 8906 -1803
rect 8935 -1816 8950 -1803
rect 8883 -1831 8910 -1823
rect 8883 -1837 8888 -1831
rect 8715 -1848 8888 -1837
rect 8905 -1848 8910 -1831
rect 8715 -1852 8910 -1848
rect 2779 -1857 2806 -1852
rect 8883 -1857 8910 -1852
<< polycont >>
rect 2740 -1548 2757 -1531
rect 8932 -1548 8949 -1531
rect 2680 -1670 2697 -1653
rect 8992 -1670 9009 -1653
rect 2680 -1726 2697 -1709
rect 8992 -1726 9009 -1709
rect 2784 -1848 2801 -1831
rect 8888 -1848 8905 -1831
<< locali >>
rect 2798 -1326 2828 -1319
rect 2798 -1344 2804 -1326
rect 2822 -1344 2828 -1326
rect 2798 -1351 2828 -1344
rect 2736 -1531 2761 -1523
rect 2736 -1548 2740 -1531
rect 2757 -1548 2761 -1531
rect 2736 -1557 2761 -1548
rect 2804 -1587 2821 -1351
rect 3613 -1385 3636 -1382
rect 3613 -1402 3616 -1385
rect 3633 -1402 3636 -1385
rect 3613 -1408 3636 -1402
rect 3035 -1426 3052 -1423
rect 2977 -1486 3000 -1480
rect 2977 -1503 2980 -1486
rect 2997 -1503 3000 -1486
rect 2977 -1509 3000 -1503
rect 2980 -1587 2997 -1509
rect 3035 -1583 3052 -1443
rect 3616 -1572 3633 -1408
rect 3660 -1514 3677 -1362
rect 3776 -1564 3793 -1281
rect 2715 -1591 2735 -1587
rect 2714 -1595 2735 -1591
rect 2714 -1612 2716 -1595
rect 2733 -1612 2735 -1595
rect 2714 -1620 2735 -1612
rect 2758 -1595 2779 -1587
rect 2758 -1612 2760 -1595
rect 2777 -1612 2779 -1595
rect 2758 -1620 2779 -1612
rect 2802 -1595 2823 -1587
rect 2802 -1612 2804 -1595
rect 2821 -1612 2823 -1595
rect 2802 -1620 2823 -1612
rect 2846 -1595 2867 -1587
rect 2846 -1612 2848 -1595
rect 2865 -1612 2867 -1595
rect 2846 -1620 2867 -1612
rect 2890 -1595 2911 -1587
rect 2890 -1612 2892 -1595
rect 2909 -1612 2911 -1595
rect 2890 -1620 2911 -1612
rect 2934 -1595 2955 -1587
rect 2934 -1612 2936 -1595
rect 2953 -1612 2955 -1595
rect 2934 -1620 2955 -1612
rect 2978 -1595 2999 -1587
rect 2978 -1612 2980 -1595
rect 2997 -1612 2999 -1595
rect 2978 -1620 2999 -1612
rect 3029 -1596 3056 -1583
rect 3616 -1589 3705 -1572
rect 3029 -1613 3034 -1596
rect 3051 -1613 3056 -1596
rect 2676 -1653 2701 -1645
rect 2676 -1670 2680 -1653
rect 2697 -1670 2701 -1653
rect 2676 -1679 2701 -1670
rect 2676 -1709 2701 -1701
rect 2676 -1726 2680 -1709
rect 2697 -1726 2701 -1709
rect 2676 -1735 2701 -1726
rect 2718 -1765 2735 -1620
rect 2760 -1765 2777 -1620
rect 2804 -1765 2821 -1620
rect 2848 -1765 2865 -1620
rect 2892 -1765 2909 -1620
rect 2936 -1765 2953 -1620
rect 2980 -1765 2997 -1620
rect 3029 -1625 3056 -1613
rect 2714 -1773 2735 -1765
rect 2714 -1790 2716 -1773
rect 2733 -1790 2735 -1773
rect 2714 -1798 2735 -1790
rect 2758 -1773 2779 -1765
rect 2758 -1790 2760 -1773
rect 2777 -1790 2779 -1773
rect 2758 -1798 2779 -1790
rect 2802 -1773 2823 -1765
rect 2802 -1790 2804 -1773
rect 2821 -1790 2823 -1773
rect 2802 -1798 2823 -1790
rect 2846 -1773 2867 -1765
rect 2846 -1790 2848 -1773
rect 2865 -1790 2867 -1773
rect 2846 -1798 2867 -1790
rect 2890 -1773 2911 -1765
rect 2890 -1790 2892 -1773
rect 2909 -1790 2911 -1773
rect 2890 -1798 2911 -1790
rect 2934 -1772 2955 -1765
rect 2934 -1790 2936 -1772
rect 2954 -1790 2955 -1772
rect 2934 -1798 2955 -1790
rect 2978 -1773 2999 -1765
rect 2978 -1790 2980 -1773
rect 2997 -1778 2999 -1773
rect 2997 -1790 3137 -1778
rect 2978 -1795 3137 -1790
rect 2978 -1798 2999 -1795
rect 2717 -1942 2734 -1798
rect 2780 -1831 2805 -1823
rect 2780 -1848 2784 -1831
rect 2801 -1848 2805 -1831
rect 2780 -1857 2805 -1848
rect 2841 -1879 2868 -1866
rect 2841 -1896 2846 -1879
rect 2863 -1896 2868 -1879
rect 2841 -1908 2868 -1896
rect 2892 -1976 2909 -1798
rect 3120 -1976 3137 -1795
rect 2885 -1983 2915 -1976
rect 2885 -2001 2891 -1983
rect 2909 -2001 2915 -1983
rect 2885 -2008 2915 -2001
rect 3113 -1983 3143 -1976
rect 3113 -2001 3119 -1983
rect 3137 -2001 3143 -1983
rect 3113 -2008 3143 -2001
rect 3620 -2003 3637 -1635
rect 3832 -1767 3849 -1322
rect 8861 -1326 8891 -1319
rect 8861 -1344 8867 -1326
rect 8885 -1344 8891 -1326
rect 8861 -1351 8891 -1344
rect 5218 -1428 5242 -1424
rect 5218 -1445 5221 -1428
rect 5238 -1445 5242 -1428
rect 5218 -1447 5242 -1445
rect 8637 -1426 8654 -1423
rect 5098 -1590 5104 -1573
rect 5121 -1590 5126 -1573
rect 5221 -1662 5238 -1447
rect 8637 -1583 8654 -1443
rect 8689 -1486 8712 -1480
rect 8689 -1503 8692 -1486
rect 8709 -1503 8712 -1486
rect 8689 -1509 8712 -1503
rect 8633 -1596 8660 -1583
rect 8692 -1587 8709 -1509
rect 8868 -1587 8885 -1351
rect 8928 -1531 8953 -1523
rect 8928 -1548 8932 -1531
rect 8949 -1548 8953 -1531
rect 8928 -1557 8953 -1548
rect 8633 -1613 8638 -1596
rect 8655 -1613 8660 -1596
rect 8633 -1625 8660 -1613
rect 8690 -1595 8711 -1587
rect 8690 -1612 8692 -1595
rect 8709 -1612 8711 -1595
rect 8690 -1620 8711 -1612
rect 8734 -1595 8755 -1587
rect 8734 -1612 8736 -1595
rect 8753 -1612 8755 -1595
rect 8734 -1620 8755 -1612
rect 8778 -1595 8799 -1587
rect 8778 -1612 8780 -1595
rect 8797 -1612 8799 -1595
rect 8778 -1620 8799 -1612
rect 8822 -1595 8843 -1587
rect 8822 -1612 8824 -1595
rect 8841 -1612 8843 -1595
rect 8822 -1620 8843 -1612
rect 8866 -1595 8887 -1587
rect 8866 -1612 8868 -1595
rect 8885 -1612 8887 -1595
rect 8866 -1620 8887 -1612
rect 8910 -1595 8931 -1587
rect 8910 -1612 8912 -1595
rect 8929 -1612 8931 -1595
rect 8910 -1620 8931 -1612
rect 8954 -1595 8975 -1587
rect 8954 -1612 8956 -1595
rect 8973 -1612 8975 -1595
rect 8954 -1620 8975 -1612
rect 3766 -1784 3849 -1767
rect 8692 -1765 8709 -1620
rect 8736 -1765 8753 -1620
rect 8780 -1765 8797 -1620
rect 8824 -1765 8841 -1620
rect 8868 -1765 8885 -1620
rect 8912 -1765 8929 -1620
rect 8954 -1765 8971 -1620
rect 8988 -1653 9013 -1645
rect 8988 -1670 8992 -1653
rect 9009 -1670 9013 -1653
rect 8988 -1679 9013 -1670
rect 8988 -1709 9013 -1701
rect 8988 -1726 8992 -1709
rect 9009 -1726 9013 -1709
rect 8988 -1735 9013 -1726
rect 8690 -1773 8711 -1765
rect 8690 -1778 8692 -1773
rect 8552 -1790 8692 -1778
rect 8709 -1790 8711 -1773
rect 8552 -1795 8711 -1790
rect 4912 -1830 4926 -1829
rect 4912 -1940 4929 -1830
rect 5230 -1879 5247 -1829
rect 5230 -1898 5247 -1896
rect 5340 -1940 5357 -1813
rect 8552 -1976 8569 -1795
rect 8690 -1798 8711 -1795
rect 8734 -1772 8755 -1765
rect 8734 -1790 8735 -1772
rect 8753 -1790 8755 -1772
rect 8734 -1798 8755 -1790
rect 8778 -1773 8799 -1765
rect 8778 -1790 8780 -1773
rect 8797 -1790 8799 -1773
rect 8778 -1798 8799 -1790
rect 8822 -1773 8843 -1765
rect 8822 -1790 8824 -1773
rect 8841 -1790 8843 -1773
rect 8822 -1798 8843 -1790
rect 8866 -1773 8887 -1765
rect 8866 -1790 8868 -1773
rect 8885 -1790 8887 -1773
rect 8866 -1798 8887 -1790
rect 8910 -1773 8931 -1765
rect 8910 -1790 8912 -1773
rect 8929 -1790 8931 -1773
rect 8910 -1798 8931 -1790
rect 8954 -1773 8975 -1765
rect 8954 -1790 8956 -1773
rect 8973 -1790 8975 -1773
rect 8954 -1798 8975 -1790
rect 8780 -1976 8797 -1798
rect 8884 -1831 8909 -1823
rect 8884 -1848 8888 -1831
rect 8905 -1848 8909 -1831
rect 8884 -1857 8909 -1848
rect 8821 -1879 8848 -1866
rect 8821 -1896 8826 -1879
rect 8843 -1896 8848 -1879
rect 8821 -1908 8848 -1896
rect 8958 -1940 8975 -1798
rect 8546 -1983 8576 -1976
rect 8546 -2001 8552 -1983
rect 8570 -2001 8576 -1983
rect 8546 -2008 8576 -2001
rect 8774 -1983 8804 -1976
rect 8774 -2001 8780 -1983
rect 8798 -2001 8804 -1983
rect 8774 -2008 8804 -2001
rect 3620 -2031 3637 -2020
<< viali >>
rect 3776 -1281 3793 -1264
rect 2804 -1344 2822 -1326
rect 2740 -1548 2757 -1531
rect 3660 -1362 3677 -1345
rect 3616 -1402 3633 -1385
rect 3035 -1443 3052 -1426
rect 2980 -1503 2997 -1486
rect 3832 -1322 3849 -1305
rect 2760 -1612 2777 -1595
rect 2680 -1670 2697 -1653
rect 2680 -1726 2697 -1709
rect 3620 -1635 3637 -1618
rect 3728 -1632 3745 -1615
rect 2848 -1790 2865 -1773
rect 2936 -1773 2954 -1772
rect 2936 -1790 2953 -1773
rect 2953 -1790 2954 -1773
rect 2784 -1848 2801 -1831
rect 2846 -1896 2863 -1879
rect 2717 -1959 2734 -1942
rect 2891 -2001 2909 -1983
rect 3119 -2001 3137 -1983
rect 8867 -1344 8885 -1326
rect 5221 -1445 5238 -1428
rect 8637 -1443 8654 -1426
rect 5104 -1590 5121 -1573
rect 4999 -1632 5016 -1615
rect 8692 -1503 8709 -1486
rect 8932 -1548 8949 -1531
rect 8912 -1612 8929 -1595
rect 5019 -1776 5036 -1759
rect 8992 -1670 9009 -1653
rect 8992 -1726 9009 -1709
rect 5066 -1813 5083 -1796
rect 5340 -1813 5357 -1796
rect 5230 -1896 5247 -1879
rect 4912 -1957 4929 -1940
rect 5340 -1957 5357 -1940
rect 8735 -1773 8753 -1772
rect 8735 -1790 8736 -1773
rect 8736 -1790 8753 -1773
rect 8824 -1790 8841 -1773
rect 8888 -1848 8905 -1831
rect 8826 -1896 8843 -1879
rect 8958 -1957 8975 -1940
rect 3620 -2020 3637 -2003
rect 8552 -2001 8570 -1983
rect 8780 -2001 8798 -1983
<< metal1 >>
rect 5766 -1258 5792 -1255
rect 3768 -1264 3803 -1261
rect 3768 -1265 3776 -1264
rect 3765 -1279 3776 -1265
rect 3768 -1281 3776 -1279
rect 3793 -1265 3803 -1264
rect 3793 -1279 5766 -1265
rect 3793 -1281 3803 -1279
rect 3768 -1284 3803 -1281
rect 5766 -1287 5792 -1284
rect 5836 -1291 5862 -1288
rect 3828 -1305 3852 -1301
rect 3825 -1319 3832 -1305
rect 2798 -1322 2828 -1319
rect 2798 -1348 2800 -1322
rect 2826 -1348 2828 -1322
rect 3828 -1322 3832 -1319
rect 3849 -1317 5836 -1305
rect 3849 -1319 5862 -1317
rect 3849 -1322 3852 -1319
rect 5836 -1320 5862 -1319
rect 3828 -1328 3852 -1322
rect 8861 -1322 8891 -1319
rect 5800 -1337 5826 -1334
rect 3656 -1345 3680 -1341
rect 2798 -1351 2828 -1348
rect 3654 -1359 3660 -1345
rect 3656 -1362 3660 -1359
rect 3677 -1359 5800 -1345
rect 3677 -1362 3680 -1359
rect 3656 -1368 3680 -1362
rect 8861 -1348 8863 -1322
rect 8889 -1348 8891 -1322
rect 8861 -1351 8891 -1348
rect 5800 -1366 5826 -1363
rect 5729 -1378 5755 -1375
rect 3613 -1385 3636 -1382
rect 3609 -1399 3616 -1385
rect 3613 -1402 3616 -1399
rect 3633 -1399 5729 -1385
rect 3633 -1402 3636 -1399
rect 3613 -1408 3636 -1402
rect 5729 -1407 5755 -1404
rect 5625 -1420 5651 -1417
rect 3029 -1426 3056 -1423
rect 5218 -1426 5242 -1424
rect 3029 -1443 3035 -1426
rect 3052 -1428 5625 -1426
rect 3052 -1443 5221 -1428
rect 3029 -1445 5221 -1443
rect 5238 -1445 5625 -1428
rect 3029 -1446 5625 -1445
rect 8633 -1426 8660 -1423
rect 5651 -1443 8637 -1426
rect 8654 -1443 8660 -1426
rect 5651 -1446 8660 -1443
rect 5218 -1448 5242 -1446
rect 5625 -1449 5651 -1446
rect 2977 -1486 3000 -1480
rect 8689 -1486 8712 -1480
rect 2977 -1503 2980 -1486
rect 2997 -1500 3062 -1486
rect 8631 -1500 8692 -1486
rect 2997 -1503 3000 -1500
rect 2977 -1509 3000 -1503
rect 8689 -1503 8692 -1500
rect 8709 -1503 8712 -1486
rect 8689 -1509 8712 -1503
rect 5906 -1523 5932 -1520
rect 2734 -1531 2763 -1526
rect 2734 -1548 2740 -1531
rect 2757 -1532 2763 -1531
rect 2757 -1546 5906 -1532
rect 2757 -1548 2763 -1546
rect 2734 -1552 2763 -1548
rect 8926 -1531 8955 -1526
rect 8926 -1532 8932 -1531
rect 5932 -1546 8932 -1532
rect 5906 -1552 5932 -1549
rect 8926 -1548 8932 -1546
rect 8949 -1548 8955 -1531
rect 8926 -1552 8955 -1548
rect 5661 -1568 5687 -1565
rect 5098 -1573 5127 -1570
rect 2636 -1587 2679 -1578
rect 2636 -1613 2641 -1587
rect 2667 -1591 2679 -1587
rect 5098 -1590 5104 -1573
rect 5121 -1575 5127 -1573
rect 5121 -1589 5661 -1575
rect 5121 -1590 5127 -1589
rect 2757 -1591 2783 -1590
rect 2667 -1595 2783 -1591
rect 5098 -1593 5127 -1590
rect 2667 -1612 2760 -1595
rect 2777 -1612 2783 -1595
rect 9010 -1587 9053 -1578
rect 5661 -1597 5687 -1594
rect 8906 -1591 8932 -1590
rect 9010 -1591 9022 -1587
rect 8906 -1595 9022 -1591
rect 6011 -1601 6037 -1598
rect 2667 -1613 2783 -1612
rect 2636 -1615 2783 -1613
rect 3725 -1615 3748 -1608
rect 2639 -1616 2669 -1615
rect 2757 -1616 2783 -1615
rect 3614 -1618 3643 -1615
rect 3725 -1618 3728 -1615
rect 3614 -1635 3620 -1618
rect 3637 -1632 3728 -1618
rect 3745 -1632 3748 -1615
rect 3637 -1635 3643 -1632
rect 3614 -1638 3643 -1635
rect 3725 -1638 3748 -1632
rect 4995 -1615 5020 -1607
rect 4995 -1632 4999 -1615
rect 5016 -1616 5020 -1615
rect 5016 -1627 6011 -1616
rect 8906 -1612 8912 -1595
rect 8929 -1612 9022 -1595
rect 8906 -1613 9022 -1612
rect 9048 -1613 9053 -1587
rect 8906 -1615 9053 -1613
rect 8906 -1616 8932 -1615
rect 9020 -1616 9050 -1615
rect 5016 -1630 6037 -1627
rect 5016 -1632 5020 -1630
rect 4995 -1639 5020 -1632
rect 5975 -1648 6001 -1645
rect 2674 -1653 2703 -1649
rect 2674 -1670 2680 -1653
rect 2697 -1654 2703 -1653
rect 2697 -1668 5975 -1654
rect 2697 -1670 2703 -1668
rect 2674 -1675 2703 -1670
rect 8986 -1653 9015 -1649
rect 8986 -1654 8992 -1653
rect 6001 -1668 8992 -1654
rect 5975 -1677 6001 -1674
rect 8986 -1670 8992 -1668
rect 9009 -1670 9015 -1653
rect 8986 -1675 9015 -1670
rect 5871 -1702 5897 -1699
rect 2674 -1709 2703 -1706
rect 2674 -1726 2680 -1709
rect 2697 -1710 2703 -1709
rect 2697 -1724 5871 -1710
rect 2697 -1726 2703 -1724
rect 2674 -1732 2703 -1726
rect 8986 -1709 9015 -1706
rect 8986 -1710 8992 -1709
rect 5897 -1724 8992 -1710
rect 5871 -1731 5897 -1728
rect 8986 -1726 8992 -1724
rect 9009 -1726 9015 -1709
rect 8986 -1732 9015 -1726
rect 5696 -1753 5722 -1750
rect 5013 -1759 5042 -1754
rect 3172 -1766 3202 -1763
rect 2845 -1771 2871 -1769
rect 2636 -1773 2871 -1771
rect 2636 -1780 2848 -1773
rect 2636 -1806 2641 -1780
rect 2667 -1790 2848 -1780
rect 2865 -1790 2871 -1773
rect 2667 -1792 2871 -1790
rect 2667 -1806 2672 -1792
rect 2845 -1794 2871 -1792
rect 2930 -1771 2959 -1769
rect 3172 -1771 3174 -1766
rect 2930 -1772 3174 -1771
rect 2930 -1790 2936 -1772
rect 2954 -1790 3174 -1772
rect 2930 -1792 3174 -1790
rect 3200 -1771 3202 -1766
rect 3200 -1792 3205 -1771
rect 5013 -1776 5019 -1759
rect 5036 -1762 5042 -1759
rect 5036 -1776 5696 -1762
rect 5013 -1780 5042 -1776
rect 8487 -1766 8517 -1763
rect 8487 -1771 8489 -1766
rect 5696 -1782 5722 -1779
rect 2930 -1793 2959 -1792
rect 3172 -1795 3202 -1792
rect 5060 -1796 5089 -1790
rect 8484 -1792 8489 -1771
rect 8515 -1771 8517 -1766
rect 8730 -1771 8759 -1769
rect 8515 -1772 8759 -1771
rect 8515 -1790 8735 -1772
rect 8753 -1790 8759 -1772
rect 8515 -1792 8759 -1790
rect 5337 -1796 5361 -1793
rect 8487 -1795 8517 -1792
rect 8730 -1793 8759 -1792
rect 8818 -1771 8844 -1769
rect 8818 -1773 9053 -1771
rect 8818 -1790 8824 -1773
rect 8841 -1780 9053 -1773
rect 8841 -1790 9022 -1780
rect 8818 -1792 9022 -1790
rect 8818 -1794 8844 -1792
rect 2639 -1809 2669 -1806
rect 5060 -1813 5066 -1796
rect 5083 -1798 5089 -1796
rect 5334 -1798 5340 -1796
rect 5083 -1812 5340 -1798
rect 5083 -1813 5089 -1812
rect 5334 -1813 5340 -1812
rect 5357 -1813 5363 -1796
rect 9017 -1806 9022 -1792
rect 9048 -1806 9053 -1780
rect 9020 -1809 9050 -1806
rect 5060 -1817 5089 -1813
rect 5337 -1816 5361 -1813
rect 5940 -1823 5966 -1820
rect 2778 -1831 2807 -1826
rect 2778 -1848 2784 -1831
rect 2801 -1832 2807 -1831
rect 2801 -1846 5940 -1832
rect 2801 -1848 2807 -1846
rect 2778 -1852 2807 -1848
rect 8882 -1831 8911 -1826
rect 8882 -1832 8888 -1831
rect 5966 -1846 8888 -1832
rect 5940 -1852 5966 -1849
rect 8882 -1848 8888 -1846
rect 8905 -1848 8911 -1831
rect 8882 -1852 8911 -1848
rect 6047 -1875 6073 -1872
rect -2059 -1895 -1892 -1877
rect 2843 -1878 2866 -1876
rect 5227 -1878 5250 -1875
rect -2059 -1954 -2005 -1895
rect -1940 -1954 -1892 -1895
rect 2840 -1879 6047 -1878
rect 2840 -1896 2846 -1879
rect 2863 -1896 5230 -1879
rect 5247 -1896 6047 -1879
rect 2840 -1898 6047 -1896
rect 2843 -1899 2866 -1898
rect 5227 -1901 5250 -1898
rect 8823 -1878 8846 -1876
rect 6073 -1879 8853 -1878
rect 6073 -1896 8826 -1879
rect 8843 -1896 8853 -1879
rect 6073 -1898 8853 -1896
rect 13581 -1895 13748 -1877
rect 8823 -1899 8846 -1898
rect 6047 -1904 6073 -1901
rect 2714 -1942 2737 -1939
rect 4909 -1940 4932 -1934
rect 5334 -1940 5360 -1937
rect 8955 -1940 8978 -1937
rect -2059 -1984 -1892 -1954
rect 2710 -1959 2717 -1942
rect 2734 -1943 2740 -1942
rect 4909 -1943 4912 -1940
rect 2734 -1957 4912 -1943
rect 4929 -1957 4935 -1940
rect 2734 -1959 2740 -1957
rect 2714 -1962 2737 -1959
rect 4909 -1960 4935 -1957
rect 5334 -1957 5340 -1940
rect 5357 -1943 5363 -1940
rect 8952 -1943 8958 -1940
rect 5357 -1957 8958 -1943
rect 8975 -1957 8981 -1940
rect 13581 -1954 13629 -1895
rect 13694 -1954 13748 -1895
rect 5334 -1960 5360 -1957
rect 8955 -1960 8978 -1957
rect 4909 -1961 4932 -1960
rect 2885 -1979 2915 -1976
rect 2885 -2005 2887 -1979
rect 2913 -2005 2915 -1979
rect 2885 -2008 2915 -2005
rect 3113 -1979 3143 -1976
rect 3113 -2005 3115 -1979
rect 3141 -2005 3143 -1979
rect 8546 -1979 8576 -1976
rect 3113 -2008 3143 -2005
rect 3614 -1998 3642 -1995
rect 3614 -2024 3616 -1998
rect 8546 -2005 8548 -1979
rect 8574 -2005 8576 -1979
rect 8546 -2008 8576 -2005
rect 8774 -1979 8804 -1976
rect 8774 -2005 8776 -1979
rect 8802 -2005 8804 -1979
rect 13581 -1984 13748 -1954
rect 8774 -2008 8804 -2005
rect 3614 -2028 3642 -2024
<< via1 >>
rect 5766 -1284 5792 -1258
rect 2800 -1326 2826 -1322
rect 2800 -1344 2804 -1326
rect 2804 -1344 2822 -1326
rect 2822 -1344 2826 -1326
rect 2800 -1348 2826 -1344
rect 5836 -1317 5862 -1291
rect 5800 -1363 5826 -1337
rect 8863 -1326 8889 -1322
rect 8863 -1344 8867 -1326
rect 8867 -1344 8885 -1326
rect 8885 -1344 8889 -1326
rect 8863 -1348 8889 -1344
rect 5729 -1404 5755 -1378
rect 5625 -1446 5651 -1420
rect 5906 -1549 5932 -1523
rect 2641 -1613 2667 -1587
rect 5661 -1594 5687 -1568
rect 6011 -1627 6037 -1601
rect 9022 -1613 9048 -1587
rect 5975 -1674 6001 -1648
rect 5871 -1728 5897 -1702
rect 2641 -1806 2667 -1780
rect 3174 -1792 3200 -1766
rect 5696 -1779 5722 -1753
rect 8489 -1792 8515 -1766
rect 9022 -1806 9048 -1780
rect 5940 -1849 5966 -1823
rect -2005 -1954 -1940 -1895
rect 6047 -1901 6073 -1875
rect 13629 -1954 13694 -1895
rect 2887 -1983 2913 -1979
rect 2887 -2001 2891 -1983
rect 2891 -2001 2909 -1983
rect 2909 -2001 2913 -1983
rect 2887 -2005 2913 -2001
rect 3115 -1983 3141 -1979
rect 3115 -2001 3119 -1983
rect 3119 -2001 3137 -1983
rect 3137 -2001 3141 -1983
rect 3115 -2005 3141 -2001
rect 3616 -2003 3642 -1998
rect 3616 -2020 3620 -2003
rect 3620 -2020 3637 -2003
rect 3637 -2020 3642 -2003
rect 8548 -1983 8574 -1979
rect 8548 -2001 8552 -1983
rect 8552 -2001 8570 -1983
rect 8570 -2001 8574 -1983
rect 8548 -2005 8574 -2001
rect 8776 -1983 8802 -1979
rect 8776 -2001 8780 -1983
rect 8780 -2001 8798 -1983
rect 8798 -2001 8802 -1983
rect 8776 -2005 8802 -2001
rect 3616 -2024 3642 -2020
<< metal2 >>
rect 2795 -1321 2831 -1316
rect 2795 -1349 2799 -1321
rect 2827 -1349 2831 -1321
rect 2795 -1354 2831 -1349
rect 5631 -1417 5645 2887
rect 5625 -1420 5651 -1417
rect 5625 -1449 5651 -1446
rect 2636 -1586 2672 -1581
rect 2636 -1614 2640 -1586
rect 2668 -1614 2672 -1586
rect 2636 -1619 2672 -1614
rect 3169 -1765 3205 -1760
rect 2636 -1779 2672 -1774
rect 2636 -1807 2640 -1779
rect 2668 -1807 2672 -1779
rect 3169 -1793 3173 -1765
rect 3201 -1793 3205 -1765
rect 3169 -1798 3205 -1793
rect 2636 -1812 2672 -1807
rect -2011 -1895 -1934 -1888
rect -2011 -1954 -2005 -1895
rect -1940 -1954 -1934 -1895
rect -2011 -1961 -1934 -1954
rect 2882 -1978 2918 -1973
rect 2882 -2006 2886 -1978
rect 2914 -2006 2918 -1978
rect 2882 -2011 2918 -2006
rect 3110 -1978 3146 -1973
rect 3110 -2006 3114 -1978
rect 3142 -2006 3146 -1978
rect 3110 -2011 3146 -2006
rect 3613 -1997 3645 -1992
rect 3613 -2025 3615 -1997
rect 3643 -2025 3645 -1997
rect 3613 -2030 3645 -2025
rect 5631 -5158 5645 -1449
rect 5666 -1565 5680 2887
rect 5661 -1568 5687 -1565
rect 5661 -1597 5687 -1594
rect 5666 -5158 5680 -1597
rect 5701 -1750 5715 2887
rect 5736 -1375 5750 2887
rect 5771 -1255 5785 2887
rect 5766 -1258 5792 -1255
rect 5766 -1287 5792 -1284
rect 5729 -1378 5755 -1375
rect 5729 -1407 5755 -1404
rect 5696 -1753 5722 -1750
rect 5696 -1782 5722 -1779
rect 5701 -5158 5715 -1782
rect 5736 -5158 5750 -1407
rect 5771 -5158 5785 -1287
rect 5806 -1334 5820 2887
rect 5841 -1288 5855 2887
rect 5836 -1291 5862 -1288
rect 5836 -1320 5862 -1317
rect 5800 -1337 5826 -1334
rect 5800 -1366 5826 -1363
rect 5806 -5158 5820 -1366
rect 5841 -5158 5855 -1320
rect 5876 -1699 5890 2887
rect 5911 -1520 5925 2887
rect 5906 -1523 5932 -1520
rect 5906 -1552 5932 -1549
rect 5871 -1702 5897 -1699
rect 5871 -1731 5897 -1728
rect 5876 -5158 5890 -1731
rect 5911 -5158 5925 -1552
rect 5946 -1820 5960 2887
rect 5981 -1645 5995 2887
rect 6016 -1598 6030 2887
rect 6011 -1601 6037 -1598
rect 6011 -1630 6037 -1627
rect 5975 -1648 6001 -1645
rect 5975 -1677 6001 -1674
rect 5940 -1823 5966 -1820
rect 5940 -1852 5966 -1849
rect 5946 -5158 5960 -1852
rect 5981 -5158 5995 -1677
rect 6016 -5158 6030 -1630
rect 6051 -1872 6065 2887
rect 8858 -1321 8894 -1316
rect 8858 -1349 8862 -1321
rect 8890 -1349 8894 -1321
rect 8858 -1354 8894 -1349
rect 9017 -1586 9053 -1581
rect 9017 -1614 9021 -1586
rect 9049 -1614 9053 -1586
rect 9017 -1619 9053 -1614
rect 8484 -1765 8520 -1760
rect 8484 -1793 8488 -1765
rect 8516 -1793 8520 -1765
rect 8484 -1798 8520 -1793
rect 9017 -1779 9053 -1774
rect 9017 -1807 9021 -1779
rect 9049 -1807 9053 -1779
rect 9017 -1812 9053 -1807
rect 6047 -1875 6073 -1872
rect 6047 -1904 6073 -1901
rect 13623 -1895 13700 -1888
rect 6051 -5158 6065 -1904
rect 13623 -1954 13629 -1895
rect 13694 -1954 13700 -1895
rect 13623 -1961 13700 -1954
rect 8543 -1978 8579 -1973
rect 8543 -2006 8547 -1978
rect 8575 -2006 8579 -1978
rect 8543 -2011 8579 -2006
rect 8771 -1978 8807 -1973
rect 8771 -2006 8775 -1978
rect 8803 -2006 8807 -1978
rect 8771 -2011 8807 -2006
<< via2 >>
rect 2799 -1322 2827 -1321
rect 2799 -1348 2800 -1322
rect 2800 -1348 2826 -1322
rect 2826 -1348 2827 -1322
rect 2799 -1349 2827 -1348
rect 2640 -1587 2668 -1586
rect 2640 -1613 2641 -1587
rect 2641 -1613 2667 -1587
rect 2667 -1613 2668 -1587
rect 2640 -1614 2668 -1613
rect 2640 -1780 2668 -1779
rect 2640 -1806 2641 -1780
rect 2641 -1806 2667 -1780
rect 2667 -1806 2668 -1780
rect 2640 -1807 2668 -1806
rect 3173 -1766 3201 -1765
rect 3173 -1792 3174 -1766
rect 3174 -1792 3200 -1766
rect 3200 -1792 3201 -1766
rect 3173 -1793 3201 -1792
rect -2005 -1954 -1940 -1895
rect 2886 -1979 2914 -1978
rect 2886 -2005 2887 -1979
rect 2887 -2005 2913 -1979
rect 2913 -2005 2914 -1979
rect 2886 -2006 2914 -2005
rect 3114 -1979 3142 -1978
rect 3114 -2005 3115 -1979
rect 3115 -2005 3141 -1979
rect 3141 -2005 3142 -1979
rect 3114 -2006 3142 -2005
rect 3615 -1998 3643 -1997
rect 3615 -2024 3616 -1998
rect 3616 -2024 3642 -1998
rect 3642 -2024 3643 -1998
rect 3615 -2025 3643 -2024
rect 8862 -1322 8890 -1321
rect 8862 -1348 8863 -1322
rect 8863 -1348 8889 -1322
rect 8889 -1348 8890 -1322
rect 8862 -1349 8890 -1348
rect 9021 -1587 9049 -1586
rect 9021 -1613 9022 -1587
rect 9022 -1613 9048 -1587
rect 9048 -1613 9049 -1587
rect 9021 -1614 9049 -1613
rect 8488 -1766 8516 -1765
rect 8488 -1792 8489 -1766
rect 8489 -1792 8515 -1766
rect 8515 -1792 8516 -1766
rect 8488 -1793 8516 -1792
rect 9021 -1780 9049 -1779
rect 9021 -1806 9022 -1780
rect 9022 -1806 9048 -1780
rect 9048 -1806 9049 -1780
rect 9021 -1807 9049 -1806
rect 13629 -1954 13694 -1895
rect 8547 -1979 8575 -1978
rect 8547 -2005 8548 -1979
rect 8548 -2005 8574 -1979
rect 8574 -2005 8575 -1979
rect 8547 -2006 8575 -2005
rect 8775 -1979 8803 -1978
rect 8775 -2005 8776 -1979
rect 8776 -2005 8802 -1979
rect 8802 -2005 8803 -1979
rect 8775 -2006 8803 -2005
<< metal3 >>
rect -2092 -1250 5604 2862
rect 6085 -1250 13781 2862
rect -2059 -1895 -1892 -1250
rect 2057 -1306 2090 -1250
rect 9599 -1306 9632 -1250
rect 2057 -1734 2585 -1306
rect 2788 -1319 2837 -1309
rect 2788 -1351 2797 -1319
rect 2829 -1351 2837 -1319
rect 2788 -1361 2837 -1351
rect 8852 -1319 8901 -1309
rect 8852 -1351 8860 -1319
rect 8892 -1351 8901 -1319
rect 8852 -1361 8901 -1351
rect 2630 -1584 2679 -1574
rect 2630 -1616 2638 -1584
rect 2670 -1616 2679 -1584
rect 2630 -1626 2679 -1616
rect 9010 -1584 9059 -1574
rect 9010 -1616 9019 -1584
rect 9051 -1616 9059 -1584
rect 9010 -1626 9059 -1616
rect 9104 -1734 9632 -1306
rect 3163 -1763 3212 -1753
rect 2630 -1777 2679 -1767
rect -2059 -1954 -2005 -1895
rect -1940 -1954 -1892 -1895
rect -2059 -2077 -1892 -1954
rect 2057 -2021 2585 -1793
rect 2630 -1809 2638 -1777
rect 2670 -1809 2679 -1777
rect 3163 -1795 3171 -1763
rect 3203 -1795 3212 -1763
rect 8477 -1763 8526 -1753
rect 3163 -1805 3212 -1795
rect 2630 -1819 2679 -1809
rect 2876 -1976 2925 -1966
rect 2876 -2008 2884 -1976
rect 2916 -2008 2925 -1976
rect 2876 -2018 2925 -2008
rect 3104 -1976 3153 -1966
rect 3104 -2008 3112 -1976
rect 3144 -2008 3153 -1976
rect 3104 -2018 3153 -2008
rect 3243 -2021 3521 -1793
rect 3602 -1995 3651 -1989
rect 2057 -2077 2090 -2021
rect 3602 -2027 3614 -1995
rect 3646 -2027 3651 -1995
rect 8168 -2021 8446 -1793
rect 8477 -1795 8486 -1763
rect 8518 -1795 8526 -1763
rect 8477 -1805 8526 -1795
rect 9010 -1777 9059 -1767
rect 9010 -1809 9019 -1777
rect 9051 -1809 9059 -1777
rect 9010 -1819 9059 -1809
rect 8536 -1976 8585 -1966
rect 8536 -2008 8545 -1976
rect 8577 -2008 8585 -1976
rect 8536 -2018 8585 -2008
rect 8764 -1976 8813 -1966
rect 8764 -2008 8773 -1976
rect 8805 -2008 8813 -1976
rect 8764 -2018 8813 -2008
rect 9104 -2021 9632 -1793
rect 3602 -2077 3651 -2027
rect 8413 -2077 8446 -2021
rect 9599 -2077 9632 -2021
rect 13581 -1895 13748 -1250
rect 13581 -1954 13629 -1895
rect 13694 -1954 13748 -1895
rect 13581 -2077 13748 -1954
rect -2093 -5105 3019 -2077
rect 3075 -5105 5604 -2077
rect 6085 -2675 8614 -2077
rect 8670 -2675 13782 -2077
rect 6085 -3034 13782 -2675
rect 6085 -5105 8614 -3034
rect 8670 -5105 13782 -3034
<< via3 >>
rect 2797 -1321 2829 -1319
rect 2797 -1349 2799 -1321
rect 2799 -1349 2827 -1321
rect 2827 -1349 2829 -1321
rect 2797 -1351 2829 -1349
rect 8860 -1321 8892 -1319
rect 8860 -1349 8862 -1321
rect 8862 -1349 8890 -1321
rect 8890 -1349 8892 -1321
rect 8860 -1351 8892 -1349
rect 2638 -1586 2670 -1584
rect 2638 -1614 2640 -1586
rect 2640 -1614 2668 -1586
rect 2668 -1614 2670 -1586
rect 2638 -1616 2670 -1614
rect 9019 -1586 9051 -1584
rect 9019 -1614 9021 -1586
rect 9021 -1614 9049 -1586
rect 9049 -1614 9051 -1586
rect 9019 -1616 9051 -1614
rect -2005 -1954 -1940 -1895
rect 2638 -1779 2670 -1777
rect 2638 -1807 2640 -1779
rect 2640 -1807 2668 -1779
rect 2668 -1807 2670 -1779
rect 2638 -1809 2670 -1807
rect 3171 -1765 3203 -1763
rect 3171 -1793 3173 -1765
rect 3173 -1793 3201 -1765
rect 3201 -1793 3203 -1765
rect 3171 -1795 3203 -1793
rect 2884 -1978 2916 -1976
rect 2884 -2006 2886 -1978
rect 2886 -2006 2914 -1978
rect 2914 -2006 2916 -1978
rect 2884 -2008 2916 -2006
rect 3112 -1978 3144 -1976
rect 3112 -2006 3114 -1978
rect 3114 -2006 3142 -1978
rect 3142 -2006 3144 -1978
rect 3112 -2008 3144 -2006
rect 3614 -1997 3646 -1995
rect 3614 -2025 3615 -1997
rect 3615 -2025 3643 -1997
rect 3643 -2025 3646 -1997
rect 3614 -2027 3646 -2025
rect 8486 -1765 8518 -1763
rect 8486 -1793 8488 -1765
rect 8488 -1793 8516 -1765
rect 8516 -1793 8518 -1765
rect 8486 -1795 8518 -1793
rect 9019 -1779 9051 -1777
rect 9019 -1807 9021 -1779
rect 9021 -1807 9049 -1779
rect 9049 -1807 9051 -1779
rect 9019 -1809 9051 -1807
rect 8545 -1978 8577 -1976
rect 8545 -2006 8547 -1978
rect 8547 -2006 8575 -1978
rect 8575 -2006 8577 -1978
rect 8545 -2008 8577 -2006
rect 8773 -1978 8805 -1976
rect 8773 -2006 8775 -1978
rect 8775 -2006 8803 -1978
rect 8803 -2006 8805 -1978
rect 8773 -2008 8805 -2006
rect 13629 -1954 13694 -1895
<< mimcap >>
rect -2078 1187 922 2848
rect -2078 1069 757 1187
rect 875 1069 922 1187
rect -2078 848 922 1069
rect 1006 1184 4006 2848
rect 1006 1066 1059 1184
rect 1177 1161 4006 1184
rect 1177 1066 3847 1161
rect 1006 1043 3847 1066
rect 3965 1043 4006 1161
rect 1006 848 4006 1043
rect 4090 1194 5590 2848
rect 4090 1076 4143 1194
rect 4261 1076 5590 1194
rect 4090 848 5590 1076
rect 6099 1194 7599 2848
rect 6099 1076 7428 1194
rect 7546 1076 7599 1194
rect 6099 848 7599 1076
rect 7683 1184 10683 2848
rect 7683 1161 10512 1184
rect 7683 1043 7724 1161
rect 7842 1066 10512 1161
rect 10630 1066 10683 1184
rect 7842 1043 10683 1066
rect 7683 848 10683 1043
rect 10767 1187 13767 2848
rect 10767 1069 10814 1187
rect 10932 1069 13767 1187
rect 10767 848 13767 1069
rect -2078 540 922 764
rect -2078 422 767 540
rect 885 422 922 540
rect -2078 -1071 922 422
rect -2078 -1189 -1858 -1071
rect -1740 -1189 922 -1071
rect -2078 -1236 922 -1189
rect 1006 547 4006 764
rect 1006 429 1040 547
rect 1158 505 4006 547
rect 1158 429 3825 505
rect 1006 387 3825 429
rect 3943 387 4006 505
rect 1006 -1236 4006 387
rect 4090 488 5590 764
rect 4090 370 4133 488
rect 4251 370 5590 488
rect 4090 -1236 5590 370
rect 6099 488 7599 764
rect 6099 370 7438 488
rect 7556 370 7599 488
rect 6099 -1236 7599 370
rect 7683 547 10683 764
rect 7683 505 10531 547
rect 7683 387 7746 505
rect 7864 429 10531 505
rect 10649 429 10683 547
rect 7864 387 10683 429
rect 7683 -1236 10683 387
rect 10767 540 13767 764
rect 10767 422 10804 540
rect 10922 422 13767 540
rect 10767 -1071 13767 422
rect 10767 -1189 13429 -1071
rect 13547 -1189 13767 -1071
rect 10767 -1236 13767 -1189
rect 2071 -1584 2571 -1320
rect 2071 -1618 2529 -1584
rect 2563 -1618 2571 -1584
rect 2071 -1720 2571 -1618
rect 9118 -1584 9618 -1320
rect 9118 -1618 9126 -1584
rect 9160 -1618 9618 -1584
rect 9118 -1720 9618 -1618
rect 2071 -1841 2571 -1807
rect 2071 -1875 2527 -1841
rect 2561 -1875 2571 -1841
rect 2071 -2007 2571 -1875
rect 3257 -1828 3507 -1807
rect 3257 -1860 3265 -1828
rect 3297 -1860 3507 -1828
rect 3257 -2007 3507 -1860
rect 8182 -1828 8432 -1807
rect 8182 -1860 8392 -1828
rect 8424 -1860 8432 -1828
rect 8182 -2007 8432 -1860
rect 9118 -1841 9618 -1807
rect 9118 -1875 9128 -1841
rect 9162 -1875 9618 -1841
rect 9118 -2007 9618 -1875
rect -2079 -2144 421 -2091
rect -2079 -2262 -1843 -2144
rect -1725 -2262 421 -2144
rect -2079 -5091 421 -2262
rect 505 -2127 3005 -2091
rect 505 -2245 725 -2127
rect 843 -2245 3005 -2127
rect 505 -5091 3005 -2245
rect 3089 -2144 5590 -2091
rect 3089 -2262 3327 -2144
rect 3445 -2262 5590 -2144
rect 3089 -5091 5590 -2262
rect 6099 -2144 8600 -2091
rect 6099 -2262 8244 -2144
rect 8362 -2262 8600 -2144
rect 6099 -5091 8600 -2262
rect 8684 -2127 11184 -2091
rect 8684 -2245 10846 -2127
rect 10964 -2245 11184 -2127
rect 8684 -5091 11184 -2245
rect 11268 -2144 13768 -2091
rect 11268 -2262 13414 -2144
rect 13532 -2262 13768 -2144
rect 11268 -5091 13768 -2262
<< mimcapcontact >>
rect 757 1069 875 1187
rect 1059 1066 1177 1184
rect 3847 1043 3965 1161
rect 4143 1076 4261 1194
rect 7428 1076 7546 1194
rect 7724 1043 7842 1161
rect 10512 1066 10630 1184
rect 10814 1069 10932 1187
rect 767 422 885 540
rect -1858 -1189 -1740 -1071
rect 1040 429 1158 547
rect 3825 387 3943 505
rect 4133 370 4251 488
rect 7438 370 7556 488
rect 7746 387 7864 505
rect 10531 429 10649 547
rect 10804 422 10922 540
rect 13429 -1189 13547 -1071
rect 2529 -1618 2563 -1584
rect 9126 -1618 9160 -1584
rect 2527 -1875 2561 -1841
rect 3265 -1860 3297 -1828
rect 8392 -1860 8424 -1828
rect 9128 -1875 9162 -1841
rect -1843 -2262 -1725 -2144
rect 725 -2245 843 -2127
rect 3327 -2262 3445 -2144
rect 8244 -2262 8362 -2144
rect 10846 -2245 10964 -2127
rect 13414 -2262 13532 -2144
<< metal4 >>
rect -2092 1194 5604 2862
rect -2092 1187 4143 1194
rect -2092 1069 757 1187
rect 875 1184 4143 1187
rect 875 1069 1059 1184
rect -2092 1066 1059 1069
rect 1177 1161 4143 1184
rect 1177 1066 3847 1161
rect -2092 1043 3847 1066
rect 3965 1076 4143 1161
rect 4261 1076 5604 1194
rect 3965 1043 5604 1076
rect -2092 547 5604 1043
rect -2092 540 1040 547
rect -2092 422 767 540
rect 885 429 1040 540
rect 1158 505 5604 547
rect 1158 429 3825 505
rect 885 422 3825 429
rect -2092 387 3825 422
rect 3943 488 5604 505
rect 3943 387 4133 488
rect -2092 370 4133 387
rect 4251 370 5604 488
rect -2092 -1071 5604 370
rect -2092 -1189 -1858 -1071
rect -1740 -1189 5604 -1071
rect -2092 -1250 5604 -1189
rect 6085 1194 13781 2862
rect 6085 1076 7428 1194
rect 7546 1187 13781 1194
rect 7546 1184 10814 1187
rect 7546 1161 10512 1184
rect 7546 1076 7724 1161
rect 6085 1043 7724 1076
rect 7842 1066 10512 1161
rect 10630 1069 10814 1184
rect 10932 1069 13781 1187
rect 10630 1066 13781 1069
rect 7842 1043 13781 1066
rect 6085 547 13781 1043
rect 6085 505 10531 547
rect 6085 488 7746 505
rect 6085 370 7438 488
rect 7556 387 7746 488
rect 7864 429 10531 505
rect 10649 540 13781 547
rect 10649 429 10804 540
rect 7864 422 10804 429
rect 10922 422 13781 540
rect 7864 387 13781 422
rect 7556 370 13781 387
rect 6085 -1071 13781 370
rect 6085 -1189 13429 -1071
rect 13547 -1189 13781 -1071
rect 6085 -1250 13781 -1189
rect 2798 -1315 2828 -1250
rect 8861 -1315 8891 -1250
rect 2796 -1319 2830 -1315
rect 2796 -1351 2797 -1319
rect 2829 -1351 2830 -1319
rect 2796 -1352 2830 -1351
rect 8859 -1319 8893 -1315
rect 8859 -1351 8860 -1319
rect 8892 -1351 8893 -1319
rect 8859 -1352 8893 -1351
rect 2528 -1584 2671 -1583
rect 2528 -1618 2529 -1584
rect 2563 -1616 2638 -1584
rect 2670 -1616 2671 -1584
rect 2563 -1618 2671 -1616
rect 2528 -1619 2671 -1618
rect 9018 -1584 9161 -1583
rect 9018 -1616 9019 -1584
rect 9051 -1616 9126 -1584
rect 9018 -1618 9126 -1616
rect 9160 -1618 9161 -1584
rect 9018 -1619 9161 -1618
rect 3170 -1763 3204 -1762
rect 2637 -1777 2671 -1776
rect 2637 -1809 2638 -1777
rect 2670 -1809 2671 -1777
rect 3170 -1795 3171 -1763
rect 3203 -1795 3204 -1763
rect 3170 -1799 3204 -1795
rect 8485 -1763 8519 -1762
rect 8485 -1795 8486 -1763
rect 8518 -1795 8519 -1763
rect 8485 -1799 8519 -1795
rect 9018 -1777 9052 -1776
rect 2637 -1813 2671 -1809
rect 2526 -1841 2562 -1840
rect 2526 -1875 2527 -1841
rect 2561 -1843 2562 -1841
rect 2639 -1843 2669 -1813
rect 2561 -1873 2669 -1843
rect 3172 -1829 3202 -1799
rect 3262 -1828 3298 -1827
rect 3262 -1829 3265 -1828
rect 3172 -1859 3265 -1829
rect 3262 -1860 3265 -1859
rect 3297 -1860 3298 -1828
rect 3262 -1861 3298 -1860
rect 8391 -1828 8427 -1827
rect 8391 -1860 8392 -1828
rect 8424 -1829 8427 -1828
rect 8487 -1829 8517 -1799
rect 9018 -1809 9019 -1777
rect 9051 -1809 9052 -1777
rect 9018 -1813 9052 -1809
rect 8424 -1859 8517 -1829
rect 9020 -1843 9050 -1813
rect 9127 -1841 9163 -1840
rect 9127 -1843 9128 -1841
rect 8424 -1860 8427 -1859
rect 8391 -1861 8427 -1860
rect 9020 -1873 9128 -1843
rect 2561 -1875 2562 -1873
rect 2526 -1876 2562 -1875
rect 9127 -1875 9128 -1873
rect 9162 -1875 9163 -1841
rect 9127 -1876 9163 -1875
rect 2883 -1976 2917 -1975
rect 2883 -2008 2884 -1976
rect 2916 -2008 2917 -1976
rect 2883 -2012 2917 -2008
rect 3111 -1976 3145 -1975
rect 3111 -2008 3112 -1976
rect 3144 -2008 3145 -1976
rect 3111 -2012 3145 -2008
rect 2885 -2077 2915 -2012
rect 3113 -2077 3143 -2012
rect 8544 -1976 8578 -1975
rect 8544 -2008 8545 -1976
rect 8577 -2008 8578 -1976
rect 8544 -2012 8578 -2008
rect 8772 -1976 8806 -1975
rect 8772 -2008 8773 -1976
rect 8805 -2008 8806 -1976
rect 8772 -2012 8806 -2008
rect 8546 -2077 8576 -2012
rect 8774 -2077 8804 -2012
rect -2093 -2127 3019 -2077
rect -2093 -2144 725 -2127
rect -2093 -2262 -1843 -2144
rect -1725 -2245 725 -2144
rect 843 -2245 3019 -2127
rect -1725 -2262 3019 -2245
rect -2093 -5105 3019 -2262
rect 3075 -2144 5604 -2077
rect 3075 -2262 3327 -2144
rect 3445 -2262 5604 -2144
rect 3075 -5105 5604 -2262
rect 6085 -2144 8614 -2077
rect 6085 -2262 8244 -2144
rect 8362 -2262 8614 -2144
rect 6085 -5105 8614 -2262
rect 8670 -2127 13782 -2077
rect 8670 -2245 10846 -2127
rect 10964 -2144 13782 -2127
rect 10964 -2245 13414 -2144
rect 8670 -2262 13414 -2245
rect 13532 -2262 13782 -2144
rect 8670 -5105 13782 -2262
<< via4 >>
rect -2030 -1895 -1908 -1853
rect -2030 -1954 -2005 -1895
rect -2005 -1954 -1940 -1895
rect -1940 -1954 -1908 -1895
rect 13597 -1895 13719 -1853
rect -2030 -1976 -1908 -1954
rect 3570 -1995 3689 -1919
rect 13597 -1954 13629 -1895
rect 13629 -1954 13694 -1895
rect 13694 -1954 13719 -1895
rect 3570 -2027 3614 -1995
rect 3614 -2027 3646 -1995
rect 3646 -2027 3689 -1995
rect 13597 -1976 13719 -1954
rect 3570 -2037 3689 -2027
<< mimcap2 >>
rect -2078 1003 922 2848
rect -2078 885 763 1003
rect 881 885 922 1003
rect -2078 848 922 885
rect 1006 1005 4006 2848
rect 1006 887 1047 1005
rect 1165 987 4006 1005
rect 1165 887 3833 987
rect 1006 869 3833 887
rect 3951 869 4006 987
rect 1006 848 4006 869
rect 4090 992 5590 2848
rect 4090 874 4124 992
rect 4242 874 5590 992
rect 4090 848 5590 874
rect 6099 992 7599 2848
rect 6099 874 7447 992
rect 7565 874 7599 992
rect 6099 848 7599 874
rect 7683 1005 10683 2848
rect 7683 987 10524 1005
rect 7683 869 7738 987
rect 7856 887 10524 987
rect 10642 887 10683 1005
rect 7856 869 10683 887
rect 7683 848 10683 869
rect 10767 1003 13767 2848
rect 10767 885 10808 1003
rect 10926 885 13767 1003
rect 10767 848 13767 885
rect -2078 726 922 764
rect -2078 608 762 726
rect 880 608 922 726
rect -2078 -1070 922 608
rect -2078 -1188 -2022 -1070
rect -1904 -1188 922 -1070
rect -2078 -1236 922 -1188
rect 1006 729 4006 764
rect 1006 611 1044 729
rect 1162 708 4006 729
rect 1162 611 3830 708
rect 1006 590 3830 611
rect 3948 590 4006 708
rect 1006 -1236 4006 590
rect 4090 706 5590 764
rect 4090 588 4122 706
rect 4240 588 5590 706
rect 4090 -1236 5590 588
rect 6099 706 7599 764
rect 6099 588 7449 706
rect 7567 588 7599 706
rect 6099 -1236 7599 588
rect 7683 729 10683 764
rect 7683 708 10527 729
rect 7683 590 7741 708
rect 7859 611 10527 708
rect 10645 611 10683 729
rect 7859 590 10683 611
rect 7683 -1236 10683 590
rect 10767 726 13767 764
rect 10767 608 10809 726
rect 10927 608 13767 726
rect 10767 -1070 13767 608
rect 10767 -1188 13593 -1070
rect 13711 -1188 13767 -1070
rect 10767 -1236 13767 -1188
rect -2079 -2122 421 -2091
rect -2079 -2240 -2037 -2122
rect -1919 -2145 421 -2122
rect -1919 -2240 241 -2145
rect -2079 -2263 241 -2240
rect 359 -2263 421 -2145
rect -2079 -5091 421 -2263
rect 505 -2145 3005 -2091
rect 505 -2263 554 -2145
rect 672 -2263 3005 -2145
rect 505 -5091 3005 -2263
rect 3089 -2127 5590 -2091
rect 3089 -2138 5438 -2127
rect 3089 -2256 3571 -2138
rect 3689 -2245 5438 -2138
rect 5556 -2245 5590 -2127
rect 3689 -2256 5590 -2245
rect 3089 -5091 5590 -2256
rect 6099 -2132 8600 -2091
rect 6099 -2135 8437 -2132
rect 6099 -2253 6126 -2135
rect 6244 -2250 8437 -2135
rect 8555 -2250 8600 -2132
rect 6244 -2253 8600 -2250
rect 6099 -5091 8600 -2253
rect 8684 -2133 11184 -2091
rect 8684 -2251 8730 -2133
rect 8848 -2145 11184 -2133
rect 8848 -2251 11017 -2145
rect 8684 -2263 11017 -2251
rect 11135 -2263 11184 -2145
rect 8684 -5091 11184 -2263
rect 11268 -2122 13768 -2091
rect 11268 -2145 13608 -2122
rect 11268 -2263 11330 -2145
rect 11448 -2240 13608 -2145
rect 13726 -2240 13768 -2122
rect 11448 -2263 13768 -2240
rect 11268 -5091 13768 -2263
<< mimcap2contact >>
rect 763 885 881 1003
rect 1047 887 1165 1005
rect 3833 869 3951 987
rect 4124 874 4242 992
rect 7447 874 7565 992
rect 7738 869 7856 987
rect 10524 887 10642 1005
rect 10808 885 10926 1003
rect 762 608 880 726
rect -2022 -1188 -1904 -1070
rect 1044 611 1162 729
rect 3830 590 3948 708
rect 4122 588 4240 706
rect 7449 588 7567 706
rect 7741 590 7859 708
rect 10527 611 10645 729
rect 10809 608 10927 726
rect 13593 -1188 13711 -1070
rect -2037 -2240 -1919 -2122
rect 241 -2263 359 -2145
rect 554 -2263 672 -2145
rect 3571 -2256 3689 -2138
rect 5438 -2245 5556 -2127
rect 6126 -2253 6244 -2135
rect 8437 -2250 8555 -2132
rect 8730 -2251 8848 -2133
rect 11017 -2263 11135 -2145
rect 11330 -2263 11448 -2145
rect 13608 -2240 13726 -2122
<< metal5 >>
rect 730 1005 1188 1029
rect 730 1003 1047 1005
rect 730 885 763 1003
rect 881 887 1047 1003
rect 1165 887 1188 1005
rect 881 885 1188 887
rect 730 729 1188 885
rect 730 726 1044 729
rect 730 608 762 726
rect 880 611 1044 726
rect 1162 611 1188 729
rect 880 608 1188 611
rect 730 592 1188 608
rect 3809 992 4266 1013
rect 3809 987 4124 992
rect 3809 869 3833 987
rect 3951 874 4124 987
rect 4242 874 4266 992
rect 3951 869 4266 874
rect 3809 708 4266 869
rect 3809 590 3830 708
rect 3948 706 4266 708
rect 3948 590 4122 706
rect 3809 588 4122 590
rect 4240 588 4266 706
rect 3809 569 4266 588
rect 7423 992 7880 1013
rect 7423 874 7447 992
rect 7565 987 7880 992
rect 7565 874 7738 987
rect 7423 869 7738 874
rect 7856 869 7880 987
rect 7423 708 7880 869
rect 7423 706 7741 708
rect 7423 588 7449 706
rect 7567 590 7741 706
rect 7859 590 7880 708
rect 10501 1005 10959 1029
rect 10501 887 10524 1005
rect 10642 1003 10959 1005
rect 10642 887 10808 1003
rect 10501 885 10808 887
rect 10926 885 10959 1003
rect 10501 729 10959 885
rect 10501 611 10527 729
rect 10645 726 10959 729
rect 10645 611 10809 726
rect 10501 608 10809 611
rect 10927 608 10959 726
rect 10501 592 10959 608
rect 7567 588 7880 590
rect 7423 569 7880 588
rect -2059 -1070 -1892 -1058
rect -2059 -1188 -2022 -1070
rect -1904 -1188 -1892 -1070
rect -2059 -1853 -1892 -1188
rect -2059 -1976 -2030 -1853
rect -1908 -1976 -1892 -1853
rect 13581 -1070 13748 -1058
rect 13581 -1188 13593 -1070
rect 13711 -1188 13748 -1070
rect 13581 -1853 13748 -1188
rect -2059 -2122 -1892 -1976
rect 3555 -1919 3719 -1906
rect 3555 -2037 3570 -1919
rect 3689 -2037 3719 -1919
rect 3555 -2116 3719 -2037
rect 13581 -1976 13597 -1853
rect 13719 -1976 13748 -1853
rect -2059 -2240 -2037 -2122
rect -1919 -2240 -1892 -2122
rect -2059 -2263 -1892 -2240
rect 218 -2145 700 -2119
rect 218 -2263 241 -2145
rect 359 -2263 554 -2145
rect 672 -2263 700 -2145
rect 218 -2280 700 -2263
rect 3555 -2138 3716 -2116
rect 3555 -2256 3571 -2138
rect 3689 -2256 3716 -2138
rect 3555 -2274 3716 -2256
rect 5403 -2127 6277 -2103
rect 5403 -2245 5438 -2127
rect 5556 -2135 6277 -2127
rect 5556 -2245 6126 -2135
rect 5403 -2253 6126 -2245
rect 6244 -2253 6277 -2135
rect 5403 -2272 6277 -2253
rect 8414 -2132 8870 -2104
rect 8414 -2250 8437 -2132
rect 8555 -2133 8870 -2132
rect 8555 -2250 8730 -2133
rect 8414 -2251 8730 -2250
rect 8848 -2251 8870 -2133
rect 8414 -2279 8870 -2251
rect 10989 -2145 11471 -2119
rect 10989 -2263 11017 -2145
rect 11135 -2263 11330 -2145
rect 11448 -2263 11471 -2145
rect 13581 -2122 13748 -1976
rect 13581 -2240 13608 -2122
rect 13726 -2240 13748 -2122
rect 13581 -2263 13748 -2240
rect 10989 -2280 11471 -2263
use mux  mux_0
timestamp 1647510647
transform 1 0 3708 0 1 -1719
box -59 -76 110 211
use multiplier  multiplier_0
timestamp 1647558825
transform 1 0 5046 0 1 -1813
box -213 -76 236 240
<< labels >>
rlabel metal4 2614 -1619 2614 -1619 5 cs1
rlabel metal4 2639 -1825 2639 -1825 7 cs2
rlabel metal4 3214 -1859 3214 -1859 5 cs3
rlabel locali 2821 -1388 2821 -1388 3 c1
rlabel locali 2909 -1946 2909 -1946 3 c2
rlabel locali 3120 -1946 3120 -1946 7 c3
rlabel metal2 5638 2887 5638 2887 1 VDD
rlabel metal2 5673 2887 5673 2887 1 inp_i
rlabel metal2 5708 2887 5708 2887 1 inm_i
rlabel metal2 5743 2887 5743 2887 1 thresh1
rlabel metal2 5778 2887 5778 2887 1 thresh2
rlabel metal2 5813 2887 5813 2887 1 cclk
rlabel metal2 5848 2887 5848 2887 1 cclkb
rlabel metal2 5883 2887 5883 2887 1 phi1
rlabel metal2 5918 2887 5918 2887 1 phi1b
rlabel metal2 5953 2887 5953 2887 1 phi2
rlabel metal2 5988 2887 5988 2887 1 phi2b
rlabel metal1 5948 -1890 5948 -1890 7 GND
rlabel via1 5948 -1839 5948 -1839 7 PHI2
rlabel metal1 5948 -1717 5948 -1717 7 PHI1
rlabel metal1 5948 -1662 5948 -1662 7 PHI2b
rlabel metal1 5948 -1540 5948 -1540 7 PHI1b
rlabel metal1 5948 -1436 5948 -1436 7 VDD
rlabel locali 8569 -1946 8569 -1946 3 c3
rlabel locali 8780 -1946 8780 -1946 7 c2
rlabel locali 8868 -1388 8868 -1388 7 c1
rlabel metal4 8475 -1859 8475 -1859 5 cs3
rlabel metal4 9050 -1825 9050 -1825 3 cs2
rlabel metal4 9075 -1619 9075 -1619 5 cs1
rlabel via1 6055 -1891 6055 -1891 7 PHI2
rlabel metal2 6058 2887 6058 2887 1 GND
rlabel metal2 6023 2887 6023 2887 1 sin
flabel metal4 1885 -36 2909 887 0 FreeSans 800 0 0 0 C1
flabel metal4 -82 -4020 942 -3097 0 FreeSans 800 0 0 0 C2
flabel mimcap2 3912 -3769 4936 -2846 0 FreeSans 800 0 0 0 C3
flabel mimcap2 6772 -3719 7796 -2796 0 FreeSans 800 0 0 0 C3
flabel metal4 10556 -3940 11580 -3017 0 FreeSans 800 0 0 0 C2
flabel mimcap2 9352 -417 10376 506 0 FreeSans 800 0 0 0 C1
flabel space 4635 -1551 5016 -1331 0 FreeSans 800 0 0 0 Multiplier
flabel mimcap 2256 -1622 2447 -1471 0 FreeSans 800 0 0 0 Cs1
flabel mimcap 2236 -1983 2427 -1832 0 FreeSans 800 0 0 0 Cs2
flabel mimcap 3300 -1963 3491 -1812 0 FreeSans 800 0 0 0 Cs3
flabel space 3871 -1679 4423 -1533 0 FreeSans 400 0 0 0 Mux_level_crossing
flabel space 2612 -1754 3046 -1673 0 FreeSans 400 0 0 0 Filter_switches
<< end >>
