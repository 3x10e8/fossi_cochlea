magic
tech sky130A
magscale 1 2
timestamp 1648937575
<< metal1 >>
rect 11566 -2518 11618 -2512
rect 11192 -2570 11566 -2546
rect 11618 -2570 11724 -2546
rect 11192 -2574 11724 -2570
rect 11566 -2576 11618 -2574
rect 11494 -2608 11546 -2604
rect 11194 -2610 11744 -2608
rect 11194 -2636 11494 -2610
rect 11546 -2636 11744 -2610
rect 11494 -2668 11546 -2662
rect 11200 -2694 11252 -2688
rect 10316 -2734 11200 -2700
rect 11252 -2734 11744 -2700
rect 11200 -2752 11252 -2746
rect 11426 -3162 11478 -3156
rect 11194 -3198 11426 -3170
rect 11426 -3220 11478 -3214
rect 11634 -3162 11686 -3156
rect 11686 -3198 11722 -3170
rect 11634 -3220 11686 -3214
rect 11285 -3436 11337 -3430
rect 11192 -3488 11285 -3468
rect 11337 -3488 11718 -3468
rect 11192 -3496 11718 -3488
rect 11366 -3530 11418 -3524
rect 11194 -3560 11366 -3532
rect 11418 -3560 11722 -3532
rect 11366 -3588 11418 -3582
rect 11208 -9720 11308 -9704
rect 11208 -9772 11215 -9720
rect 11267 -9772 11308 -9720
rect 11208 -9802 11308 -9772
rect 21487 -9947 27164 -9907
rect 13450 -10116 13508 -10101
rect 13450 -10168 13453 -10116
rect 13505 -10168 13508 -10116
rect 13450 -10182 13508 -10168
rect 21494 -10262 27166 -10222
rect 19471 -10439 19472 -10387
rect 19524 -10439 19525 -10387
<< via1 >>
rect 11566 -2570 11618 -2518
rect 11494 -2662 11546 -2610
rect 11200 -2746 11252 -2694
rect 11426 -3214 11478 -3162
rect 11634 -3214 11686 -3162
rect 11285 -3488 11337 -3436
rect 11366 -3582 11418 -3530
rect 11215 -9772 11267 -9720
rect 13453 -10168 13505 -10116
rect 19472 -10439 19524 -10387
<< metal2 >>
rect 8930 6502 11396 6542
rect 7336 6278 11326 6318
rect 5626 6088 11256 6128
rect 11226 -2688 11256 6088
rect 11200 -2694 11256 -2688
rect 11252 -2746 11256 -2694
rect 11200 -2752 11256 -2746
rect 11226 -9704 11256 -2752
rect 11296 -3430 11326 6278
rect 11285 -3436 11337 -3430
rect 11285 -3494 11337 -3488
rect 11295 -3496 11337 -3494
rect 11296 -3497 11337 -3496
rect 11296 -9682 11326 -3497
rect 11366 -3524 11396 6502
rect 11436 -3156 11466 7440
rect 11506 6504 14192 6544
rect 11506 -2604 11536 6504
rect 11576 6276 15768 6316
rect 11576 -2512 11606 6276
rect 11646 6088 17002 6128
rect 11566 -2518 11618 -2512
rect 11566 -2576 11618 -2570
rect 11494 -2610 11546 -2604
rect 11494 -2668 11546 -2662
rect 11426 -3162 11478 -3156
rect 11426 -3220 11478 -3214
rect 11366 -3530 11418 -3524
rect 11366 -3588 11418 -3582
rect 11506 -9680 11536 -2668
rect 11646 -3156 11676 6088
rect 11634 -3162 11686 -3156
rect 11634 -3220 11686 -3214
rect 11208 -9720 11268 -9704
rect 11208 -9772 11215 -9720
rect 11267 -9772 11268 -9720
rect 11208 -9802 11268 -9772
rect 13450 -10116 13508 -10096
rect 13450 -10168 13453 -10116
rect 13505 -10168 13508 -10116
rect 13450 -10551 13508 -10168
rect 19459 -10387 19536 -10378
rect 19459 -10443 19469 -10387
rect 19525 -10443 19536 -10387
rect 19459 -10453 19536 -10443
<< via2 >>
rect 19469 -10439 19472 -10387
rect 19472 -10439 19524 -10387
rect 19524 -10439 19525 -10387
rect 19469 -10443 19525 -10439
<< metal3 >>
rect -5284 5705 -5096 6012
rect 11120 5512 11761 5675
rect 11139 4857 11780 5020
rect 10991 3273 11899 3546
rect 11015 2017 11923 2290
rect 10976 820 11884 1093
rect 11049 -308 11957 -35
rect 10991 -1407 11899 -1134
rect 19415 -10387 19583 -9532
rect 19415 -10443 19469 -10387
rect 19525 -10443 19583 -10387
rect 19415 -10468 19583 -10443
<< metal4 >>
rect 11126 -9630 11184 -9628
rect 11126 -10112 11186 -9630
rect 11614 -9650 11720 -9552
rect 11614 -10048 11674 -9650
rect 11596 -10088 11674 -10048
rect 11126 -10172 11357 -10112
use ../comparator/comparator_final  comparator_final_0
timestamp 1647895372
transform 1 0 11870 0 1 -10038
box -574 -430 9642 401
use fitler_cell  fitler_cell_0
timestamp 1647840975
transform 1 0 4 0 1 0
box -5288 -9650 11208 6206
use fitler_cell  fitler_cell_1
timestamp 1647840975
transform -1 0 22898 0 1 0
box -5288 -9650 11208 6206
<< labels >>
rlabel metal2 s 13477 -10551 13477 -10551 4 compout
port 1 nsew
rlabel metal3 s -5197 6012 -5197 6012 4 vssa1
port 8 nsew
rlabel space 27695 6206 27695 6206 1 inm
port 12 n
rlabel space -4792 6206 -4792 6206 1 inp
port 13 n
rlabel metal2 14192 6526 14192 6526 3 phi1b
port 14 e
rlabel metal2 15768 6294 15768 6294 3 phi2b
port 15 e
rlabel metal2 17002 6108 17002 6108 3 vbotm
port 16 e
rlabel metal2 11452 7440 11452 7440 1 vbotp
port 17 n
rlabel metal2 5626 6108 5626 6108 7 vdda1
port 18 w
rlabel metal2 7336 6298 7336 6298 7 phi1
port 19 w
rlabel metal2 8930 6524 8930 6524 7 phi2
port 20 w
rlabel metal1 27166 -10244 27166 -10244 3 events
port 21 e
rlabel metal1 27164 -9928 27164 -9928 3 polxevent
port 22 e
<< end >>
