VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO analog_core_Q
  CLASS BLOCK ;
  FOREIGN analog_core_Q ;
  ORIGIN 0.000 2.450 ;
  SIZE 2038.520 BY 187.340 ;
  PIN fb1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.390 184.885 25.670 184.895 ;
    END
  END fb1[0]
  PIN fb1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 279.310 184.885 279.590 184.895 ;
    END
  END fb1[1]
  PIN fb1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 533.230 184.885 533.510 184.895 ;
    END
  END fb1[2]
  PIN fb1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.150 184.885 787.430 184.895 ;
    END
  END fb1[3]
  PIN fb1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1041.070 184.885 1041.350 184.895 ;
    END
  END fb1[4]
  PIN fb1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1294.990 184.885 1295.270 184.895 ;
    END
  END fb1[5]
  PIN fb1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1548.910 184.885 1549.190 184.895 ;
    END
  END fb1[6]
  PIN fb1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1802.830 184.885 1803.110 184.895 ;
    END
  END fb1[7]
  PIN cclk[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.710 184.885 67.990 184.895 ;
    END
  END cclk[0]
  PIN cclk[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 321.630 184.885 321.910 184.895 ;
    END
  END cclk[1]
  PIN cclk[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 575.550 184.885 575.830 184.895 ;
    END
  END cclk[2]
  PIN cclk[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.470 184.885 829.750 184.895 ;
    END
  END cclk[3]
  PIN cclk[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1083.390 184.885 1083.670 184.895 ;
    END
  END cclk[4]
  PIN cclk[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1337.310 184.885 1337.590 184.895 ;
    END
  END cclk[5]
  PIN cclk[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1591.230 184.885 1591.510 184.895 ;
    END
  END cclk[6]
  PIN cclk[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.150 184.885 1845.430 184.895 ;
    END
  END cclk[7]
  PIN div2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.030 184.885 110.310 184.895 ;
    END
  END div2[0]
  PIN div2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 363.950 184.885 364.230 184.895 ;
    END
  END div2[1]
  PIN div2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 617.870 184.885 618.150 184.895 ;
    END
  END div2[2]
  PIN div2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 871.790 184.885 872.070 184.895 ;
    END
  END div2[3]
  PIN div2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1125.710 184.885 1125.990 184.895 ;
    END
  END div2[4]
  PIN div2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1379.630 184.885 1379.910 184.895 ;
    END
  END div2[5]
  PIN div2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1633.550 184.885 1633.830 184.895 ;
    END
  END div2[6]
  PIN div2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1887.470 184.885 1887.750 184.895 ;
    END
  END div2[7]
  PIN high_buf[0]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 152.350 184.885 152.630 184.895 ;
    END
  END high_buf[0]
  PIN high_buf[1]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 406.270 184.885 406.550 184.895 ;
    END
  END high_buf[1]
  PIN high_buf[2]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 660.190 184.885 660.470 184.895 ;
    END
  END high_buf[2]
  PIN high_buf[3]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 914.110 184.885 914.390 184.895 ;
    END
  END high_buf[3]
  PIN high_buf[4]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.030 184.885 1168.310 184.895 ;
    END
  END high_buf[4]
  PIN high_buf[5]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 1421.950 184.885 1422.230 184.895 ;
    END
  END high_buf[5]
  PIN high_buf[6]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 1675.870 184.885 1676.150 184.895 ;
    END
  END high_buf[6]
  PIN high_buf[7]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.790 184.885 1930.070 184.895 ;
    END
  END high_buf[7]
  PIN phi1b_dig[0]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 194.670 184.885 194.950 184.895 ;
    END
  END phi1b_dig[0]
  PIN phi1b_dig[1]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 448.590 184.885 448.870 184.895 ;
    END
  END phi1b_dig[1]
  PIN phi1b_dig[2]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 702.510 184.885 702.790 184.895 ;
    END
  END phi1b_dig[2]
  PIN phi1b_dig[3]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 956.430 184.885 956.710 184.895 ;
    END
  END phi1b_dig[3]
  PIN phi1b_dig[4]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 1210.350 184.885 1210.630 184.895 ;
    END
  END phi1b_dig[4]
  PIN phi1b_dig[5]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 1464.270 184.885 1464.550 184.895 ;
    END
  END phi1b_dig[5]
  PIN phi1b_dig[6]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 1718.190 184.885 1718.470 184.895 ;
    END
  END phi1b_dig[6]
  PIN phi1b_dig[7]
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 1972.110 184.885 1972.390 184.895 ;
    END
  END phi1b_dig[7]
  PIN lo[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.990 184.885 237.270 184.895 ;
    END
  END lo[0]
  PIN lo[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.910 184.885 491.190 184.895 ;
    END
  END lo[1]
  PIN lo[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 744.830 184.885 745.110 184.895 ;
    END
  END lo[2]
  PIN lo[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 998.750 184.885 999.030 184.895 ;
    END
  END lo[3]
  PIN lo[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1252.670 184.885 1252.950 184.895 ;
    END
  END lo[4]
  PIN lo[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.590 184.885 1506.870 184.895 ;
    END
  END lo[5]
  PIN lo[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1760.510 184.885 1760.790 184.895 ;
    END
  END lo[6]
  PIN lo[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2014.430 184.885 2014.710 184.895 ;
    END
  END lo[7]
  PIN vnb
    DIRECTION INOUT ;
    PORT
      LAYER met1 ;
        RECT 2038.515 184.360 2038.525 184.860 ;
    END
  END vnb
  PIN vpb
    DIRECTION INOUT ;
    PORT
      LAYER met1 ;
        RECT 2038.515 164.465 2038.525 164.970 ;
    END
  END vpb
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 2038.515 144.500 2038.525 145.000 ;
    END
  END vccd1
  PIN th1
    DIRECTION INOUT ;
    PORT
      LAYER met1 ;
        RECT 2038.515 124.500 2038.525 125.000 ;
    END
  END th1
  PIN th2
    DIRECTION INOUT ;
    PORT
      LAYER met1 ;
        RECT 2038.515 104.500 2038.525 105.000 ;
    END
  END th2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 2038.515 84.500 2038.525 85.000 ;
    END
  END vssd1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 2038.515 64.500 2038.525 65.000 ;
    END
  END vdda1
  OBS
      LAYER li1 ;
        RECT 3.230 124.330 2014.850 175.040 ;
      LAYER met1 ;
        RECT 2.565 184.080 2038.235 184.890 ;
        RECT 2.565 165.250 2038.515 184.080 ;
        RECT 2.565 164.185 2038.235 165.250 ;
        RECT 2.565 145.280 2038.515 164.185 ;
        RECT 2.565 144.220 2038.235 145.280 ;
        RECT 2.565 125.280 2038.515 144.220 ;
        RECT 2.565 124.220 2038.235 125.280 ;
        RECT 2.565 105.280 2038.515 124.220 ;
        RECT 2.565 104.220 2038.235 105.280 ;
        RECT 2.565 85.280 2038.515 104.220 ;
        RECT 2.565 84.220 2038.235 85.280 ;
        RECT 2.565 65.280 2038.515 84.220 ;
        RECT 2.565 64.500 2038.235 65.280 ;
      LAYER met2 ;
        RECT 2.590 184.605 25.110 184.890 ;
        RECT 25.950 184.605 67.430 184.890 ;
        RECT 68.270 184.605 109.750 184.890 ;
        RECT 110.590 184.605 152.070 184.890 ;
        RECT 152.910 184.605 194.390 184.890 ;
        RECT 195.230 184.605 236.710 184.890 ;
        RECT 237.550 184.605 279.030 184.890 ;
        RECT 279.870 184.605 321.350 184.890 ;
        RECT 322.190 184.605 363.670 184.890 ;
        RECT 364.510 184.605 405.990 184.890 ;
        RECT 406.830 184.605 448.310 184.890 ;
        RECT 449.150 184.605 490.630 184.890 ;
        RECT 491.470 184.605 532.950 184.890 ;
        RECT 533.790 184.605 575.270 184.890 ;
        RECT 576.110 184.605 617.590 184.890 ;
        RECT 618.430 184.605 659.910 184.890 ;
        RECT 660.750 184.605 702.230 184.890 ;
        RECT 703.070 184.605 744.550 184.890 ;
        RECT 745.390 184.605 786.870 184.890 ;
        RECT 787.710 184.605 829.190 184.890 ;
        RECT 830.030 184.605 871.510 184.890 ;
        RECT 872.350 184.605 913.830 184.890 ;
        RECT 914.670 184.605 956.150 184.890 ;
        RECT 956.990 184.605 998.470 184.890 ;
        RECT 999.310 184.605 1040.790 184.890 ;
        RECT 1041.630 184.605 1083.110 184.890 ;
        RECT 1083.950 184.605 1125.430 184.890 ;
        RECT 1126.270 184.605 1167.750 184.890 ;
        RECT 1168.590 184.605 1210.070 184.890 ;
        RECT 1210.910 184.605 1252.390 184.890 ;
        RECT 1253.230 184.605 1294.710 184.890 ;
        RECT 1295.550 184.605 1337.030 184.890 ;
        RECT 1337.870 184.605 1379.350 184.890 ;
        RECT 1380.190 184.605 1421.670 184.890 ;
        RECT 1422.510 184.605 1463.990 184.890 ;
        RECT 1464.830 184.605 1506.310 184.890 ;
        RECT 1507.150 184.605 1548.630 184.890 ;
        RECT 1549.470 184.605 1590.950 184.890 ;
        RECT 1591.790 184.605 1633.270 184.890 ;
        RECT 1634.110 184.605 1675.590 184.890 ;
        RECT 1676.430 184.605 1717.910 184.890 ;
        RECT 1718.750 184.605 1760.230 184.890 ;
        RECT 1761.070 184.605 1802.550 184.890 ;
        RECT 1803.390 184.605 1844.870 184.890 ;
        RECT 1845.710 184.605 1887.190 184.890 ;
        RECT 1888.030 184.605 1929.510 184.890 ;
        RECT 1930.350 184.605 1971.830 184.890 ;
        RECT 1972.670 184.605 2014.150 184.890 ;
        RECT 2014.990 184.605 2037.360 184.890 ;
        RECT 2.590 64.470 2037.360 184.605 ;
      LAYER met3 ;
        RECT 0.000 -0.810 2037.360 176.620 ;
      LAYER met4 ;
        RECT 0.000 -2.450 2031.360 176.620 ;
      LAYER met5 ;
        RECT 0.000 -2.450 2031.360 139.505 ;
  END
END analog_core_Q
END LIBRARY

