* NGSPICE file created from comparator.ext - technology: sky130B

.subckt inv_LV A w_987_322# a_1138_96# a_1032_466# a_1136_466# VSUBS
X0 a_1136_466# A a_1032_466# w_987_322# sky130_fd_pr__pfet_01v8 ad=1.554e+11p pd=1.58e+06u as=1.554e+11p ps=1.58e+06u w=420000u l=150000u
X1 a_1138_96# A a_1032_466# VSUBS sky130_fd_pr__nfet_01v8 ad=1.554e+11p pd=1.58e+06u as=1.554e+11p ps=1.58e+06u w=420000u l=150000u
.ends

.subckt comparator
Xinv_LV_2 inv_LV_2/A w_n359_n11# inv_LV_7/VSUBS inv_LV_3/A w_n359_n11# inv_LV_7/VSUBS
+ inv_LV
Xinv_LV_3 inv_LV_3/A w_n359_n11# inv_LV_7/VSUBS li_1873_504# w_n359_n11# inv_LV_7/VSUBS
+ inv_LV
Xinv_LV_4 inv_LV_4/A w_n359_n11# inv_LV_7/VSUBS inv_LV_4/a_1032_466# w_n359_n11# inv_LV_7/VSUBS
+ inv_LV
Xinv_LV_5 inv_LV_5/A w_n359_n11# inv_LV_7/VSUBS inv_LV_4/A w_n359_n11# inv_LV_7/VSUBS
+ inv_LV
Xinv_LV_6 inv_LV_6/A w_n359_n11# inv_LV_7/VSUBS inv_LV_5/A w_n359_n11# inv_LV_7/VSUBS
+ inv_LV
Xinv_LV_7 low w_n359_n11# inv_LV_7/VSUBS inv_LV_6/A w_n359_n11# inv_LV_7/VSUBS inv_LV
Xinv_LV_0 low w_n359_n11# inv_LV_7/VSUBS inv_LV_1/A w_n359_n11# inv_LV_7/VSUBS inv_LV
Xinv_LV_1 inv_LV_1/A w_n359_n11# inv_LV_7/VSUBS inv_LV_2/A w_n359_n11# inv_LV_7/VSUBS
+ inv_LV
X0 tail a_10_n824# inv_LV_7/VSUBS inv_LV_7/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.197e+11p pd=1.41e+06u as=1.9131e+12p ps=2.003e+07u w=420000u l=2e+06u
X1 inv_LV_7/VSUBS a_n618_473# low inv_LV_7/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.394e+11p ps=2.82e+06u w=420000u l=2e+06u
X2 low FP pfetw w_n359_n11# sky130_fd_pr__pfet_01v8 ad=5.9e+11p pd=5.18e+06u as=2.815e+11p ps=2.65e+06u w=1e+06u l=150000u
X3 inv_LV_7/VSUBS a_n618_473# low inv_LV_7/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=2e+06u
X4 pfetw low w_n359_n11# w_n359_n11# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.5981e+12p ps=1.685e+07u w=420000u l=150000u
X5 FN a_10_n824# w_n359_n11# w_n359_n11# sky130_fd_pr__pfet_01v8 ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X6 FP inp tail inv_LV_7/VSUBS sky130_fd_pr__nfet_03v3_nvt ad=2.85e+11p pd=2.57e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=500000u
X7 pfete FN low w_n359_n11# sky130_fd_pr__pfet_01v8 ad=2.815e+11p pd=2.65e+06u as=0p ps=0u w=1e+06u l=150000u
X8 w_n359_n11# low pfete w_n359_n11# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 low low inv_LV_7/VSUBS inv_LV_7/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=2e+06u
X10 FN a_280_n337# tail inv_LV_7/VSUBS sky130_fd_pr__nfet_03v3_nvt ad=2.85e+11p pd=2.57e+06u as=0p ps=0u w=1e+06u l=500000u
X11 low low inv_LV_7/VSUBS inv_LV_7/VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=2e+06u
X12 w_n359_n11# a_10_n824# FP w_n359_n11# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
.ends

