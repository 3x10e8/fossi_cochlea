* NGSPICE file created from /local_disk/fossi_cochlea/mag/final_designs/caps/cap_3pF.ext - technology: sky130B

.subckt cap_10_10_center_x2 m3_n710_n366# c1_n16_n6#
X0 m3_n710_n366# c1_n16_n6# sky130_fd_pr__cap_mim_m3_2 l=1e+07u w=1e+07u
X1 c1_n16_n6# m3_n710_n366# sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
.ends

.subckt cap_10_10_side2_x2 m3_n710_n366# c1_n16_n6#
X0 m3_n710_n366# c1_n16_n6# sky130_fd_pr__cap_mim_m3_2 l=1e+07u w=1e+07u
X1 c1_n16_n6# m3_n710_n366# sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
.ends

.subckt cap_3pF ref sig
Xcap_10_10_center_x2_0[0] ref sig cap_10_10_center_x2
Xcap_10_10_center_x2_0[1] ref sig cap_10_10_center_x2
Xcap_10_10_center_x2_0[2] ref sig cap_10_10_center_x2
Xcap_10_10_center_x2_0[3] ref sig cap_10_10_center_x2
Xcap_10_10_center_x2_0[4] ref sig cap_10_10_center_x2
Xcap_10_10_center_x2_0[5] ref sig cap_10_10_center_x2
Xcap_10_10_side2_x2_0 ref sig cap_10_10_side2_x2
Xcap_10_10_side2_x2_1 ref sig cap_10_10_side2_x2
.ends

