magic
tech sky130A
timestamp 1647558825
<< nwell >>
rect -213 95 236 182
<< nmos >>
rect -155 -21 -140 21
rect -111 -21 -96 21
rect -1 -21 14 21
rect 43 -21 58 21
rect 144 -21 159 21
<< pmos >>
rect -155 114 -140 156
rect -111 114 -96 156
rect -1 114 14 156
rect 43 114 58 156
rect 144 114 159 156
<< ndiff >>
rect -184 9 -155 21
rect -184 -8 -178 9
rect -161 -8 -155 9
rect -184 -21 -155 -8
rect -140 9 -111 21
rect -140 -8 -134 9
rect -117 -8 -111 9
rect -140 -21 -111 -8
rect -96 9 -67 21
rect -96 -8 -90 9
rect -73 -8 -67 9
rect -96 -21 -67 -8
rect -30 9 -1 21
rect -30 -8 -24 9
rect -7 -8 -1 9
rect -30 -21 -1 -8
rect 14 9 43 21
rect 14 -8 20 9
rect 37 -8 43 9
rect 14 -21 43 -8
rect 58 9 87 21
rect 58 -8 64 9
rect 81 -8 87 9
rect 58 -21 87 -8
rect 117 8 144 21
rect 117 -9 121 8
rect 138 -9 144 8
rect 117 -21 144 -9
rect 159 8 190 21
rect 159 -9 165 8
rect 182 -9 190 8
rect 159 -21 190 -9
<< pdiff >>
rect -184 144 -155 156
rect -184 127 -178 144
rect -161 127 -155 144
rect -184 114 -155 127
rect -140 144 -111 156
rect -140 127 -134 144
rect -117 127 -111 144
rect -140 114 -111 127
rect -96 144 -67 156
rect -96 127 -90 144
rect -73 127 -67 144
rect -96 114 -67 127
rect -30 144 -1 156
rect -30 127 -24 144
rect -7 127 -1 144
rect -30 114 -1 127
rect 14 144 43 156
rect 14 127 20 144
rect 37 127 43 144
rect 14 114 43 127
rect 58 144 87 156
rect 58 127 64 144
rect 81 127 87 144
rect 58 114 87 127
rect 117 143 144 156
rect 117 126 121 143
rect 138 126 144 143
rect 117 114 144 126
rect 159 143 189 156
rect 159 126 165 143
rect 182 126 189 143
rect 159 114 189 126
<< ndiffc >>
rect -178 -8 -161 9
rect -134 -8 -117 9
rect -90 -8 -73 9
rect -24 -8 -7 9
rect 20 -8 37 9
rect 64 -8 81 9
rect 121 -9 138 8
rect 165 -9 182 8
<< pdiffc >>
rect -178 127 -161 144
rect -134 127 -117 144
rect -90 127 -73 144
rect -24 127 -7 144
rect 20 127 37 144
rect 64 127 81 144
rect 121 126 138 143
rect 165 126 182 143
<< psubdiff >>
rect 190 8 221 21
rect 190 -9 199 8
rect 216 -9 221 8
rect 190 -21 221 -9
<< nsubdiff >>
rect 189 143 218 156
rect 189 126 199 143
rect 216 126 218 143
rect 189 114 218 126
<< psubdiffcont >>
rect 199 -9 216 8
<< nsubdiffcont >>
rect 199 126 216 143
<< poly >>
rect -206 205 -179 206
rect -111 205 -25 206
rect -206 198 159 205
rect -206 190 -47 198
rect -206 189 -176 190
rect -213 173 -176 189
rect -111 189 -47 190
rect -213 44 -195 173
rect -155 156 -140 169
rect -111 156 -96 189
rect -59 181 -47 189
rect -30 190 159 198
rect -30 181 -22 190
rect -59 173 -22 181
rect -155 80 -140 114
rect -111 101 -96 114
rect -155 65 -96 80
rect -213 29 -140 44
rect -155 21 -140 29
rect -111 21 -96 65
rect -59 44 -41 173
rect -1 156 14 169
rect 43 156 58 190
rect 144 156 159 190
rect -1 80 14 114
rect 43 101 58 114
rect -1 65 58 80
rect -59 29 14 44
rect -1 21 14 29
rect 43 21 58 65
rect 144 21 159 114
rect -155 -34 -140 -21
rect -111 -56 -96 -21
rect -1 -34 14 -21
rect 43 -38 58 -21
rect 144 -34 159 -21
rect 37 -46 64 -38
rect 37 -56 42 -46
rect -111 -63 42 -56
rect 59 -63 64 -46
rect -111 -71 64 -63
<< polycont >>
rect -47 181 -30 198
rect 42 -63 59 -46
<< locali >>
rect -180 223 82 240
rect -180 156 -163 223
rect -50 198 -27 206
rect -50 181 -47 198
rect -30 181 -27 198
rect -50 173 -27 181
rect 65 156 82 223
rect -182 144 -157 156
rect -182 127 -178 144
rect -161 127 -157 144
rect -182 114 -157 127
rect -138 144 -113 156
rect -138 127 -134 144
rect -117 127 -113 144
rect -138 114 -113 127
rect -94 144 -69 156
rect -94 127 -90 144
rect -73 127 -69 144
rect -94 114 -69 127
rect -28 144 -3 156
rect -28 127 -24 144
rect -7 127 -3 144
rect -28 114 -3 127
rect 16 144 41 156
rect 16 127 20 144
rect 37 127 41 144
rect 16 114 41 127
rect 60 144 85 156
rect 60 127 64 144
rect 81 127 85 144
rect 60 114 85 127
rect 117 143 142 156
rect 117 126 121 143
rect 138 126 142 143
rect 117 114 142 126
rect 161 143 218 156
rect 161 126 165 143
rect 182 126 199 143
rect 216 126 218 143
rect 161 114 218 126
rect -181 21 -164 114
rect -134 21 -117 114
rect -89 21 -72 114
rect -27 21 -10 114
rect 20 21 37 114
rect 65 21 82 114
rect 117 21 134 114
rect -182 9 -157 21
rect -182 -8 -178 9
rect -161 -8 -157 9
rect -182 -21 -157 -8
rect -138 9 -113 21
rect -138 -8 -134 9
rect -117 -8 -113 9
rect -138 -21 -113 -8
rect -94 9 -69 21
rect -94 -8 -90 9
rect -73 8 -69 9
rect -28 9 -3 21
rect -28 8 -24 9
rect -73 -8 -24 8
rect -7 -8 -3 9
rect -94 -9 -3 -8
rect -94 -21 -69 -9
rect -28 -21 -3 -9
rect 16 9 41 21
rect 16 -8 20 9
rect 37 -8 41 9
rect 16 -21 41 -8
rect 60 9 85 21
rect 60 -8 64 9
rect 81 -8 85 9
rect 60 -21 85 -8
rect 117 8 142 21
rect 117 -9 121 8
rect 138 -9 142 8
rect 117 -21 142 -9
rect 161 8 221 21
rect 161 -9 165 8
rect 182 -9 199 8
rect 216 -9 221 8
rect 161 -21 221 -9
rect 39 -40 62 -38
rect 117 -40 134 -21
rect 39 -46 134 -40
rect 39 -63 42 -46
rect 59 -57 134 -46
rect 59 -63 62 -57
rect 39 -71 62 -63
<< labels >>
flabel locali -26 -20 -4 -9 0 FreeSans 80 0 0 0 Vref1
flabel locali 61 -21 83 -10 0 FreeSans 80 0 0 0 Vref2
flabel locali 18 -20 40 -9 0 FreeSans 80 0 0 0 Out
flabel space -51 200 -29 211 0 FreeSans 80 0 0 0 C
flabel space 39 -76 61 -65 0 FreeSans 80 0 0 0 Cbar
flabel locali -180 -20 -158 -9 0 FreeSans 80 0 0 0 Vref1
flabel locali -93 -21 -71 -10 0 FreeSans 80 0 0 0 Vref2
flabel locali -136 -20 -114 -9 0 FreeSans 80 0 0 0 Out
flabel space -205 200 -183 211 0 FreeSans 80 0 0 0 C
flabel space -115 -76 -93 -65 0 FreeSans 80 0 0 0 Cbar
flabel nwell 165 125 183 143 0 FreeSans 40 0 0 0 VDD
flabel locali 165 -10 183 8 0 FreeSans 40 0 0 0 GND
<< end >>
