magic
tech sky130B
magscale 1 2
timestamp 1662788822
<< viali >>
rect 4629 17289 4663 17323
rect 5273 17289 5307 17323
rect 12633 17289 12667 17323
rect 20361 17289 20395 17323
rect 28273 17289 28307 17323
rect 43637 17289 43671 17323
rect 52101 17289 52135 17323
rect 59921 17289 59955 17323
rect 68569 17289 68603 17323
rect 76297 17289 76331 17323
rect 91569 17289 91603 17323
rect 34345 17221 34379 17255
rect 55965 17221 55999 17255
rect 83289 17221 83323 17255
rect 85589 17221 85623 17255
rect 1685 17153 1719 17187
rect 4813 17153 4847 17187
rect 5457 17153 5491 17187
rect 12449 17153 12483 17187
rect 20545 17153 20579 17187
rect 28457 17153 28491 17187
rect 44281 17153 44315 17187
rect 52285 17153 52319 17187
rect 58817 17153 58851 17187
rect 60105 17153 60139 17187
rect 61301 17153 61335 17187
rect 62313 17153 62347 17187
rect 68385 17153 68419 17187
rect 76113 17153 76147 17187
rect 91753 17153 91787 17187
rect 92213 17153 92247 17187
rect 34897 17085 34931 17119
rect 36645 17085 36679 17119
rect 36921 17085 36955 17119
rect 37565 17085 37599 17119
rect 61117 17085 61151 17119
rect 63233 17085 63267 17119
rect 64337 17085 64371 17119
rect 65809 17085 65843 17119
rect 83841 17085 83875 17119
rect 85865 17085 85899 17119
rect 86417 17085 86451 17119
rect 44097 17017 44131 17051
rect 57069 17017 57103 17051
rect 63877 17017 63911 17051
rect 64981 17017 65015 17051
rect 67741 17017 67775 17051
rect 1961 16949 1995 16983
rect 42625 16949 42659 16983
rect 45937 16949 45971 16983
rect 46489 16949 46523 16983
rect 47041 16949 47075 16983
rect 56609 16949 56643 16983
rect 59369 16949 59403 16983
rect 61761 16949 61795 16983
rect 36369 16745 36403 16779
rect 38761 16745 38795 16779
rect 50353 16745 50387 16779
rect 60657 16745 60691 16779
rect 83841 16745 83875 16779
rect 94237 16745 94271 16779
rect 1593 16677 1627 16711
rect 54953 16677 54987 16711
rect 68109 16677 68143 16711
rect 68661 16677 68695 16711
rect 20361 16609 20395 16643
rect 31769 16609 31803 16643
rect 35725 16609 35759 16643
rect 41061 16609 41095 16643
rect 41705 16609 41739 16643
rect 42349 16609 42383 16643
rect 42809 16609 42843 16643
rect 45293 16609 45327 16643
rect 46213 16609 46247 16643
rect 46673 16609 46707 16643
rect 47501 16609 47535 16643
rect 56057 16609 56091 16643
rect 56793 16609 56827 16643
rect 57345 16609 57379 16643
rect 58725 16609 58759 16643
rect 62129 16609 62163 16643
rect 65809 16609 65843 16643
rect 67281 16609 67315 16643
rect 77033 16609 77067 16643
rect 93225 16609 93259 16643
rect 19717 16541 19751 16575
rect 36277 16541 36311 16575
rect 47317 16541 47351 16575
rect 59921 16541 59955 16575
rect 62405 16541 62439 16575
rect 62865 16541 62899 16575
rect 67557 16541 67591 16575
rect 83197 16541 83231 16575
rect 83749 16541 83783 16575
rect 92581 16541 92615 16575
rect 94053 16541 94087 16575
rect 53113 16473 53147 16507
rect 55505 16473 55539 16507
rect 63141 16473 63175 16507
rect 19625 16405 19659 16439
rect 32229 16405 32263 16439
rect 32873 16405 32907 16439
rect 43545 16405 43579 16439
rect 48237 16405 48271 16439
rect 52469 16405 52503 16439
rect 54401 16405 54435 16439
rect 58173 16405 58207 16439
rect 59185 16405 59219 16439
rect 60013 16405 60047 16439
rect 64613 16405 64647 16439
rect 65073 16405 65107 16439
rect 71973 16405 72007 16439
rect 92765 16405 92799 16439
rect 20085 16201 20119 16235
rect 44925 16201 44959 16235
rect 46765 16201 46799 16235
rect 52193 16201 52227 16235
rect 72525 16201 72559 16235
rect 31125 16133 31159 16167
rect 53573 16133 53607 16167
rect 55597 16133 55631 16167
rect 59737 16133 59771 16167
rect 65533 16133 65567 16167
rect 20821 16065 20855 16099
rect 29009 16065 29043 16099
rect 40877 16065 40911 16099
rect 41521 16065 41555 16099
rect 45385 16065 45419 16099
rect 46029 16065 46063 16099
rect 46673 16065 46707 16099
rect 50353 16065 50387 16099
rect 52377 16065 52411 16099
rect 53113 16065 53147 16099
rect 54217 16065 54251 16099
rect 56425 16065 56459 16099
rect 64337 16065 64371 16099
rect 65073 16065 65107 16099
rect 67373 16065 67407 16099
rect 71145 16065 71179 16099
rect 78873 16065 78907 16099
rect 18337 15997 18371 16031
rect 18613 15997 18647 16031
rect 39589 15997 39623 16031
rect 40141 15997 40175 16031
rect 40785 15997 40819 16031
rect 41981 15997 42015 16031
rect 49341 15997 49375 16031
rect 50537 15997 50571 16031
rect 61485 15997 61519 16031
rect 61761 15997 61795 16031
rect 63785 15997 63819 16031
rect 66453 15997 66487 16031
rect 76573 15997 76607 16031
rect 31585 15929 31619 15963
rect 34805 15929 34839 15963
rect 35357 15929 35391 15963
rect 65809 15929 65843 15963
rect 66729 15929 66763 15963
rect 70409 15929 70443 15963
rect 76021 15929 76055 15963
rect 79333 15929 79367 15963
rect 79977 15929 80011 15963
rect 20729 15861 20763 15895
rect 28917 15861 28951 15895
rect 29561 15861 29595 15895
rect 32689 15861 32723 15895
rect 33701 15861 33735 15895
rect 34253 15861 34287 15895
rect 35909 15861 35943 15895
rect 38761 15861 38795 15895
rect 42809 15861 42843 15895
rect 43453 15861 43487 15895
rect 44281 15861 44315 15895
rect 45477 15861 45511 15895
rect 46121 15861 46155 15895
rect 47777 15861 47811 15895
rect 48789 15861 48823 15895
rect 53021 15861 53055 15895
rect 55045 15861 55079 15895
rect 56517 15861 56551 15895
rect 57161 15861 57195 15895
rect 58081 15861 58115 15895
rect 58633 15861 58667 15895
rect 59185 15861 59219 15895
rect 62221 15861 62255 15895
rect 63233 15861 63267 15895
rect 65993 15861 66027 15895
rect 66913 15861 66947 15895
rect 68385 15861 68419 15895
rect 69029 15861 69063 15895
rect 69673 15861 69707 15895
rect 71053 15861 71087 15895
rect 72065 15861 72099 15895
rect 77033 15861 77067 15895
rect 77585 15861 77619 15895
rect 78781 15861 78815 15895
rect 80529 15861 80563 15895
rect 83197 15861 83231 15895
rect 83933 15861 83967 15895
rect 30113 15657 30147 15691
rect 38393 15657 38427 15691
rect 43821 15657 43855 15691
rect 68109 15657 68143 15691
rect 31585 15589 31619 15623
rect 44649 15589 44683 15623
rect 59369 15589 59403 15623
rect 67281 15589 67315 15623
rect 69673 15589 69707 15623
rect 72525 15589 72559 15623
rect 73169 15589 73203 15623
rect 73721 15589 73755 15623
rect 34989 15521 35023 15555
rect 36829 15521 36863 15555
rect 48973 15521 49007 15555
rect 61117 15521 61151 15555
rect 64705 15521 64739 15555
rect 64981 15521 65015 15555
rect 78873 15521 78907 15555
rect 79701 15521 79735 15555
rect 20177 15453 20211 15487
rect 20821 15453 20855 15487
rect 22661 15453 22695 15487
rect 28549 15453 28583 15487
rect 29193 15453 29227 15487
rect 31677 15453 31711 15487
rect 33425 15453 33459 15487
rect 33885 15453 33919 15487
rect 35081 15453 35115 15487
rect 38301 15453 38335 15487
rect 40325 15453 40359 15487
rect 40785 15453 40819 15487
rect 43729 15453 43763 15487
rect 45753 15453 45787 15487
rect 46673 15453 46707 15487
rect 48881 15453 48915 15487
rect 49525 15453 49559 15487
rect 51181 15453 51215 15487
rect 53849 15453 53883 15487
rect 56149 15453 56183 15487
rect 57069 15453 57103 15487
rect 60105 15453 60139 15487
rect 65809 15453 65843 15487
rect 65993 15453 66027 15487
rect 66821 15453 66855 15487
rect 67465 15453 67499 15487
rect 67925 15453 67959 15487
rect 69213 15453 69247 15487
rect 71513 15453 71547 15487
rect 72157 15453 72191 15487
rect 74181 15453 74215 15487
rect 75469 15453 75503 15487
rect 76297 15453 76331 15487
rect 79149 15453 79183 15487
rect 82921 15453 82955 15487
rect 30665 15385 30699 15419
rect 32505 15385 32539 15419
rect 43177 15385 43211 15419
rect 46949 15385 46983 15419
rect 51457 15385 51491 15419
rect 57345 15385 57379 15419
rect 61393 15385 61427 15419
rect 64889 15385 64923 15419
rect 66177 15385 66211 15419
rect 75101 15385 75135 15419
rect 75285 15385 75319 15419
rect 20085 15317 20119 15351
rect 20729 15317 20763 15351
rect 22753 15317 22787 15351
rect 23673 15317 23707 15351
rect 24869 15317 24903 15351
rect 28457 15317 28491 15351
rect 29101 15317 29135 15351
rect 33057 15317 33091 15351
rect 35541 15317 35575 15351
rect 36277 15317 36311 15351
rect 37657 15317 37691 15351
rect 39221 15317 39255 15351
rect 41153 15317 41187 15351
rect 41797 15317 41831 15351
rect 42349 15317 42383 15351
rect 45661 15317 45695 15351
rect 48421 15317 48455 15351
rect 50629 15317 50663 15351
rect 52929 15317 52963 15351
rect 53757 15317 53791 15351
rect 54401 15317 54435 15351
rect 54861 15317 54895 15351
rect 56057 15317 56091 15351
rect 58817 15317 58851 15351
rect 60013 15317 60047 15351
rect 62865 15317 62899 15351
rect 63417 15317 63451 15351
rect 66729 15317 66763 15351
rect 68661 15317 68695 15351
rect 70225 15317 70259 15351
rect 70961 15317 70995 15351
rect 71605 15317 71639 15351
rect 72617 15317 72651 15351
rect 74365 15317 74399 15351
rect 76481 15317 76515 15351
rect 77401 15317 77435 15351
rect 80161 15317 80195 15351
rect 81357 15317 81391 15351
rect 83749 15317 83783 15351
rect 84393 15317 84427 15351
rect 86509 15317 86543 15351
rect 88073 15317 88107 15351
rect 88901 15317 88935 15351
rect 28181 15113 28215 15147
rect 36829 15113 36863 15147
rect 53021 15113 53055 15147
rect 62313 15113 62347 15147
rect 67373 15113 67407 15147
rect 71513 15113 71547 15147
rect 72617 15113 72651 15147
rect 82185 15113 82219 15147
rect 19349 15045 19383 15079
rect 21097 15045 21131 15079
rect 29653 15045 29687 15079
rect 49433 15045 49467 15079
rect 59093 15045 59127 15079
rect 60841 15045 60875 15079
rect 63233 15045 63267 15079
rect 69213 15045 69247 15079
rect 70041 15045 70075 15079
rect 73721 15045 73755 15079
rect 77217 15045 77251 15079
rect 77309 15045 77343 15079
rect 77861 15045 77895 15079
rect 84025 15045 84059 15079
rect 22201 14977 22235 15011
rect 22845 14977 22879 15011
rect 23489 14977 23523 15011
rect 24317 14977 24351 15011
rect 31033 14977 31067 15011
rect 31401 14977 31435 15011
rect 32873 14977 32907 15011
rect 33149 14977 33183 15011
rect 33885 14977 33919 15011
rect 34989 14977 35023 15011
rect 36093 14977 36127 15011
rect 36921 14977 36955 15011
rect 38117 14977 38151 15011
rect 38485 14977 38519 15011
rect 39221 14977 39255 15011
rect 39313 14977 39347 15011
rect 40325 14977 40359 15011
rect 40877 14977 40911 15011
rect 41705 14977 41739 15011
rect 43453 14977 43487 15011
rect 45937 14977 45971 15011
rect 48053 14977 48087 15011
rect 49157 14977 49191 15011
rect 54769 14977 54803 15011
rect 61117 14977 61151 15011
rect 61577 14977 61611 15011
rect 64337 14977 64371 15011
rect 67189 14977 67223 15011
rect 68569 14977 68603 15011
rect 69121 14977 69155 15011
rect 72157 14977 72191 15011
rect 75837 14977 75871 15011
rect 78873 14977 78907 15011
rect 80621 14977 80655 15011
rect 82553 14977 82587 15011
rect 82921 14977 82955 15011
rect 86877 14977 86911 15011
rect 19073 14909 19107 14943
rect 25881 14909 25915 14943
rect 29929 14909 29963 14943
rect 30481 14909 30515 14943
rect 34345 14909 34379 14943
rect 34897 14909 34931 14943
rect 37473 14909 37507 14943
rect 45845 14909 45879 14943
rect 46673 14909 46707 14943
rect 48329 14909 48363 14943
rect 54493 14909 54527 14943
rect 55229 14909 55263 14943
rect 55505 14909 55539 14943
rect 56977 14909 57011 14943
rect 64889 14909 64923 14943
rect 65165 14909 65199 14943
rect 69765 14909 69799 14943
rect 73629 14909 73663 14943
rect 80713 14909 80747 14943
rect 83933 14909 83967 14943
rect 85681 14909 85715 14943
rect 87981 14909 88015 14943
rect 12725 14841 12759 14875
rect 23397 14841 23431 14875
rect 72433 14841 72467 14875
rect 74181 14841 74215 14875
rect 75285 14841 75319 14875
rect 84485 14841 84519 14875
rect 14657 14773 14691 14807
rect 22661 14773 22695 14807
rect 36001 14773 36035 14807
rect 40233 14773 40267 14807
rect 40969 14773 41003 14807
rect 41613 14773 41647 14807
rect 42901 14773 42935 14807
rect 44741 14773 44775 14807
rect 50905 14773 50939 14807
rect 51549 14773 51583 14807
rect 52009 14773 52043 14807
rect 58173 14773 58207 14807
rect 61669 14773 61703 14807
rect 63877 14773 63911 14807
rect 66637 14773 66671 14807
rect 68477 14773 68511 14807
rect 74733 14773 74767 14807
rect 76389 14773 76423 14807
rect 78781 14773 78815 14807
rect 79333 14773 79367 14807
rect 80345 14773 80379 14807
rect 81357 14773 81391 14807
rect 85221 14773 85255 14807
rect 86417 14773 86451 14807
rect 87429 14773 87463 14807
rect 89085 14773 89119 14807
rect 89545 14773 89579 14807
rect 90097 14773 90131 14807
rect 90741 14773 90775 14807
rect 24593 14569 24627 14603
rect 46305 14569 46339 14603
rect 56241 14569 56275 14603
rect 81265 14569 81299 14603
rect 92673 14569 92707 14603
rect 11805 14501 11839 14535
rect 28917 14501 28951 14535
rect 63233 14501 63267 14535
rect 71513 14501 71547 14535
rect 83841 14501 83875 14535
rect 11345 14433 11379 14467
rect 12449 14433 12483 14467
rect 19441 14433 19475 14467
rect 19717 14433 19751 14467
rect 21465 14433 21499 14467
rect 27445 14433 27479 14467
rect 31861 14433 31895 14467
rect 32045 14433 32079 14467
rect 40601 14433 40635 14467
rect 44097 14433 44131 14467
rect 48605 14433 48639 14467
rect 55873 14433 55907 14467
rect 60657 14433 60691 14467
rect 71053 14433 71087 14467
rect 76941 14433 76975 14467
rect 78965 14433 78999 14467
rect 83565 14433 83599 14467
rect 88441 14433 88475 14467
rect 7297 14365 7331 14399
rect 8033 14365 8067 14399
rect 11437 14365 11471 14399
rect 12541 14365 12575 14399
rect 15669 14365 15703 14399
rect 23765 14365 23799 14399
rect 24777 14365 24811 14399
rect 25697 14365 25731 14399
rect 27169 14365 27203 14399
rect 29837 14365 29871 14399
rect 30481 14365 30515 14399
rect 35173 14365 35207 14399
rect 37105 14365 37139 14399
rect 37381 14365 37415 14399
rect 38301 14365 38335 14399
rect 38853 14365 38887 14399
rect 40325 14365 40359 14399
rect 42625 14365 42659 14399
rect 43821 14365 43855 14399
rect 45477 14365 45511 14399
rect 46213 14365 46247 14399
rect 49249 14365 49283 14399
rect 50997 14365 51031 14399
rect 51549 14365 51583 14399
rect 54033 14365 54067 14399
rect 55965 14365 55999 14399
rect 59921 14365 59955 14399
rect 62681 14365 62715 14399
rect 65257 14365 65291 14399
rect 66085 14365 66119 14399
rect 66637 14365 66671 14399
rect 67741 14365 67775 14399
rect 68201 14365 68235 14399
rect 71145 14365 71179 14399
rect 72157 14365 72191 14399
rect 79609 14365 79643 14399
rect 80069 14365 80103 14399
rect 82369 14365 82403 14399
rect 83473 14365 83507 14399
rect 84945 14365 84979 14399
rect 86785 14365 86819 14399
rect 87061 14365 87095 14399
rect 88533 14365 88567 14399
rect 89361 14365 89395 14399
rect 9229 14297 9263 14331
rect 13093 14297 13127 14331
rect 23489 14297 23523 14331
rect 33701 14297 33735 14331
rect 36001 14297 36035 14331
rect 38209 14297 38243 14331
rect 39129 14297 39163 14331
rect 46857 14297 46891 14331
rect 51825 14297 51859 14331
rect 53941 14297 53975 14331
rect 57253 14297 57287 14331
rect 58817 14297 58851 14331
rect 59369 14297 59403 14331
rect 62405 14297 62439 14331
rect 67649 14297 67683 14331
rect 68477 14297 68511 14331
rect 72709 14297 72743 14331
rect 78689 14297 78723 14331
rect 84393 14297 84427 14331
rect 89269 14297 89303 14331
rect 14565 14229 14599 14263
rect 15577 14229 15611 14263
rect 16221 14229 16255 14263
rect 22017 14229 22051 14263
rect 25605 14229 25639 14263
rect 26617 14229 26651 14263
rect 29929 14229 29963 14263
rect 30573 14229 30607 14263
rect 31401 14229 31435 14263
rect 34253 14229 34287 14263
rect 35081 14229 35115 14263
rect 36553 14229 36587 14263
rect 42073 14229 42107 14263
rect 42717 14229 42751 14263
rect 44649 14229 44683 14263
rect 45385 14229 45419 14263
rect 49157 14229 49191 14263
rect 49709 14229 49743 14263
rect 50353 14229 50387 14263
rect 53297 14229 53331 14263
rect 54585 14229 54619 14263
rect 60013 14229 60047 14263
rect 63693 14229 63727 14263
rect 64245 14229 64279 14263
rect 65165 14229 65199 14263
rect 65901 14229 65935 14263
rect 69949 14229 69983 14263
rect 72065 14229 72099 14263
rect 73997 14229 74031 14263
rect 75009 14229 75043 14263
rect 75561 14229 75595 14263
rect 76205 14229 76239 14263
rect 79517 14229 79551 14263
rect 80161 14229 80195 14263
rect 81817 14229 81851 14263
rect 85037 14229 85071 14263
rect 85589 14229 85623 14263
rect 86417 14229 86451 14263
rect 88165 14229 88199 14263
rect 90005 14229 90039 14263
rect 90557 14229 90591 14263
rect 91569 14229 91603 14263
rect 92213 14229 92247 14263
rect 20545 14025 20579 14059
rect 22477 14025 22511 14059
rect 27721 14025 27755 14059
rect 47225 14025 47259 14059
rect 58265 14025 58299 14059
rect 67465 14025 67499 14059
rect 74825 14025 74859 14059
rect 76205 14025 76239 14059
rect 80989 14025 81023 14059
rect 82645 14025 82679 14059
rect 88257 14025 88291 14059
rect 92765 14025 92799 14059
rect 7757 13957 7791 13991
rect 9321 13957 9355 13991
rect 16957 13957 16991 13991
rect 23765 13957 23799 13991
rect 24593 13957 24627 13991
rect 35449 13957 35483 13991
rect 39221 13957 39255 13991
rect 43729 13957 43763 13991
rect 49985 13957 50019 13991
rect 51089 13957 51123 13991
rect 53021 13957 53055 13991
rect 59277 13957 59311 13991
rect 61025 13957 61059 13991
rect 62405 13957 62439 13991
rect 75561 13957 75595 13991
rect 78965 13957 78999 13991
rect 89269 13957 89303 13991
rect 2973 13889 3007 13923
rect 3893 13889 3927 13923
rect 8585 13889 8619 13923
rect 11897 13889 11931 13923
rect 13277 13889 13311 13923
rect 13921 13889 13955 13923
rect 14933 13889 14967 13923
rect 15945 13889 15979 13923
rect 21281 13889 21315 13923
rect 27629 13889 27663 13923
rect 30113 13889 30147 13923
rect 30849 13889 30883 13923
rect 31769 13889 31803 13923
rect 32505 13889 32539 13923
rect 33149 13889 33183 13923
rect 36369 13889 36403 13923
rect 38485 13889 38519 13923
rect 38945 13889 38979 13923
rect 40969 13889 41003 13923
rect 41691 13889 41725 13923
rect 42717 13889 42751 13923
rect 42901 13889 42935 13923
rect 44557 13889 44591 13923
rect 45477 13889 45511 13923
rect 47777 13889 47811 13923
rect 52929 13889 52963 13923
rect 53757 13889 53791 13923
rect 55045 13889 55079 13923
rect 57069 13889 57103 13923
rect 58081 13889 58115 13923
rect 61301 13889 61335 13923
rect 63601 13889 63635 13923
rect 68937 13889 68971 13923
rect 69305 13889 69339 13923
rect 72617 13889 72651 13923
rect 73537 13889 73571 13923
rect 75653 13889 75687 13923
rect 76113 13889 76147 13923
rect 76941 13889 76975 13923
rect 77401 13889 77435 13923
rect 77493 13889 77527 13923
rect 78689 13889 78723 13923
rect 83197 13889 83231 13923
rect 85313 13889 85347 13923
rect 86233 13889 86267 13923
rect 87153 13889 87187 13923
rect 91845 13889 91879 13923
rect 92581 13889 92615 13923
rect 8217 13821 8251 13855
rect 8493 13821 8527 13855
rect 11161 13821 11195 13855
rect 11989 13821 12023 13855
rect 14013 13821 14047 13855
rect 15025 13821 15059 13855
rect 15853 13821 15887 13855
rect 18797 13821 18831 13855
rect 19073 13821 19107 13855
rect 21373 13821 21407 13855
rect 26341 13821 26375 13855
rect 26617 13821 26651 13855
rect 28365 13821 28399 13855
rect 32413 13821 32447 13855
rect 33977 13821 34011 13855
rect 35633 13821 35667 13855
rect 36921 13821 36955 13855
rect 37749 13821 37783 13855
rect 38393 13821 38427 13855
rect 41613 13821 41647 13855
rect 44833 13821 44867 13855
rect 45753 13821 45787 13855
rect 49525 13821 49559 13855
rect 54217 13821 54251 13855
rect 61761 13821 61795 13855
rect 64061 13821 64095 13855
rect 66453 13821 66487 13855
rect 66913 13821 66947 13855
rect 70869 13821 70903 13855
rect 73629 13821 73663 13855
rect 78137 13821 78171 13855
rect 83841 13821 83875 13855
rect 84945 13821 84979 13855
rect 87705 13821 87739 13855
rect 88993 13821 89027 13855
rect 91293 13821 91327 13855
rect 12265 13753 12299 13787
rect 14289 13753 14323 13787
rect 15301 13753 15335 13787
rect 41981 13753 42015 13787
rect 58817 13753 58851 13787
rect 74273 13753 74307 13787
rect 81541 13753 81575 13787
rect 4813 13685 4847 13719
rect 6653 13685 6687 13719
rect 17417 13685 17451 13719
rect 29855 13685 29889 13719
rect 30757 13685 30791 13719
rect 33241 13685 33275 13719
rect 48034 13685 48068 13719
rect 50537 13685 50571 13719
rect 51641 13685 51675 13719
rect 52193 13685 52227 13719
rect 53665 13685 53699 13719
rect 56805 13685 56839 13719
rect 63509 13685 63543 13719
rect 64705 13685 64739 13719
rect 66195 13685 66229 13719
rect 68385 13685 68419 13719
rect 72353 13685 72387 13719
rect 76849 13685 76883 13719
rect 80437 13685 80471 13719
rect 82093 13685 82127 13719
rect 90741 13685 90775 13719
rect 93225 13685 93259 13719
rect 94145 13685 94179 13719
rect 5089 13481 5123 13515
rect 21189 13481 21223 13515
rect 27537 13481 27571 13515
rect 28457 13481 28491 13515
rect 31493 13481 31527 13515
rect 36001 13481 36035 13515
rect 37289 13481 37323 13515
rect 38209 13481 38243 13515
rect 44373 13481 44407 13515
rect 52837 13481 52871 13515
rect 65165 13481 65199 13515
rect 69949 13481 69983 13515
rect 71053 13481 71087 13515
rect 76113 13481 76147 13515
rect 79425 13481 79459 13515
rect 81817 13481 81851 13515
rect 85221 13481 85255 13515
rect 89177 13481 89211 13515
rect 89821 13481 89855 13515
rect 5733 13413 5767 13447
rect 7481 13413 7515 13447
rect 13461 13413 13495 13447
rect 41153 13413 41187 13447
rect 66637 13413 66671 13447
rect 73353 13413 73387 13447
rect 78781 13413 78815 13447
rect 85681 13413 85715 13447
rect 86693 13413 86727 13447
rect 2973 13345 3007 13379
rect 4077 13345 4111 13379
rect 8125 13345 8159 13379
rect 9781 13345 9815 13379
rect 12081 13345 12115 13379
rect 14565 13345 14599 13379
rect 16313 13345 16347 13379
rect 23949 13345 23983 13379
rect 25421 13345 25455 13379
rect 32689 13345 32723 13379
rect 45201 13345 45235 13379
rect 47409 13345 47443 13379
rect 49709 13345 49743 13379
rect 50445 13345 50479 13379
rect 54309 13345 54343 13379
rect 59001 13345 59035 13379
rect 75561 13345 75595 13379
rect 80069 13345 80103 13379
rect 82921 13345 82955 13379
rect 84669 13345 84703 13379
rect 87705 13345 87739 13379
rect 90465 13345 90499 13379
rect 93593 13345 93627 13379
rect 3065 13277 3099 13311
rect 4169 13277 4203 13311
rect 5825 13277 5859 13311
rect 6009 13277 6043 13311
rect 8217 13277 8251 13311
rect 10149 13277 10183 13311
rect 10517 13277 10551 13311
rect 12633 13277 12667 13311
rect 14289 13277 14323 13311
rect 17049 13277 17083 13311
rect 18245 13277 18279 13311
rect 18889 13277 18923 13311
rect 19441 13277 19475 13311
rect 22201 13277 22235 13311
rect 25145 13277 25179 13311
rect 26065 13277 26099 13311
rect 28273 13277 28307 13311
rect 29745 13277 29779 13311
rect 32505 13277 32539 13311
rect 35449 13277 35483 13311
rect 36093 13277 36127 13311
rect 36737 13277 36771 13311
rect 40233 13277 40267 13311
rect 42441 13277 42475 13311
rect 49617 13277 49651 13311
rect 51825 13277 51859 13311
rect 54585 13277 54619 13311
rect 56149 13277 56183 13311
rect 56425 13277 56459 13311
rect 59645 13277 59679 13311
rect 60657 13277 60691 13311
rect 61577 13277 61611 13311
rect 62221 13277 62255 13311
rect 64705 13277 64739 13311
rect 65993 13277 66027 13311
rect 66453 13277 66487 13311
rect 69397 13277 69431 13311
rect 69857 13277 69891 13311
rect 71145 13277 71179 13311
rect 71605 13277 71639 13311
rect 73813 13277 73847 13311
rect 76297 13277 76331 13311
rect 77033 13277 77067 13311
rect 79517 13277 79551 13311
rect 79969 13277 80003 13311
rect 86693 13277 86727 13311
rect 87429 13277 87463 13311
rect 89729 13277 89763 13311
rect 90557 13277 90591 13311
rect 18153 13209 18187 13243
rect 19717 13209 19751 13243
rect 22477 13209 22511 13243
rect 24593 13209 24627 13243
rect 30021 13209 30055 13243
rect 34345 13209 34379 13243
rect 39497 13209 39531 13243
rect 42901 13209 42935 13243
rect 45477 13209 45511 13243
rect 47685 13209 47719 13243
rect 52101 13209 52135 13243
rect 57253 13209 57287 13243
rect 62497 13209 62531 13243
rect 67833 13209 67867 13243
rect 71881 13209 71915 13243
rect 77309 13209 77343 13243
rect 82369 13209 82403 13243
rect 83197 13209 83231 13243
rect 93317 13209 93351 13243
rect 3433 13141 3467 13175
rect 4537 13141 4571 13175
rect 6929 13141 6963 13175
rect 8585 13141 8619 13175
rect 16865 13141 16899 13175
rect 17601 13141 17635 13175
rect 18797 13141 18831 13175
rect 29193 13141 29227 13175
rect 32045 13141 32079 13175
rect 35357 13141 35391 13175
rect 40141 13141 40175 13175
rect 46949 13141 46983 13175
rect 49157 13141 49191 13175
rect 50997 13141 51031 13175
rect 56793 13141 56827 13175
rect 59553 13141 59587 13175
rect 60749 13141 60783 13175
rect 61669 13141 61703 13175
rect 63969 13141 64003 13175
rect 64613 13141 64647 13175
rect 65901 13141 65935 13175
rect 67097 13141 67131 13175
rect 80621 13141 80655 13175
rect 81357 13141 81391 13175
rect 91845 13141 91879 13175
rect 94053 13141 94087 13175
rect 4445 12937 4479 12971
rect 6561 12937 6595 12971
rect 9965 12937 9999 12971
rect 11897 12937 11931 12971
rect 30481 12937 30515 12971
rect 45477 12937 45511 12971
rect 47777 12937 47811 12971
rect 53389 12937 53423 12971
rect 56793 12937 56827 12971
rect 61577 12937 61611 12971
rect 64981 12937 65015 12971
rect 66545 12937 66579 12971
rect 76941 12937 76975 12971
rect 83933 12937 83967 12971
rect 84669 12937 84703 12971
rect 87797 12937 87831 12971
rect 93317 12937 93351 12971
rect 14749 12869 14783 12903
rect 16957 12869 16991 12903
rect 21097 12869 21131 12903
rect 24501 12869 24535 12903
rect 29285 12869 29319 12903
rect 32873 12869 32907 12903
rect 38669 12869 38703 12903
rect 44189 12869 44223 12903
rect 54677 12869 54711 12903
rect 63509 12869 63543 12903
rect 70777 12869 70811 12903
rect 75745 12869 75779 12903
rect 77769 12869 77803 12903
rect 94237 12869 94271 12903
rect 3801 12801 3835 12835
rect 4997 12801 5031 12835
rect 6929 12801 6963 12835
rect 7757 12801 7791 12835
rect 8585 12801 8619 12835
rect 9597 12801 9631 12835
rect 11713 12801 11747 12835
rect 13921 12801 13955 12835
rect 17969 12801 18003 12835
rect 18521 12801 18555 12835
rect 22569 12801 22603 12835
rect 25237 12807 25271 12841
rect 26249 12801 26283 12835
rect 30389 12801 30423 12835
rect 31585 12801 31619 12835
rect 32597 12801 32631 12835
rect 34989 12801 35023 12835
rect 35173 12801 35207 12835
rect 35909 12801 35943 12835
rect 37749 12801 37783 12835
rect 41705 12801 41739 12835
rect 42809 12801 42843 12835
rect 46765 12801 46799 12835
rect 48145 12801 48179 12835
rect 48973 12801 49007 12835
rect 49341 12801 49375 12835
rect 50905 12801 50939 12835
rect 51825 12801 51859 12835
rect 55413 12801 55447 12835
rect 58081 12801 58115 12835
rect 59093 12801 59127 12835
rect 61117 12801 61151 12835
rect 63233 12801 63267 12835
rect 65533 12801 65567 12835
rect 66453 12801 66487 12835
rect 67557 12801 67591 12835
rect 67649 12801 67683 12835
rect 68385 12801 68419 12835
rect 68661 12801 68695 12835
rect 69765 12801 69799 12835
rect 70501 12801 70535 12835
rect 73629 12801 73663 12835
rect 75193 12801 75227 12835
rect 75653 12801 75687 12835
rect 76757 12801 76791 12835
rect 77493 12801 77527 12835
rect 81909 12801 81943 12835
rect 82277 12801 82311 12835
rect 84117 12801 84151 12835
rect 84761 12801 84795 12835
rect 85497 12801 85531 12835
rect 86233 12801 86267 12835
rect 86877 12801 86911 12835
rect 87705 12801 87739 12835
rect 89453 12801 89487 12835
rect 89545 12801 89579 12835
rect 90741 12801 90775 12835
rect 91109 12801 91143 12835
rect 92581 12801 92615 12835
rect 92765 12801 92799 12835
rect 93225 12801 93259 12835
rect 94145 12801 94179 12835
rect 3893 12733 3927 12767
rect 7021 12733 7055 12767
rect 7849 12733 7883 12767
rect 8125 12733 8159 12767
rect 9505 12733 9539 12767
rect 14473 12733 14507 12767
rect 24777 12733 24811 12767
rect 25329 12733 25363 12767
rect 26341 12733 26375 12767
rect 26617 12733 26651 12767
rect 27445 12733 27479 12767
rect 27629 12733 27663 12767
rect 29837 12733 29871 12767
rect 31677 12733 31711 12767
rect 36185 12733 36219 12767
rect 38393 12733 38427 12767
rect 40141 12733 40175 12767
rect 41797 12733 41831 12767
rect 42901 12733 42935 12767
rect 47041 12733 47075 12767
rect 48053 12733 48087 12767
rect 50077 12733 50111 12767
rect 50997 12733 51031 12767
rect 51917 12733 51951 12767
rect 55321 12733 55355 12767
rect 56241 12733 56275 12767
rect 58173 12733 58207 12767
rect 59369 12733 59403 12767
rect 62129 12733 62163 12767
rect 69305 12733 69339 12767
rect 72525 12733 72559 12767
rect 80161 12733 80195 12767
rect 80437 12733 80471 12767
rect 86785 12733 86819 12767
rect 88349 12733 88383 12767
rect 35173 12665 35207 12699
rect 43177 12665 43211 12699
rect 65717 12665 65751 12699
rect 68661 12665 68695 12699
rect 87245 12665 87279 12699
rect 5273 12597 5307 12631
rect 6009 12597 6043 12631
rect 13185 12597 13219 12631
rect 13829 12597 13863 12631
rect 16221 12597 16255 12631
rect 17049 12597 17083 12631
rect 17877 12597 17911 12631
rect 18613 12597 18647 12631
rect 19625 12597 19659 12631
rect 22477 12597 22511 12631
rect 23029 12597 23063 12631
rect 31309 12597 31343 12631
rect 34345 12597 34379 12631
rect 36921 12597 36955 12631
rect 37841 12597 37875 12631
rect 41061 12597 41095 12631
rect 41981 12597 42015 12631
rect 43729 12597 43763 12631
rect 52193 12597 52227 12631
rect 57345 12597 57379 12631
rect 69949 12597 69983 12631
rect 73721 12597 73755 12631
rect 74273 12597 74307 12631
rect 75009 12597 75043 12631
rect 78689 12597 78723 12631
rect 81541 12597 81575 12631
rect 85405 12597 85439 12631
rect 86141 12597 86175 12631
rect 90189 12597 90223 12631
rect 92765 12597 92799 12631
rect 21189 12393 21223 12427
rect 21833 12393 21867 12427
rect 24869 12393 24903 12427
rect 29929 12393 29963 12427
rect 30849 12393 30883 12427
rect 34989 12393 35023 12427
rect 37749 12393 37783 12427
rect 40325 12393 40359 12427
rect 42717 12393 42751 12427
rect 49617 12393 49651 12427
rect 53389 12393 53423 12427
rect 59369 12393 59403 12427
rect 61577 12393 61611 12427
rect 80253 12393 80287 12427
rect 84117 12393 84151 12427
rect 89729 12393 89763 12427
rect 93317 12393 93351 12427
rect 94237 12393 94271 12427
rect 24041 12325 24075 12359
rect 29193 12325 29227 12359
rect 33425 12325 33459 12359
rect 54677 12325 54711 12359
rect 58817 12325 58851 12359
rect 66545 12325 66579 12359
rect 78045 12325 78079 12359
rect 79609 12325 79643 12359
rect 81265 12325 81299 12359
rect 3341 12257 3375 12291
rect 8033 12257 8067 12291
rect 13737 12257 13771 12291
rect 15853 12257 15887 12291
rect 18521 12257 18555 12291
rect 19441 12257 19475 12291
rect 19717 12257 19751 12291
rect 22293 12257 22327 12291
rect 22569 12257 22603 12291
rect 26341 12257 26375 12291
rect 28181 12257 28215 12291
rect 30297 12257 30331 12291
rect 31125 12257 31159 12291
rect 33701 12257 33735 12291
rect 37013 12257 37047 12291
rect 39221 12257 39255 12291
rect 39497 12257 39531 12291
rect 42073 12257 42107 12291
rect 46213 12257 46247 12291
rect 46489 12257 46523 12291
rect 54033 12257 54067 12291
rect 56517 12257 56551 12291
rect 62681 12257 62715 12291
rect 62957 12257 62991 12291
rect 73537 12257 73571 12291
rect 75561 12257 75595 12291
rect 77125 12257 77159 12291
rect 78505 12257 78539 12291
rect 81725 12257 81759 12291
rect 85589 12257 85623 12291
rect 85865 12257 85899 12291
rect 87613 12257 87647 12291
rect 91845 12257 91879 12291
rect 3249 12189 3283 12223
rect 5089 12189 5123 12223
rect 8493 12189 8527 12223
rect 16129 12189 16163 12223
rect 21649 12189 21683 12223
rect 26249 12189 26283 12223
rect 27077 12189 27111 12223
rect 27997 12189 28031 12223
rect 30205 12189 30239 12223
rect 31217 12189 31251 12223
rect 31953 12189 31987 12223
rect 32137 12189 32171 12223
rect 33793 12189 33827 12223
rect 35081 12189 35115 12223
rect 37289 12189 37323 12223
rect 42533 12189 42567 12223
rect 43821 12189 43855 12223
rect 44005 12189 44039 12223
rect 45377 12189 45411 12223
rect 46029 12189 46063 12223
rect 48513 12189 48547 12223
rect 49433 12189 49467 12223
rect 49525 12189 49559 12223
rect 50629 12189 50663 12223
rect 51181 12189 51215 12223
rect 56425 12189 56459 12223
rect 57161 12189 57195 12223
rect 57345 12189 57379 12223
rect 57805 12189 57839 12223
rect 57989 12189 58023 12223
rect 58909 12189 58943 12223
rect 60657 12189 60691 12223
rect 65993 12189 66027 12223
rect 66637 12189 66671 12223
rect 67281 12189 67315 12223
rect 67373 12189 67407 12223
rect 67925 12189 67959 12223
rect 70409 12189 70443 12223
rect 73077 12189 73111 12223
rect 76297 12189 76331 12223
rect 76389 12189 76423 12223
rect 77033 12189 77067 12223
rect 77217 12189 77251 12223
rect 77309 12189 77343 12223
rect 77953 12189 77987 12223
rect 78321 12189 78355 12223
rect 78965 12189 78999 12223
rect 81633 12189 81667 12223
rect 82277 12189 82311 12223
rect 83013 12189 83047 12223
rect 86601 12189 86635 12223
rect 87705 12189 87739 12223
rect 90373 12189 90407 12223
rect 90649 12189 90683 12223
rect 91569 12189 91603 12223
rect 94053 12189 94087 12223
rect 4353 12121 4387 12155
rect 6101 12121 6135 12155
rect 13461 12121 13495 12155
rect 18245 12121 18279 12155
rect 27353 12121 27387 12155
rect 41797 12121 41831 12155
rect 44557 12121 44591 12155
rect 48789 12121 48823 12155
rect 53757 12121 53791 12155
rect 57253 12121 57287 12155
rect 57897 12121 57931 12155
rect 61853 12121 61887 12155
rect 62037 12121 62071 12155
rect 62129 12121 62163 12155
rect 64705 12121 64739 12155
rect 68201 12121 68235 12155
rect 72801 12121 72835 12155
rect 73813 12121 73847 12155
rect 79057 12121 79091 12155
rect 83565 12121 83599 12155
rect 87061 12121 87095 12155
rect 2881 12053 2915 12087
rect 6009 12053 6043 12087
rect 6837 12053 6871 12087
rect 7297 12053 7331 12087
rect 11989 12053 12023 12087
rect 14381 12053 14415 12087
rect 16773 12053 16807 12087
rect 25421 12053 25455 12087
rect 25881 12053 25915 12087
rect 32965 12053 32999 12087
rect 35541 12053 35575 12087
rect 45477 12053 45511 12087
rect 49801 12053 49835 12087
rect 53849 12053 53883 12087
rect 55597 12053 55631 12087
rect 59921 12053 59955 12087
rect 60749 12053 60783 12087
rect 65165 12053 65199 12087
rect 65901 12053 65935 12087
rect 69673 12053 69707 12087
rect 70317 12053 70351 12087
rect 71329 12053 71363 12087
rect 77493 12053 77527 12087
rect 82369 12053 82403 12087
rect 86509 12053 86543 12087
rect 88625 12053 88659 12087
rect 89177 12053 89211 12087
rect 4537 11849 4571 11883
rect 9689 11849 9723 11883
rect 14013 11849 14047 11883
rect 16313 11849 16347 11883
rect 29101 11849 29135 11883
rect 36553 11849 36587 11883
rect 41061 11849 41095 11883
rect 41429 11849 41463 11883
rect 42625 11849 42659 11883
rect 43821 11849 43855 11883
rect 52009 11849 52043 11883
rect 53021 11849 53055 11883
rect 61577 11849 61611 11883
rect 65625 11849 65659 11883
rect 73629 11849 73663 11883
rect 78781 11849 78815 11883
rect 85221 11849 85255 11883
rect 94237 11849 94271 11883
rect 3065 11781 3099 11815
rect 8217 11781 8251 11815
rect 21465 11781 21499 11815
rect 22293 11781 22327 11815
rect 24317 11781 24351 11815
rect 26433 11781 26467 11815
rect 30665 11781 30699 11815
rect 39037 11781 39071 11815
rect 40601 11781 40635 11815
rect 41521 11781 41555 11815
rect 46581 11781 46615 11815
rect 51273 11781 51307 11815
rect 57529 11781 57563 11815
rect 63601 11781 63635 11815
rect 68385 11781 68419 11815
rect 74181 11781 74215 11815
rect 75469 11781 75503 11815
rect 79609 11781 79643 11815
rect 80161 11781 80195 11815
rect 80529 11781 80563 11815
rect 81817 11781 81851 11815
rect 89085 11781 89119 11815
rect 90097 11781 90131 11815
rect 6745 11713 6779 11747
rect 10149 11713 10183 11747
rect 13093 11713 13127 11747
rect 13921 11713 13955 11747
rect 17141 11713 17175 11747
rect 17693 11713 17727 11747
rect 20177 11713 20211 11747
rect 20453 11713 20487 11747
rect 27537 11713 27571 11747
rect 29469 11713 29503 11747
rect 30399 11713 30433 11747
rect 33977 11713 34011 11747
rect 34161 11713 34195 11747
rect 35265 11713 35299 11747
rect 35541 11713 35575 11747
rect 36645 11713 36679 11747
rect 38025 11713 38059 11747
rect 42993 11713 43027 11747
rect 52193 11713 52227 11747
rect 52377 11713 52411 11747
rect 52929 11713 52963 11747
rect 53113 11713 53147 11747
rect 54401 11713 54435 11747
rect 55045 11713 55079 11747
rect 56149 11713 56183 11747
rect 56701 11713 56735 11747
rect 57345 11713 57379 11747
rect 58265 11713 58299 11747
rect 58428 11713 58462 11747
rect 58541 11713 58575 11747
rect 58679 11713 58713 11747
rect 61945 11713 61979 11747
rect 62405 11713 62439 11747
rect 63325 11713 63359 11747
rect 67373 11713 67407 11747
rect 67557 11713 67591 11747
rect 71145 11713 71179 11747
rect 71237 11713 71271 11747
rect 72157 11713 72191 11747
rect 72341 11713 72375 11747
rect 72433 11713 72467 11747
rect 72709 11713 72743 11747
rect 73537 11713 73571 11747
rect 75377 11713 75411 11747
rect 75561 11713 75595 11747
rect 76021 11713 76055 11747
rect 76757 11713 76791 11747
rect 76941 11713 76975 11747
rect 77217 11713 77251 11747
rect 77401 11713 77435 11747
rect 77861 11713 77895 11747
rect 78045 11713 78079 11747
rect 79057 11713 79091 11747
rect 80621 11713 80655 11747
rect 80713 11713 80747 11747
rect 84209 11713 84243 11747
rect 84945 11713 84979 11747
rect 89177 11713 89211 11747
rect 92121 11713 92155 11747
rect 92305 11713 92339 11747
rect 94145 11713 94179 11747
rect 2789 11645 2823 11679
rect 6653 11645 6687 11679
rect 7941 11645 7975 11679
rect 10425 11645 10459 11679
rect 12265 11645 12299 11679
rect 13185 11645 13219 11679
rect 14565 11645 14599 11679
rect 14841 11645 14875 11679
rect 17233 11645 17267 11679
rect 17969 11645 18003 11679
rect 19717 11645 19751 11679
rect 22017 11645 22051 11679
rect 25053 11645 25087 11679
rect 26617 11645 26651 11679
rect 27445 11645 27479 11679
rect 28549 11645 28583 11679
rect 29377 11645 29411 11679
rect 33241 11645 33275 11679
rect 35817 11645 35851 11679
rect 39773 11645 39807 11679
rect 41613 11645 41647 11679
rect 43085 11645 43119 11679
rect 44373 11645 44407 11679
rect 44925 11645 44959 11679
rect 46765 11645 46799 11679
rect 48513 11645 48547 11679
rect 49341 11645 49375 11679
rect 50445 11645 50479 11679
rect 53757 11645 53791 11679
rect 57161 11645 57195 11679
rect 65073 11645 65107 11679
rect 66545 11645 66579 11679
rect 70593 11645 70627 11679
rect 72525 11645 72559 11679
rect 74733 11645 74767 11679
rect 80897 11645 80931 11679
rect 81541 11645 81575 11679
rect 83841 11645 83875 11679
rect 84301 11645 84335 11679
rect 87705 11645 87739 11679
rect 87981 11645 88015 11679
rect 89821 11645 89855 11679
rect 91569 11645 91603 11679
rect 93133 11645 93167 11679
rect 7113 11577 7147 11611
rect 27169 11577 27203 11611
rect 56609 11577 56643 11611
rect 59921 11577 59955 11611
rect 61025 11577 61059 11611
rect 77033 11577 77067 11611
rect 77125 11577 77159 11611
rect 1593 11509 1627 11543
rect 5089 11509 5123 11543
rect 5549 11509 5583 11543
rect 12817 11509 12851 11543
rect 23765 11509 23799 11543
rect 31769 11509 31803 11543
rect 32597 11509 32631 11543
rect 52377 11509 52411 11543
rect 58909 11509 58943 11543
rect 59369 11509 59403 11543
rect 60565 11509 60599 11543
rect 69673 11509 69707 11543
rect 72893 11509 72927 11543
rect 76205 11509 76239 11543
rect 78045 11509 78079 11543
rect 83289 11509 83323 11543
rect 86233 11509 86267 11543
rect 1777 11305 1811 11339
rect 9137 11305 9171 11339
rect 9597 11305 9631 11339
rect 11253 11305 11287 11339
rect 11989 11305 12023 11339
rect 13553 11305 13587 11339
rect 20269 11305 20303 11339
rect 27721 11305 27755 11339
rect 28549 11305 28583 11339
rect 30021 11305 30055 11339
rect 31493 11305 31527 11339
rect 39497 11305 39531 11339
rect 41981 11305 42015 11339
rect 43085 11305 43119 11339
rect 54493 11305 54527 11339
rect 56333 11305 56367 11339
rect 63601 11305 63635 11339
rect 64889 11305 64923 11339
rect 74089 11305 74123 11339
rect 76941 11305 76975 11339
rect 77401 11305 77435 11339
rect 78873 11305 78907 11339
rect 79517 11305 79551 11339
rect 84623 11305 84657 11339
rect 85221 11305 85255 11339
rect 87981 11305 88015 11339
rect 90557 11305 90591 11339
rect 93317 11305 93351 11339
rect 19533 11237 19567 11271
rect 30665 11237 30699 11271
rect 54677 11237 54711 11271
rect 55873 11237 55907 11271
rect 56977 11237 57011 11271
rect 58725 11237 58759 11271
rect 66361 11237 66395 11271
rect 70041 11237 70075 11271
rect 74365 11237 74399 11271
rect 76205 11237 76239 11271
rect 84485 11237 84519 11271
rect 85773 11237 85807 11271
rect 88717 11237 88751 11271
rect 5181 11169 5215 11203
rect 7573 11169 7607 11203
rect 8493 11169 8527 11203
rect 9413 11169 9447 11203
rect 10701 11169 10735 11203
rect 13185 11169 13219 11203
rect 21649 11169 21683 11203
rect 23121 11169 23155 11203
rect 26249 11169 26283 11203
rect 34253 11169 34287 11203
rect 38025 11169 38059 11203
rect 38301 11169 38335 11203
rect 44005 11169 44039 11203
rect 44649 11169 44683 11203
rect 48973 11169 49007 11203
rect 58633 11169 58667 11203
rect 58854 11169 58888 11203
rect 60749 11169 60783 11203
rect 60933 11169 60967 11203
rect 61853 11169 61887 11203
rect 62129 11169 62163 11203
rect 65901 11169 65935 11203
rect 69765 11169 69799 11203
rect 76665 11169 76699 11203
rect 76757 11169 76791 11203
rect 77666 11169 77700 11203
rect 77861 11169 77895 11203
rect 84393 11169 84427 11203
rect 86601 11169 86635 11203
rect 89269 11169 89303 11203
rect 91845 11169 91879 11203
rect 93869 11169 93903 11203
rect 2237 11101 2271 11135
rect 2513 11101 2547 11135
rect 3249 11101 3283 11135
rect 3985 11101 4019 11135
rect 4261 11101 4295 11135
rect 4905 11101 4939 11135
rect 6377 11101 6411 11135
rect 8401 11101 8435 11135
rect 9689 11101 9723 11135
rect 13277 11101 13311 11135
rect 15393 11101 15427 11135
rect 16589 11101 16623 11135
rect 17141 11101 17175 11135
rect 18797 11101 18831 11135
rect 19441 11101 19475 11135
rect 19625 11101 19659 11135
rect 20085 11101 20119 11135
rect 21373 11101 21407 11135
rect 24961 11101 24995 11135
rect 25973 11101 26007 11135
rect 32505 11101 32539 11135
rect 35357 11101 35391 11135
rect 38393 11101 38427 11135
rect 40509 11101 40543 11135
rect 41429 11101 41463 11135
rect 42441 11101 42475 11135
rect 43821 11101 43855 11135
rect 45569 11101 45603 11135
rect 46765 11101 46799 11135
rect 47501 11101 47535 11135
rect 49433 11101 49467 11135
rect 49617 11101 49651 11135
rect 49709 11101 49743 11135
rect 50353 11101 50387 11135
rect 50629 11101 50663 11135
rect 51273 11101 51307 11135
rect 51457 11101 51491 11135
rect 52009 11101 52043 11135
rect 52837 11101 52871 11135
rect 56057 11101 56091 11135
rect 56149 11101 56183 11135
rect 56333 11101 56367 11135
rect 57345 11101 57379 11135
rect 59461 11101 59495 11135
rect 59645 11101 59679 11135
rect 61025 11101 61059 11135
rect 64337 11101 64371 11135
rect 65993 11101 66027 11135
rect 68569 11101 68603 11135
rect 68937 11101 68971 11135
rect 69673 11101 69707 11135
rect 71145 11101 71179 11135
rect 71237 11101 71271 11135
rect 72341 11101 72375 11135
rect 72709 11101 72743 11135
rect 73537 11101 73571 11135
rect 74273 11101 74307 11135
rect 74457 11101 74491 11135
rect 74549 11101 74583 11135
rect 75101 11101 75135 11135
rect 75285 11101 75319 11135
rect 75571 11101 75605 11135
rect 77585 11101 77619 11135
rect 77769 11101 77803 11135
rect 78413 11101 78447 11135
rect 78505 11101 78539 11135
rect 78689 11101 78723 11135
rect 79609 11101 79643 11135
rect 80529 11101 80563 11135
rect 81725 11101 81759 11135
rect 82553 11101 82587 11135
rect 86693 11101 86727 11135
rect 87981 11101 88015 11135
rect 90005 11101 90039 11135
rect 90465 11101 90499 11135
rect 91569 11101 91603 11135
rect 93777 11101 93811 11135
rect 6929 11033 6963 11067
rect 10241 11033 10275 11067
rect 12633 11033 12667 11067
rect 14565 11033 14599 11067
rect 25237 11033 25271 11067
rect 31217 11033 31251 11067
rect 32781 11033 32815 11067
rect 35541 11033 35575 11067
rect 37197 11033 37231 11067
rect 51365 11033 51399 11067
rect 54309 11033 54343 11067
rect 57161 11033 57195 11067
rect 58265 11033 58299 11067
rect 59001 11033 59035 11067
rect 59553 11033 59587 11067
rect 64245 11033 64279 11067
rect 67097 11033 67131 11067
rect 71881 11033 71915 11067
rect 75469 11033 75503 11067
rect 76205 11033 76239 11067
rect 84025 11033 84059 11067
rect 84761 11033 84795 11067
rect 87521 11033 87555 11067
rect 3433 10965 3467 10999
rect 5825 10965 5859 10999
rect 8033 10965 8067 10999
rect 15301 10965 15335 10999
rect 20821 10965 20855 10999
rect 24041 10965 24075 10999
rect 29193 10965 29227 10999
rect 50445 10965 50479 10999
rect 50813 10965 50847 10999
rect 54509 10965 54543 10999
rect 61393 10965 61427 10999
rect 71145 10965 71179 10999
rect 80437 10965 80471 10999
rect 89913 10965 89947 10999
rect 1777 10761 1811 10795
rect 4077 10761 4111 10795
rect 9229 10761 9263 10795
rect 11161 10761 11195 10795
rect 12265 10761 12299 10795
rect 15230 10761 15264 10795
rect 15393 10761 15427 10795
rect 18705 10761 18739 10795
rect 31217 10761 31251 10795
rect 37473 10761 37507 10795
rect 42073 10761 42107 10795
rect 48329 10761 48363 10795
rect 88441 10761 88475 10795
rect 91661 10761 91695 10795
rect 94237 10761 94271 10795
rect 7757 10693 7791 10727
rect 13001 10693 13035 10727
rect 15025 10693 15059 10727
rect 21281 10693 21315 10727
rect 26617 10693 26651 10727
rect 27997 10693 28031 10727
rect 30665 10693 30699 10727
rect 33885 10693 33919 10727
rect 35541 10693 35575 10727
rect 41337 10693 41371 10727
rect 44925 10693 44959 10727
rect 54217 10693 54251 10727
rect 55873 10693 55907 10727
rect 65441 10693 65475 10727
rect 67189 10693 67223 10727
rect 70593 10693 70627 10727
rect 72341 10693 72375 10727
rect 79609 10693 79643 10727
rect 86141 10693 86175 10727
rect 86969 10693 87003 10727
rect 89085 10693 89119 10727
rect 90189 10693 90223 10727
rect 4537 10625 4571 10659
rect 6745 10625 6779 10659
rect 7481 10625 7515 10659
rect 10057 10625 10091 10659
rect 11989 10625 12023 10659
rect 15853 10625 15887 10659
rect 17049 10625 17083 10659
rect 18061 10625 18095 10659
rect 18245 10625 18279 10659
rect 19073 10625 19107 10659
rect 19717 10625 19751 10659
rect 27261 10625 27295 10659
rect 27721 10625 27755 10659
rect 29745 10625 29779 10659
rect 31769 10625 31803 10659
rect 32597 10625 32631 10659
rect 33701 10625 33735 10659
rect 36277 10625 36311 10659
rect 36435 10625 36469 10659
rect 36645 10625 36679 10659
rect 36921 10625 36955 10659
rect 38117 10625 38151 10659
rect 38867 10625 38901 10659
rect 41521 10625 41555 10659
rect 42809 10625 42843 10659
rect 44005 10625 44039 10659
rect 44741 10625 44775 10659
rect 48513 10625 48547 10659
rect 48605 10625 48639 10659
rect 49525 10625 49559 10659
rect 49617 10625 49651 10659
rect 49893 10625 49927 10659
rect 53205 10625 53239 10659
rect 53297 10625 53331 10659
rect 53481 10625 53515 10659
rect 53665 10625 53699 10659
rect 54125 10625 54159 10659
rect 54309 10625 54343 10659
rect 54953 10625 54987 10659
rect 55781 10625 55815 10659
rect 55965 10625 55999 10659
rect 56517 10625 56551 10659
rect 57345 10625 57379 10659
rect 60749 10625 60783 10659
rect 62313 10625 62347 10659
rect 63233 10625 63267 10659
rect 67833 10625 67867 10659
rect 72985 10625 73019 10659
rect 73721 10625 73755 10659
rect 77585 10625 77619 10659
rect 78689 10625 78723 10659
rect 78781 10625 78815 10659
rect 82001 10625 82035 10659
rect 82277 10625 82311 10659
rect 83289 10625 83323 10659
rect 83841 10625 83875 10659
rect 83933 10625 83967 10659
rect 84209 10625 84243 10659
rect 84669 10625 84703 10659
rect 86049 10625 86083 10659
rect 89177 10625 89211 10659
rect 92581 10625 92615 10659
rect 94145 10625 94179 10659
rect 2329 10557 2363 10591
rect 2605 10557 2639 10591
rect 4813 10557 4847 10591
rect 10149 10557 10183 10591
rect 12265 10557 12299 10591
rect 12725 10557 12759 10591
rect 14473 10557 14507 10591
rect 16037 10557 16071 10591
rect 16957 10557 16991 10591
rect 19165 10557 19199 10591
rect 22017 10557 22051 10591
rect 22293 10557 22327 10591
rect 24593 10557 24627 10591
rect 24869 10557 24903 10591
rect 32689 10557 32723 10591
rect 39037 10557 39071 10591
rect 39681 10557 39715 10591
rect 42901 10557 42935 10591
rect 43177 10557 43211 10591
rect 43913 10557 43947 10591
rect 45201 10557 45235 10591
rect 47225 10557 47259 10591
rect 48881 10557 48915 10591
rect 50445 10557 50479 10591
rect 50721 10557 50755 10591
rect 54861 10557 54895 10591
rect 57437 10557 57471 10591
rect 58081 10557 58115 10591
rect 58357 10557 58391 10591
rect 60657 10557 60691 10591
rect 61577 10557 61611 10591
rect 62129 10557 62163 10591
rect 64981 10557 65015 10591
rect 68385 10557 68419 10591
rect 68661 10557 68695 10591
rect 75193 10557 75227 10591
rect 75469 10557 75503 10591
rect 79333 10557 79367 10591
rect 81081 10557 81115 10591
rect 82645 10557 82679 10591
rect 86693 10557 86727 10591
rect 89913 10557 89947 10591
rect 92489 10557 92523 10591
rect 93225 10557 93259 10591
rect 5549 10489 5583 10523
rect 10425 10489 10459 10523
rect 12081 10489 12115 10523
rect 17417 10489 17451 10523
rect 32965 10489 32999 10523
rect 38577 10489 38611 10523
rect 43637 10489 43671 10523
rect 48789 10489 48823 10523
rect 53021 10489 53055 10523
rect 53389 10489 53423 10523
rect 56977 10489 57011 10523
rect 59829 10489 59863 10523
rect 83197 10489 83231 10523
rect 6653 10421 6687 10455
rect 15209 10421 15243 10455
rect 18245 10421 18279 10455
rect 23765 10421 23799 10455
rect 36645 10421 36679 10455
rect 49341 10421 49375 10455
rect 49801 10421 49835 10455
rect 52193 10421 52227 10455
rect 55321 10421 55355 10455
rect 63490 10421 63524 10455
rect 67741 10421 67775 10455
rect 70133 10421 70167 10455
rect 72893 10421 72927 10455
rect 73629 10421 73663 10455
rect 74181 10421 74215 10455
rect 76941 10421 76975 10455
rect 77677 10421 77711 10455
rect 84761 10421 84795 10455
rect 85313 10421 85347 10455
rect 1777 10217 1811 10251
rect 11805 10217 11839 10251
rect 18797 10217 18831 10251
rect 22569 10217 22603 10251
rect 32551 10217 32585 10251
rect 36553 10217 36587 10251
rect 41981 10217 42015 10251
rect 42809 10217 42843 10251
rect 44465 10217 44499 10251
rect 47041 10217 47075 10251
rect 48053 10217 48087 10251
rect 48605 10217 48639 10251
rect 49801 10217 49835 10251
rect 53481 10217 53515 10251
rect 53757 10217 53791 10251
rect 54401 10217 54435 10251
rect 59185 10217 59219 10251
rect 62681 10217 62715 10251
rect 63325 10217 63359 10251
rect 67465 10217 67499 10251
rect 68109 10217 68143 10251
rect 75469 10217 75503 10251
rect 81357 10217 81391 10251
rect 82001 10217 82035 10251
rect 88625 10217 88659 10251
rect 89913 10217 89947 10251
rect 3433 10149 3467 10183
rect 4077 10149 4111 10183
rect 19441 10149 19475 10183
rect 29101 10149 29135 10183
rect 38209 10149 38243 10183
rect 40141 10149 40175 10183
rect 90465 10149 90499 10183
rect 4905 10081 4939 10115
rect 10793 10081 10827 10115
rect 13553 10081 13587 10115
rect 15117 10081 15151 10115
rect 18245 10081 18279 10115
rect 19993 10081 20027 10115
rect 20269 10081 20303 10115
rect 22017 10081 22051 10115
rect 25421 10081 25455 10115
rect 30573 10081 30607 10115
rect 34345 10081 34379 10115
rect 36921 10081 36955 10115
rect 38485 10081 38519 10115
rect 40049 10051 40083 10085
rect 41245 10081 41279 10115
rect 42717 10081 42751 10115
rect 42901 10081 42935 10115
rect 45845 10081 45879 10115
rect 47225 10081 47259 10115
rect 48973 10081 49007 10115
rect 53573 10081 53607 10115
rect 55781 10081 55815 10115
rect 56977 10081 57011 10115
rect 59369 10081 59403 10115
rect 71237 10081 71271 10115
rect 72709 10081 72743 10115
rect 76389 10081 76423 10115
rect 79057 10081 79091 10115
rect 79793 10081 79827 10115
rect 82461 10081 82495 10115
rect 83933 10081 83967 10115
rect 89177 10081 89211 10115
rect 91569 10081 91603 10115
rect 93317 10081 93351 10115
rect 1593 10013 1627 10047
rect 2237 10013 2271 10047
rect 2513 10013 2547 10047
rect 3249 10013 3283 10047
rect 3985 10013 4019 10047
rect 4169 10013 4203 10047
rect 4629 10013 4663 10047
rect 7297 10013 7331 10047
rect 8033 10013 8067 10047
rect 8309 10013 8343 10047
rect 10885 10013 10919 10047
rect 15025 10013 15059 10047
rect 17417 10013 17451 10047
rect 27445 10013 27479 10047
rect 30205 10013 30239 10047
rect 31999 10013 32033 10047
rect 33977 10013 34011 10047
rect 36751 10013 36785 10047
rect 38577 10013 38611 10047
rect 40233 10013 40267 10047
rect 40325 10013 40359 10047
rect 41153 10013 41187 10047
rect 41331 10013 41365 10047
rect 42625 10013 42659 10047
rect 43545 10013 43579 10047
rect 43821 10013 43855 10047
rect 44465 10013 44499 10047
rect 44649 10013 44683 10047
rect 45385 10013 45419 10047
rect 45661 10013 45695 10047
rect 46305 10013 46339 10047
rect 46489 10013 46523 10047
rect 47317 10013 47351 10047
rect 48789 10013 48823 10047
rect 49065 10013 49099 10047
rect 49801 10013 49835 10047
rect 50353 10013 50387 10047
rect 52745 10013 52779 10047
rect 53481 10013 53515 10047
rect 53849 10013 53883 10047
rect 54493 10013 54527 10047
rect 55873 10013 55907 10047
rect 56793 10013 56827 10047
rect 59461 10013 59495 10047
rect 60749 10013 60783 10047
rect 61117 10013 61151 10047
rect 62589 10013 62623 10047
rect 63509 10013 63543 10047
rect 64429 10013 64463 10047
rect 66177 10013 66211 10047
rect 66545 10013 66579 10047
rect 67925 10013 67959 10047
rect 70409 10013 70443 10047
rect 70961 10013 70995 10047
rect 73169 10013 73203 10047
rect 75377 10013 75411 10047
rect 76113 10013 76147 10047
rect 78321 10013 78355 10047
rect 79149 10013 79183 10047
rect 79963 10013 79997 10047
rect 81449 10013 81483 10047
rect 84209 10013 84243 10047
rect 84853 10013 84887 10047
rect 85773 10013 85807 10047
rect 86417 10013 86451 10047
rect 89821 10013 89855 10047
rect 93961 10013 93995 10047
rect 6653 9945 6687 9979
rect 13277 9945 13311 9979
rect 15669 9945 15703 9979
rect 18429 9945 18463 9979
rect 23949 9945 23983 9979
rect 24685 9945 24719 9979
rect 24869 9945 24903 9979
rect 25697 9945 25731 9979
rect 27997 9945 28031 9979
rect 35265 9945 35299 9979
rect 41797 9945 41831 9979
rect 45477 9945 45511 9979
rect 46397 9945 46431 9979
rect 50905 9945 50939 9979
rect 52561 9945 52595 9979
rect 58633 9945 58667 9979
rect 61761 9945 61795 9979
rect 64705 9945 64739 9979
rect 66913 9945 66947 9979
rect 70133 9945 70167 9979
rect 73445 9945 73479 9979
rect 85865 9945 85899 9979
rect 86693 9945 86727 9979
rect 90649 9945 90683 9979
rect 91845 9945 91879 9979
rect 7113 9877 7147 9911
rect 9229 9877 9263 9911
rect 9781 9877 9815 9911
rect 10517 9877 10551 9911
rect 14657 9877 14691 9911
rect 18521 9877 18555 9911
rect 18613 9877 18647 9911
rect 23121 9877 23155 9911
rect 23857 9877 23891 9911
rect 28089 9877 28123 9911
rect 34989 9877 35023 9911
rect 36001 9877 36035 9911
rect 37657 9877 37691 9911
rect 39497 9877 39531 9911
rect 41997 9877 42031 9911
rect 42165 9877 42199 9911
rect 43361 9877 43395 9911
rect 43729 9877 43763 9911
rect 44281 9877 44315 9911
rect 55505 9877 55539 9911
rect 65257 9877 65291 9911
rect 68661 9877 68695 9911
rect 74917 9877 74951 9911
rect 77861 9877 77895 9911
rect 78413 9877 78447 9911
rect 80253 9877 80287 9911
rect 84761 9877 84795 9911
rect 88165 9877 88199 9911
rect 93869 9877 93903 9911
rect 17877 9673 17911 9707
rect 21097 9673 21131 9707
rect 39313 9673 39347 9707
rect 40325 9673 40359 9707
rect 49157 9673 49191 9707
rect 9505 9605 9539 9639
rect 11161 9605 11195 9639
rect 12633 9605 12667 9639
rect 13553 9605 13587 9639
rect 15853 9605 15887 9639
rect 19809 9605 19843 9639
rect 23213 9605 23247 9639
rect 30205 9605 30239 9639
rect 33248 9605 33282 9639
rect 35357 9605 35391 9639
rect 35541 9605 35575 9639
rect 39865 9605 39899 9639
rect 43637 9605 43671 9639
rect 47133 9605 47167 9639
rect 48329 9605 48363 9639
rect 48513 9605 48547 9639
rect 49985 9605 50019 9639
rect 52929 9605 52963 9639
rect 53113 9605 53147 9639
rect 53849 9605 53883 9639
rect 63325 9605 63359 9639
rect 64797 9605 64831 9639
rect 67741 9605 67775 9639
rect 72985 9605 73019 9639
rect 75377 9605 75411 9639
rect 76021 9605 76055 9639
rect 82461 9605 82495 9639
rect 87797 9605 87831 9639
rect 94237 9605 94271 9639
rect 2145 9537 2179 9571
rect 2605 9537 2639 9571
rect 2881 9537 2915 9571
rect 3617 9537 3651 9571
rect 4353 9537 4387 9571
rect 5089 9537 5123 9571
rect 5825 9537 5859 9571
rect 6653 9537 6687 9571
rect 6929 9537 6963 9571
rect 7665 9537 7699 9571
rect 8585 9537 8619 9571
rect 9321 9537 9355 9571
rect 11713 9537 11747 9571
rect 12909 9537 12943 9571
rect 14197 9537 14231 9571
rect 16037 9537 16071 9571
rect 16221 9537 16255 9571
rect 16313 9537 16347 9571
rect 17509 9537 17543 9571
rect 18889 9537 18923 9571
rect 19165 9537 19199 9571
rect 19993 9537 20027 9571
rect 20085 9537 20119 9571
rect 20729 9537 20763 9571
rect 24593 9537 24627 9571
rect 26617 9537 26651 9571
rect 27169 9537 27203 9571
rect 32965 9537 32999 9571
rect 36185 9537 36219 9571
rect 36377 9537 36411 9571
rect 36829 9537 36863 9571
rect 37749 9537 37783 9571
rect 38853 9537 38887 9571
rect 39129 9537 39163 9571
rect 41153 9537 41187 9571
rect 41981 9537 42015 9571
rect 43177 9537 43211 9571
rect 43821 9537 43855 9571
rect 43913 9537 43947 9571
rect 44097 9537 44131 9571
rect 44189 9537 44223 9571
rect 45385 9537 45419 9571
rect 49249 9537 49283 9571
rect 49341 9537 49375 9571
rect 52193 9537 52227 9571
rect 52377 9537 52411 9571
rect 53297 9537 53331 9571
rect 57345 9537 57379 9571
rect 58081 9537 58115 9571
rect 58173 9537 58207 9571
rect 58909 9537 58943 9571
rect 61945 9537 61979 9571
rect 62405 9537 62439 9571
rect 62589 9537 62623 9571
rect 63233 9537 63267 9571
rect 63447 9537 63481 9571
rect 67557 9537 67591 9571
rect 67833 9537 67867 9571
rect 71593 9543 71627 9577
rect 71697 9537 71731 9571
rect 72709 9537 72743 9571
rect 73905 9537 73939 9571
rect 74825 9537 74859 9571
rect 75469 9537 75503 9571
rect 75929 9537 75963 9571
rect 76665 9537 76699 9571
rect 78137 9537 78171 9571
rect 79517 9537 79551 9571
rect 83105 9537 83139 9571
rect 84209 9537 84243 9571
rect 84485 9537 84519 9571
rect 87889 9537 87923 9571
rect 88993 9537 89027 9571
rect 90189 9537 90223 9571
rect 93225 9537 93259 9571
rect 94145 9537 94179 9571
rect 4813 9469 4847 9503
rect 8309 9469 8343 9503
rect 9965 9469 9999 9503
rect 12633 9469 12667 9503
rect 14289 9469 14323 9503
rect 17417 9469 17451 9503
rect 18981 9469 19015 9503
rect 19073 9469 19107 9503
rect 19349 9469 19383 9503
rect 20821 9469 20855 9503
rect 22109 9469 22143 9503
rect 24869 9469 24903 9503
rect 27445 9469 27479 9503
rect 29929 9469 29963 9503
rect 32413 9469 32447 9503
rect 38945 9469 38979 9503
rect 41245 9469 41279 9503
rect 45477 9469 45511 9503
rect 46581 9469 46615 9503
rect 48973 9469 49007 9503
rect 49801 9469 49835 9503
rect 51641 9469 51675 9503
rect 55781 9469 55815 9503
rect 56057 9469 56091 9503
rect 56241 9469 56275 9503
rect 60657 9469 60691 9503
rect 61117 9469 61151 9503
rect 61301 9469 61335 9503
rect 63601 9469 63635 9503
rect 64521 9469 64555 9503
rect 68845 9469 68879 9503
rect 69121 9469 69155 9503
rect 70593 9469 70627 9503
rect 74733 9469 74767 9503
rect 76941 9469 76975 9503
rect 77861 9469 77895 9503
rect 79425 9469 79459 9503
rect 80345 9469 80379 9503
rect 80805 9469 80839 9503
rect 82645 9469 82679 9503
rect 83841 9469 83875 9503
rect 86969 9469 87003 9503
rect 87245 9469 87279 9503
rect 90649 9469 90683 9503
rect 90925 9469 90959 9503
rect 3801 9401 3835 9435
rect 7849 9401 7883 9435
rect 10609 9401 10643 9435
rect 12817 9401 12851 9435
rect 14565 9401 14599 9435
rect 15393 9401 15427 9435
rect 20085 9401 20119 9435
rect 34713 9401 34747 9435
rect 40141 9401 40175 9435
rect 40785 9401 40819 9435
rect 45017 9401 45051 9435
rect 48145 9401 48179 9435
rect 63509 9401 63543 9435
rect 83197 9401 83231 9435
rect 89085 9401 89119 9435
rect 1961 9333 1995 9367
rect 6009 9333 6043 9367
rect 11897 9333 11931 9367
rect 22661 9333 22695 9367
rect 28917 9333 28951 9367
rect 31677 9333 31711 9367
rect 35725 9333 35759 9367
rect 36277 9333 36311 9367
rect 38301 9333 38335 9367
rect 38853 9333 38887 9367
rect 46029 9333 46063 9367
rect 49065 9333 49099 9367
rect 57161 9333 57195 9367
rect 58817 9333 58851 9367
rect 61853 9333 61887 9367
rect 62589 9333 62623 9367
rect 66269 9333 66303 9367
rect 66729 9333 66763 9367
rect 67373 9333 67407 9367
rect 71053 9333 71087 9367
rect 71789 9333 71823 9367
rect 71973 9333 72007 9367
rect 74089 9333 74123 9367
rect 78781 9333 78815 9367
rect 85497 9333 85531 9367
rect 88349 9333 88383 9367
rect 90189 9333 90223 9367
rect 92397 9333 92431 9367
rect 92949 9333 92983 9367
rect 1777 9129 1811 9163
rect 3433 9129 3467 9163
rect 14657 9129 14691 9163
rect 15669 9129 15703 9163
rect 16221 9129 16255 9163
rect 16957 9129 16991 9163
rect 17693 9129 17727 9163
rect 18153 9129 18187 9163
rect 19717 9129 19751 9163
rect 19901 9129 19935 9163
rect 20913 9129 20947 9163
rect 21833 9129 21867 9163
rect 29837 9129 29871 9163
rect 44373 9129 44407 9163
rect 45201 9129 45235 9163
rect 46213 9129 46247 9163
rect 49801 9129 49835 9163
rect 59921 9129 59955 9163
rect 71697 9129 71731 9163
rect 77033 9129 77067 9163
rect 79333 9129 79367 9163
rect 93961 9129 93995 9163
rect 8401 9061 8435 9095
rect 21465 9061 21499 9095
rect 24777 9061 24811 9095
rect 25329 9061 25363 9095
rect 31033 9061 31067 9095
rect 36645 9061 36679 9095
rect 64705 9061 64739 9095
rect 2237 8993 2271 9027
rect 4261 8993 4295 9027
rect 5089 8993 5123 9027
rect 7757 8993 7791 9027
rect 9413 8993 9447 9027
rect 12265 8993 12299 9027
rect 13737 8993 13771 9027
rect 17049 8993 17083 9027
rect 19533 8993 19567 9027
rect 20545 8993 20579 9027
rect 25789 8993 25823 9027
rect 26065 8993 26099 9027
rect 28549 8993 28583 9027
rect 31585 8993 31619 9027
rect 34897 8993 34931 9027
rect 37657 8993 37691 9027
rect 38301 8993 38335 9027
rect 39313 8993 39347 9027
rect 43361 8993 43395 9027
rect 43637 8993 43671 9027
rect 44281 8993 44315 9027
rect 51641 8993 51675 9027
rect 53757 8993 53791 9027
rect 53941 8993 53975 9027
rect 57345 8993 57379 9027
rect 60657 8993 60691 9027
rect 62313 8993 62347 9027
rect 63509 8993 63543 9027
rect 66177 8993 66211 9027
rect 66453 8993 66487 9027
rect 68477 8993 68511 9027
rect 71053 8993 71087 9027
rect 73169 8993 73203 9027
rect 74089 8993 74123 9027
rect 77861 8993 77895 9027
rect 84025 8993 84059 9027
rect 88165 8993 88199 9027
rect 88441 8993 88475 9027
rect 90833 8993 90867 9027
rect 93225 8993 93259 9027
rect 2513 8925 2547 8959
rect 3249 8925 3283 8959
rect 4445 8925 4479 8959
rect 6009 8925 6043 8959
rect 9505 8925 9539 8959
rect 12725 8925 12759 8959
rect 13001 8925 13035 8959
rect 14565 8925 14599 8959
rect 14749 8925 14783 8959
rect 16129 8925 16163 8959
rect 16313 8925 16347 8959
rect 16773 8925 16807 8959
rect 16865 8925 16899 8959
rect 17509 8925 17543 8959
rect 17693 8925 17727 8959
rect 19441 8925 19475 8959
rect 19717 8925 19751 8959
rect 20637 8925 20671 8959
rect 21649 8925 21683 8959
rect 21741 8925 21775 8959
rect 22385 8925 22419 8959
rect 22569 8925 22603 8959
rect 28457 8925 28491 8959
rect 34069 8925 34103 8959
rect 34345 8925 34379 8959
rect 37565 8925 37599 8959
rect 38209 8925 38243 8959
rect 38393 8925 38427 8959
rect 39221 8925 39255 8959
rect 40509 8925 40543 8959
rect 40693 8925 40727 8959
rect 43821 8925 43855 8959
rect 44557 8925 44591 8959
rect 44649 8925 44683 8959
rect 45385 8925 45419 8959
rect 45477 8925 45511 8959
rect 45661 8925 45695 8959
rect 45753 8925 45787 8959
rect 46397 8925 46431 8959
rect 46673 8925 46707 8959
rect 47409 8925 47443 8959
rect 50813 8925 50847 8959
rect 51273 8925 51307 8959
rect 52101 8925 52135 8959
rect 54585 8925 54619 8959
rect 57805 8925 57839 8959
rect 58357 8925 58391 8959
rect 58909 8925 58943 8959
rect 59001 8925 59035 8959
rect 62497 8925 62531 8959
rect 63601 8925 63635 8959
rect 64245 8925 64279 8959
rect 65993 8925 66027 8959
rect 68293 8925 68327 8959
rect 71145 8925 71179 8959
rect 71789 8925 71823 8959
rect 72893 8925 72927 8959
rect 73813 8925 73847 8959
rect 76389 8925 76423 8959
rect 76941 8925 76975 8959
rect 77585 8925 77619 8959
rect 79977 8925 80011 8959
rect 80529 8927 80563 8961
rect 81265 8925 81299 8959
rect 86509 8925 86543 8959
rect 86877 8925 86911 8959
rect 87981 8925 88015 8959
rect 91017 8925 91051 8959
rect 93409 8925 93443 8959
rect 93869 8925 93903 8959
rect 6285 8857 6319 8891
rect 11989 8857 12023 8891
rect 18337 8857 18371 8891
rect 18705 8857 18739 8891
rect 21925 8857 21959 8891
rect 27813 8857 27847 8891
rect 31861 8857 31895 8891
rect 35173 8857 35207 8891
rect 47593 8857 47627 8891
rect 49249 8857 49283 8891
rect 57621 8857 57655 8891
rect 60105 8857 60139 8891
rect 70133 8857 70167 8891
rect 72249 8857 72283 8891
rect 79885 8857 79919 8891
rect 81541 8857 81575 8891
rect 84209 8857 84243 8891
rect 85865 8857 85899 8891
rect 91569 8857 91603 8891
rect 9137 8789 9171 8823
rect 10517 8789 10551 8823
rect 18429 8789 18463 8823
rect 18521 8789 18555 8823
rect 22385 8789 22419 8823
rect 23121 8789 23155 8823
rect 28825 8789 28859 8823
rect 30481 8789 30515 8823
rect 33333 8789 33367 8823
rect 33885 8789 33919 8823
rect 34253 8789 34287 8823
rect 37197 8789 37231 8823
rect 38853 8789 38887 8823
rect 40693 8789 40727 8823
rect 41429 8789 41463 8823
rect 44465 8789 44499 8823
rect 46581 8789 46615 8823
rect 54493 8789 54527 8823
rect 59737 8789 59771 8823
rect 59905 8789 59939 8823
rect 75561 8789 75595 8823
rect 76205 8789 76239 8823
rect 80621 8789 80655 8823
rect 83013 8789 83047 8823
rect 87521 8789 87555 8823
rect 2145 8585 2179 8619
rect 4721 8585 4755 8619
rect 8493 8585 8527 8619
rect 16313 8585 16347 8619
rect 17049 8585 17083 8619
rect 20637 8585 20671 8619
rect 22569 8585 22603 8619
rect 27629 8585 27663 8619
rect 36461 8585 36495 8619
rect 37841 8585 37875 8619
rect 40325 8585 40359 8619
rect 42993 8585 43027 8619
rect 45201 8585 45235 8619
rect 47869 8585 47903 8619
rect 49525 8585 49559 8619
rect 50629 8585 50663 8619
rect 53481 8585 53515 8619
rect 54585 8585 54619 8619
rect 57437 8585 57471 8619
rect 64061 8585 64095 8619
rect 75193 8585 75227 8619
rect 78137 8585 78171 8619
rect 82185 8585 82219 8619
rect 86877 8585 86911 8619
rect 13461 8517 13495 8551
rect 15853 8517 15887 8551
rect 20269 8517 20303 8551
rect 21465 8517 21499 8551
rect 26249 8517 26283 8551
rect 28917 8517 28951 8551
rect 48513 8517 48547 8551
rect 52101 8517 52135 8551
rect 69029 8517 69063 8551
rect 77539 8517 77573 8551
rect 78873 8517 78907 8551
rect 87889 8517 87923 8551
rect 93409 8517 93443 8551
rect 2973 8449 3007 8483
rect 4353 8449 4387 8483
rect 5365 8449 5399 8483
rect 6653 8449 6687 8483
rect 6929 8449 6963 8483
rect 7573 8449 7607 8483
rect 8585 8449 8619 8483
rect 9137 8449 9171 8483
rect 9505 8449 9539 8483
rect 13737 8449 13771 8483
rect 14749 8449 14783 8483
rect 17694 8449 17728 8483
rect 17877 8449 17911 8483
rect 19165 8449 19199 8483
rect 20177 8449 20211 8483
rect 20453 8449 20487 8483
rect 21373 8449 21407 8483
rect 22201 8449 22235 8483
rect 23029 8449 23063 8483
rect 23765 8449 23799 8483
rect 26525 8449 26559 8483
rect 29929 8449 29963 8483
rect 33609 8449 33643 8483
rect 36277 8449 36311 8483
rect 36553 8449 36587 8483
rect 37473 8449 37507 8483
rect 37657 8449 37691 8483
rect 39313 8449 39347 8483
rect 40509 8449 40543 8483
rect 40785 8449 40819 8483
rect 41705 8449 41739 8483
rect 42809 8449 42843 8483
rect 42901 8449 42935 8483
rect 43913 8449 43947 8483
rect 46213 8449 46247 8483
rect 47777 8449 47811 8483
rect 47961 8449 47995 8483
rect 48789 8449 48823 8483
rect 49893 8449 49927 8483
rect 53205 8449 53239 8483
rect 53941 8449 53975 8483
rect 54125 8449 54159 8483
rect 58081 8449 58115 8483
rect 59369 8449 59403 8483
rect 62221 8449 62255 8483
rect 63693 8449 63727 8483
rect 64521 8449 64555 8483
rect 73629 8449 73663 8483
rect 73813 8449 73847 8483
rect 75285 8449 75319 8483
rect 75745 8449 75779 8483
rect 81265 8449 81299 8483
rect 82277 8449 82311 8483
rect 82921 8449 82955 8483
rect 84117 8449 84151 8483
rect 87521 8449 87555 8483
rect 89269 8449 89303 8483
rect 89913 8449 89947 8483
rect 90833 8449 90867 8483
rect 3065 8381 3099 8415
rect 3709 8381 3743 8415
rect 4261 8381 4295 8415
rect 5917 8381 5951 8415
rect 7849 8381 7883 8415
rect 10885 8381 10919 8415
rect 11713 8381 11747 8415
rect 14841 8381 14875 8415
rect 17785 8381 17819 8415
rect 17969 8381 18003 8415
rect 19073 8381 19107 8415
rect 22293 8381 22327 8415
rect 23121 8381 23155 8415
rect 23305 8381 23339 8415
rect 24777 8381 24811 8415
rect 30205 8381 30239 8415
rect 33885 8381 33919 8415
rect 35633 8381 35667 8415
rect 40601 8381 40635 8415
rect 40693 8381 40727 8415
rect 41613 8381 41647 8415
rect 42073 8381 42107 8415
rect 42625 8381 42659 8415
rect 44005 8381 44039 8415
rect 44281 8381 44315 8415
rect 46765 8381 46799 8415
rect 47225 8381 47259 8415
rect 48697 8381 48731 8415
rect 49985 8381 50019 8415
rect 52377 8381 52411 8415
rect 53481 8381 53515 8415
rect 55229 8381 55263 8415
rect 55505 8381 55539 8415
rect 59093 8381 59127 8415
rect 59277 8381 59311 8415
rect 59829 8381 59863 8415
rect 60105 8381 60139 8415
rect 63785 8381 63819 8415
rect 64797 8381 64831 8415
rect 67557 8381 67591 8415
rect 67833 8381 67867 8415
rect 68845 8381 68879 8415
rect 70685 8381 70719 8415
rect 72525 8381 72559 8415
rect 72801 8381 72835 8415
rect 72985 8381 73019 8415
rect 74641 8381 74675 8415
rect 76113 8381 76147 8415
rect 78689 8381 78723 8415
rect 79149 8381 79183 8415
rect 83013 8381 83047 8415
rect 85129 8381 85163 8415
rect 85405 8381 85439 8415
rect 90189 8381 90223 8415
rect 90741 8381 90775 8415
rect 91753 8381 91787 8415
rect 93593 8381 93627 8415
rect 2605 8313 2639 8347
rect 15117 8313 15151 8347
rect 16221 8313 16255 8347
rect 17509 8313 17543 8347
rect 19533 8313 19567 8347
rect 23213 8313 23247 8347
rect 29469 8313 29503 8347
rect 32597 8313 32631 8347
rect 39773 8313 39807 8347
rect 43177 8313 43211 8347
rect 46949 8313 46983 8347
rect 53297 8313 53331 8347
rect 58173 8313 58207 8347
rect 62497 8313 62531 8347
rect 81265 8313 81299 8347
rect 83289 8313 83323 8347
rect 91201 8313 91235 8347
rect 94145 8313 94179 8347
rect 5273 8245 5307 8279
rect 31677 8245 31711 8279
rect 33057 8245 33091 8279
rect 36093 8245 36127 8279
rect 38761 8245 38795 8279
rect 45753 8245 45787 8279
rect 48789 8245 48823 8279
rect 48973 8245 49007 8279
rect 53941 8245 53975 8279
rect 56977 8245 57011 8279
rect 59185 8245 59219 8279
rect 61577 8245 61611 8279
rect 65441 8245 65475 8279
rect 66085 8245 66119 8279
rect 84209 8245 84243 8279
rect 88993 8245 89027 8279
rect 2881 8041 2915 8075
rect 3433 8041 3467 8075
rect 15577 8041 15611 8075
rect 17417 8041 17451 8075
rect 18613 8041 18647 8075
rect 20637 8041 20671 8075
rect 21649 8041 21683 8075
rect 21833 8041 21867 8075
rect 28549 8041 28583 8075
rect 33333 8041 33367 8075
rect 40417 8041 40451 8075
rect 42993 8041 43027 8075
rect 47961 8041 47995 8075
rect 48237 8041 48271 8075
rect 49249 8041 49283 8075
rect 49709 8041 49743 8075
rect 50997 8041 51031 8075
rect 52193 8041 52227 8075
rect 52377 8041 52411 8075
rect 54861 8041 54895 8075
rect 58081 8041 58115 8075
rect 62405 8041 62439 8075
rect 66361 8041 66395 8075
rect 79149 8041 79183 8075
rect 93547 8041 93581 8075
rect 7665 7973 7699 8007
rect 13645 7973 13679 8007
rect 27813 7973 27847 8007
rect 34253 7973 34287 8007
rect 37289 7973 37323 8007
rect 45293 7973 45327 8007
rect 46949 7973 46983 8007
rect 47041 7973 47075 8007
rect 54033 7973 54067 8007
rect 59921 7973 59955 8007
rect 69121 7973 69155 8007
rect 71329 7973 71363 8007
rect 75377 7973 75411 8007
rect 79977 7973 80011 8007
rect 80529 7973 80563 8007
rect 86693 7973 86727 8007
rect 4997 7905 5031 7939
rect 5273 7905 5307 7939
rect 7021 7905 7055 7939
rect 18521 7905 18555 7939
rect 20085 7905 20119 7939
rect 20913 7905 20947 7939
rect 27169 7905 27203 7939
rect 36645 7905 36679 7939
rect 40785 7905 40819 7939
rect 42901 7905 42935 7939
rect 45753 7905 45787 7939
rect 46857 7905 46891 7939
rect 53481 7905 53515 7939
rect 56333 7905 56367 7939
rect 56609 7905 56643 7939
rect 59461 7905 59495 7939
rect 60933 7905 60967 7939
rect 63325 7905 63359 7939
rect 66085 7905 66119 7939
rect 67373 7905 67407 7939
rect 67649 7905 67683 7939
rect 69673 7905 69707 7939
rect 74733 7905 74767 7939
rect 76205 7905 76239 7939
rect 78045 7905 78079 7939
rect 78781 7905 78815 7939
rect 80713 7905 80747 7939
rect 81449 7905 81483 7939
rect 83841 7905 83875 7939
rect 84117 7905 84151 7939
rect 88717 7905 88751 7939
rect 88993 7905 89027 7939
rect 89453 7905 89487 7939
rect 92121 7905 92155 7939
rect 3985 7837 4019 7871
rect 8401 7837 8435 7871
rect 9413 7837 9447 7871
rect 10057 7837 10091 7871
rect 10333 7837 10367 7871
rect 11345 7837 11379 7871
rect 11713 7837 11747 7871
rect 18061 7837 18095 7871
rect 18705 7837 18739 7871
rect 18797 7837 18831 7871
rect 21005 7837 21039 7871
rect 28733 7837 28767 7871
rect 29101 7837 29135 7871
rect 31585 7837 31619 7871
rect 34897 7837 34931 7871
rect 39405 7837 39439 7871
rect 40693 7837 40727 7871
rect 41337 7837 41371 7871
rect 41613 7837 41647 7871
rect 42993 7837 43027 7871
rect 45661 7837 45695 7871
rect 47133 7837 47167 7871
rect 48237 7837 48271 7871
rect 48329 7837 48363 7871
rect 51200 7837 51234 7871
rect 51457 7837 51491 7871
rect 53021 7837 53055 7871
rect 54953 7837 54987 7871
rect 55873 7837 55907 7871
rect 59553 7837 59587 7871
rect 60657 7837 60691 7871
rect 65165 7837 65199 7871
rect 65993 7837 66027 7871
rect 69765 7837 69799 7871
rect 70409 7837 70443 7871
rect 71513 7837 71547 7871
rect 72065 7837 72099 7871
rect 72171 7837 72205 7871
rect 72341 7837 72375 7871
rect 72433 7837 72467 7871
rect 73077 7837 73111 7871
rect 74917 7837 74951 7871
rect 78873 7837 78907 7871
rect 79793 7837 79827 7871
rect 79977 7837 80011 7871
rect 80437 7837 80471 7871
rect 82645 7837 82679 7871
rect 82921 7837 82955 7871
rect 83657 7837 83691 7871
rect 86509 7837 86543 7871
rect 89729 7837 89763 7871
rect 90465 7837 90499 7871
rect 91753 7837 91787 7871
rect 94053 7837 94087 7871
rect 8309 7769 8343 7803
rect 13185 7769 13219 7803
rect 14289 7769 14323 7803
rect 19809 7769 19843 7803
rect 19901 7769 19935 7803
rect 21812 7769 21846 7803
rect 22017 7769 22051 7803
rect 26893 7769 26927 7803
rect 29837 7769 29871 7803
rect 32045 7769 32079 7803
rect 35173 7769 35207 7803
rect 38301 7769 38335 7803
rect 41429 7769 41463 7803
rect 42717 7769 42751 7803
rect 50445 7769 50479 7803
rect 51365 7769 51399 7803
rect 52009 7769 52043 7803
rect 64981 7769 65015 7803
rect 70317 7769 70351 7803
rect 77861 7769 77895 7803
rect 4169 7701 4203 7735
rect 9137 7701 9171 7735
rect 16957 7701 16991 7735
rect 19441 7701 19475 7735
rect 22937 7701 22971 7735
rect 25421 7701 25455 7735
rect 28825 7701 28859 7735
rect 28917 7701 28951 7735
rect 37749 7701 37783 7735
rect 38945 7701 38979 7735
rect 41797 7701 41831 7735
rect 43177 7701 43211 7735
rect 44097 7701 44131 7735
rect 44649 7701 44683 7735
rect 46397 7701 46431 7735
rect 52209 7701 52243 7735
rect 52929 7701 52963 7735
rect 55781 7701 55815 7735
rect 58541 7701 58575 7735
rect 66913 7701 66947 7735
rect 72617 7701 72651 7735
rect 80713 7701 80747 7735
rect 87245 7701 87279 7735
rect 90649 7701 90683 7735
rect 94237 7701 94271 7735
rect 5917 7497 5951 7531
rect 18337 7497 18371 7531
rect 18981 7497 19015 7531
rect 24685 7497 24719 7531
rect 27537 7497 27571 7531
rect 28457 7497 28491 7531
rect 35449 7497 35483 7531
rect 39773 7497 39807 7531
rect 42625 7497 42659 7531
rect 42993 7497 43027 7531
rect 44189 7497 44223 7531
rect 45477 7497 45511 7531
rect 46581 7497 46615 7531
rect 47225 7497 47259 7531
rect 49249 7497 49283 7531
rect 52193 7497 52227 7531
rect 60565 7497 60599 7531
rect 60841 7497 60875 7531
rect 64797 7497 64831 7531
rect 66821 7497 66855 7531
rect 67833 7497 67867 7531
rect 75101 7497 75135 7531
rect 76481 7497 76515 7531
rect 76941 7497 76975 7531
rect 78137 7497 78171 7531
rect 85313 7497 85347 7531
rect 86049 7497 86083 7531
rect 86601 7497 86635 7531
rect 93133 7497 93167 7531
rect 2237 7429 2271 7463
rect 4445 7429 4479 7463
rect 9597 7429 9631 7463
rect 13737 7429 13771 7463
rect 14473 7429 14507 7463
rect 16865 7429 16899 7463
rect 17693 7429 17727 7463
rect 26157 7429 26191 7463
rect 27997 7429 28031 7463
rect 29929 7429 29963 7463
rect 32413 7429 32447 7463
rect 33149 7429 33183 7463
rect 34897 7429 34931 7463
rect 49985 7429 50019 7463
rect 52929 7429 52963 7463
rect 57529 7429 57563 7463
rect 58357 7429 58391 7463
rect 62589 7429 62623 7463
rect 63509 7429 63543 7463
rect 70501 7429 70535 7463
rect 77769 7429 77803 7463
rect 78781 7429 78815 7463
rect 79701 7429 79735 7463
rect 80713 7429 80747 7463
rect 83197 7429 83231 7463
rect 84761 7429 84795 7463
rect 89177 7429 89211 7463
rect 79931 7395 79965 7429
rect 1961 7361 1995 7395
rect 6653 7361 6687 7395
rect 7205 7361 7239 7395
rect 10057 7361 10091 7395
rect 11989 7361 12023 7395
rect 18245 7361 18279 7395
rect 18429 7361 18463 7395
rect 19073 7361 19107 7395
rect 19625 7361 19659 7395
rect 20453 7361 20487 7395
rect 22109 7361 22143 7395
rect 27721 7361 27755 7395
rect 35817 7361 35851 7395
rect 36829 7361 36863 7395
rect 38209 7361 38243 7395
rect 39129 7361 39163 7395
rect 40141 7361 40175 7395
rect 41061 7361 41095 7395
rect 42073 7361 42107 7395
rect 42809 7361 42843 7395
rect 42901 7361 42935 7395
rect 49157 7361 49191 7395
rect 49801 7361 49835 7395
rect 52101 7361 52135 7395
rect 52285 7361 52319 7395
rect 53573 7361 53607 7395
rect 57253 7361 57287 7395
rect 58081 7361 58115 7395
rect 60749 7361 60783 7395
rect 60933 7361 60967 7395
rect 62681 7361 62715 7395
rect 63877 7361 63911 7395
rect 64337 7361 64371 7395
rect 64613 7361 64647 7395
rect 65533 7361 65567 7395
rect 65625 7361 65659 7395
rect 65809 7361 65843 7395
rect 66453 7361 66487 7395
rect 66637 7361 66671 7395
rect 67511 7361 67545 7395
rect 68753 7361 68787 7395
rect 69581 7361 69615 7395
rect 72985 7361 73019 7395
rect 74733 7361 74767 7395
rect 76021 7361 76055 7395
rect 76297 7361 76331 7395
rect 77677 7361 77711 7395
rect 77953 7361 77987 7395
rect 78689 7361 78723 7395
rect 78873 7361 78907 7395
rect 83013 7361 83047 7395
rect 83289 7361 83323 7395
rect 84209 7361 84243 7395
rect 84301 7361 84335 7395
rect 84485 7361 84519 7395
rect 84577 7361 84611 7395
rect 85957 7361 85991 7395
rect 87521 7361 87555 7395
rect 88257 7361 88291 7395
rect 91569 7361 91603 7395
rect 92305 7361 92339 7395
rect 92949 7361 92983 7395
rect 3709 7293 3743 7327
rect 4169 7293 4203 7327
rect 14197 7293 14231 7327
rect 16221 7293 16255 7327
rect 23121 7293 23155 7327
rect 26433 7293 26467 7327
rect 27905 7293 27939 7327
rect 30205 7293 30239 7327
rect 32873 7293 32907 7327
rect 35725 7293 35759 7327
rect 39037 7293 39071 7327
rect 40233 7293 40267 7327
rect 40877 7293 40911 7327
rect 40969 7293 41003 7327
rect 41153 7293 41187 7327
rect 41793 7293 41827 7327
rect 46121 7293 46155 7327
rect 51641 7293 51675 7327
rect 53757 7293 53791 7327
rect 54585 7293 54619 7327
rect 54861 7293 54895 7327
rect 61577 7293 61611 7327
rect 64429 7293 64463 7327
rect 67373 7293 67407 7327
rect 68661 7293 68695 7327
rect 69489 7293 69523 7327
rect 72709 7293 72743 7327
rect 73537 7293 73571 7327
rect 74641 7293 74675 7327
rect 76113 7293 76147 7327
rect 80529 7293 80563 7327
rect 81725 7293 81759 7327
rect 87245 7293 87279 7327
rect 88993 7293 89027 7327
rect 89453 7293 89487 7327
rect 91293 7293 91327 7327
rect 94145 7293 94179 7327
rect 38761 7225 38795 7259
rect 41889 7225 41923 7259
rect 43177 7225 43211 7259
rect 47869 7225 47903 7259
rect 48513 7225 48547 7259
rect 61117 7225 61151 7259
rect 61945 7225 61979 7259
rect 65993 7225 66027 7259
rect 69949 7225 69983 7259
rect 8309 7157 8343 7191
rect 10241 7157 10275 7191
rect 11069 7157 11103 7191
rect 23673 7157 23707 7191
rect 24225 7157 24259 7191
rect 27997 7157 28031 7191
rect 30665 7157 30699 7191
rect 37749 7157 37783 7191
rect 41337 7157 41371 7191
rect 41981 7157 42015 7191
rect 44925 7157 44959 7191
rect 56333 7157 56367 7191
rect 59829 7157 59863 7191
rect 62037 7157 62071 7191
rect 64613 7157 64647 7191
rect 66637 7157 66671 7191
rect 68477 7157 68511 7191
rect 71237 7157 71271 7191
rect 76297 7157 76331 7191
rect 79885 7157 79919 7191
rect 80069 7157 80103 7191
rect 82829 7157 82863 7191
rect 88441 7157 88475 7191
rect 92489 7157 92523 7191
rect 21465 6953 21499 6987
rect 22109 6953 22143 6987
rect 28089 6953 28123 6987
rect 28733 6953 28767 6987
rect 32247 6953 32281 6987
rect 35160 6953 35194 6987
rect 37841 6953 37875 6987
rect 38945 6953 38979 6987
rect 41061 6953 41095 6987
rect 49249 6953 49283 6987
rect 50616 6953 50650 6987
rect 52653 6953 52687 6987
rect 53757 6953 53791 6987
rect 54585 6953 54619 6987
rect 58541 6953 58575 6987
rect 65257 6953 65291 6987
rect 67943 6953 67977 6987
rect 81541 6953 81575 6987
rect 84393 6953 84427 6987
rect 84761 6953 84795 6987
rect 88165 6953 88199 6987
rect 93409 6953 93443 6987
rect 16681 6885 16715 6919
rect 22937 6885 22971 6919
rect 34161 6885 34195 6919
rect 40417 6885 40451 6919
rect 74181 6885 74215 6919
rect 80713 6885 80747 6919
rect 87061 6885 87095 6919
rect 89913 6885 89947 6919
rect 4261 6817 4295 6851
rect 10057 6817 10091 6851
rect 12906 6817 12940 6851
rect 13461 6817 13495 6851
rect 14565 6817 14599 6851
rect 20177 6817 20211 6851
rect 23581 6817 23615 6851
rect 24869 6817 24903 6851
rect 25329 6817 25363 6851
rect 29929 6817 29963 6851
rect 32505 6817 32539 6851
rect 32965 6817 32999 6851
rect 33425 6817 33459 6851
rect 34897 6817 34931 6851
rect 36645 6817 36679 6851
rect 37289 6817 37323 6851
rect 38485 6817 38519 6851
rect 40049 6817 40083 6851
rect 40509 6817 40543 6851
rect 42901 6817 42935 6851
rect 44649 6817 44683 6851
rect 45477 6817 45511 6851
rect 48789 6817 48823 6851
rect 49433 6817 49467 6851
rect 50353 6817 50387 6851
rect 53205 6817 53239 6851
rect 56425 6817 56459 6851
rect 57989 6817 58023 6851
rect 60749 6817 60783 6851
rect 61853 6817 61887 6851
rect 62037 6817 62071 6851
rect 62773 6817 62807 6851
rect 62957 6817 62991 6851
rect 69305 6817 69339 6851
rect 71605 6817 71639 6851
rect 74641 6817 74675 6851
rect 75285 6817 75319 6851
rect 80437 6817 80471 6851
rect 82461 6817 82495 6851
rect 84485 6817 84519 6851
rect 88717 6817 88751 6851
rect 90925 6817 90959 6851
rect 92397 6817 92431 6851
rect 3065 6749 3099 6783
rect 4169 6749 4203 6783
rect 7205 6749 7239 6783
rect 7481 6749 7515 6783
rect 8125 6749 8159 6783
rect 10333 6749 10367 6783
rect 10977 6749 11011 6783
rect 11897 6749 11931 6783
rect 12633 6749 12667 6783
rect 14657 6749 14691 6783
rect 15301 6749 15335 6783
rect 18797 6749 18831 6783
rect 19993 6749 20027 6783
rect 23029 6749 23063 6783
rect 23673 6749 23707 6783
rect 27353 6749 27387 6783
rect 33333 6749 33367 6783
rect 34343 6727 34377 6761
rect 39129 6749 39163 6783
rect 39405 6749 39439 6783
rect 40969 6749 41003 6783
rect 41153 6749 41187 6783
rect 42809 6749 42843 6783
rect 45201 6749 45235 6783
rect 45293 6749 45327 6783
rect 46029 6749 46063 6783
rect 47869 6749 47903 6783
rect 49525 6749 49559 6783
rect 52745 6749 52779 6783
rect 54401 6749 54435 6783
rect 56333 6749 56367 6783
rect 59553 6749 59587 6783
rect 59829 6749 59863 6783
rect 60841 6749 60875 6783
rect 61945 6749 61979 6783
rect 62129 6749 62163 6783
rect 62681 6749 62715 6783
rect 63509 6749 63543 6783
rect 68201 6749 68235 6783
rect 71329 6749 71363 6783
rect 74549 6749 74583 6783
rect 75469 6749 75503 6783
rect 75561 6749 75595 6783
rect 76205 6749 76239 6783
rect 76389 6749 76423 6783
rect 77309 6749 77343 6783
rect 78321 6749 78355 6783
rect 79425 6749 79459 6783
rect 80345 6749 80379 6783
rect 81265 6759 81299 6793
rect 81633 6749 81667 6783
rect 82185 6749 82219 6783
rect 84393 6749 84427 6783
rect 85221 6749 85255 6783
rect 86877 6749 86911 6783
rect 87981 6749 88015 6783
rect 88993 6749 89027 6783
rect 89637 6749 89671 6783
rect 90465 6749 90499 6783
rect 92673 6749 92707 6783
rect 8401 6681 8435 6715
rect 19441 6681 19475 6715
rect 21005 6681 21039 6715
rect 22753 6681 22787 6715
rect 25605 6681 25639 6715
rect 28549 6681 28583 6715
rect 30481 6681 30515 6715
rect 34069 6681 34103 6715
rect 34253 6681 34287 6715
rect 41981 6681 42015 6715
rect 43545 6681 43579 6715
rect 46213 6681 46247 6715
rect 49249 6681 49283 6715
rect 56977 6681 57011 6715
rect 63785 6681 63819 6715
rect 66177 6681 66211 6715
rect 69765 6681 69799 6715
rect 73629 6681 73663 6715
rect 75285 6681 75319 6715
rect 76757 6681 76791 6715
rect 78873 6681 78907 6715
rect 81357 6681 81391 6715
rect 91845 6681 91879 6715
rect 93961 6681 93995 6715
rect 3249 6613 3283 6647
rect 4537 6613 4571 6647
rect 5089 6613 5123 6647
rect 6653 6613 6687 6647
rect 9597 6613 9631 6647
rect 11253 6613 11287 6647
rect 11713 6613 11747 6647
rect 14289 6613 14323 6647
rect 18245 6613 18279 6647
rect 23029 6613 23063 6647
rect 24041 6613 24075 6647
rect 28749 6613 28783 6647
rect 28917 6613 28951 6647
rect 39313 6613 39347 6647
rect 42441 6613 42475 6647
rect 43637 6613 43671 6647
rect 45477 6613 45511 6647
rect 49709 6613 49743 6647
rect 52101 6613 52135 6647
rect 57437 6613 57471 6647
rect 59645 6613 59679 6647
rect 60013 6613 60047 6647
rect 61209 6613 61243 6647
rect 61669 6613 61703 6647
rect 62957 6613 62991 6647
rect 68753 6613 68787 6647
rect 70409 6613 70443 6647
rect 73077 6613 73111 6647
rect 76481 6613 76515 6647
rect 76573 6613 76607 6647
rect 77769 6613 77803 6647
rect 81449 6613 81483 6647
rect 83933 6613 83967 6647
rect 85865 6613 85899 6647
rect 4721 6409 4755 6443
rect 15025 6409 15059 6443
rect 17969 6409 18003 6443
rect 19441 6409 19475 6443
rect 20545 6409 20579 6443
rect 26617 6409 26651 6443
rect 32413 6409 32447 6443
rect 39313 6409 39347 6443
rect 40233 6409 40267 6443
rect 43729 6409 43763 6443
rect 45201 6409 45235 6443
rect 46949 6409 46983 6443
rect 49801 6409 49835 6443
rect 49985 6409 50019 6443
rect 52101 6409 52135 6443
rect 58173 6409 58207 6443
rect 59553 6409 59587 6443
rect 60657 6409 60691 6443
rect 64613 6409 64647 6443
rect 65349 6409 65383 6443
rect 67373 6409 67407 6443
rect 68569 6409 68603 6443
rect 71605 6409 71639 6443
rect 72157 6409 72191 6443
rect 74733 6409 74767 6443
rect 76297 6409 76331 6443
rect 83289 6409 83323 6443
rect 94145 6409 94179 6443
rect 6009 6341 6043 6375
rect 22937 6341 22971 6375
rect 33149 6341 33183 6375
rect 34897 6341 34931 6375
rect 49893 6341 49927 6375
rect 50629 6341 50663 6375
rect 53849 6341 53883 6375
rect 56517 6341 56551 6375
rect 58725 6341 58759 6375
rect 70041 6341 70075 6375
rect 78781 6341 78815 6375
rect 79241 6341 79275 6375
rect 90557 6341 90591 6375
rect 6837 6273 6871 6307
rect 7481 6273 7515 6307
rect 8217 6273 8251 6307
rect 8493 6273 8527 6307
rect 9229 6273 9263 6307
rect 9873 6273 9907 6307
rect 10149 6273 10183 6307
rect 10793 6273 10827 6307
rect 14289 6273 14323 6307
rect 18705 6273 18739 6307
rect 19533 6273 19567 6307
rect 20361 6273 20395 6307
rect 20545 6273 20579 6307
rect 21005 6273 21039 6307
rect 23489 6273 23523 6307
rect 23765 6273 23799 6307
rect 27537 6273 27571 6307
rect 30113 6273 30147 6307
rect 32873 6273 32907 6307
rect 36001 6273 36035 6307
rect 36277 6273 36311 6307
rect 38025 6273 38059 6307
rect 39129 6273 39163 6307
rect 39313 6273 39347 6307
rect 40141 6273 40175 6307
rect 40325 6273 40359 6307
rect 40969 6273 41003 6307
rect 42073 6273 42107 6307
rect 44557 6273 44591 6307
rect 45569 6273 45603 6307
rect 46213 6273 46247 6307
rect 46397 6273 46431 6307
rect 48145 6273 48179 6307
rect 48414 6273 48448 6307
rect 48973 6273 49007 6307
rect 49151 6273 49185 6307
rect 51733 6273 51767 6307
rect 54493 6273 54527 6307
rect 56977 6273 57011 6307
rect 57161 6273 57195 6307
rect 59369 6273 59403 6307
rect 59553 6273 59587 6307
rect 60565 6273 60599 6307
rect 60749 6273 60783 6307
rect 61853 6273 61887 6307
rect 63785 6273 63819 6307
rect 64521 6273 64555 6307
rect 64705 6273 64739 6307
rect 65165 6273 65199 6307
rect 65349 6273 65383 6307
rect 66729 6273 66763 6307
rect 70317 6273 70351 6307
rect 71421 6273 71455 6307
rect 71697 6273 71731 6307
rect 72525 6273 72559 6307
rect 73537 6273 73571 6307
rect 73721 6273 73755 6307
rect 74549 6273 74583 6307
rect 74825 6273 74859 6307
rect 75561 6273 75595 6307
rect 77217 6273 77251 6307
rect 77401 6273 77435 6307
rect 79977 6273 80011 6307
rect 82921 6273 82955 6307
rect 83933 6273 83967 6307
rect 84761 6273 84795 6307
rect 85037 6273 85071 6307
rect 85773 6273 85807 6307
rect 86680 6273 86714 6307
rect 87429 6273 87463 6307
rect 88349 6273 88383 6307
rect 90833 6273 90867 6307
rect 92121 6273 92155 6307
rect 92397 6273 92431 6307
rect 93041 6273 93075 6307
rect 6561 6205 6595 6239
rect 18429 6205 18463 6239
rect 18613 6205 18647 6239
rect 19349 6205 19383 6239
rect 23673 6205 23707 6239
rect 24869 6205 24903 6239
rect 25145 6205 25179 6239
rect 27445 6205 27479 6239
rect 29837 6205 29871 6239
rect 37933 6205 37967 6239
rect 40877 6205 40911 6239
rect 43177 6205 43211 6239
rect 44649 6205 44683 6239
rect 45477 6205 45511 6239
rect 47961 6205 47995 6239
rect 48237 6205 48271 6239
rect 48330 6205 48364 6239
rect 51641 6205 51675 6239
rect 53665 6205 53699 6239
rect 53941 6205 53975 6239
rect 54769 6205 54803 6239
rect 61761 6205 61795 6239
rect 66821 6205 66855 6239
rect 72617 6205 72651 6239
rect 73629 6205 73663 6239
rect 75285 6205 75319 6239
rect 75469 6205 75503 6239
rect 75644 6205 75678 6239
rect 75745 6205 75779 6239
rect 76757 6205 76791 6239
rect 80253 6205 80287 6239
rect 82001 6205 82035 6239
rect 82829 6205 82863 6239
rect 86417 6205 86451 6239
rect 89085 6205 89119 6239
rect 11713 6137 11747 6171
rect 14381 6137 14415 6171
rect 19901 6137 19935 6171
rect 27169 6137 27203 6171
rect 35357 6137 35391 6171
rect 41337 6137 41371 6171
rect 46305 6137 46339 6171
rect 49617 6137 49651 6171
rect 50905 6137 50939 6171
rect 60105 6137 60139 6171
rect 74365 6137 74399 6171
rect 76389 6137 76423 6171
rect 77217 6137 77251 6171
rect 7757 6069 7791 6103
rect 9413 6069 9447 6103
rect 11069 6069 11103 6103
rect 18521 6069 18555 6103
rect 22477 6069 22511 6103
rect 23765 6069 23799 6103
rect 23949 6069 23983 6103
rect 28365 6069 28399 6103
rect 37657 6069 37691 6103
rect 44281 6069 44315 6103
rect 49157 6069 49191 6103
rect 50169 6069 50203 6103
rect 51089 6069 51123 6103
rect 57069 6069 57103 6103
rect 62129 6069 62163 6103
rect 63325 6069 63359 6103
rect 63969 6069 64003 6103
rect 65901 6069 65935 6103
rect 66453 6069 66487 6103
rect 71237 6069 71271 6103
rect 77861 6069 77895 6103
rect 84025 6069 84059 6103
rect 85957 6069 85991 6103
rect 87613 6069 87647 6103
rect 88165 6069 88199 6103
rect 91385 6069 91419 6103
rect 93317 6069 93351 6103
rect 10333 5865 10367 5899
rect 19901 5865 19935 5899
rect 23121 5865 23155 5899
rect 25881 5865 25915 5899
rect 34253 5865 34287 5899
rect 40785 5865 40819 5899
rect 42993 5865 43027 5899
rect 47777 5865 47811 5899
rect 49801 5865 49835 5899
rect 50813 5865 50847 5899
rect 51457 5865 51491 5899
rect 52009 5865 52043 5899
rect 52837 5865 52871 5899
rect 53389 5865 53423 5899
rect 53941 5865 53975 5899
rect 54493 5865 54527 5899
rect 60105 5865 60139 5899
rect 62116 5865 62150 5899
rect 65073 5865 65107 5899
rect 68109 5865 68143 5899
rect 68661 5865 68695 5899
rect 69213 5865 69247 5899
rect 70409 5865 70443 5899
rect 70961 5865 70995 5899
rect 75285 5865 75319 5899
rect 79057 5865 79091 5899
rect 82921 5865 82955 5899
rect 83473 5865 83507 5899
rect 85865 5865 85899 5899
rect 88441 5865 88475 5899
rect 93409 5865 93443 5899
rect 93869 5865 93903 5899
rect 8585 5797 8619 5831
rect 22661 5797 22695 5831
rect 28457 5797 28491 5831
rect 36829 5797 36863 5831
rect 38117 5797 38151 5831
rect 38853 5797 38887 5831
rect 39405 5797 39439 5831
rect 44005 5797 44039 5831
rect 46581 5797 46615 5831
rect 51365 5797 51399 5831
rect 67557 5797 67591 5831
rect 75101 5797 75135 5831
rect 77401 5797 77435 5831
rect 81265 5797 81299 5831
rect 85129 5797 85163 5831
rect 92765 5797 92799 5831
rect 3985 5729 4019 5763
rect 6377 5729 6411 5763
rect 6837 5729 6871 5763
rect 7113 5729 7147 5763
rect 9229 5729 9263 5763
rect 16313 5729 16347 5763
rect 19533 5729 19567 5763
rect 20545 5729 20579 5763
rect 23029 5729 23063 5763
rect 26985 5729 27019 5763
rect 32045 5729 32079 5763
rect 32505 5729 32539 5763
rect 35449 5729 35483 5763
rect 36001 5729 36035 5763
rect 40141 5729 40175 5763
rect 41521 5729 41555 5763
rect 45201 5729 45235 5763
rect 48789 5729 48823 5763
rect 51549 5729 51583 5763
rect 55597 5729 55631 5763
rect 56609 5729 56643 5763
rect 60749 5729 60783 5763
rect 61853 5729 61887 5763
rect 63877 5729 63911 5763
rect 64613 5729 64647 5763
rect 66085 5729 66119 5763
rect 71973 5729 72007 5763
rect 73169 5729 73203 5763
rect 78781 5729 78815 5763
rect 80713 5729 80747 5763
rect 84025 5729 84059 5763
rect 87981 5729 88015 5763
rect 89637 5729 89671 5763
rect 91569 5729 91603 5763
rect 9321 5661 9355 5695
rect 14289 5661 14323 5695
rect 15301 5661 15335 5695
rect 15485 5661 15519 5695
rect 19625 5661 19659 5695
rect 20637 5661 20671 5695
rect 21833 5661 21867 5695
rect 22845 5661 22879 5695
rect 24041 5661 24075 5695
rect 24777 5661 24811 5695
rect 24961 5661 24995 5695
rect 25421 5661 25455 5695
rect 25697 5661 25731 5695
rect 26709 5661 26743 5695
rect 41245 5661 41279 5695
rect 44465 5661 44499 5695
rect 44649 5661 44683 5695
rect 48697 5661 48731 5695
rect 48881 5661 48915 5695
rect 49525 5661 49559 5695
rect 49617 5661 49651 5695
rect 50353 5661 50387 5695
rect 50445 5661 50479 5695
rect 50629 5661 50663 5695
rect 51273 5661 51307 5695
rect 55689 5661 55723 5695
rect 56793 5661 56827 5695
rect 56977 5661 57011 5695
rect 57069 5661 57103 5695
rect 57529 5661 57563 5695
rect 58909 5661 58943 5695
rect 60841 5661 60875 5695
rect 64705 5661 64739 5695
rect 65809 5661 65843 5695
rect 69857 5661 69891 5695
rect 71789 5661 71823 5695
rect 75285 5661 75319 5695
rect 75377 5661 75411 5695
rect 75561 5661 75595 5695
rect 76389 5661 76423 5695
rect 77125 5661 77159 5695
rect 78689 5661 78723 5695
rect 79701 5661 79735 5695
rect 80437 5661 80471 5695
rect 86969 5661 87003 5695
rect 87705 5661 87739 5695
rect 88625 5661 88659 5695
rect 89361 5661 89395 5695
rect 91845 5661 91879 5695
rect 92489 5661 92523 5695
rect 93225 5661 93259 5695
rect 4261 5593 4295 5627
rect 14565 5593 14599 5627
rect 21649 5593 21683 5627
rect 21925 5593 21959 5627
rect 22201 5593 22235 5627
rect 23121 5593 23155 5627
rect 25513 5593 25547 5627
rect 30297 5593 30331 5627
rect 32781 5593 32815 5627
rect 37565 5593 37599 5627
rect 46029 5593 46063 5627
rect 47317 5593 47351 5627
rect 49801 5593 49835 5627
rect 57713 5593 57747 5627
rect 57897 5593 57931 5627
rect 76113 5593 76147 5627
rect 81817 5593 81851 5627
rect 84577 5593 84611 5627
rect 5733 5525 5767 5559
rect 9873 5525 9907 5559
rect 11161 5525 11195 5559
rect 22017 5525 22051 5559
rect 24961 5525 24995 5559
rect 44465 5525 44499 5559
rect 49341 5525 49375 5559
rect 56057 5525 56091 5559
rect 58357 5525 58391 5559
rect 59461 5525 59495 5559
rect 61209 5525 61243 5559
rect 74089 5525 74123 5559
rect 76297 5525 76331 5559
rect 76481 5525 76515 5559
rect 76665 5525 76699 5559
rect 77585 5525 77619 5559
rect 79517 5525 79551 5559
rect 82461 5525 82495 5559
rect 86785 5525 86819 5559
rect 90189 5525 90223 5559
rect 90649 5525 90683 5559
rect 4261 5321 4295 5355
rect 8309 5321 8343 5355
rect 22109 5321 22143 5355
rect 22845 5321 22879 5355
rect 34437 5321 34471 5355
rect 37933 5321 37967 5355
rect 39681 5321 39715 5355
rect 40141 5321 40175 5355
rect 40877 5321 40911 5355
rect 90649 5321 90683 5355
rect 91293 5321 91327 5355
rect 94145 5321 94179 5355
rect 9597 5253 9631 5287
rect 13001 5253 13035 5287
rect 23305 5253 23339 5287
rect 26157 5253 26191 5287
rect 27353 5253 27387 5287
rect 28273 5253 28307 5287
rect 41521 5253 41555 5287
rect 44281 5253 44315 5287
rect 46305 5253 46339 5287
rect 48237 5253 48271 5287
rect 49417 5253 49451 5287
rect 49617 5253 49651 5287
rect 52193 5253 52227 5287
rect 53573 5253 53607 5287
rect 55873 5253 55907 5287
rect 58173 5253 58207 5287
rect 62405 5253 62439 5287
rect 63785 5253 63819 5287
rect 64889 5253 64923 5287
rect 66361 5253 66395 5287
rect 68385 5253 68419 5287
rect 73629 5253 73663 5287
rect 76757 5253 76791 5287
rect 84669 5253 84703 5287
rect 4353 5185 4387 5219
rect 6837 5185 6871 5219
rect 22569 5185 22603 5219
rect 22753 5185 22787 5219
rect 22845 5185 22879 5219
rect 23489 5185 23523 5219
rect 28733 5185 28767 5219
rect 31769 5185 31803 5219
rect 32689 5185 32723 5219
rect 36369 5185 36403 5219
rect 37657 5185 37691 5219
rect 42993 5185 43027 5219
rect 48145 5185 48179 5219
rect 50077 5185 50111 5219
rect 50905 5185 50939 5219
rect 53205 5185 53239 5219
rect 53389 5185 53423 5219
rect 53481 5185 53515 5219
rect 56793 5185 56827 5219
rect 56977 5185 57011 5219
rect 57069 5185 57103 5219
rect 58081 5185 58115 5219
rect 58357 5185 58391 5219
rect 62681 5185 62715 5219
rect 64429 5185 64463 5219
rect 69765 5185 69799 5219
rect 72433 5185 72467 5219
rect 73529 5175 73563 5209
rect 73721 5185 73755 5219
rect 74181 5185 74215 5219
rect 74365 5185 74399 5219
rect 75285 5185 75319 5219
rect 75469 5185 75503 5219
rect 76021 5185 76055 5219
rect 76205 5185 76239 5219
rect 76665 5185 76699 5219
rect 76849 5185 76883 5219
rect 77585 5185 77619 5219
rect 77677 5185 77711 5219
rect 79241 5185 79275 5219
rect 84393 5185 84427 5219
rect 85405 5185 85439 5219
rect 86049 5185 86083 5219
rect 87061 5185 87095 5219
rect 87705 5185 87739 5219
rect 90189 5185 90223 5219
rect 92397 5185 92431 5219
rect 93041 5185 93075 5219
rect 14749 5117 14783 5151
rect 26433 5117 26467 5151
rect 27261 5117 27295 5151
rect 31493 5117 31527 5151
rect 32597 5117 32631 5151
rect 36921 5117 36955 5151
rect 41981 5117 42015 5151
rect 43085 5117 43119 5151
rect 44005 5117 44039 5151
rect 48329 5117 48363 5151
rect 50353 5117 50387 5151
rect 51181 5117 51215 5151
rect 56149 5117 56183 5151
rect 66913 5117 66947 5151
rect 69213 5117 69247 5151
rect 70041 5117 70075 5151
rect 72341 5117 72375 5151
rect 75009 5117 75043 5151
rect 75193 5117 75227 5151
rect 75377 5117 75411 5151
rect 77861 5117 77895 5151
rect 79149 5117 79183 5151
rect 80713 5117 80747 5151
rect 80989 5117 81023 5151
rect 84577 5117 84611 5151
rect 86325 5117 86359 5151
rect 86785 5117 86819 5151
rect 92121 5117 92155 5151
rect 32321 5049 32355 5083
rect 33793 5049 33827 5083
rect 45753 5049 45787 5083
rect 47777 5049 47811 5083
rect 49249 5049 49283 5083
rect 50169 5049 50203 5083
rect 51089 5049 51123 5083
rect 53757 5049 53791 5083
rect 54401 5049 54435 5083
rect 58081 5049 58115 5083
rect 58817 5049 58851 5083
rect 59921 5049 59955 5083
rect 63233 5049 63267 5083
rect 65441 5049 65475 5083
rect 71513 5049 71547 5083
rect 72065 5049 72099 5083
rect 76113 5049 76147 5083
rect 77769 5049 77803 5083
rect 79609 5049 79643 5083
rect 82461 5049 82495 5083
rect 6929 4981 6963 5015
rect 23673 4981 23707 5015
rect 24225 4981 24259 5015
rect 24685 4981 24719 5015
rect 28917 4981 28951 5015
rect 30021 4981 30055 5015
rect 38485 4981 38519 5015
rect 39037 4981 39071 5015
rect 42717 4981 42751 5015
rect 46949 4981 46983 5015
rect 49433 4981 49467 5015
rect 50261 4981 50295 5015
rect 50997 4981 51031 5015
rect 51733 4981 51767 5015
rect 56609 4981 56643 5015
rect 59461 4981 59495 5015
rect 60933 4981 60967 5015
rect 74273 4981 74307 5015
rect 80161 4981 80195 5015
rect 83105 4981 83139 5015
rect 84209 4981 84243 5015
rect 84669 4981 84703 5015
rect 85129 4981 85163 5015
rect 87981 4981 88015 5015
rect 88993 4981 89027 5015
rect 89545 4981 89579 5015
rect 93317 4981 93351 5015
rect 8493 4777 8527 4811
rect 22845 4777 22879 4811
rect 26525 4777 26559 4811
rect 29745 4777 29779 4811
rect 38117 4777 38151 4811
rect 47685 4777 47719 4811
rect 49157 4777 49191 4811
rect 50905 4777 50939 4811
rect 52469 4777 52503 4811
rect 53757 4777 53791 4811
rect 54769 4777 54803 4811
rect 56885 4777 56919 4811
rect 59185 4777 59219 4811
rect 60749 4777 60783 4811
rect 62405 4777 62439 4811
rect 65901 4777 65935 4811
rect 73261 4777 73295 4811
rect 73629 4777 73663 4811
rect 74365 4777 74399 4811
rect 76205 4777 76239 4811
rect 77953 4777 77987 4811
rect 82461 4777 82495 4811
rect 85037 4777 85071 4811
rect 87981 4777 88015 4811
rect 22385 4709 22419 4743
rect 23489 4709 23523 4743
rect 25513 4709 25547 4743
rect 33701 4709 33735 4743
rect 34989 4709 35023 4743
rect 39037 4709 39071 4743
rect 43361 4709 43395 4743
rect 44373 4709 44407 4743
rect 45201 4709 45235 4743
rect 46949 4709 46983 4743
rect 53389 4709 53423 4743
rect 58081 4709 58115 4743
rect 61209 4709 61243 4743
rect 62957 4709 62991 4743
rect 65165 4709 65199 4743
rect 72249 4709 72283 4743
rect 74549 4709 74583 4743
rect 77861 4709 77895 4743
rect 93225 4709 93259 4743
rect 6745 4641 6779 4675
rect 7021 4641 7055 4675
rect 31309 4641 31343 4675
rect 33977 4641 34011 4675
rect 36645 4641 36679 4675
rect 45937 4641 45971 4675
rect 47501 4641 47535 4675
rect 50445 4641 50479 4675
rect 53665 4641 53699 4675
rect 56149 4641 56183 4675
rect 61761 4641 61795 4675
rect 63509 4641 63543 4675
rect 64061 4641 64095 4675
rect 64521 4641 64555 4675
rect 67373 4641 67407 4675
rect 67649 4641 67683 4675
rect 68109 4641 68143 4675
rect 68385 4641 68419 4675
rect 69857 4641 69891 4675
rect 71697 4641 71731 4675
rect 72709 4641 72743 4675
rect 75101 4641 75135 4675
rect 77033 4641 77067 4675
rect 77769 4641 77803 4675
rect 79793 4641 79827 4675
rect 86785 4641 86819 4675
rect 88533 4641 88567 4675
rect 91017 4641 91051 4675
rect 91937 4641 91971 4675
rect 9137 4573 9171 4607
rect 9413 4573 9447 4607
rect 10149 4573 10183 4607
rect 14381 4573 14415 4607
rect 14565 4573 14599 4607
rect 25053 4573 25087 4607
rect 25145 4573 25179 4607
rect 25329 4573 25363 4607
rect 27813 4573 27847 4607
rect 29929 4573 29963 4607
rect 36369 4573 36403 4607
rect 40417 4573 40451 4607
rect 46029 4573 46063 4607
rect 47777 4573 47811 4607
rect 49249 4573 49283 4607
rect 52009 4573 52043 4607
rect 53573 4573 53607 4607
rect 54953 4573 54987 4607
rect 56030 4573 56064 4607
rect 57253 4573 57287 4607
rect 58725 4573 58759 4607
rect 59737 4573 59771 4607
rect 71527 4573 71561 4607
rect 72617 4573 72651 4607
rect 73445 4573 73479 4607
rect 73537 4573 73571 4607
rect 76941 4573 76975 4607
rect 78045 4573 78079 4607
rect 78505 4573 78539 4607
rect 78689 4573 78723 4607
rect 79517 4573 79551 4607
rect 81265 4573 81299 4607
rect 81541 4573 81575 4607
rect 82277 4573 82311 4607
rect 83381 4573 83415 4607
rect 83657 4573 83691 4607
rect 84393 4573 84427 4607
rect 85681 4573 85715 4607
rect 85865 4573 85899 4607
rect 87061 4573 87095 4607
rect 87705 4573 87739 4607
rect 88625 4573 88659 4607
rect 90557 4573 90591 4607
rect 90833 4573 90867 4607
rect 92029 4573 92063 4607
rect 93041 4573 93075 4607
rect 31401 4505 31435 4539
rect 32321 4505 32355 4539
rect 35357 4505 35391 4539
rect 40693 4505 40727 4539
rect 42625 4505 42659 4539
rect 49801 4505 49835 4539
rect 53849 4505 53883 4539
rect 57069 4505 57103 4539
rect 57713 4505 57747 4539
rect 57897 4505 57931 4539
rect 73721 4505 73755 4539
rect 74181 4505 74215 4539
rect 74397 4505 74431 4539
rect 79609 4505 79643 4539
rect 80345 4505 80379 4539
rect 89453 4505 89487 4539
rect 89637 4505 89671 4539
rect 89821 4505 89855 4539
rect 92857 4505 92891 4539
rect 10333 4437 10367 4471
rect 10793 4437 10827 4471
rect 15393 4437 15427 4471
rect 23949 4437 23983 4471
rect 33517 4437 33551 4471
rect 34897 4437 34931 4471
rect 42165 4437 42199 4471
rect 46397 4437 46431 4471
rect 47501 4437 47535 4471
rect 56425 4437 56459 4471
rect 58541 4437 58575 4471
rect 71237 4437 71271 4471
rect 77309 4437 77343 4471
rect 78597 4437 78631 4471
rect 79149 4437 79183 4471
rect 84577 4437 84611 4471
rect 85865 4437 85899 4471
rect 88993 4437 89027 4471
rect 90649 4437 90683 4471
rect 92397 4437 92431 4471
rect 93685 4437 93719 4471
rect 94237 4437 94271 4471
rect 34437 4233 34471 4267
rect 43269 4233 43303 4267
rect 51457 4233 51491 4267
rect 56609 4233 56643 4267
rect 59369 4233 59403 4267
rect 64337 4233 64371 4267
rect 75929 4233 75963 4267
rect 77493 4233 77527 4267
rect 84025 4233 84059 4267
rect 84209 4233 84243 4267
rect 86785 4233 86819 4267
rect 90281 4233 90315 4267
rect 91753 4233 91787 4267
rect 23029 4165 23063 4199
rect 25973 4165 26007 4199
rect 26157 4165 26191 4199
rect 33425 4165 33459 4199
rect 33609 4165 33643 4199
rect 53757 4165 53791 4199
rect 55505 4165 55539 4199
rect 71513 4165 71547 4199
rect 73537 4165 73571 4199
rect 78965 4165 78999 4199
rect 84117 4165 84151 4199
rect 90189 4165 90223 4199
rect 9597 4097 9631 4131
rect 9873 4097 9907 4131
rect 10609 4097 10643 4131
rect 14841 4097 14875 4131
rect 25513 4097 25547 4131
rect 33241 4097 33275 4131
rect 34621 4097 34655 4131
rect 39773 4097 39807 4131
rect 40325 4097 40359 4131
rect 41429 4097 41463 4131
rect 43821 4097 43855 4131
rect 52285 4097 52319 4131
rect 53205 4097 53239 4131
rect 58633 4097 58667 4131
rect 62037 4097 62071 4131
rect 62589 4097 62623 4131
rect 63785 4097 63819 4131
rect 65441 4097 65475 4131
rect 71237 4097 71271 4131
rect 73813 4097 73847 4131
rect 77401 4097 77435 4131
rect 80897 4097 80931 4131
rect 81541 4097 81575 4131
rect 83289 4097 83323 4131
rect 83841 4097 83875 4131
rect 84853 4097 84887 4131
rect 85497 4097 85531 4131
rect 86233 4097 86267 4131
rect 86969 4097 87003 4131
rect 87705 4097 87739 4131
rect 87981 4097 88015 4131
rect 90005 4097 90039 4131
rect 90281 4097 90315 4131
rect 90741 4097 90775 4131
rect 13093 4029 13127 4063
rect 14565 4029 14599 4063
rect 26341 4029 26375 4063
rect 37473 4029 37507 4063
rect 37749 4029 37783 4063
rect 39221 4029 39255 4063
rect 40785 4029 40819 4063
rect 49157 4029 49191 4063
rect 49433 4029 49467 4063
rect 50905 4029 50939 4063
rect 55137 4029 55171 4063
rect 55597 4029 55631 4063
rect 56149 4029 56183 4063
rect 57069 4029 57103 4063
rect 57529 4029 57563 4063
rect 60841 4029 60875 4063
rect 61117 4029 61151 4063
rect 72985 4029 73019 4063
rect 74365 4029 74399 4063
rect 75193 4029 75227 4063
rect 78689 4029 78723 4063
rect 80437 4029 80471 4063
rect 82185 4029 82219 4063
rect 93225 4029 93259 4063
rect 93501 4029 93535 4063
rect 94145 4029 94179 4063
rect 10793 3961 10827 3995
rect 56425 3961 56459 3995
rect 57345 3961 57379 3995
rect 64981 3961 65015 3995
rect 73721 3961 73755 3995
rect 84393 3961 84427 3995
rect 11805 3893 11839 3927
rect 36921 3893 36955 3927
rect 58173 3893 58207 3927
rect 63233 3893 63267 3927
rect 65993 3893 66027 3927
rect 68385 3893 68419 3927
rect 73629 3893 73663 3927
rect 76481 3893 76515 3927
rect 78045 3893 78079 3927
rect 82645 3893 82679 3927
rect 88993 3893 89027 3927
rect 14289 3689 14323 3723
rect 59277 3689 59311 3723
rect 61485 3689 61519 3723
rect 68569 3689 68603 3723
rect 86417 3689 86451 3723
rect 87429 3689 87463 3723
rect 90833 3689 90867 3723
rect 93225 3689 93259 3723
rect 40049 3621 40083 3655
rect 51089 3621 51123 3655
rect 54217 3621 54251 3655
rect 54677 3621 54711 3655
rect 60749 3621 60783 3655
rect 64521 3621 64555 3655
rect 72065 3621 72099 3655
rect 72157 3621 72191 3655
rect 76113 3621 76147 3655
rect 76849 3621 76883 3655
rect 80713 3621 80747 3655
rect 83473 3621 83507 3655
rect 87889 3621 87923 3655
rect 88441 3621 88475 3655
rect 92673 3621 92707 3655
rect 39405 3553 39439 3587
rect 51917 3553 51951 3587
rect 55965 3553 55999 3587
rect 64061 3553 64095 3587
rect 71513 3553 71547 3587
rect 71973 3553 72007 3587
rect 80069 3553 80103 3587
rect 83933 3553 83967 3587
rect 85313 3553 85347 3587
rect 89361 3553 89395 3587
rect 14473 3485 14507 3519
rect 15209 3485 15243 3519
rect 15485 3485 15519 3519
rect 53665 3485 53699 3519
rect 55689 3485 55723 3519
rect 57897 3485 57931 3519
rect 62037 3485 62071 3519
rect 65165 3485 65199 3519
rect 67925 3485 67959 3519
rect 72249 3485 72283 3519
rect 79609 3485 79643 3519
rect 81725 3485 81759 3519
rect 82001 3485 82035 3519
rect 82737 3485 82771 3519
rect 84853 3485 84887 3519
rect 86969 3485 87003 3519
rect 87061 3485 87095 3519
rect 87245 3485 87279 3519
rect 89085 3485 89119 3519
rect 91937 3485 91971 3519
rect 94053 3485 94087 3519
rect 15945 3417 15979 3451
rect 39129 3417 39163 3451
rect 53389 3417 53423 3451
rect 58449 3417 58483 3451
rect 63785 3417 63819 3451
rect 65809 3417 65843 3451
rect 73353 3417 73387 3451
rect 79333 3417 79367 3451
rect 82921 3417 82955 3451
rect 37657 3349 37691 3383
rect 57437 3349 57471 3383
rect 68109 3349 68143 3383
rect 72893 3349 72927 3383
rect 73997 3349 74031 3383
rect 77861 3349 77895 3383
rect 92121 3349 92155 3383
rect 94237 3349 94271 3383
rect 37565 3145 37599 3179
rect 53849 3145 53883 3179
rect 54401 3145 54435 3179
rect 54953 3145 54987 3179
rect 55505 3145 55539 3179
rect 56241 3145 56275 3179
rect 57161 3145 57195 3179
rect 79241 3145 79275 3179
rect 80621 3145 80655 3179
rect 81541 3145 81575 3179
rect 85221 3145 85255 3179
rect 85957 3145 85991 3179
rect 90465 3145 90499 3179
rect 91017 3145 91051 3179
rect 92029 3145 92063 3179
rect 39037 3077 39071 3111
rect 39773 3077 39807 3111
rect 53021 3077 53055 3111
rect 61301 3077 61335 3111
rect 64705 3077 64739 3111
rect 76297 3077 76331 3111
rect 77493 3077 77527 3111
rect 78045 3077 78079 3111
rect 89821 3077 89855 3111
rect 39313 3009 39347 3043
rect 51273 3009 51307 3043
rect 51825 3009 51859 3043
rect 78873 3009 78907 3043
rect 79885 3009 79919 3043
rect 86601 3009 86635 3043
rect 87153 3009 87187 3043
rect 64981 2941 65015 2975
rect 65441 2941 65475 2975
rect 78781 2941 78815 2975
rect 82645 2941 82679 2975
rect 83197 2941 83231 2975
rect 84761 2941 84795 2975
rect 63233 2873 63267 2907
rect 92489 2873 92523 2907
rect 79701 2805 79735 2839
rect 36369 2601 36403 2635
rect 39405 2601 39439 2635
rect 44097 2601 44131 2635
rect 54401 2601 54435 2635
rect 64337 2601 64371 2635
rect 78781 2601 78815 2635
rect 86877 2601 86911 2635
rect 90925 2601 90959 2635
rect 53389 2533 53423 2567
rect 83841 2465 83875 2499
rect 91845 2465 91879 2499
rect 4537 2397 4571 2431
rect 12725 2397 12759 2431
rect 13369 2397 13403 2431
rect 20085 2397 20119 2431
rect 21005 2397 21039 2431
rect 28457 2397 28491 2431
rect 36185 2397 36219 2431
rect 36829 2397 36863 2431
rect 44281 2397 44315 2431
rect 52285 2397 52319 2431
rect 53573 2397 53607 2431
rect 60933 2397 60967 2431
rect 68385 2397 68419 2431
rect 75193 2397 75227 2431
rect 76113 2397 76147 2431
rect 91569 2397 91603 2431
rect 92857 2397 92891 2431
rect 61485 2329 61519 2363
rect 84025 2329 84059 2363
rect 4721 2261 4755 2295
rect 12541 2261 12575 2295
rect 13185 2261 13219 2295
rect 20269 2261 20303 2295
rect 20821 2261 20855 2295
rect 28273 2261 28307 2295
rect 43637 2261 43671 2295
rect 52101 2261 52135 2295
rect 60749 2261 60783 2295
rect 68569 2261 68603 2295
rect 75377 2261 75411 2295
rect 76297 2261 76331 2295
rect 83289 2261 83323 2295
<< metal1 >>
rect 20898 17484 20904 17536
rect 20956 17524 20962 17536
rect 69658 17524 69664 17536
rect 20956 17496 69664 17524
rect 20956 17484 20962 17496
rect 69658 17484 69664 17496
rect 69716 17484 69722 17536
rect 1104 17434 95011 17456
rect 1104 17382 24386 17434
rect 24438 17382 24450 17434
rect 24502 17382 24514 17434
rect 24566 17382 24578 17434
rect 24630 17382 24642 17434
rect 24694 17382 47823 17434
rect 47875 17382 47887 17434
rect 47939 17382 47951 17434
rect 48003 17382 48015 17434
rect 48067 17382 48079 17434
rect 48131 17382 71260 17434
rect 71312 17382 71324 17434
rect 71376 17382 71388 17434
rect 71440 17382 71452 17434
rect 71504 17382 71516 17434
rect 71568 17382 94697 17434
rect 94749 17382 94761 17434
rect 94813 17382 94825 17434
rect 94877 17382 94889 17434
rect 94941 17382 94953 17434
rect 95005 17382 95011 17434
rect 1104 17360 95011 17382
rect 4430 17280 4436 17332
rect 4488 17320 4494 17332
rect 4617 17323 4675 17329
rect 4617 17320 4629 17323
rect 4488 17292 4629 17320
rect 4488 17280 4494 17292
rect 4617 17289 4629 17292
rect 4663 17289 4675 17323
rect 4617 17283 4675 17289
rect 5261 17323 5319 17329
rect 5261 17289 5273 17323
rect 5307 17289 5319 17323
rect 5261 17283 5319 17289
rect 1578 17144 1584 17196
rect 1636 17184 1642 17196
rect 1673 17187 1731 17193
rect 1673 17184 1685 17187
rect 1636 17156 1685 17184
rect 1636 17144 1642 17156
rect 1673 17153 1685 17156
rect 1719 17153 1731 17187
rect 1673 17147 1731 17153
rect 4801 17187 4859 17193
rect 4801 17153 4813 17187
rect 4847 17184 4859 17187
rect 5276 17184 5304 17283
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 12621 17323 12679 17329
rect 12621 17320 12633 17323
rect 12492 17292 12633 17320
rect 12492 17280 12498 17292
rect 12621 17289 12633 17292
rect 12667 17289 12679 17323
rect 12621 17283 12679 17289
rect 20254 17280 20260 17332
rect 20312 17320 20318 17332
rect 20349 17323 20407 17329
rect 20349 17320 20361 17323
rect 20312 17292 20361 17320
rect 20312 17280 20318 17292
rect 20349 17289 20361 17292
rect 20395 17289 20407 17323
rect 20349 17283 20407 17289
rect 28166 17280 28172 17332
rect 28224 17320 28230 17332
rect 28261 17323 28319 17329
rect 28261 17320 28273 17323
rect 28224 17292 28273 17320
rect 28224 17280 28230 17292
rect 28261 17289 28273 17292
rect 28307 17289 28319 17323
rect 43625 17323 43683 17329
rect 28261 17283 28319 17289
rect 31726 17292 41414 17320
rect 31726 17252 31754 17292
rect 34330 17252 34336 17264
rect 6656 17224 31754 17252
rect 34243 17224 34336 17252
rect 4847 17156 5304 17184
rect 5445 17187 5503 17193
rect 4847 17153 4859 17156
rect 4801 17147 4859 17153
rect 5445 17153 5457 17187
rect 5491 17184 5503 17187
rect 6546 17184 6552 17196
rect 5491 17156 6552 17184
rect 5491 17153 5503 17156
rect 5445 17147 5503 17153
rect 6546 17144 6552 17156
rect 6604 17144 6610 17196
rect 1949 16983 2007 16989
rect 1949 16949 1961 16983
rect 1995 16980 2007 16983
rect 5074 16980 5080 16992
rect 1995 16952 5080 16980
rect 1995 16949 2007 16952
rect 1949 16943 2007 16949
rect 5074 16940 5080 16952
rect 5132 16980 5138 16992
rect 6656 16980 6684 17224
rect 34330 17212 34336 17224
rect 34388 17252 34394 17264
rect 41386 17252 41414 17292
rect 43625 17289 43637 17323
rect 43671 17320 43683 17323
rect 43990 17320 43996 17332
rect 43671 17292 43996 17320
rect 43671 17289 43683 17292
rect 43625 17283 43683 17289
rect 43990 17280 43996 17292
rect 44048 17280 44054 17332
rect 50338 17320 50344 17332
rect 46032 17292 50344 17320
rect 46032 17252 46060 17292
rect 50338 17280 50344 17292
rect 50396 17280 50402 17332
rect 51902 17280 51908 17332
rect 51960 17320 51966 17332
rect 52089 17323 52147 17329
rect 52089 17320 52101 17323
rect 51960 17292 52101 17320
rect 51960 17280 51966 17292
rect 52089 17289 52101 17292
rect 52135 17289 52147 17323
rect 52089 17283 52147 17289
rect 59814 17280 59820 17332
rect 59872 17320 59878 17332
rect 59909 17323 59967 17329
rect 59909 17320 59921 17323
rect 59872 17292 59921 17320
rect 59872 17280 59878 17292
rect 59909 17289 59921 17292
rect 59955 17289 59967 17323
rect 59909 17283 59967 17289
rect 67726 17280 67732 17332
rect 67784 17320 67790 17332
rect 68557 17323 68615 17329
rect 68557 17320 68569 17323
rect 67784 17292 68569 17320
rect 67784 17280 67790 17292
rect 68557 17289 68569 17292
rect 68603 17289 68615 17323
rect 68557 17283 68615 17289
rect 75638 17280 75644 17332
rect 75696 17320 75702 17332
rect 76285 17323 76343 17329
rect 76285 17320 76297 17323
rect 75696 17292 76297 17320
rect 75696 17280 75702 17292
rect 76285 17289 76297 17292
rect 76331 17289 76343 17323
rect 91557 17323 91615 17329
rect 91557 17320 91569 17323
rect 76285 17283 76343 17289
rect 89686 17292 91569 17320
rect 49510 17252 49516 17264
rect 34388 17224 35466 17252
rect 41386 17224 46060 17252
rect 46124 17224 49516 17252
rect 34388 17212 34394 17224
rect 11882 17144 11888 17196
rect 11940 17184 11946 17196
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 11940 17156 12449 17184
rect 11940 17144 11946 17156
rect 12437 17153 12449 17156
rect 12483 17153 12495 17187
rect 20530 17184 20536 17196
rect 20491 17156 20536 17184
rect 12437 17147 12495 17153
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 28442 17184 28448 17196
rect 28403 17156 28448 17184
rect 28442 17144 28448 17156
rect 28500 17144 28506 17196
rect 43990 17144 43996 17196
rect 44048 17184 44054 17196
rect 44269 17187 44327 17193
rect 44269 17184 44281 17187
rect 44048 17156 44281 17184
rect 44048 17144 44054 17156
rect 44269 17153 44281 17156
rect 44315 17153 44327 17187
rect 44269 17147 44327 17153
rect 34882 17116 34888 17128
rect 34843 17088 34888 17116
rect 34882 17076 34888 17088
rect 34940 17076 34946 17128
rect 36633 17119 36691 17125
rect 36633 17085 36645 17119
rect 36679 17116 36691 17119
rect 36679 17088 36860 17116
rect 36679 17085 36691 17088
rect 36633 17079 36691 17085
rect 36832 17048 36860 17088
rect 36906 17076 36912 17128
rect 36964 17116 36970 17128
rect 37553 17119 37611 17125
rect 37553 17116 37565 17119
rect 36964 17088 37565 17116
rect 36964 17076 36970 17088
rect 37553 17085 37565 17088
rect 37599 17116 37611 17119
rect 46124 17116 46152 17224
rect 49510 17212 49516 17224
rect 49568 17252 49574 17264
rect 55953 17255 56011 17261
rect 55953 17252 55965 17255
rect 49568 17224 55965 17252
rect 49568 17212 49574 17224
rect 55953 17221 55965 17224
rect 55999 17252 56011 17255
rect 57054 17252 57060 17264
rect 55999 17224 57060 17252
rect 55999 17221 56011 17224
rect 55953 17215 56011 17221
rect 57054 17212 57060 17224
rect 57112 17212 57118 17264
rect 65886 17252 65892 17264
rect 60108 17224 65892 17252
rect 52270 17184 52276 17196
rect 52231 17156 52276 17184
rect 52270 17144 52276 17156
rect 52328 17144 52334 17196
rect 60108 17193 60136 17224
rect 65886 17212 65892 17224
rect 65944 17212 65950 17264
rect 83277 17255 83335 17261
rect 83277 17221 83289 17255
rect 83323 17252 83335 17255
rect 84010 17252 84016 17264
rect 83323 17224 84016 17252
rect 83323 17221 83335 17224
rect 83277 17215 83335 17221
rect 84010 17212 84016 17224
rect 84068 17252 84074 17264
rect 85577 17255 85635 17261
rect 84068 17224 84410 17252
rect 84068 17212 84074 17224
rect 85577 17221 85589 17255
rect 85623 17252 85635 17255
rect 89686 17252 89714 17292
rect 91557 17289 91569 17292
rect 91603 17289 91615 17323
rect 91557 17283 91615 17289
rect 85623 17224 89714 17252
rect 85623 17221 85635 17224
rect 85577 17215 85635 17221
rect 58805 17187 58863 17193
rect 58805 17153 58817 17187
rect 58851 17184 58863 17187
rect 60093 17187 60151 17193
rect 60093 17184 60105 17187
rect 58851 17156 60105 17184
rect 58851 17153 58863 17156
rect 58805 17147 58863 17153
rect 60093 17153 60105 17156
rect 60139 17153 60151 17187
rect 61289 17187 61347 17193
rect 61289 17184 61301 17187
rect 60093 17147 60151 17153
rect 60706 17156 61301 17184
rect 37599 17088 46152 17116
rect 37599 17085 37611 17088
rect 37553 17079 37611 17085
rect 46198 17076 46204 17128
rect 46256 17116 46262 17128
rect 59354 17116 59360 17128
rect 46256 17088 59360 17116
rect 46256 17076 46262 17088
rect 59354 17076 59360 17088
rect 59412 17076 59418 17128
rect 44085 17051 44143 17057
rect 44085 17048 44097 17051
rect 36832 17020 44097 17048
rect 44085 17017 44097 17020
rect 44131 17017 44143 17051
rect 44085 17011 44143 17017
rect 55122 17008 55128 17060
rect 55180 17048 55186 17060
rect 57057 17051 57115 17057
rect 57057 17048 57069 17051
rect 55180 17020 57069 17048
rect 55180 17008 55186 17020
rect 57057 17017 57069 17020
rect 57103 17048 57115 17051
rect 57974 17048 57980 17060
rect 57103 17020 57980 17048
rect 57103 17017 57115 17020
rect 57057 17011 57115 17017
rect 57974 17008 57980 17020
rect 58032 17048 58038 17060
rect 60706 17048 60734 17156
rect 61289 17153 61301 17156
rect 61335 17184 61347 17187
rect 62301 17187 62359 17193
rect 62301 17184 62313 17187
rect 61335 17156 62313 17184
rect 61335 17153 61347 17156
rect 61289 17147 61347 17153
rect 62301 17153 62313 17156
rect 62347 17153 62359 17187
rect 68370 17184 68376 17196
rect 68331 17156 68376 17184
rect 62301 17147 62359 17153
rect 68370 17144 68376 17156
rect 68428 17144 68434 17196
rect 76098 17184 76104 17196
rect 76059 17156 76104 17184
rect 76098 17144 76104 17156
rect 76156 17144 76162 17196
rect 91462 17144 91468 17196
rect 91520 17184 91526 17196
rect 91741 17187 91799 17193
rect 91741 17184 91753 17187
rect 91520 17156 91753 17184
rect 91520 17144 91526 17156
rect 91741 17153 91753 17156
rect 91787 17184 91799 17187
rect 92201 17187 92259 17193
rect 92201 17184 92213 17187
rect 91787 17156 92213 17184
rect 91787 17153 91799 17156
rect 91741 17147 91799 17153
rect 92201 17153 92213 17156
rect 92247 17153 92259 17187
rect 92201 17147 92259 17153
rect 61105 17119 61163 17125
rect 61105 17085 61117 17119
rect 61151 17116 61163 17119
rect 61838 17116 61844 17128
rect 61151 17088 61844 17116
rect 61151 17085 61163 17088
rect 61105 17079 61163 17085
rect 61838 17076 61844 17088
rect 61896 17116 61902 17128
rect 63221 17119 63279 17125
rect 63221 17116 63233 17119
rect 61896 17088 63233 17116
rect 61896 17076 61902 17088
rect 63221 17085 63233 17088
rect 63267 17116 63279 17119
rect 63586 17116 63592 17128
rect 63267 17088 63592 17116
rect 63267 17085 63279 17088
rect 63221 17079 63279 17085
rect 63586 17076 63592 17088
rect 63644 17116 63650 17128
rect 64325 17119 64383 17125
rect 64325 17116 64337 17119
rect 63644 17088 64337 17116
rect 63644 17076 63650 17088
rect 64325 17085 64337 17088
rect 64371 17116 64383 17119
rect 65794 17116 65800 17128
rect 64371 17088 65800 17116
rect 64371 17085 64383 17088
rect 64325 17079 64383 17085
rect 65794 17076 65800 17088
rect 65852 17076 65858 17128
rect 83366 17076 83372 17128
rect 83424 17116 83430 17128
rect 83829 17119 83887 17125
rect 83829 17116 83841 17119
rect 83424 17088 83841 17116
rect 83424 17076 83430 17088
rect 83829 17085 83841 17088
rect 83875 17085 83887 17119
rect 85853 17119 85911 17125
rect 85853 17116 85865 17119
rect 83829 17079 83887 17085
rect 84028 17088 85865 17116
rect 58032 17020 60734 17048
rect 58032 17008 58038 17020
rect 62850 17008 62856 17060
rect 62908 17048 62914 17060
rect 63865 17051 63923 17057
rect 63865 17048 63877 17051
rect 62908 17020 63877 17048
rect 62908 17008 62914 17020
rect 63865 17017 63877 17020
rect 63911 17048 63923 17051
rect 64969 17051 65027 17057
rect 64969 17048 64981 17051
rect 63911 17020 64981 17048
rect 63911 17017 63923 17020
rect 63865 17011 63923 17017
rect 64969 17017 64981 17020
rect 65015 17048 65027 17051
rect 67542 17048 67548 17060
rect 65015 17020 67548 17048
rect 65015 17017 65027 17020
rect 64969 17011 65027 17017
rect 67542 17008 67548 17020
rect 67600 17048 67606 17060
rect 67729 17051 67787 17057
rect 67729 17048 67741 17051
rect 67600 17020 67741 17048
rect 67600 17008 67606 17020
rect 67729 17017 67741 17020
rect 67775 17048 67787 17051
rect 83734 17048 83740 17060
rect 67775 17020 83740 17048
rect 67775 17017 67787 17020
rect 67729 17011 67787 17017
rect 83734 17008 83740 17020
rect 83792 17048 83798 17060
rect 84028 17048 84056 17088
rect 85853 17085 85865 17088
rect 85899 17116 85911 17119
rect 86405 17119 86463 17125
rect 86405 17116 86417 17119
rect 85899 17088 86417 17116
rect 85899 17085 85911 17088
rect 85853 17079 85911 17085
rect 86405 17085 86417 17088
rect 86451 17085 86463 17119
rect 86405 17079 86463 17085
rect 83792 17020 84056 17048
rect 83792 17008 83798 17020
rect 5132 16952 6684 16980
rect 5132 16940 5138 16952
rect 32214 16940 32220 16992
rect 32272 16980 32278 16992
rect 38654 16980 38660 16992
rect 32272 16952 38660 16980
rect 32272 16940 32278 16952
rect 38654 16940 38660 16952
rect 38712 16940 38718 16992
rect 40586 16940 40592 16992
rect 40644 16980 40650 16992
rect 42613 16983 42671 16989
rect 42613 16980 42625 16983
rect 40644 16952 42625 16980
rect 40644 16940 40650 16952
rect 42613 16949 42625 16952
rect 42659 16949 42671 16983
rect 42613 16943 42671 16949
rect 45925 16983 45983 16989
rect 45925 16949 45937 16983
rect 45971 16980 45983 16983
rect 46014 16980 46020 16992
rect 45971 16952 46020 16980
rect 45971 16949 45983 16952
rect 45925 16943 45983 16949
rect 46014 16940 46020 16952
rect 46072 16940 46078 16992
rect 46474 16980 46480 16992
rect 46435 16952 46480 16980
rect 46474 16940 46480 16952
rect 46532 16940 46538 16992
rect 47026 16980 47032 16992
rect 46987 16952 47032 16980
rect 47026 16940 47032 16952
rect 47084 16940 47090 16992
rect 56597 16983 56655 16989
rect 56597 16949 56609 16983
rect 56643 16980 56655 16983
rect 56686 16980 56692 16992
rect 56643 16952 56692 16980
rect 56643 16949 56655 16952
rect 56597 16943 56655 16949
rect 56686 16940 56692 16952
rect 56744 16940 56750 16992
rect 59357 16983 59415 16989
rect 59357 16949 59369 16983
rect 59403 16980 59415 16983
rect 60734 16980 60740 16992
rect 59403 16952 60740 16980
rect 59403 16949 59415 16952
rect 59357 16943 59415 16949
rect 60734 16940 60740 16952
rect 60792 16940 60798 16992
rect 61102 16940 61108 16992
rect 61160 16980 61166 16992
rect 61749 16983 61807 16989
rect 61749 16980 61761 16983
rect 61160 16952 61761 16980
rect 61160 16940 61166 16952
rect 61749 16949 61761 16952
rect 61795 16949 61807 16983
rect 61749 16943 61807 16949
rect 1104 16890 94852 16912
rect 1104 16838 12668 16890
rect 12720 16838 12732 16890
rect 12784 16838 12796 16890
rect 12848 16838 12860 16890
rect 12912 16838 12924 16890
rect 12976 16838 36105 16890
rect 36157 16838 36169 16890
rect 36221 16838 36233 16890
rect 36285 16838 36297 16890
rect 36349 16838 36361 16890
rect 36413 16838 59542 16890
rect 59594 16838 59606 16890
rect 59658 16838 59670 16890
rect 59722 16838 59734 16890
rect 59786 16838 59798 16890
rect 59850 16838 82979 16890
rect 83031 16838 83043 16890
rect 83095 16838 83107 16890
rect 83159 16838 83171 16890
rect 83223 16838 83235 16890
rect 83287 16838 94852 16890
rect 1104 16816 94852 16838
rect 36357 16779 36415 16785
rect 36357 16745 36369 16779
rect 36403 16776 36415 16779
rect 36906 16776 36912 16788
rect 36403 16748 36912 16776
rect 36403 16745 36415 16748
rect 36357 16739 36415 16745
rect 36906 16736 36912 16748
rect 36964 16736 36970 16788
rect 38654 16736 38660 16788
rect 38712 16776 38718 16788
rect 38749 16779 38807 16785
rect 38749 16776 38761 16779
rect 38712 16748 38761 16776
rect 38712 16736 38718 16748
rect 38749 16745 38761 16748
rect 38795 16776 38807 16779
rect 46198 16776 46204 16788
rect 38795 16748 46204 16776
rect 38795 16745 38807 16748
rect 38749 16739 38807 16745
rect 46198 16736 46204 16748
rect 46256 16736 46262 16788
rect 50338 16776 50344 16788
rect 50299 16748 50344 16776
rect 50338 16736 50344 16748
rect 50396 16736 50402 16788
rect 50522 16736 50528 16788
rect 50580 16776 50586 16788
rect 55122 16776 55128 16788
rect 50580 16748 55128 16776
rect 50580 16736 50586 16748
rect 55122 16736 55128 16748
rect 55180 16736 55186 16788
rect 57054 16736 57060 16788
rect 57112 16776 57118 16788
rect 60645 16779 60703 16785
rect 57112 16748 59216 16776
rect 57112 16736 57118 16748
rect 1578 16708 1584 16720
rect 1539 16680 1584 16708
rect 1578 16668 1584 16680
rect 1636 16668 1642 16720
rect 24302 16668 24308 16720
rect 24360 16708 24366 16720
rect 47026 16708 47032 16720
rect 24360 16680 47032 16708
rect 24360 16668 24366 16680
rect 47026 16668 47032 16680
rect 47084 16708 47090 16720
rect 54938 16708 54944 16720
rect 47084 16680 47532 16708
rect 54899 16680 54944 16708
rect 47084 16668 47090 16680
rect 20346 16640 20352 16652
rect 20307 16612 20352 16640
rect 20346 16600 20352 16612
rect 20404 16600 20410 16652
rect 31757 16643 31815 16649
rect 31757 16609 31769 16643
rect 31803 16640 31815 16643
rect 31846 16640 31852 16652
rect 31803 16612 31852 16640
rect 31803 16609 31815 16612
rect 31757 16603 31815 16609
rect 31846 16600 31852 16612
rect 31904 16600 31910 16652
rect 35713 16643 35771 16649
rect 35713 16609 35725 16643
rect 35759 16640 35771 16643
rect 35759 16612 36032 16640
rect 35759 16609 35771 16612
rect 35713 16603 35771 16609
rect 36004 16584 36032 16612
rect 40126 16600 40132 16652
rect 40184 16640 40190 16652
rect 41049 16643 41107 16649
rect 41049 16640 41061 16643
rect 40184 16612 41061 16640
rect 40184 16600 40190 16612
rect 41049 16609 41061 16612
rect 41095 16640 41107 16643
rect 41693 16643 41751 16649
rect 41693 16640 41705 16643
rect 41095 16612 41705 16640
rect 41095 16609 41107 16612
rect 41049 16603 41107 16609
rect 41693 16609 41705 16612
rect 41739 16609 41751 16643
rect 42334 16640 42340 16652
rect 42295 16612 42340 16640
rect 41693 16603 41751 16609
rect 42334 16600 42340 16612
rect 42392 16600 42398 16652
rect 42426 16600 42432 16652
rect 42484 16640 42490 16652
rect 42797 16643 42855 16649
rect 42797 16640 42809 16643
rect 42484 16612 42809 16640
rect 42484 16600 42490 16612
rect 42797 16609 42809 16612
rect 42843 16609 42855 16643
rect 42797 16603 42855 16609
rect 45281 16643 45339 16649
rect 45281 16609 45293 16643
rect 45327 16640 45339 16643
rect 45830 16640 45836 16652
rect 45327 16612 45836 16640
rect 45327 16609 45339 16612
rect 45281 16603 45339 16609
rect 45830 16600 45836 16612
rect 45888 16600 45894 16652
rect 46201 16643 46259 16649
rect 46201 16609 46213 16643
rect 46247 16640 46259 16643
rect 46382 16640 46388 16652
rect 46247 16612 46388 16640
rect 46247 16609 46259 16612
rect 46201 16603 46259 16609
rect 46382 16600 46388 16612
rect 46440 16600 46446 16652
rect 46566 16600 46572 16652
rect 46624 16640 46630 16652
rect 47504 16649 47532 16680
rect 54938 16668 54944 16680
rect 54996 16668 55002 16720
rect 59188 16708 59216 16748
rect 60645 16745 60657 16779
rect 60691 16776 60703 16779
rect 62022 16776 62028 16788
rect 60691 16748 62028 16776
rect 60691 16745 60703 16748
rect 60645 16739 60703 16745
rect 62022 16736 62028 16748
rect 62080 16736 62086 16788
rect 65886 16736 65892 16788
rect 65944 16776 65950 16788
rect 65944 16748 83688 16776
rect 65944 16736 65950 16748
rect 61102 16708 61108 16720
rect 59188 16680 61108 16708
rect 61102 16668 61108 16680
rect 61160 16668 61166 16720
rect 68097 16711 68155 16717
rect 68097 16677 68109 16711
rect 68143 16708 68155 16711
rect 68186 16708 68192 16720
rect 68143 16680 68192 16708
rect 68143 16677 68155 16680
rect 68097 16671 68155 16677
rect 68186 16668 68192 16680
rect 68244 16668 68250 16720
rect 68649 16711 68707 16717
rect 68649 16677 68661 16711
rect 68695 16708 68707 16711
rect 83366 16708 83372 16720
rect 68695 16680 83372 16708
rect 68695 16677 68707 16680
rect 68649 16671 68707 16677
rect 46661 16643 46719 16649
rect 46661 16640 46673 16643
rect 46624 16612 46673 16640
rect 46624 16600 46630 16612
rect 46661 16609 46673 16612
rect 46707 16609 46719 16643
rect 47489 16643 47547 16649
rect 46661 16603 46719 16609
rect 47136 16612 47440 16640
rect 19705 16575 19763 16581
rect 19705 16541 19717 16575
rect 19751 16572 19763 16575
rect 20622 16572 20628 16584
rect 19751 16544 20628 16572
rect 19751 16541 19763 16544
rect 19705 16535 19763 16541
rect 20622 16532 20628 16544
rect 20680 16532 20686 16584
rect 35986 16572 35992 16584
rect 35899 16544 35992 16572
rect 35986 16532 35992 16544
rect 36044 16572 36050 16584
rect 36265 16575 36323 16581
rect 36265 16572 36277 16575
rect 36044 16544 36277 16572
rect 36044 16532 36050 16544
rect 36265 16541 36277 16544
rect 36311 16541 36323 16575
rect 47136 16572 47164 16612
rect 36265 16535 36323 16541
rect 40696 16544 47164 16572
rect 47305 16575 47363 16581
rect 29362 16464 29368 16516
rect 29420 16504 29426 16516
rect 40696 16504 40724 16544
rect 47305 16541 47317 16575
rect 47351 16541 47363 16575
rect 47412 16572 47440 16612
rect 47489 16609 47501 16643
rect 47535 16640 47547 16643
rect 53558 16640 53564 16652
rect 47535 16612 53564 16640
rect 47535 16609 47547 16612
rect 47489 16603 47547 16609
rect 53558 16600 53564 16612
rect 53616 16600 53622 16652
rect 55950 16600 55956 16652
rect 56008 16640 56014 16652
rect 56045 16643 56103 16649
rect 56045 16640 56057 16643
rect 56008 16612 56057 16640
rect 56008 16600 56014 16612
rect 56045 16609 56057 16612
rect 56091 16609 56103 16643
rect 56778 16640 56784 16652
rect 56739 16612 56784 16640
rect 56045 16603 56103 16609
rect 56778 16600 56784 16612
rect 56836 16600 56842 16652
rect 57330 16640 57336 16652
rect 57291 16612 57336 16640
rect 57330 16600 57336 16612
rect 57388 16600 57394 16652
rect 58713 16643 58771 16649
rect 58713 16609 58725 16643
rect 58759 16640 58771 16643
rect 59446 16640 59452 16652
rect 58759 16612 59452 16640
rect 58759 16609 58771 16612
rect 58713 16603 58771 16609
rect 59446 16600 59452 16612
rect 59504 16600 59510 16652
rect 62117 16643 62175 16649
rect 60016 16612 60320 16640
rect 59906 16572 59912 16584
rect 47412 16544 55904 16572
rect 59867 16544 59912 16572
rect 47305 16535 47363 16541
rect 29420 16476 40724 16504
rect 29420 16464 29426 16476
rect 40770 16464 40776 16516
rect 40828 16504 40834 16516
rect 47118 16504 47124 16516
rect 40828 16476 47124 16504
rect 40828 16464 40834 16476
rect 47118 16464 47124 16476
rect 47176 16464 47182 16516
rect 19610 16436 19616 16448
rect 19571 16408 19616 16436
rect 19610 16396 19616 16408
rect 19668 16396 19674 16448
rect 32214 16436 32220 16448
rect 32175 16408 32220 16436
rect 32214 16396 32220 16408
rect 32272 16396 32278 16448
rect 32858 16436 32864 16448
rect 32819 16408 32864 16436
rect 32858 16396 32864 16408
rect 32916 16396 32922 16448
rect 39574 16396 39580 16448
rect 39632 16436 39638 16448
rect 43533 16439 43591 16445
rect 43533 16436 43545 16439
rect 39632 16408 43545 16436
rect 39632 16396 39638 16408
rect 43533 16405 43545 16408
rect 43579 16436 43591 16439
rect 43714 16436 43720 16448
rect 43579 16408 43720 16436
rect 43579 16405 43591 16408
rect 43533 16399 43591 16405
rect 43714 16396 43720 16408
rect 43772 16396 43778 16448
rect 44818 16396 44824 16448
rect 44876 16436 44882 16448
rect 47320 16436 47348 16535
rect 47394 16464 47400 16516
rect 47452 16504 47458 16516
rect 51810 16504 51816 16516
rect 47452 16476 51816 16504
rect 47452 16464 47458 16476
rect 51810 16464 51816 16476
rect 51868 16464 51874 16516
rect 53101 16507 53159 16513
rect 53101 16504 53113 16507
rect 51920 16476 53113 16504
rect 48225 16439 48283 16445
rect 48225 16436 48237 16439
rect 44876 16408 48237 16436
rect 44876 16396 44882 16408
rect 48225 16405 48237 16408
rect 48271 16436 48283 16439
rect 48866 16436 48872 16448
rect 48271 16408 48872 16436
rect 48271 16405 48283 16408
rect 48225 16399 48283 16405
rect 48866 16396 48872 16408
rect 48924 16396 48930 16448
rect 51166 16396 51172 16448
rect 51224 16436 51230 16448
rect 51920 16436 51948 16476
rect 53101 16473 53113 16476
rect 53147 16473 53159 16507
rect 53101 16467 53159 16473
rect 54846 16464 54852 16516
rect 54904 16504 54910 16516
rect 55493 16507 55551 16513
rect 55493 16504 55505 16507
rect 54904 16476 55505 16504
rect 54904 16464 54910 16476
rect 55493 16473 55505 16476
rect 55539 16473 55551 16507
rect 55876 16504 55904 16544
rect 59906 16532 59912 16544
rect 59964 16532 59970 16584
rect 60016 16504 60044 16612
rect 60292 16572 60320 16612
rect 62117 16609 62129 16643
rect 62163 16640 62175 16643
rect 65518 16640 65524 16652
rect 62163 16612 65524 16640
rect 62163 16609 62175 16612
rect 62117 16603 62175 16609
rect 65518 16600 65524 16612
rect 65576 16640 65582 16652
rect 65797 16643 65855 16649
rect 65797 16640 65809 16643
rect 65576 16612 65809 16640
rect 65576 16600 65582 16612
rect 65797 16609 65809 16612
rect 65843 16609 65855 16643
rect 65797 16603 65855 16609
rect 67269 16643 67327 16649
rect 67269 16609 67281 16643
rect 67315 16640 67327 16643
rect 68664 16640 68692 16671
rect 83366 16668 83372 16680
rect 83424 16668 83430 16720
rect 83660 16708 83688 16748
rect 83734 16736 83740 16788
rect 83792 16776 83798 16788
rect 83829 16779 83887 16785
rect 83829 16776 83841 16779
rect 83792 16748 83841 16776
rect 83792 16736 83798 16748
rect 83829 16745 83841 16748
rect 83875 16745 83887 16779
rect 94222 16776 94228 16788
rect 94183 16748 94228 16776
rect 83829 16739 83887 16745
rect 94222 16736 94228 16748
rect 94280 16736 94286 16788
rect 87874 16708 87880 16720
rect 83660 16680 87880 16708
rect 87874 16668 87880 16680
rect 87932 16668 87938 16720
rect 67315 16612 68692 16640
rect 77021 16643 77079 16649
rect 67315 16609 67327 16612
rect 67269 16603 67327 16609
rect 77021 16609 77033 16643
rect 77067 16640 77079 16643
rect 77294 16640 77300 16652
rect 77067 16612 77300 16640
rect 77067 16609 77079 16612
rect 77021 16603 77079 16609
rect 77294 16600 77300 16612
rect 77352 16600 77358 16652
rect 93213 16643 93271 16649
rect 93213 16640 93225 16643
rect 92584 16612 93225 16640
rect 92584 16584 92612 16612
rect 93213 16609 93225 16612
rect 93259 16609 93271 16643
rect 93213 16603 93271 16609
rect 60826 16572 60832 16584
rect 60292 16544 60832 16572
rect 60826 16532 60832 16544
rect 60884 16532 60890 16584
rect 62393 16575 62451 16581
rect 62393 16541 62405 16575
rect 62439 16572 62451 16575
rect 62850 16572 62856 16584
rect 62439 16544 62856 16572
rect 62439 16541 62451 16544
rect 62393 16535 62451 16541
rect 62850 16532 62856 16544
rect 62908 16532 62914 16584
rect 67542 16532 67548 16584
rect 67600 16572 67606 16584
rect 83185 16575 83243 16581
rect 67600 16544 67645 16572
rect 67600 16532 67606 16544
rect 83185 16541 83197 16575
rect 83231 16572 83243 16575
rect 83550 16572 83556 16584
rect 83231 16544 83556 16572
rect 83231 16541 83243 16544
rect 83185 16535 83243 16541
rect 83550 16532 83556 16544
rect 83608 16572 83614 16584
rect 83737 16575 83795 16581
rect 83737 16572 83749 16575
rect 83608 16544 83749 16572
rect 83608 16532 83614 16544
rect 83737 16541 83749 16544
rect 83783 16541 83795 16575
rect 92566 16572 92572 16584
rect 92479 16544 92572 16572
rect 83737 16535 83795 16541
rect 92566 16532 92572 16544
rect 92624 16532 92630 16584
rect 94041 16575 94099 16581
rect 94041 16572 94053 16575
rect 92768 16544 94053 16572
rect 61838 16504 61844 16516
rect 55876 16476 60044 16504
rect 61686 16476 61844 16504
rect 55493 16467 55551 16473
rect 61838 16464 61844 16476
rect 61896 16464 61902 16516
rect 63129 16507 63187 16513
rect 63129 16473 63141 16507
rect 63175 16473 63187 16507
rect 63129 16467 63187 16473
rect 51224 16408 51948 16436
rect 51224 16396 51230 16408
rect 52362 16396 52368 16448
rect 52420 16436 52426 16448
rect 52457 16439 52515 16445
rect 52457 16436 52469 16439
rect 52420 16408 52469 16436
rect 52420 16396 52426 16408
rect 52457 16405 52469 16408
rect 52503 16405 52515 16439
rect 52457 16399 52515 16405
rect 54389 16439 54447 16445
rect 54389 16405 54401 16439
rect 54435 16436 54447 16439
rect 55214 16436 55220 16448
rect 54435 16408 55220 16436
rect 54435 16405 54447 16408
rect 54389 16399 54447 16405
rect 55214 16396 55220 16408
rect 55272 16396 55278 16448
rect 58158 16436 58164 16448
rect 58119 16408 58164 16436
rect 58158 16396 58164 16408
rect 58216 16396 58222 16448
rect 59170 16436 59176 16448
rect 59131 16408 59176 16436
rect 59170 16396 59176 16408
rect 59228 16396 59234 16448
rect 59998 16436 60004 16448
rect 59959 16408 60004 16436
rect 59998 16396 60004 16408
rect 60056 16396 60062 16448
rect 60090 16396 60096 16448
rect 60148 16436 60154 16448
rect 61930 16436 61936 16448
rect 60148 16408 61936 16436
rect 60148 16396 60154 16408
rect 61930 16396 61936 16408
rect 61988 16396 61994 16448
rect 62022 16396 62028 16448
rect 62080 16436 62086 16448
rect 63144 16436 63172 16467
rect 63586 16464 63592 16516
rect 63644 16464 63650 16516
rect 65794 16464 65800 16516
rect 65852 16504 65858 16516
rect 68738 16504 68744 16516
rect 65852 16476 66102 16504
rect 67606 16476 68744 16504
rect 65852 16464 65858 16476
rect 64598 16436 64604 16448
rect 62080 16408 63172 16436
rect 64559 16408 64604 16436
rect 62080 16396 62086 16408
rect 64598 16396 64604 16408
rect 64656 16396 64662 16448
rect 64966 16396 64972 16448
rect 65024 16436 65030 16448
rect 65061 16439 65119 16445
rect 65061 16436 65073 16439
rect 65024 16408 65073 16436
rect 65024 16396 65030 16408
rect 65061 16405 65073 16408
rect 65107 16405 65119 16439
rect 65996 16436 66024 16476
rect 67606 16436 67634 16476
rect 68738 16464 68744 16476
rect 68796 16464 68802 16516
rect 71958 16436 71964 16448
rect 65996 16408 67634 16436
rect 71919 16408 71964 16436
rect 65061 16399 65119 16405
rect 71958 16396 71964 16408
rect 72016 16396 72022 16448
rect 92768 16445 92796 16544
rect 94041 16541 94053 16544
rect 94087 16541 94099 16575
rect 94041 16535 94099 16541
rect 92753 16439 92811 16445
rect 92753 16405 92765 16439
rect 92799 16405 92811 16439
rect 92753 16399 92811 16405
rect 1104 16346 95011 16368
rect 1104 16294 24386 16346
rect 24438 16294 24450 16346
rect 24502 16294 24514 16346
rect 24566 16294 24578 16346
rect 24630 16294 24642 16346
rect 24694 16294 47823 16346
rect 47875 16294 47887 16346
rect 47939 16294 47951 16346
rect 48003 16294 48015 16346
rect 48067 16294 48079 16346
rect 48131 16294 71260 16346
rect 71312 16294 71324 16346
rect 71376 16294 71388 16346
rect 71440 16294 71452 16346
rect 71504 16294 71516 16346
rect 71568 16294 94697 16346
rect 94749 16294 94761 16346
rect 94813 16294 94825 16346
rect 94877 16294 94889 16346
rect 94941 16294 94953 16346
rect 95005 16294 95011 16346
rect 1104 16272 95011 16294
rect 20073 16235 20131 16241
rect 20073 16201 20085 16235
rect 20119 16232 20131 16235
rect 20119 16204 22094 16232
rect 20119 16201 20131 16204
rect 20073 16195 20131 16201
rect 19610 16124 19616 16176
rect 19668 16124 19674 16176
rect 20622 16056 20628 16108
rect 20680 16096 20686 16108
rect 20809 16099 20867 16105
rect 20809 16096 20821 16099
rect 20680 16068 20821 16096
rect 20680 16056 20686 16068
rect 20809 16065 20821 16068
rect 20855 16065 20867 16099
rect 20809 16059 20867 16065
rect 15378 15988 15384 16040
rect 15436 16028 15442 16040
rect 18325 16031 18383 16037
rect 18325 16028 18337 16031
rect 15436 16000 18337 16028
rect 15436 15988 15442 16000
rect 18325 15997 18337 16000
rect 18371 15997 18383 16031
rect 18325 15991 18383 15997
rect 18601 16031 18659 16037
rect 18601 15997 18613 16031
rect 18647 16028 18659 16031
rect 20346 16028 20352 16040
rect 18647 16000 20352 16028
rect 18647 15997 18659 16000
rect 18601 15991 18659 15997
rect 20346 15988 20352 16000
rect 20404 15988 20410 16040
rect 22066 16028 22094 16204
rect 32858 16192 32864 16244
rect 32916 16232 32922 16244
rect 39574 16232 39580 16244
rect 32916 16204 39580 16232
rect 32916 16192 32922 16204
rect 39574 16192 39580 16204
rect 39632 16192 39638 16244
rect 39684 16204 41414 16232
rect 31113 16167 31171 16173
rect 31113 16133 31125 16167
rect 31159 16164 31171 16167
rect 31386 16164 31392 16176
rect 31159 16136 31392 16164
rect 31159 16133 31171 16136
rect 31113 16127 31171 16133
rect 31386 16124 31392 16136
rect 31444 16124 31450 16176
rect 28997 16099 29055 16105
rect 28997 16065 29009 16099
rect 29043 16096 29055 16099
rect 29546 16096 29552 16108
rect 29043 16068 29552 16096
rect 29043 16065 29055 16068
rect 28997 16059 29055 16065
rect 29546 16056 29552 16068
rect 29604 16056 29610 16108
rect 30098 16056 30104 16108
rect 30156 16096 30162 16108
rect 30156 16094 39620 16096
rect 39684 16094 39712 16204
rect 39758 16124 39764 16176
rect 39816 16164 39822 16176
rect 40770 16164 40776 16176
rect 39816 16136 40776 16164
rect 39816 16124 39822 16136
rect 40770 16124 40776 16136
rect 40828 16124 40834 16176
rect 41386 16164 41414 16204
rect 41598 16192 41604 16244
rect 41656 16232 41662 16244
rect 44818 16232 44824 16244
rect 41656 16204 44824 16232
rect 41656 16192 41662 16204
rect 44818 16192 44824 16204
rect 44876 16192 44882 16244
rect 44913 16235 44971 16241
rect 44913 16201 44925 16235
rect 44959 16232 44971 16235
rect 46382 16232 46388 16244
rect 44959 16204 46388 16232
rect 44959 16201 44971 16204
rect 44913 16195 44971 16201
rect 46382 16192 46388 16204
rect 46440 16192 46446 16244
rect 46753 16235 46811 16241
rect 46753 16201 46765 16235
rect 46799 16232 46811 16235
rect 52086 16232 52092 16244
rect 46799 16204 52092 16232
rect 46799 16201 46811 16204
rect 46753 16195 46811 16201
rect 52086 16192 52092 16204
rect 52144 16192 52150 16244
rect 52181 16235 52239 16241
rect 52181 16201 52193 16235
rect 52227 16232 52239 16235
rect 52270 16232 52276 16244
rect 52227 16204 52276 16232
rect 52227 16201 52239 16204
rect 52181 16195 52239 16201
rect 52270 16192 52276 16204
rect 52328 16192 52334 16244
rect 52932 16204 61884 16232
rect 46474 16164 46480 16176
rect 41386 16136 46480 16164
rect 46474 16124 46480 16136
rect 46532 16164 46538 16176
rect 51442 16164 51448 16176
rect 46532 16136 46704 16164
rect 46532 16124 46538 16136
rect 40862 16096 40868 16108
rect 30156 16068 39712 16094
rect 40823 16068 40868 16096
rect 30156 16056 30162 16068
rect 39592 16066 39712 16068
rect 40862 16056 40868 16068
rect 40920 16056 40926 16108
rect 41509 16099 41567 16105
rect 41509 16065 41521 16099
rect 41555 16096 41567 16099
rect 42794 16096 42800 16108
rect 41555 16068 42800 16096
rect 41555 16065 41567 16068
rect 41509 16059 41567 16065
rect 39577 16031 39635 16037
rect 39577 16028 39589 16031
rect 22066 16000 39589 16028
rect 39577 15997 39589 16000
rect 39623 16028 39635 16031
rect 40129 16031 40187 16037
rect 40129 16028 40141 16031
rect 39623 16000 40141 16028
rect 39623 15997 39635 16000
rect 39577 15991 39635 15997
rect 40129 15997 40141 16000
rect 40175 16028 40187 16031
rect 40310 16028 40316 16040
rect 40175 16000 40316 16028
rect 40175 15997 40187 16000
rect 40129 15991 40187 15997
rect 40310 15988 40316 16000
rect 40368 15988 40374 16040
rect 40770 16028 40776 16040
rect 40731 16000 40776 16028
rect 40770 15988 40776 16000
rect 40828 15988 40834 16040
rect 40954 15988 40960 16040
rect 41012 16028 41018 16040
rect 41969 16031 42027 16037
rect 41969 16028 41981 16031
rect 41012 16000 41981 16028
rect 41012 15988 41018 16000
rect 41969 15997 41981 16000
rect 42015 15997 42027 16031
rect 41969 15991 42027 15997
rect 22094 15920 22100 15972
rect 22152 15960 22158 15972
rect 22152 15932 29684 15960
rect 22152 15920 22158 15932
rect 20714 15892 20720 15904
rect 20675 15864 20720 15892
rect 20714 15852 20720 15864
rect 20772 15852 20778 15904
rect 27706 15852 27712 15904
rect 27764 15892 27770 15904
rect 28905 15895 28963 15901
rect 28905 15892 28917 15895
rect 27764 15864 28917 15892
rect 27764 15852 27770 15864
rect 28905 15861 28917 15864
rect 28951 15861 28963 15895
rect 29546 15892 29552 15904
rect 29507 15864 29552 15892
rect 28905 15855 28963 15861
rect 29546 15852 29552 15864
rect 29604 15852 29610 15904
rect 29656 15892 29684 15932
rect 29730 15920 29736 15972
rect 29788 15960 29794 15972
rect 31573 15963 31631 15969
rect 31573 15960 31585 15963
rect 29788 15932 31585 15960
rect 29788 15920 29794 15932
rect 31573 15929 31585 15932
rect 31619 15929 31631 15963
rect 32858 15960 32864 15972
rect 31573 15923 31631 15929
rect 31726 15932 32864 15960
rect 31726 15892 31754 15932
rect 32858 15920 32864 15932
rect 32916 15920 32922 15972
rect 34790 15960 34796 15972
rect 34703 15932 34796 15960
rect 34790 15920 34796 15932
rect 34848 15960 34854 15972
rect 35345 15963 35403 15969
rect 35345 15960 35357 15963
rect 34848 15932 35357 15960
rect 34848 15920 34854 15932
rect 35345 15929 35357 15932
rect 35391 15960 35403 15963
rect 41874 15960 41880 15972
rect 35391 15932 41880 15960
rect 35391 15929 35403 15932
rect 35345 15923 35403 15929
rect 41874 15920 41880 15932
rect 41932 15920 41938 15972
rect 29656 15864 31754 15892
rect 32677 15895 32735 15901
rect 32677 15861 32689 15895
rect 32723 15892 32735 15895
rect 32766 15892 32772 15904
rect 32723 15864 32772 15892
rect 32723 15861 32735 15864
rect 32677 15855 32735 15861
rect 32766 15852 32772 15864
rect 32824 15852 32830 15904
rect 33689 15895 33747 15901
rect 33689 15861 33701 15895
rect 33735 15892 33747 15895
rect 34054 15892 34060 15904
rect 33735 15864 34060 15892
rect 33735 15861 33747 15864
rect 33689 15855 33747 15861
rect 34054 15852 34060 15864
rect 34112 15852 34118 15904
rect 34241 15895 34299 15901
rect 34241 15861 34253 15895
rect 34287 15892 34299 15895
rect 34514 15892 34520 15904
rect 34287 15864 34520 15892
rect 34287 15861 34299 15864
rect 34241 15855 34299 15861
rect 34514 15852 34520 15864
rect 34572 15852 34578 15904
rect 35802 15852 35808 15904
rect 35860 15892 35866 15904
rect 35897 15895 35955 15901
rect 35897 15892 35909 15895
rect 35860 15864 35909 15892
rect 35860 15852 35866 15864
rect 35897 15861 35909 15864
rect 35943 15861 35955 15895
rect 35897 15855 35955 15861
rect 38749 15895 38807 15901
rect 38749 15861 38761 15895
rect 38795 15892 38807 15895
rect 38838 15892 38844 15904
rect 38795 15864 38844 15892
rect 38795 15861 38807 15864
rect 38749 15855 38807 15861
rect 38838 15852 38844 15864
rect 38896 15892 38902 15904
rect 42076 15892 42104 16068
rect 42794 16056 42800 16068
rect 42852 16056 42858 16108
rect 44266 16056 44272 16108
rect 44324 16096 44330 16108
rect 45373 16099 45431 16105
rect 45373 16096 45385 16099
rect 44324 16068 45385 16096
rect 44324 16056 44330 16068
rect 45373 16065 45385 16068
rect 45419 16065 45431 16099
rect 46014 16096 46020 16108
rect 45975 16068 46020 16096
rect 45373 16059 45431 16065
rect 46014 16056 46020 16068
rect 46072 16056 46078 16108
rect 46676 16105 46704 16136
rect 46768 16136 51448 16164
rect 46661 16099 46719 16105
rect 46661 16065 46673 16099
rect 46707 16065 46719 16099
rect 46661 16059 46719 16065
rect 44358 15988 44364 16040
rect 44416 16028 44422 16040
rect 46768 16028 46796 16136
rect 51442 16124 51448 16136
rect 51500 16124 51506 16176
rect 52932 16164 52960 16204
rect 53558 16164 53564 16176
rect 52288 16136 52960 16164
rect 53519 16136 53564 16164
rect 47026 16056 47032 16108
rect 47084 16096 47090 16108
rect 49050 16096 49056 16108
rect 47084 16068 49056 16096
rect 47084 16056 47090 16068
rect 49050 16056 49056 16068
rect 49108 16056 49114 16108
rect 50338 16096 50344 16108
rect 50299 16068 50344 16096
rect 50338 16056 50344 16068
rect 50396 16056 50402 16108
rect 50430 16056 50436 16108
rect 50488 16096 50494 16108
rect 52288 16096 52316 16136
rect 53558 16124 53564 16136
rect 53616 16124 53622 16176
rect 55585 16167 55643 16173
rect 55585 16133 55597 16167
rect 55631 16164 55643 16167
rect 55858 16164 55864 16176
rect 55631 16136 55864 16164
rect 55631 16133 55643 16136
rect 55585 16127 55643 16133
rect 55858 16124 55864 16136
rect 55916 16164 55922 16176
rect 59170 16164 59176 16176
rect 55916 16136 59176 16164
rect 55916 16124 55922 16136
rect 59170 16124 59176 16136
rect 59228 16124 59234 16176
rect 59354 16124 59360 16176
rect 59412 16164 59418 16176
rect 59725 16167 59783 16173
rect 59725 16164 59737 16167
rect 59412 16136 59737 16164
rect 59412 16124 59418 16136
rect 59725 16133 59737 16136
rect 59771 16133 59783 16167
rect 59725 16127 59783 16133
rect 59998 16124 60004 16176
rect 60056 16164 60062 16176
rect 61856 16164 61884 16204
rect 61930 16192 61936 16244
rect 61988 16232 61994 16244
rect 71958 16232 71964 16244
rect 61988 16204 71964 16232
rect 61988 16192 61994 16204
rect 71958 16192 71964 16204
rect 72016 16232 72022 16244
rect 72142 16232 72148 16244
rect 72016 16204 72148 16232
rect 72016 16192 72022 16204
rect 72142 16192 72148 16204
rect 72200 16232 72206 16244
rect 72513 16235 72571 16241
rect 72513 16232 72525 16235
rect 72200 16204 72525 16232
rect 72200 16192 72206 16204
rect 72513 16201 72525 16204
rect 72559 16201 72571 16235
rect 72513 16195 72571 16201
rect 77846 16192 77852 16244
rect 77904 16232 77910 16244
rect 92566 16232 92572 16244
rect 77904 16204 92572 16232
rect 77904 16192 77910 16204
rect 92566 16192 92572 16204
rect 92624 16192 92630 16244
rect 64966 16164 64972 16176
rect 60056 16136 60306 16164
rect 61856 16136 64972 16164
rect 60056 16124 60062 16136
rect 64966 16124 64972 16136
rect 65024 16124 65030 16176
rect 65518 16164 65524 16176
rect 65479 16136 65524 16164
rect 65518 16124 65524 16136
rect 65576 16164 65582 16176
rect 66070 16164 66076 16176
rect 65576 16136 66076 16164
rect 65576 16124 65582 16136
rect 66070 16124 66076 16136
rect 66128 16124 66134 16176
rect 72050 16164 72056 16176
rect 66180 16136 66668 16164
rect 66180 16108 66208 16136
rect 50488 16068 52316 16096
rect 50488 16056 50494 16068
rect 52362 16056 52368 16108
rect 52420 16096 52426 16108
rect 53101 16099 53159 16105
rect 52420 16068 52465 16096
rect 52420 16056 52426 16068
rect 53101 16065 53113 16099
rect 53147 16096 53159 16099
rect 53650 16096 53656 16108
rect 53147 16068 53656 16096
rect 53147 16065 53159 16068
rect 53101 16059 53159 16065
rect 53650 16056 53656 16068
rect 53708 16056 53714 16108
rect 54202 16096 54208 16108
rect 54115 16068 54208 16096
rect 54202 16056 54208 16068
rect 54260 16096 54266 16108
rect 56410 16096 56416 16108
rect 54260 16068 55996 16096
rect 56371 16068 56416 16096
rect 54260 16056 54266 16068
rect 44416 16000 46796 16028
rect 44416 15988 44422 16000
rect 48682 15988 48688 16040
rect 48740 16028 48746 16040
rect 49329 16031 49387 16037
rect 49329 16028 49341 16031
rect 48740 16000 49341 16028
rect 48740 15988 48746 16000
rect 49329 15997 49341 16000
rect 49375 15997 49387 16031
rect 50522 16028 50528 16040
rect 50483 16000 50528 16028
rect 49329 15991 49387 15997
rect 50522 15988 50528 16000
rect 50580 15988 50586 16040
rect 55968 16028 55996 16068
rect 56410 16056 56416 16068
rect 56468 16056 56474 16108
rect 56686 16056 56692 16108
rect 56744 16096 56750 16108
rect 60090 16096 60096 16108
rect 56744 16068 60096 16096
rect 56744 16056 56750 16068
rect 60090 16056 60096 16068
rect 60148 16056 60154 16108
rect 63586 16056 63592 16108
rect 63644 16096 63650 16108
rect 64325 16099 64383 16105
rect 64325 16096 64337 16099
rect 63644 16068 64337 16096
rect 63644 16056 63650 16068
rect 64325 16065 64337 16068
rect 64371 16065 64383 16099
rect 64325 16059 64383 16065
rect 65061 16099 65119 16105
rect 65061 16065 65073 16099
rect 65107 16096 65119 16099
rect 66162 16096 66168 16108
rect 65107 16068 66168 16096
rect 65107 16065 65119 16068
rect 65061 16059 65119 16065
rect 66162 16056 66168 16068
rect 66220 16056 66226 16108
rect 66640 16096 66668 16136
rect 70366 16136 72056 16164
rect 67361 16099 67419 16105
rect 67361 16096 67373 16099
rect 66640 16068 67373 16096
rect 67361 16065 67373 16068
rect 67407 16065 67419 16099
rect 67361 16059 67419 16065
rect 56318 16028 56324 16040
rect 50632 16000 55904 16028
rect 55968 16000 56324 16028
rect 46014 15960 46020 15972
rect 43824 15932 46020 15960
rect 43824 15904 43852 15932
rect 46014 15920 46020 15932
rect 46072 15920 46078 15972
rect 46198 15920 46204 15972
rect 46256 15960 46262 15972
rect 50632 15960 50660 16000
rect 55306 15960 55312 15972
rect 46256 15932 50660 15960
rect 51046 15932 55312 15960
rect 46256 15920 46262 15932
rect 38896 15864 42104 15892
rect 42797 15895 42855 15901
rect 38896 15852 38902 15864
rect 42797 15861 42809 15895
rect 42843 15892 42855 15895
rect 42886 15892 42892 15904
rect 42843 15864 42892 15892
rect 42843 15861 42855 15864
rect 42797 15855 42855 15861
rect 42886 15852 42892 15864
rect 42944 15852 42950 15904
rect 43441 15895 43499 15901
rect 43441 15861 43453 15895
rect 43487 15892 43499 15895
rect 43806 15892 43812 15904
rect 43487 15864 43812 15892
rect 43487 15861 43499 15864
rect 43441 15855 43499 15861
rect 43806 15852 43812 15864
rect 43864 15852 43870 15904
rect 44266 15892 44272 15904
rect 44227 15864 44272 15892
rect 44266 15852 44272 15864
rect 44324 15852 44330 15904
rect 45462 15892 45468 15904
rect 45423 15864 45468 15892
rect 45462 15852 45468 15864
rect 45520 15852 45526 15904
rect 46109 15895 46167 15901
rect 46109 15861 46121 15895
rect 46155 15892 46167 15895
rect 47026 15892 47032 15904
rect 46155 15864 47032 15892
rect 46155 15861 46167 15864
rect 46109 15855 46167 15861
rect 47026 15852 47032 15864
rect 47084 15852 47090 15904
rect 47118 15852 47124 15904
rect 47176 15892 47182 15904
rect 47765 15895 47823 15901
rect 47765 15892 47777 15895
rect 47176 15864 47777 15892
rect 47176 15852 47182 15864
rect 47765 15861 47777 15864
rect 47811 15861 47823 15895
rect 48774 15892 48780 15904
rect 48735 15864 48780 15892
rect 47765 15855 47823 15861
rect 48774 15852 48780 15864
rect 48832 15852 48838 15904
rect 48866 15852 48872 15904
rect 48924 15892 48930 15904
rect 51046 15892 51074 15932
rect 55306 15920 55312 15932
rect 55364 15920 55370 15972
rect 55876 15960 55904 16000
rect 56318 15988 56324 16000
rect 56376 15988 56382 16040
rect 60734 16028 60740 16040
rect 59832 16000 60740 16028
rect 59832 15960 59860 16000
rect 60734 15988 60740 16000
rect 60792 16028 60798 16040
rect 61473 16031 61531 16037
rect 61473 16028 61485 16031
rect 60792 16000 61485 16028
rect 60792 15988 60798 16000
rect 61473 15997 61485 16000
rect 61519 15997 61531 16031
rect 61473 15991 61531 15997
rect 61749 16031 61807 16037
rect 61749 15997 61761 16031
rect 61795 16028 61807 16031
rect 61838 16028 61844 16040
rect 61795 16000 61844 16028
rect 61795 15997 61807 16000
rect 61749 15991 61807 15997
rect 61838 15988 61844 16000
rect 61896 16028 61902 16040
rect 63773 16031 63831 16037
rect 63773 16028 63785 16031
rect 61896 16000 63785 16028
rect 61896 15988 61902 16000
rect 63773 15997 63785 16000
rect 63819 16028 63831 16031
rect 66346 16028 66352 16040
rect 63819 16000 66352 16028
rect 63819 15997 63831 16000
rect 63773 15991 63831 15997
rect 66346 15988 66352 16000
rect 66404 15988 66410 16040
rect 66441 16031 66499 16037
rect 66441 15997 66453 16031
rect 66487 15997 66499 16031
rect 66441 15991 66499 15997
rect 55876 15932 59860 15960
rect 64598 15920 64604 15972
rect 64656 15960 64662 15972
rect 65797 15963 65855 15969
rect 65797 15960 65809 15963
rect 64656 15932 65809 15960
rect 64656 15920 64662 15932
rect 65797 15929 65809 15932
rect 65843 15960 65855 15963
rect 66456 15960 66484 15991
rect 66530 15988 66536 16040
rect 66588 16028 66594 16040
rect 70366 16028 70394 16136
rect 72050 16124 72056 16136
rect 72108 16124 72114 16176
rect 71130 16096 71136 16108
rect 71091 16068 71136 16096
rect 71130 16056 71136 16068
rect 71188 16056 71194 16108
rect 78858 16096 78864 16108
rect 78819 16068 78864 16096
rect 78858 16056 78864 16068
rect 78916 16056 78922 16108
rect 66588 16000 70394 16028
rect 76561 16031 76619 16037
rect 66588 15988 66594 16000
rect 76561 15997 76573 16031
rect 76607 16028 76619 16031
rect 77202 16028 77208 16040
rect 76607 16000 77208 16028
rect 76607 15997 76619 16000
rect 76561 15991 76619 15997
rect 77202 15988 77208 16000
rect 77260 15988 77266 16040
rect 65843 15932 66484 15960
rect 66717 15963 66775 15969
rect 65843 15929 65855 15932
rect 65797 15923 65855 15929
rect 66717 15929 66729 15963
rect 66763 15929 66775 15963
rect 70397 15963 70455 15969
rect 70397 15960 70409 15963
rect 66717 15923 66775 15929
rect 69032 15932 70409 15960
rect 53006 15892 53012 15904
rect 48924 15864 51074 15892
rect 52967 15864 53012 15892
rect 48924 15852 48930 15864
rect 53006 15852 53012 15864
rect 53064 15852 53070 15904
rect 55033 15895 55091 15901
rect 55033 15861 55045 15895
rect 55079 15892 55091 15895
rect 55950 15892 55956 15904
rect 55079 15864 55956 15892
rect 55079 15861 55091 15864
rect 55033 15855 55091 15861
rect 55950 15852 55956 15864
rect 56008 15852 56014 15904
rect 56505 15895 56563 15901
rect 56505 15861 56517 15895
rect 56551 15892 56563 15895
rect 56594 15892 56600 15904
rect 56551 15864 56600 15892
rect 56551 15861 56563 15864
rect 56505 15855 56563 15861
rect 56594 15852 56600 15864
rect 56652 15852 56658 15904
rect 57149 15895 57207 15901
rect 57149 15861 57161 15895
rect 57195 15892 57207 15895
rect 57882 15892 57888 15904
rect 57195 15864 57888 15892
rect 57195 15861 57207 15864
rect 57149 15855 57207 15861
rect 57882 15852 57888 15864
rect 57940 15892 57946 15904
rect 58069 15895 58127 15901
rect 58069 15892 58081 15895
rect 57940 15864 58081 15892
rect 57940 15852 57946 15864
rect 58069 15861 58081 15864
rect 58115 15861 58127 15895
rect 58618 15892 58624 15904
rect 58579 15864 58624 15892
rect 58069 15855 58127 15861
rect 58618 15852 58624 15864
rect 58676 15852 58682 15904
rect 58710 15852 58716 15904
rect 58768 15892 58774 15904
rect 59173 15895 59231 15901
rect 59173 15892 59185 15895
rect 58768 15864 59185 15892
rect 58768 15852 58774 15864
rect 59173 15861 59185 15864
rect 59219 15861 59231 15895
rect 62206 15892 62212 15904
rect 62167 15864 62212 15892
rect 59173 15855 59231 15861
rect 62206 15852 62212 15864
rect 62264 15852 62270 15904
rect 62942 15852 62948 15904
rect 63000 15892 63006 15904
rect 63221 15895 63279 15901
rect 63221 15892 63233 15895
rect 63000 15864 63233 15892
rect 63000 15852 63006 15864
rect 63221 15861 63233 15864
rect 63267 15861 63279 15895
rect 63221 15855 63279 15861
rect 65886 15852 65892 15904
rect 65944 15892 65950 15904
rect 65981 15895 66039 15901
rect 65981 15892 65993 15895
rect 65944 15864 65993 15892
rect 65944 15852 65950 15864
rect 65981 15861 65993 15864
rect 66027 15861 66039 15895
rect 65981 15855 66039 15861
rect 66070 15852 66076 15904
rect 66128 15892 66134 15904
rect 66732 15892 66760 15923
rect 69032 15904 69060 15932
rect 70397 15929 70409 15932
rect 70443 15929 70455 15963
rect 70397 15923 70455 15929
rect 76009 15963 76067 15969
rect 76009 15929 76021 15963
rect 76055 15960 76067 15963
rect 76742 15960 76748 15972
rect 76055 15932 76748 15960
rect 76055 15929 76067 15932
rect 76009 15923 76067 15929
rect 76742 15920 76748 15932
rect 76800 15920 76806 15972
rect 77110 15920 77116 15972
rect 77168 15960 77174 15972
rect 79321 15963 79379 15969
rect 79321 15960 79333 15963
rect 77168 15932 79333 15960
rect 77168 15920 77174 15932
rect 79321 15929 79333 15932
rect 79367 15929 79379 15963
rect 79321 15923 79379 15929
rect 79965 15963 80023 15969
rect 79965 15929 79977 15963
rect 80011 15960 80023 15963
rect 80698 15960 80704 15972
rect 80011 15932 80704 15960
rect 80011 15929 80023 15932
rect 79965 15923 80023 15929
rect 80698 15920 80704 15932
rect 80756 15920 80762 15972
rect 66128 15864 66760 15892
rect 66901 15895 66959 15901
rect 66128 15852 66134 15864
rect 66901 15861 66913 15895
rect 66947 15892 66959 15895
rect 67910 15892 67916 15904
rect 66947 15864 67916 15892
rect 66947 15861 66959 15864
rect 66901 15855 66959 15861
rect 67910 15852 67916 15864
rect 67968 15852 67974 15904
rect 68002 15852 68008 15904
rect 68060 15892 68066 15904
rect 68373 15895 68431 15901
rect 68373 15892 68385 15895
rect 68060 15864 68385 15892
rect 68060 15852 68066 15864
rect 68373 15861 68385 15864
rect 68419 15861 68431 15895
rect 69014 15892 69020 15904
rect 68975 15864 69020 15892
rect 68373 15855 68431 15861
rect 69014 15852 69020 15864
rect 69072 15852 69078 15904
rect 69661 15895 69719 15901
rect 69661 15861 69673 15895
rect 69707 15892 69719 15895
rect 69750 15892 69756 15904
rect 69707 15864 69756 15892
rect 69707 15861 69719 15864
rect 69661 15855 69719 15861
rect 69750 15852 69756 15864
rect 69808 15852 69814 15904
rect 71038 15892 71044 15904
rect 70999 15864 71044 15892
rect 71038 15852 71044 15864
rect 71096 15852 71102 15904
rect 72053 15895 72111 15901
rect 72053 15861 72065 15895
rect 72099 15892 72111 15895
rect 74258 15892 74264 15904
rect 72099 15864 74264 15892
rect 72099 15861 72111 15864
rect 72053 15855 72111 15861
rect 74258 15852 74264 15864
rect 74316 15852 74322 15904
rect 76558 15852 76564 15904
rect 76616 15892 76622 15904
rect 77021 15895 77079 15901
rect 77021 15892 77033 15895
rect 76616 15864 77033 15892
rect 76616 15852 76622 15864
rect 77021 15861 77033 15864
rect 77067 15861 77079 15895
rect 77021 15855 77079 15861
rect 77478 15852 77484 15904
rect 77536 15892 77542 15904
rect 77573 15895 77631 15901
rect 77573 15892 77585 15895
rect 77536 15864 77585 15892
rect 77536 15852 77542 15864
rect 77573 15861 77585 15864
rect 77619 15861 77631 15895
rect 78766 15892 78772 15904
rect 78727 15864 78772 15892
rect 77573 15855 77631 15861
rect 78766 15852 78772 15864
rect 78824 15852 78830 15904
rect 80517 15895 80575 15901
rect 80517 15861 80529 15895
rect 80563 15892 80575 15895
rect 80606 15892 80612 15904
rect 80563 15864 80612 15892
rect 80563 15861 80575 15864
rect 80517 15855 80575 15861
rect 80606 15852 80612 15864
rect 80664 15852 80670 15904
rect 83185 15895 83243 15901
rect 83185 15861 83197 15895
rect 83231 15892 83243 15895
rect 83458 15892 83464 15904
rect 83231 15864 83464 15892
rect 83231 15861 83243 15864
rect 83185 15855 83243 15861
rect 83458 15852 83464 15864
rect 83516 15852 83522 15904
rect 83918 15892 83924 15904
rect 83879 15864 83924 15892
rect 83918 15852 83924 15864
rect 83976 15852 83982 15904
rect 1104 15802 94852 15824
rect 1104 15750 12668 15802
rect 12720 15750 12732 15802
rect 12784 15750 12796 15802
rect 12848 15750 12860 15802
rect 12912 15750 12924 15802
rect 12976 15750 36105 15802
rect 36157 15750 36169 15802
rect 36221 15750 36233 15802
rect 36285 15750 36297 15802
rect 36349 15750 36361 15802
rect 36413 15750 59542 15802
rect 59594 15750 59606 15802
rect 59658 15750 59670 15802
rect 59722 15750 59734 15802
rect 59786 15750 59798 15802
rect 59850 15750 82979 15802
rect 83031 15750 83043 15802
rect 83095 15750 83107 15802
rect 83159 15750 83171 15802
rect 83223 15750 83235 15802
rect 83287 15750 94852 15802
rect 1104 15728 94852 15750
rect 28074 15648 28080 15700
rect 28132 15688 28138 15700
rect 30098 15688 30104 15700
rect 28132 15660 30104 15688
rect 28132 15648 28138 15660
rect 30098 15648 30104 15660
rect 30156 15648 30162 15700
rect 31386 15648 31392 15700
rect 31444 15688 31450 15700
rect 31444 15660 33456 15688
rect 31444 15648 31450 15660
rect 27798 15580 27804 15632
rect 27856 15620 27862 15632
rect 31573 15623 31631 15629
rect 31573 15620 31585 15623
rect 27856 15592 31585 15620
rect 27856 15580 27862 15592
rect 31573 15589 31585 15592
rect 31619 15589 31631 15623
rect 33428 15620 33456 15660
rect 34974 15648 34980 15700
rect 35032 15688 35038 15700
rect 38381 15691 38439 15697
rect 35032 15660 35894 15688
rect 35032 15648 35038 15660
rect 35866 15620 35894 15660
rect 38381 15657 38393 15691
rect 38427 15688 38439 15691
rect 39758 15688 39764 15700
rect 38427 15660 39764 15688
rect 38427 15657 38439 15660
rect 38381 15651 38439 15657
rect 39758 15648 39764 15660
rect 39816 15648 39822 15700
rect 43809 15691 43867 15697
rect 43809 15657 43821 15691
rect 43855 15688 43867 15691
rect 44358 15688 44364 15700
rect 43855 15660 44364 15688
rect 43855 15657 43867 15660
rect 43809 15651 43867 15657
rect 44358 15648 44364 15660
rect 44416 15648 44422 15700
rect 45462 15648 45468 15700
rect 45520 15688 45526 15700
rect 60826 15688 60832 15700
rect 45520 15660 60832 15688
rect 45520 15648 45526 15660
rect 60826 15648 60832 15660
rect 60884 15648 60890 15700
rect 65978 15648 65984 15700
rect 66036 15688 66042 15700
rect 68097 15691 68155 15697
rect 68097 15688 68109 15691
rect 66036 15660 68109 15688
rect 66036 15648 66042 15660
rect 68097 15657 68109 15660
rect 68143 15688 68155 15691
rect 73246 15688 73252 15700
rect 68143 15660 73252 15688
rect 68143 15657 68155 15660
rect 68097 15651 68155 15657
rect 73246 15648 73252 15660
rect 73304 15648 73310 15700
rect 73632 15660 79732 15688
rect 44266 15620 44272 15632
rect 33428 15592 35112 15620
rect 35866 15592 44272 15620
rect 31573 15583 31631 15589
rect 19610 15512 19616 15564
rect 19668 15552 19674 15564
rect 34977 15555 35035 15561
rect 34977 15552 34989 15555
rect 19668 15524 34989 15552
rect 19668 15512 19674 15524
rect 34977 15521 34989 15524
rect 35023 15521 35035 15555
rect 34977 15515 35035 15521
rect 35084 15552 35112 15592
rect 44266 15580 44272 15592
rect 44324 15580 44330 15632
rect 44637 15623 44695 15629
rect 44637 15589 44649 15623
rect 44683 15620 44695 15623
rect 44683 15592 46520 15620
rect 44683 15589 44695 15592
rect 44637 15583 44695 15589
rect 46492 15564 46520 15592
rect 47946 15580 47952 15632
rect 48004 15620 48010 15632
rect 50430 15620 50436 15632
rect 48004 15592 50436 15620
rect 48004 15580 48010 15592
rect 50430 15580 50436 15592
rect 50488 15580 50494 15632
rect 59357 15623 59415 15629
rect 59357 15589 59369 15623
rect 59403 15620 59415 15623
rect 60274 15620 60280 15632
rect 59403 15592 60280 15620
rect 59403 15589 59415 15592
rect 59357 15583 59415 15589
rect 60274 15580 60280 15592
rect 60332 15580 60338 15632
rect 67269 15623 67327 15629
rect 67269 15620 67281 15623
rect 64984 15592 67281 15620
rect 36817 15555 36875 15561
rect 36817 15552 36829 15555
rect 35084 15524 36829 15552
rect 19334 15444 19340 15496
rect 19392 15484 19398 15496
rect 20165 15487 20223 15493
rect 20165 15484 20177 15487
rect 19392 15456 20177 15484
rect 19392 15444 19398 15456
rect 20165 15453 20177 15456
rect 20211 15484 20223 15487
rect 20622 15484 20628 15496
rect 20211 15456 20628 15484
rect 20211 15453 20223 15456
rect 20165 15447 20223 15453
rect 20622 15444 20628 15456
rect 20680 15484 20686 15496
rect 20809 15487 20867 15493
rect 20809 15484 20821 15487
rect 20680 15456 20821 15484
rect 20680 15444 20686 15456
rect 20809 15453 20821 15456
rect 20855 15484 20867 15487
rect 22646 15484 22652 15496
rect 20855 15456 22652 15484
rect 20855 15453 20867 15456
rect 20809 15447 20867 15453
rect 22646 15444 22652 15456
rect 22704 15444 22710 15496
rect 27614 15444 27620 15496
rect 27672 15484 27678 15496
rect 28537 15487 28595 15493
rect 28537 15484 28549 15487
rect 27672 15456 28549 15484
rect 27672 15444 27678 15456
rect 28537 15453 28549 15456
rect 28583 15484 28595 15487
rect 29181 15487 29239 15493
rect 29181 15484 29193 15487
rect 28583 15456 29193 15484
rect 28583 15453 28595 15456
rect 28537 15447 28595 15453
rect 29181 15453 29193 15456
rect 29227 15484 29239 15487
rect 30466 15484 30472 15496
rect 29227 15456 30472 15484
rect 29227 15453 29239 15456
rect 29181 15447 29239 15453
rect 30466 15444 30472 15456
rect 30524 15444 30530 15496
rect 31665 15487 31723 15493
rect 31665 15453 31677 15487
rect 31711 15484 31723 15487
rect 32214 15484 32220 15496
rect 31711 15456 32220 15484
rect 31711 15453 31723 15456
rect 31665 15447 31723 15453
rect 32214 15444 32220 15456
rect 32272 15444 32278 15496
rect 32858 15444 32864 15496
rect 32916 15484 32922 15496
rect 33413 15487 33471 15493
rect 33413 15484 33425 15487
rect 32916 15456 33425 15484
rect 32916 15444 32922 15456
rect 33413 15453 33425 15456
rect 33459 15453 33471 15487
rect 33413 15447 33471 15453
rect 33873 15487 33931 15493
rect 33873 15453 33885 15487
rect 33919 15484 33931 15487
rect 34790 15484 34796 15496
rect 33919 15456 34796 15484
rect 33919 15453 33931 15456
rect 33873 15447 33931 15453
rect 34790 15444 34796 15456
rect 34848 15444 34854 15496
rect 35084 15493 35112 15524
rect 36817 15521 36829 15524
rect 36863 15552 36875 15555
rect 38746 15552 38752 15564
rect 36863 15524 38752 15552
rect 36863 15521 36875 15524
rect 36817 15515 36875 15521
rect 38746 15512 38752 15524
rect 38804 15512 38810 15564
rect 39298 15512 39304 15564
rect 39356 15552 39362 15564
rect 46198 15552 46204 15564
rect 39356 15524 46204 15552
rect 39356 15512 39362 15524
rect 46198 15512 46204 15524
rect 46256 15512 46262 15564
rect 46474 15512 46480 15564
rect 46532 15552 46538 15564
rect 48961 15555 49019 15561
rect 46532 15524 48084 15552
rect 46532 15512 46538 15524
rect 35069 15487 35127 15493
rect 35069 15453 35081 15487
rect 35115 15453 35127 15487
rect 35069 15447 35127 15453
rect 37090 15444 37096 15496
rect 37148 15484 37154 15496
rect 38289 15487 38347 15493
rect 38289 15484 38301 15487
rect 37148 15456 38301 15484
rect 37148 15444 37154 15456
rect 38289 15453 38301 15456
rect 38335 15453 38347 15487
rect 40310 15484 40316 15496
rect 40271 15456 40316 15484
rect 38289 15447 38347 15453
rect 40310 15444 40316 15456
rect 40368 15444 40374 15496
rect 40770 15484 40776 15496
rect 40731 15456 40776 15484
rect 40770 15444 40776 15456
rect 40828 15444 40834 15496
rect 40862 15444 40868 15496
rect 40920 15484 40926 15496
rect 43714 15484 43720 15496
rect 40920 15456 43116 15484
rect 43675 15456 43720 15484
rect 40920 15444 40926 15456
rect 43088 15428 43116 15456
rect 43714 15444 43720 15456
rect 43772 15444 43778 15496
rect 45738 15484 45744 15496
rect 45699 15456 45744 15484
rect 45738 15444 45744 15456
rect 45796 15444 45802 15496
rect 46658 15484 46664 15496
rect 46619 15456 46664 15484
rect 46658 15444 46664 15456
rect 46716 15444 46722 15496
rect 48056 15470 48084 15524
rect 48961 15521 48973 15555
rect 49007 15552 49019 15555
rect 61102 15552 61108 15564
rect 49007 15524 60734 15552
rect 61063 15524 61108 15552
rect 49007 15521 49019 15524
rect 48961 15515 49019 15521
rect 48682 15444 48688 15496
rect 48740 15484 48746 15496
rect 48869 15487 48927 15493
rect 48869 15484 48881 15487
rect 48740 15456 48881 15484
rect 48740 15444 48746 15456
rect 48869 15453 48881 15456
rect 48915 15453 48927 15487
rect 48869 15447 48927 15453
rect 49142 15444 49148 15496
rect 49200 15484 49206 15496
rect 49510 15484 49516 15496
rect 49200 15456 49516 15484
rect 49200 15444 49206 15456
rect 49510 15444 49516 15456
rect 49568 15444 49574 15496
rect 51166 15484 51172 15496
rect 51127 15456 51172 15484
rect 51166 15444 51172 15456
rect 51224 15444 51230 15496
rect 53650 15444 53656 15496
rect 53708 15484 53714 15496
rect 53837 15487 53895 15493
rect 53837 15484 53849 15487
rect 53708 15456 53849 15484
rect 53708 15444 53714 15456
rect 53837 15453 53849 15456
rect 53883 15484 53895 15487
rect 56137 15487 56195 15493
rect 56137 15484 56149 15487
rect 53883 15456 56149 15484
rect 53883 15453 53895 15456
rect 53837 15447 53895 15453
rect 56137 15453 56149 15456
rect 56183 15484 56195 15487
rect 56410 15484 56416 15496
rect 56183 15456 56416 15484
rect 56183 15453 56195 15456
rect 56137 15447 56195 15453
rect 56410 15444 56416 15456
rect 56468 15444 56474 15496
rect 57054 15484 57060 15496
rect 57015 15456 57060 15484
rect 57054 15444 57060 15456
rect 57112 15444 57118 15496
rect 59906 15444 59912 15496
rect 59964 15484 59970 15496
rect 60093 15487 60151 15493
rect 60093 15484 60105 15487
rect 59964 15456 60105 15484
rect 59964 15444 59970 15456
rect 60093 15453 60105 15456
rect 60139 15453 60151 15487
rect 60706 15484 60734 15524
rect 61102 15512 61108 15524
rect 61160 15512 61166 15564
rect 64690 15552 64696 15564
rect 64651 15524 64696 15552
rect 64690 15512 64696 15524
rect 64748 15512 64754 15564
rect 64984 15561 65012 15592
rect 67269 15589 67281 15592
rect 67315 15589 67327 15623
rect 67269 15583 67327 15589
rect 67358 15580 67364 15632
rect 67416 15620 67422 15632
rect 69661 15623 69719 15629
rect 69661 15620 69673 15623
rect 67416 15592 69673 15620
rect 67416 15580 67422 15592
rect 69661 15589 69673 15592
rect 69707 15589 69719 15623
rect 69661 15583 69719 15589
rect 70486 15580 70492 15632
rect 70544 15620 70550 15632
rect 72418 15620 72424 15632
rect 70544 15592 72424 15620
rect 70544 15580 70550 15592
rect 72418 15580 72424 15592
rect 72476 15580 72482 15632
rect 72513 15623 72571 15629
rect 72513 15589 72525 15623
rect 72559 15589 72571 15623
rect 72513 15583 72571 15589
rect 64969 15555 65027 15561
rect 64969 15521 64981 15555
rect 65015 15521 65027 15555
rect 67634 15552 67640 15564
rect 64969 15515 65027 15521
rect 66824 15524 67640 15552
rect 61010 15484 61016 15496
rect 60706 15456 61016 15484
rect 60093 15447 60151 15453
rect 61010 15444 61016 15456
rect 61068 15444 61074 15496
rect 65797 15487 65855 15493
rect 65797 15453 65809 15487
rect 65843 15484 65855 15487
rect 65886 15484 65892 15496
rect 65843 15456 65892 15484
rect 65843 15453 65855 15456
rect 65797 15447 65855 15453
rect 65886 15444 65892 15456
rect 65944 15444 65950 15496
rect 65978 15444 65984 15496
rect 66036 15484 66042 15496
rect 66824 15493 66852 15524
rect 67634 15512 67640 15524
rect 67692 15552 67698 15564
rect 70302 15552 70308 15564
rect 67692 15524 70308 15552
rect 67692 15512 67698 15524
rect 70302 15512 70308 15524
rect 70360 15552 70366 15564
rect 71130 15552 71136 15564
rect 70360 15524 71136 15552
rect 70360 15512 70366 15524
rect 71130 15512 71136 15524
rect 71188 15552 71194 15564
rect 71188 15524 71544 15552
rect 71188 15512 71194 15524
rect 66809 15487 66867 15493
rect 66036 15456 66081 15484
rect 66036 15444 66042 15456
rect 66809 15453 66821 15487
rect 66855 15453 66867 15487
rect 66809 15447 66867 15453
rect 67453 15487 67511 15493
rect 67453 15453 67465 15487
rect 67499 15453 67511 15487
rect 67910 15484 67916 15496
rect 67871 15456 67916 15484
rect 67453 15447 67511 15453
rect 30653 15419 30711 15425
rect 30653 15416 30665 15419
rect 24872 15388 30665 15416
rect 20070 15348 20076 15360
rect 20031 15320 20076 15348
rect 20070 15308 20076 15320
rect 20128 15308 20134 15360
rect 20717 15351 20775 15357
rect 20717 15317 20729 15351
rect 20763 15348 20775 15351
rect 20806 15348 20812 15360
rect 20763 15320 20812 15348
rect 20763 15317 20775 15320
rect 20717 15311 20775 15317
rect 20806 15308 20812 15320
rect 20864 15308 20870 15360
rect 22738 15348 22744 15360
rect 22699 15320 22744 15348
rect 22738 15308 22744 15320
rect 22796 15308 22802 15360
rect 23658 15348 23664 15360
rect 23619 15320 23664 15348
rect 23658 15308 23664 15320
rect 23716 15308 23722 15360
rect 24762 15308 24768 15360
rect 24820 15348 24826 15360
rect 24872 15357 24900 15388
rect 30653 15385 30665 15388
rect 30699 15416 30711 15419
rect 32398 15416 32404 15428
rect 30699 15388 32404 15416
rect 30699 15385 30711 15388
rect 30653 15379 30711 15385
rect 32398 15376 32404 15388
rect 32456 15416 32462 15428
rect 32493 15419 32551 15425
rect 32493 15416 32505 15419
rect 32456 15388 32505 15416
rect 32456 15376 32462 15388
rect 32493 15385 32505 15388
rect 32539 15385 32551 15419
rect 32493 15379 32551 15385
rect 32582 15376 32588 15428
rect 32640 15416 32646 15428
rect 32766 15416 32772 15428
rect 32640 15388 32772 15416
rect 32640 15376 32646 15388
rect 32766 15376 32772 15388
rect 32824 15416 32830 15428
rect 41598 15416 41604 15428
rect 32824 15388 41604 15416
rect 32824 15376 32830 15388
rect 41598 15376 41604 15388
rect 41656 15376 41662 15428
rect 41874 15376 41880 15428
rect 41932 15416 41938 15428
rect 41932 15388 42472 15416
rect 41932 15376 41938 15388
rect 24857 15351 24915 15357
rect 24857 15348 24869 15351
rect 24820 15320 24869 15348
rect 24820 15308 24826 15320
rect 24857 15317 24869 15320
rect 24903 15317 24915 15351
rect 24857 15311 24915 15317
rect 28445 15351 28503 15357
rect 28445 15317 28457 15351
rect 28491 15348 28503 15351
rect 28534 15348 28540 15360
rect 28491 15320 28540 15348
rect 28491 15317 28503 15320
rect 28445 15311 28503 15317
rect 28534 15308 28540 15320
rect 28592 15308 28598 15360
rect 28902 15308 28908 15360
rect 28960 15348 28966 15360
rect 29089 15351 29147 15357
rect 29089 15348 29101 15351
rect 28960 15320 29101 15348
rect 28960 15308 28966 15320
rect 29089 15317 29101 15320
rect 29135 15317 29147 15351
rect 29089 15311 29147 15317
rect 32674 15308 32680 15360
rect 32732 15348 32738 15360
rect 33045 15351 33103 15357
rect 33045 15348 33057 15351
rect 32732 15320 33057 15348
rect 32732 15308 32738 15320
rect 33045 15317 33057 15320
rect 33091 15317 33103 15351
rect 33045 15311 33103 15317
rect 33134 15308 33140 15360
rect 33192 15348 33198 15360
rect 34514 15348 34520 15360
rect 33192 15320 34520 15348
rect 33192 15308 33198 15320
rect 34514 15308 34520 15320
rect 34572 15348 34578 15360
rect 34974 15348 34980 15360
rect 34572 15320 34980 15348
rect 34572 15308 34578 15320
rect 34974 15308 34980 15320
rect 35032 15308 35038 15360
rect 35526 15348 35532 15360
rect 35487 15320 35532 15348
rect 35526 15308 35532 15320
rect 35584 15308 35590 15360
rect 36262 15348 36268 15360
rect 36223 15320 36268 15348
rect 36262 15308 36268 15320
rect 36320 15308 36326 15360
rect 37645 15351 37703 15357
rect 37645 15317 37657 15351
rect 37691 15348 37703 15351
rect 37734 15348 37740 15360
rect 37691 15320 37740 15348
rect 37691 15317 37703 15320
rect 37645 15311 37703 15317
rect 37734 15308 37740 15320
rect 37792 15308 37798 15360
rect 38102 15308 38108 15360
rect 38160 15348 38166 15360
rect 39209 15351 39267 15357
rect 39209 15348 39221 15351
rect 38160 15320 39221 15348
rect 38160 15308 38166 15320
rect 39209 15317 39221 15320
rect 39255 15348 39267 15351
rect 40862 15348 40868 15360
rect 39255 15320 40868 15348
rect 39255 15317 39267 15320
rect 39209 15311 39267 15317
rect 40862 15308 40868 15320
rect 40920 15308 40926 15360
rect 41138 15348 41144 15360
rect 41099 15320 41144 15348
rect 41138 15308 41144 15320
rect 41196 15308 41202 15360
rect 41690 15308 41696 15360
rect 41748 15348 41754 15360
rect 41785 15351 41843 15357
rect 41785 15348 41797 15351
rect 41748 15320 41797 15348
rect 41748 15308 41754 15320
rect 41785 15317 41797 15320
rect 41831 15317 41843 15351
rect 42334 15348 42340 15360
rect 42295 15320 42340 15348
rect 41785 15311 41843 15317
rect 42334 15308 42340 15320
rect 42392 15308 42398 15360
rect 42444 15348 42472 15388
rect 43070 15376 43076 15428
rect 43128 15416 43134 15428
rect 43165 15419 43223 15425
rect 43165 15416 43177 15419
rect 43128 15388 43177 15416
rect 43128 15376 43134 15388
rect 43165 15385 43177 15388
rect 43211 15385 43223 15419
rect 46934 15416 46940 15428
rect 43165 15379 43223 15385
rect 43640 15388 45784 15416
rect 46895 15388 46940 15416
rect 43640 15348 43668 15388
rect 45646 15348 45652 15360
rect 42444 15320 43668 15348
rect 45607 15320 45652 15348
rect 45646 15308 45652 15320
rect 45704 15308 45710 15360
rect 45756 15348 45784 15388
rect 46934 15376 46940 15388
rect 46992 15376 46998 15428
rect 51442 15416 51448 15428
rect 48240 15388 51074 15416
rect 51403 15388 51448 15416
rect 48240 15348 48268 15388
rect 45756 15320 48268 15348
rect 48409 15351 48467 15357
rect 48409 15317 48421 15351
rect 48455 15348 48467 15351
rect 48498 15348 48504 15360
rect 48455 15320 48504 15348
rect 48455 15317 48467 15320
rect 48409 15311 48467 15317
rect 48498 15308 48504 15320
rect 48556 15308 48562 15360
rect 49694 15308 49700 15360
rect 49752 15348 49758 15360
rect 50522 15348 50528 15360
rect 49752 15320 50528 15348
rect 49752 15308 49758 15320
rect 50522 15308 50528 15320
rect 50580 15348 50586 15360
rect 50617 15351 50675 15357
rect 50617 15348 50629 15351
rect 50580 15320 50629 15348
rect 50580 15308 50586 15320
rect 50617 15317 50629 15320
rect 50663 15317 50675 15351
rect 51046 15348 51074 15388
rect 51442 15376 51448 15388
rect 51500 15376 51506 15428
rect 53006 15416 53012 15428
rect 52670 15388 53012 15416
rect 53006 15376 53012 15388
rect 53064 15376 53070 15428
rect 56686 15376 56692 15428
rect 56744 15416 56750 15428
rect 57333 15419 57391 15425
rect 57333 15416 57345 15419
rect 56744 15388 57345 15416
rect 56744 15376 56750 15388
rect 57333 15385 57345 15388
rect 57379 15385 57391 15419
rect 57333 15379 57391 15385
rect 57974 15376 57980 15428
rect 58032 15376 58038 15428
rect 61381 15419 61439 15425
rect 61381 15416 61393 15419
rect 58820 15388 61393 15416
rect 52917 15351 52975 15357
rect 52917 15348 52929 15351
rect 51046 15320 52929 15348
rect 50617 15311 50675 15317
rect 52917 15317 52929 15320
rect 52963 15317 52975 15351
rect 53742 15348 53748 15360
rect 53703 15320 53748 15348
rect 52917 15311 52975 15317
rect 53742 15308 53748 15320
rect 53800 15308 53806 15360
rect 54389 15351 54447 15357
rect 54389 15317 54401 15351
rect 54435 15348 54447 15351
rect 54478 15348 54484 15360
rect 54435 15320 54484 15348
rect 54435 15317 54447 15320
rect 54389 15311 54447 15317
rect 54478 15308 54484 15320
rect 54536 15308 54542 15360
rect 54846 15348 54852 15360
rect 54807 15320 54852 15348
rect 54846 15308 54852 15320
rect 54904 15308 54910 15360
rect 56042 15348 56048 15360
rect 56003 15320 56048 15348
rect 56042 15308 56048 15320
rect 56100 15308 56106 15360
rect 58820 15357 58848 15388
rect 61381 15385 61393 15388
rect 61427 15385 61439 15419
rect 61381 15379 61439 15385
rect 61930 15376 61936 15428
rect 61988 15376 61994 15428
rect 64877 15419 64935 15425
rect 62868 15388 64828 15416
rect 58805 15351 58863 15357
rect 58805 15317 58817 15351
rect 58851 15317 58863 15351
rect 58805 15311 58863 15317
rect 60001 15351 60059 15357
rect 60001 15317 60013 15351
rect 60047 15348 60059 15351
rect 60090 15348 60096 15360
rect 60047 15320 60096 15348
rect 60047 15317 60059 15320
rect 60001 15311 60059 15317
rect 60090 15308 60096 15320
rect 60148 15308 60154 15360
rect 62868 15357 62896 15388
rect 62853 15351 62911 15357
rect 62853 15317 62865 15351
rect 62899 15317 62911 15351
rect 62853 15311 62911 15317
rect 63405 15351 63463 15357
rect 63405 15317 63417 15351
rect 63451 15348 63463 15351
rect 63586 15348 63592 15360
rect 63451 15320 63592 15348
rect 63451 15317 63463 15320
rect 63405 15311 63463 15317
rect 63586 15308 63592 15320
rect 63644 15308 63650 15360
rect 64800 15348 64828 15388
rect 64877 15385 64889 15419
rect 64923 15416 64935 15419
rect 64966 15416 64972 15428
rect 64923 15388 64972 15416
rect 64923 15385 64935 15388
rect 64877 15379 64935 15385
rect 64966 15376 64972 15388
rect 65024 15376 65030 15428
rect 66165 15419 66223 15425
rect 66165 15385 66177 15419
rect 66211 15416 66223 15419
rect 67468 15416 67496 15447
rect 67910 15444 67916 15456
rect 67968 15444 67974 15496
rect 69201 15487 69259 15493
rect 69201 15453 69213 15487
rect 69247 15484 69259 15487
rect 70854 15484 70860 15496
rect 69247 15456 70860 15484
rect 69247 15453 69259 15456
rect 69201 15447 69259 15453
rect 70854 15444 70860 15456
rect 70912 15444 70918 15496
rect 71516 15493 71544 15524
rect 72050 15512 72056 15564
rect 72108 15552 72114 15564
rect 72528 15552 72556 15583
rect 72602 15580 72608 15632
rect 72660 15620 72666 15632
rect 73157 15623 73215 15629
rect 73157 15620 73169 15623
rect 72660 15592 73169 15620
rect 72660 15580 72666 15592
rect 73157 15589 73169 15592
rect 73203 15620 73215 15623
rect 73632 15620 73660 15660
rect 73203 15592 73660 15620
rect 73709 15623 73767 15629
rect 73203 15589 73215 15592
rect 73157 15583 73215 15589
rect 73709 15589 73721 15623
rect 73755 15620 73767 15623
rect 74626 15620 74632 15632
rect 73755 15592 74632 15620
rect 73755 15589 73767 15592
rect 73709 15583 73767 15589
rect 74626 15580 74632 15592
rect 74684 15580 74690 15632
rect 79704 15561 79732 15660
rect 78861 15555 78919 15561
rect 78861 15552 78873 15555
rect 72108 15524 72556 15552
rect 72620 15524 78873 15552
rect 72108 15512 72114 15524
rect 71501 15487 71559 15493
rect 71501 15453 71513 15487
rect 71547 15453 71559 15487
rect 71501 15447 71559 15453
rect 72142 15444 72148 15496
rect 72200 15484 72206 15496
rect 72200 15456 72245 15484
rect 72620 15478 72648 15524
rect 78861 15521 78873 15524
rect 78907 15521 78919 15555
rect 78861 15515 78919 15521
rect 79689 15555 79747 15561
rect 79689 15521 79701 15555
rect 79735 15552 79747 15555
rect 80238 15552 80244 15564
rect 79735 15524 80244 15552
rect 79735 15521 79747 15524
rect 79689 15515 79747 15521
rect 80238 15512 80244 15524
rect 80296 15512 80302 15564
rect 74166 15484 74172 15496
rect 72200 15444 72206 15456
rect 72436 15450 72648 15478
rect 74127 15456 74172 15484
rect 66211 15388 67496 15416
rect 66211 15385 66223 15388
rect 66165 15379 66223 15385
rect 67818 15376 67824 15428
rect 67876 15416 67882 15428
rect 72436 15416 72464 15450
rect 74166 15444 74172 15456
rect 74224 15444 74230 15496
rect 75457 15487 75515 15493
rect 75457 15453 75469 15487
rect 75503 15484 75515 15487
rect 76285 15487 76343 15493
rect 76285 15484 76297 15487
rect 75503 15456 76297 15484
rect 75503 15453 75515 15456
rect 75457 15447 75515 15453
rect 76285 15453 76297 15456
rect 76331 15453 76343 15487
rect 76285 15447 76343 15453
rect 79137 15487 79195 15493
rect 79137 15453 79149 15487
rect 79183 15484 79195 15487
rect 81250 15484 81256 15496
rect 79183 15456 81256 15484
rect 79183 15453 79195 15456
rect 79137 15447 79195 15453
rect 81250 15444 81256 15456
rect 81308 15444 81314 15496
rect 82814 15444 82820 15496
rect 82872 15484 82878 15496
rect 82909 15487 82967 15493
rect 82909 15484 82921 15487
rect 82872 15456 82921 15484
rect 82872 15444 82878 15456
rect 82909 15453 82921 15456
rect 82955 15484 82967 15487
rect 82955 15456 84148 15484
rect 82955 15453 82967 15456
rect 82909 15447 82967 15453
rect 75089 15419 75147 15425
rect 75089 15416 75101 15419
rect 67876 15388 72464 15416
rect 72620 15388 75101 15416
rect 67876 15376 67882 15388
rect 66530 15348 66536 15360
rect 64800 15320 66536 15348
rect 66530 15308 66536 15320
rect 66588 15308 66594 15360
rect 66714 15348 66720 15360
rect 66675 15320 66720 15348
rect 66714 15308 66720 15320
rect 66772 15308 66778 15360
rect 68649 15351 68707 15357
rect 68649 15317 68661 15351
rect 68695 15348 68707 15351
rect 68738 15348 68744 15360
rect 68695 15320 68744 15348
rect 68695 15317 68707 15320
rect 68649 15311 68707 15317
rect 68738 15308 68744 15320
rect 68796 15308 68802 15360
rect 69842 15308 69848 15360
rect 69900 15348 69906 15360
rect 70213 15351 70271 15357
rect 70213 15348 70225 15351
rect 69900 15320 70225 15348
rect 69900 15308 69906 15320
rect 70213 15317 70225 15320
rect 70259 15317 70271 15351
rect 70213 15311 70271 15317
rect 70854 15308 70860 15360
rect 70912 15348 70918 15360
rect 70949 15351 71007 15357
rect 70949 15348 70961 15351
rect 70912 15320 70961 15348
rect 70912 15308 70918 15320
rect 70949 15317 70961 15320
rect 70995 15317 71007 15351
rect 71590 15348 71596 15360
rect 71551 15320 71596 15348
rect 70949 15311 71007 15317
rect 71590 15308 71596 15320
rect 71648 15308 71654 15360
rect 72620 15357 72648 15388
rect 75089 15385 75101 15388
rect 75135 15385 75147 15419
rect 75089 15379 75147 15385
rect 75273 15419 75331 15425
rect 75273 15385 75285 15419
rect 75319 15416 75331 15419
rect 78766 15416 78772 15428
rect 75319 15388 77524 15416
rect 78430 15388 78772 15416
rect 75319 15385 75331 15388
rect 75273 15379 75331 15385
rect 72605 15351 72663 15357
rect 72605 15317 72617 15351
rect 72651 15317 72663 15351
rect 72605 15311 72663 15317
rect 74353 15351 74411 15357
rect 74353 15317 74365 15351
rect 74399 15348 74411 15351
rect 75288 15348 75316 15379
rect 76466 15348 76472 15360
rect 74399 15320 75316 15348
rect 76427 15320 76472 15348
rect 74399 15317 74411 15320
rect 74353 15311 74411 15317
rect 76466 15308 76472 15320
rect 76524 15308 76530 15360
rect 77386 15348 77392 15360
rect 77347 15320 77392 15348
rect 77386 15308 77392 15320
rect 77444 15308 77450 15360
rect 77496 15348 77524 15388
rect 78766 15376 78772 15388
rect 78824 15376 78830 15428
rect 82998 15416 83004 15428
rect 78876 15388 83004 15416
rect 78876 15348 78904 15388
rect 82998 15376 83004 15388
rect 83056 15376 83062 15428
rect 84120 15360 84148 15456
rect 80146 15348 80152 15360
rect 77496 15320 78904 15348
rect 80107 15320 80152 15348
rect 80146 15308 80152 15320
rect 80204 15308 80210 15360
rect 81345 15351 81403 15357
rect 81345 15317 81357 15351
rect 81391 15348 81403 15351
rect 81618 15348 81624 15360
rect 81391 15320 81624 15348
rect 81391 15317 81403 15320
rect 81345 15311 81403 15317
rect 81618 15308 81624 15320
rect 81676 15308 81682 15360
rect 83734 15348 83740 15360
rect 83695 15320 83740 15348
rect 83734 15308 83740 15320
rect 83792 15308 83798 15360
rect 84102 15308 84108 15360
rect 84160 15348 84166 15360
rect 84381 15351 84439 15357
rect 84381 15348 84393 15351
rect 84160 15320 84393 15348
rect 84160 15308 84166 15320
rect 84381 15317 84393 15320
rect 84427 15317 84439 15351
rect 84381 15311 84439 15317
rect 86497 15351 86555 15357
rect 86497 15317 86509 15351
rect 86543 15348 86555 15351
rect 86770 15348 86776 15360
rect 86543 15320 86776 15348
rect 86543 15317 86555 15320
rect 86497 15311 86555 15317
rect 86770 15308 86776 15320
rect 86828 15308 86834 15360
rect 88061 15351 88119 15357
rect 88061 15317 88073 15351
rect 88107 15348 88119 15351
rect 88242 15348 88248 15360
rect 88107 15320 88248 15348
rect 88107 15317 88119 15320
rect 88061 15311 88119 15317
rect 88242 15308 88248 15320
rect 88300 15308 88306 15360
rect 88889 15351 88947 15357
rect 88889 15317 88901 15351
rect 88935 15348 88947 15351
rect 88978 15348 88984 15360
rect 88935 15320 88984 15348
rect 88935 15317 88947 15320
rect 88889 15311 88947 15317
rect 88978 15308 88984 15320
rect 89036 15308 89042 15360
rect 1104 15258 95011 15280
rect 1104 15206 24386 15258
rect 24438 15206 24450 15258
rect 24502 15206 24514 15258
rect 24566 15206 24578 15258
rect 24630 15206 24642 15258
rect 24694 15206 47823 15258
rect 47875 15206 47887 15258
rect 47939 15206 47951 15258
rect 48003 15206 48015 15258
rect 48067 15206 48079 15258
rect 48131 15206 71260 15258
rect 71312 15206 71324 15258
rect 71376 15206 71388 15258
rect 71440 15206 71452 15258
rect 71504 15206 71516 15258
rect 71568 15206 94697 15258
rect 94749 15206 94761 15258
rect 94813 15206 94825 15258
rect 94877 15206 94889 15258
rect 94941 15206 94953 15258
rect 95005 15206 95011 15258
rect 1104 15184 95011 15206
rect 16298 15104 16304 15156
rect 16356 15144 16362 15156
rect 22554 15144 22560 15156
rect 16356 15116 22560 15144
rect 16356 15104 16362 15116
rect 22554 15104 22560 15116
rect 22612 15104 22618 15156
rect 28074 15144 28080 15156
rect 22756 15116 28080 15144
rect 19337 15079 19395 15085
rect 19337 15045 19349 15079
rect 19383 15076 19395 15079
rect 19610 15076 19616 15088
rect 19383 15048 19616 15076
rect 19383 15045 19395 15048
rect 19337 15039 19395 15045
rect 19610 15036 19616 15048
rect 19668 15036 19674 15088
rect 20714 15076 20720 15088
rect 20562 15048 20720 15076
rect 20714 15036 20720 15048
rect 20772 15036 20778 15088
rect 21085 15079 21143 15085
rect 21085 15045 21097 15079
rect 21131 15076 21143 15079
rect 22756 15076 22784 15116
rect 28074 15104 28080 15116
rect 28132 15104 28138 15156
rect 28169 15147 28227 15153
rect 28169 15113 28181 15147
rect 28215 15144 28227 15147
rect 28215 15116 32076 15144
rect 28215 15113 28227 15116
rect 28169 15107 28227 15113
rect 24762 15076 24768 15088
rect 21131 15048 22784 15076
rect 22848 15048 24768 15076
rect 21131 15045 21143 15048
rect 21085 15039 21143 15045
rect 22848 15017 22876 15048
rect 24762 15036 24768 15048
rect 24820 15036 24826 15088
rect 24854 15036 24860 15088
rect 24912 15076 24918 15088
rect 27798 15076 27804 15088
rect 24912 15048 27804 15076
rect 24912 15036 24918 15048
rect 27798 15036 27804 15048
rect 27856 15036 27862 15088
rect 28902 15036 28908 15088
rect 28960 15036 28966 15088
rect 29641 15079 29699 15085
rect 29641 15045 29653 15079
rect 29687 15076 29699 15079
rect 32048 15076 32076 15116
rect 33318 15104 33324 15156
rect 33376 15144 33382 15156
rect 36817 15147 36875 15153
rect 36817 15144 36829 15147
rect 33376 15116 36829 15144
rect 33376 15104 33382 15116
rect 36817 15113 36829 15116
rect 36863 15113 36875 15147
rect 36817 15107 36875 15113
rect 38746 15104 38752 15156
rect 38804 15144 38810 15156
rect 53009 15147 53067 15153
rect 53009 15144 53021 15147
rect 38804 15116 53021 15144
rect 38804 15104 38810 15116
rect 53009 15113 53021 15116
rect 53055 15113 53067 15147
rect 53009 15107 53067 15113
rect 53208 15116 59216 15144
rect 35986 15076 35992 15088
rect 29687 15048 31156 15076
rect 32048 15048 35992 15076
rect 29687 15045 29699 15048
rect 29641 15039 29699 15045
rect 22189 15011 22247 15017
rect 22189 14977 22201 15011
rect 22235 15008 22247 15011
rect 22833 15011 22891 15017
rect 22833 15008 22845 15011
rect 22235 14980 22845 15008
rect 22235 14977 22247 14980
rect 22189 14971 22247 14977
rect 22833 14977 22845 14980
rect 22879 14977 22891 15011
rect 22833 14971 22891 14977
rect 23477 15011 23535 15017
rect 23477 14977 23489 15011
rect 23523 14977 23535 15011
rect 23477 14971 23535 14977
rect 24305 15011 24363 15017
rect 24305 14977 24317 15011
rect 24351 15008 24363 15011
rect 24578 15008 24584 15020
rect 24351 14980 24584 15008
rect 24351 14977 24363 14980
rect 24305 14971 24363 14977
rect 15746 14900 15752 14952
rect 15804 14940 15810 14952
rect 19061 14943 19119 14949
rect 19061 14940 19073 14943
rect 15804 14912 19073 14940
rect 15804 14900 15810 14912
rect 19061 14909 19073 14912
rect 19107 14909 19119 14943
rect 23492 14940 23520 14971
rect 24578 14968 24584 14980
rect 24636 14968 24642 15020
rect 24688 14980 26280 15008
rect 23658 14940 23664 14952
rect 23492 14912 23664 14940
rect 19061 14903 19119 14909
rect 23658 14900 23664 14912
rect 23716 14940 23722 14952
rect 24688 14940 24716 14980
rect 25866 14940 25872 14952
rect 23716 14912 24716 14940
rect 25827 14912 25872 14940
rect 23716 14900 23722 14912
rect 25866 14900 25872 14912
rect 25924 14900 25930 14952
rect 26252 14940 26280 14980
rect 30098 14968 30104 15020
rect 30156 15008 30162 15020
rect 31021 15011 31079 15017
rect 30156 14980 30880 15008
rect 30156 14968 30162 14980
rect 29638 14940 29644 14952
rect 26252 14912 29644 14940
rect 29638 14900 29644 14912
rect 29696 14900 29702 14952
rect 29914 14940 29920 14952
rect 29875 14912 29920 14940
rect 29914 14900 29920 14912
rect 29972 14900 29978 14952
rect 30469 14943 30527 14949
rect 30469 14909 30481 14943
rect 30515 14940 30527 14943
rect 30742 14940 30748 14952
rect 30515 14912 30748 14940
rect 30515 14909 30527 14912
rect 30469 14903 30527 14909
rect 30742 14900 30748 14912
rect 30800 14900 30806 14952
rect 30852 14940 30880 14980
rect 31021 14977 31033 15011
rect 31067 14977 31079 15011
rect 31021 14971 31079 14977
rect 31036 14940 31064 14971
rect 30852 14912 31064 14940
rect 31128 14940 31156 15048
rect 35986 15036 35992 15048
rect 36044 15036 36050 15088
rect 36262 15076 36268 15088
rect 36096 15048 36268 15076
rect 31386 15008 31392 15020
rect 31347 14980 31392 15008
rect 31386 14968 31392 14980
rect 31444 14968 31450 15020
rect 31478 14968 31484 15020
rect 31536 15008 31542 15020
rect 32861 15011 32919 15017
rect 32861 15008 32873 15011
rect 31536 14980 32873 15008
rect 31536 14968 31542 14980
rect 32861 14977 32873 14980
rect 32907 14977 32919 15011
rect 32861 14971 32919 14977
rect 32950 14968 32956 15020
rect 33008 15008 33014 15020
rect 33137 15011 33195 15017
rect 33137 15008 33149 15011
rect 33008 14980 33149 15008
rect 33008 14968 33014 14980
rect 33137 14977 33149 14980
rect 33183 14977 33195 15011
rect 33137 14971 33195 14977
rect 33873 15011 33931 15017
rect 33873 14977 33885 15011
rect 33919 15008 33931 15011
rect 34790 15008 34796 15020
rect 33919 14980 34796 15008
rect 33919 14977 33931 14980
rect 33873 14971 33931 14977
rect 34790 14968 34796 14980
rect 34848 14968 34854 15020
rect 34974 15008 34980 15020
rect 34935 14980 34980 15008
rect 34974 14968 34980 14980
rect 35032 14968 35038 15020
rect 36096 15017 36124 15048
rect 36262 15036 36268 15048
rect 36320 15076 36326 15088
rect 36320 15048 45968 15076
rect 36320 15036 36326 15048
rect 36081 15011 36139 15017
rect 36081 14977 36093 15011
rect 36127 14977 36139 15011
rect 36081 14971 36139 14977
rect 36909 15011 36967 15017
rect 36909 14977 36921 15011
rect 36955 15008 36967 15011
rect 37274 15008 37280 15020
rect 36955 14980 37280 15008
rect 36955 14977 36967 14980
rect 36909 14971 36967 14977
rect 37274 14968 37280 14980
rect 37332 14968 37338 15020
rect 38105 15011 38163 15017
rect 38105 15008 38117 15011
rect 37384 14980 38117 15008
rect 32766 14940 32772 14952
rect 31128 14912 32772 14940
rect 32766 14900 32772 14912
rect 32824 14900 32830 14952
rect 33226 14900 33232 14952
rect 33284 14940 33290 14952
rect 34333 14943 34391 14949
rect 34333 14940 34345 14943
rect 33284 14912 34345 14940
rect 33284 14900 33290 14912
rect 34333 14909 34345 14912
rect 34379 14909 34391 14943
rect 34333 14903 34391 14909
rect 34698 14900 34704 14952
rect 34756 14940 34762 14952
rect 34885 14943 34943 14949
rect 34885 14940 34897 14943
rect 34756 14912 34897 14940
rect 34756 14900 34762 14912
rect 34885 14909 34897 14912
rect 34931 14909 34943 14943
rect 34885 14903 34943 14909
rect 35066 14900 35072 14952
rect 35124 14940 35130 14952
rect 37384 14940 37412 14980
rect 38105 14977 38117 14980
rect 38151 14977 38163 15011
rect 38105 14971 38163 14977
rect 38473 15011 38531 15017
rect 38473 14977 38485 15011
rect 38519 15008 38531 15011
rect 38654 15008 38660 15020
rect 38519 14980 38660 15008
rect 38519 14977 38531 14980
rect 38473 14971 38531 14977
rect 35124 14912 37412 14940
rect 37461 14943 37519 14949
rect 35124 14900 35130 14912
rect 37461 14909 37473 14943
rect 37507 14909 37519 14943
rect 38120 14940 38148 14971
rect 38654 14968 38660 14980
rect 38712 14968 38718 15020
rect 39209 15011 39267 15017
rect 39209 14977 39221 15011
rect 39255 14977 39267 15011
rect 39209 14971 39267 14977
rect 39224 14940 39252 14971
rect 39298 14968 39304 15020
rect 39356 15008 39362 15020
rect 40310 15008 40316 15020
rect 39356 14980 39401 15008
rect 40271 14980 40316 15008
rect 39356 14968 39362 14980
rect 40310 14968 40316 14980
rect 40368 14968 40374 15020
rect 40402 14968 40408 15020
rect 40460 15008 40466 15020
rect 40865 15011 40923 15017
rect 40865 15008 40877 15011
rect 40460 14980 40877 15008
rect 40460 14968 40466 14980
rect 40865 14977 40877 14980
rect 40911 14977 40923 15011
rect 40865 14971 40923 14977
rect 41693 15011 41751 15017
rect 41693 14977 41705 15011
rect 41739 14977 41751 15011
rect 43438 15008 43444 15020
rect 43399 14980 43444 15008
rect 41693 14971 41751 14977
rect 38120 14912 39252 14940
rect 37461 14903 37519 14909
rect 12526 14832 12532 14884
rect 12584 14872 12590 14884
rect 12710 14872 12716 14884
rect 12584 14844 12716 14872
rect 12584 14832 12590 14844
rect 12710 14832 12716 14844
rect 12768 14832 12774 14884
rect 23385 14875 23443 14881
rect 23385 14872 23397 14875
rect 22066 14844 23397 14872
rect 14645 14807 14703 14813
rect 14645 14773 14657 14807
rect 14691 14804 14703 14807
rect 15010 14804 15016 14816
rect 14691 14776 15016 14804
rect 14691 14773 14703 14776
rect 14645 14767 14703 14773
rect 15010 14764 15016 14776
rect 15068 14764 15074 14816
rect 16114 14764 16120 14816
rect 16172 14804 16178 14816
rect 22066 14804 22094 14844
rect 23385 14841 23397 14844
rect 23431 14841 23443 14875
rect 23385 14835 23443 14841
rect 24394 14832 24400 14884
rect 24452 14872 24458 14884
rect 27706 14872 27712 14884
rect 24452 14844 27712 14872
rect 24452 14832 24458 14844
rect 27706 14832 27712 14844
rect 27764 14832 27770 14884
rect 29840 14844 31984 14872
rect 16172 14776 22094 14804
rect 16172 14764 16178 14776
rect 22370 14764 22376 14816
rect 22428 14804 22434 14816
rect 22649 14807 22707 14813
rect 22649 14804 22661 14807
rect 22428 14776 22661 14804
rect 22428 14764 22434 14776
rect 22649 14773 22661 14776
rect 22695 14773 22707 14807
rect 22649 14767 22707 14773
rect 24486 14764 24492 14816
rect 24544 14804 24550 14816
rect 26786 14804 26792 14816
rect 24544 14776 26792 14804
rect 24544 14764 24550 14776
rect 26786 14764 26792 14776
rect 26844 14764 26850 14816
rect 26878 14764 26884 14816
rect 26936 14804 26942 14816
rect 29840 14804 29868 14844
rect 26936 14776 29868 14804
rect 31956 14804 31984 14844
rect 32030 14832 32036 14884
rect 32088 14872 32094 14884
rect 37476 14872 37504 14903
rect 41322 14900 41328 14952
rect 41380 14940 41386 14952
rect 41708 14940 41736 14971
rect 43438 14968 43444 14980
rect 43496 14968 43502 15020
rect 45940 15017 45968 15048
rect 46014 15036 46020 15088
rect 46072 15076 46078 15088
rect 48682 15076 48688 15088
rect 46072 15048 48688 15076
rect 46072 15036 46078 15048
rect 48682 15036 48688 15048
rect 48740 15036 48746 15088
rect 48774 15036 48780 15088
rect 48832 15076 48838 15088
rect 49421 15079 49479 15085
rect 49421 15076 49433 15079
rect 48832 15048 49433 15076
rect 48832 15036 48838 15048
rect 49421 15045 49433 15048
rect 49467 15045 49479 15079
rect 49421 15039 49479 15045
rect 49694 15036 49700 15088
rect 49752 15076 49758 15088
rect 49752 15048 49910 15076
rect 49752 15036 49758 15048
rect 50706 15036 50712 15088
rect 50764 15076 50770 15088
rect 53098 15076 53104 15088
rect 50764 15048 53104 15076
rect 50764 15036 50770 15048
rect 53098 15036 53104 15048
rect 53156 15036 53162 15088
rect 45925 15011 45983 15017
rect 45925 14977 45937 15011
rect 45971 15008 45983 15011
rect 47118 15008 47124 15020
rect 45971 14980 47124 15008
rect 45971 14977 45983 14980
rect 45925 14971 45983 14977
rect 47118 14968 47124 14980
rect 47176 14968 47182 15020
rect 47210 14968 47216 15020
rect 47268 15008 47274 15020
rect 48041 15011 48099 15017
rect 48041 15008 48053 15011
rect 47268 14980 48053 15008
rect 47268 14968 47274 14980
rect 48041 14977 48053 14980
rect 48087 14977 48099 15011
rect 49142 15008 49148 15020
rect 49103 14980 49148 15008
rect 48041 14971 48099 14977
rect 49142 14968 49148 14980
rect 49200 14968 49206 15020
rect 53208 15008 53236 15116
rect 53742 15036 53748 15088
rect 53800 15036 53806 15088
rect 54938 15076 54944 15088
rect 54772 15048 54944 15076
rect 54772 15017 54800 15048
rect 54938 15036 54944 15048
rect 54996 15076 55002 15088
rect 55490 15076 55496 15088
rect 54996 15048 55496 15076
rect 54996 15036 55002 15048
rect 55490 15036 55496 15048
rect 55548 15036 55554 15088
rect 59078 15076 59084 15088
rect 59039 15048 59084 15076
rect 59078 15036 59084 15048
rect 59136 15036 59142 15088
rect 51046 14980 53236 15008
rect 54757 15011 54815 15017
rect 41380 14912 41736 14940
rect 41380 14900 41386 14912
rect 42702 14900 42708 14952
rect 42760 14940 42766 14952
rect 45833 14943 45891 14949
rect 45833 14940 45845 14943
rect 42760 14912 45845 14940
rect 42760 14900 42766 14912
rect 45833 14909 45845 14912
rect 45879 14940 45891 14943
rect 46014 14940 46020 14952
rect 45879 14912 46020 14940
rect 45879 14909 45891 14912
rect 45833 14903 45891 14909
rect 46014 14900 46020 14912
rect 46072 14900 46078 14952
rect 46290 14900 46296 14952
rect 46348 14940 46354 14952
rect 46661 14943 46719 14949
rect 46661 14940 46673 14943
rect 46348 14912 46673 14940
rect 46348 14900 46354 14912
rect 46661 14909 46673 14912
rect 46707 14909 46719 14943
rect 48314 14940 48320 14952
rect 48275 14912 48320 14940
rect 46661 14903 46719 14909
rect 48314 14900 48320 14912
rect 48372 14900 48378 14952
rect 51046 14940 51074 14980
rect 54757 14977 54769 15011
rect 54803 14977 54815 15011
rect 54757 14971 54815 14977
rect 56594 14968 56600 15020
rect 56652 14968 56658 15020
rect 49252 14912 51074 14940
rect 41230 14872 41236 14884
rect 32088 14844 37504 14872
rect 37844 14844 41236 14872
rect 32088 14832 32094 14844
rect 33042 14804 33048 14816
rect 31956 14776 33048 14804
rect 26936 14764 26942 14776
rect 33042 14764 33048 14776
rect 33100 14764 33106 14816
rect 35986 14804 35992 14816
rect 35947 14776 35992 14804
rect 35986 14764 35992 14776
rect 36044 14764 36050 14816
rect 36078 14764 36084 14816
rect 36136 14804 36142 14816
rect 37844 14804 37872 14844
rect 41230 14832 41236 14844
rect 41288 14832 41294 14884
rect 48332 14872 48360 14900
rect 49252 14872 49280 14912
rect 52086 14900 52092 14952
rect 52144 14940 52150 14952
rect 54481 14943 54539 14949
rect 54481 14940 54493 14943
rect 52144 14912 54493 14940
rect 52144 14900 52150 14912
rect 54481 14909 54493 14912
rect 54527 14909 54539 14943
rect 55214 14940 55220 14952
rect 55175 14912 55220 14940
rect 54481 14903 54539 14909
rect 55214 14900 55220 14912
rect 55272 14900 55278 14952
rect 55493 14943 55551 14949
rect 55493 14940 55505 14943
rect 55324 14912 55505 14940
rect 41386 14844 46428 14872
rect 48332 14844 49280 14872
rect 50448 14844 53328 14872
rect 40218 14804 40224 14816
rect 36136 14776 37872 14804
rect 40179 14776 40224 14804
rect 36136 14764 36142 14776
rect 40218 14764 40224 14776
rect 40276 14764 40282 14816
rect 40957 14807 41015 14813
rect 40957 14773 40969 14807
rect 41003 14804 41015 14807
rect 41386 14804 41414 14844
rect 41598 14804 41604 14816
rect 41003 14776 41414 14804
rect 41559 14776 41604 14804
rect 41003 14773 41015 14776
rect 40957 14767 41015 14773
rect 41598 14764 41604 14776
rect 41656 14764 41662 14816
rect 42702 14764 42708 14816
rect 42760 14804 42766 14816
rect 42889 14807 42947 14813
rect 42889 14804 42901 14807
rect 42760 14776 42901 14804
rect 42760 14764 42766 14776
rect 42889 14773 42901 14776
rect 42935 14773 42947 14807
rect 44726 14804 44732 14816
rect 44687 14776 44732 14804
rect 42889 14767 42947 14773
rect 44726 14764 44732 14776
rect 44784 14764 44790 14816
rect 46400 14804 46428 14844
rect 50448 14804 50476 14844
rect 50890 14804 50896 14816
rect 46400 14776 50476 14804
rect 50851 14776 50896 14804
rect 50890 14764 50896 14776
rect 50948 14764 50954 14816
rect 51537 14807 51595 14813
rect 51537 14773 51549 14807
rect 51583 14804 51595 14807
rect 51718 14804 51724 14816
rect 51583 14776 51724 14804
rect 51583 14773 51595 14776
rect 51537 14767 51595 14773
rect 51718 14764 51724 14776
rect 51776 14764 51782 14816
rect 51994 14804 52000 14816
rect 51955 14776 52000 14804
rect 51994 14764 52000 14776
rect 52052 14764 52058 14816
rect 53300 14804 53328 14844
rect 55324 14804 55352 14912
rect 55493 14909 55505 14912
rect 55539 14909 55551 14943
rect 55493 14903 55551 14909
rect 55582 14900 55588 14952
rect 55640 14940 55646 14952
rect 56686 14940 56692 14952
rect 55640 14912 56692 14940
rect 55640 14900 55646 14912
rect 56686 14900 56692 14912
rect 56744 14900 56750 14952
rect 56962 14940 56968 14952
rect 56923 14912 56968 14940
rect 56962 14900 56968 14912
rect 57020 14900 57026 14952
rect 59188 14940 59216 15116
rect 59906 15104 59912 15156
rect 59964 15144 59970 15156
rect 61562 15144 61568 15156
rect 59964 15116 61568 15144
rect 59964 15104 59970 15116
rect 61562 15104 61568 15116
rect 61620 15104 61626 15156
rect 62298 15144 62304 15156
rect 62211 15116 62304 15144
rect 62298 15104 62304 15116
rect 62356 15144 62362 15156
rect 66162 15144 66168 15156
rect 62356 15116 66168 15144
rect 62356 15104 62362 15116
rect 66162 15104 66168 15116
rect 66220 15104 66226 15156
rect 67361 15147 67419 15153
rect 67361 15113 67373 15147
rect 67407 15144 67419 15147
rect 68370 15144 68376 15156
rect 67407 15116 68376 15144
rect 67407 15113 67419 15116
rect 67361 15107 67419 15113
rect 68370 15104 68376 15116
rect 68428 15104 68434 15156
rect 70946 15144 70952 15156
rect 68572 15116 70952 15144
rect 60090 15036 60096 15088
rect 60148 15036 60154 15088
rect 60826 15076 60832 15088
rect 60787 15048 60832 15076
rect 60826 15036 60832 15048
rect 60884 15036 60890 15088
rect 61470 15036 61476 15088
rect 61528 15076 61534 15088
rect 61528 15048 61884 15076
rect 61528 15036 61534 15048
rect 61105 15011 61163 15017
rect 61105 14977 61117 15011
rect 61151 15008 61163 15011
rect 61286 15008 61292 15020
rect 61151 14980 61292 15008
rect 61151 14977 61163 14980
rect 61105 14971 61163 14977
rect 61286 14968 61292 14980
rect 61344 14968 61350 15020
rect 61562 14968 61568 15020
rect 61620 15008 61626 15020
rect 61856 15008 61884 15048
rect 61930 15036 61936 15088
rect 61988 15076 61994 15088
rect 63221 15079 63279 15085
rect 63221 15076 63233 15079
rect 61988 15048 63233 15076
rect 61988 15036 61994 15048
rect 63221 15045 63233 15048
rect 63267 15045 63279 15079
rect 65426 15076 65432 15088
rect 63221 15039 63279 15045
rect 64340 15048 65432 15076
rect 63126 15008 63132 15020
rect 61620 14980 61665 15008
rect 61856 14980 63132 15008
rect 61620 14968 61626 14980
rect 63126 14968 63132 14980
rect 63184 15008 63190 15020
rect 64340 15017 64368 15048
rect 65426 15036 65432 15048
rect 65484 15036 65490 15088
rect 66714 15076 66720 15088
rect 66378 15048 66720 15076
rect 66714 15036 66720 15048
rect 66772 15036 66778 15088
rect 64325 15011 64383 15017
rect 64325 15008 64337 15011
rect 63184 14980 64337 15008
rect 63184 14968 63190 14980
rect 64325 14977 64337 14980
rect 64371 14977 64383 15011
rect 67174 15008 67180 15020
rect 67135 14980 67180 15008
rect 64325 14971 64383 14977
rect 67174 14968 67180 14980
rect 67232 14968 67238 15020
rect 68572 15017 68600 15116
rect 70946 15104 70952 15116
rect 71004 15144 71010 15156
rect 71501 15147 71559 15153
rect 71501 15144 71513 15147
rect 71004 15116 71513 15144
rect 71004 15104 71010 15116
rect 71501 15113 71513 15116
rect 71547 15113 71559 15147
rect 71501 15107 71559 15113
rect 72605 15147 72663 15153
rect 72605 15113 72617 15147
rect 72651 15144 72663 15147
rect 74166 15144 74172 15156
rect 72651 15116 74172 15144
rect 72651 15113 72663 15116
rect 72605 15107 72663 15113
rect 74166 15104 74172 15116
rect 74224 15104 74230 15156
rect 74534 15104 74540 15156
rect 74592 15144 74598 15156
rect 80606 15144 80612 15156
rect 74592 15116 80612 15144
rect 74592 15104 74598 15116
rect 80606 15104 80612 15116
rect 80664 15104 80670 15156
rect 82170 15144 82176 15156
rect 82131 15116 82176 15144
rect 82170 15104 82176 15116
rect 82228 15104 82234 15156
rect 84930 15144 84936 15156
rect 82924 15116 84936 15144
rect 69201 15079 69259 15085
rect 69201 15045 69213 15079
rect 69247 15076 69259 15079
rect 70029 15079 70087 15085
rect 70029 15076 70041 15079
rect 69247 15048 70041 15076
rect 69247 15045 69259 15048
rect 69201 15039 69259 15045
rect 70029 15045 70041 15048
rect 70075 15045 70087 15079
rect 70029 15039 70087 15045
rect 71038 15036 71044 15088
rect 71096 15036 71102 15088
rect 73709 15079 73767 15085
rect 73709 15076 73721 15079
rect 71516 15048 73721 15076
rect 71516 15020 71544 15048
rect 73709 15045 73721 15048
rect 73755 15045 73767 15079
rect 73709 15039 73767 15045
rect 76466 15036 76472 15088
rect 76524 15076 76530 15088
rect 77205 15079 77263 15085
rect 77205 15076 77217 15079
rect 76524 15048 77217 15076
rect 76524 15036 76530 15048
rect 77205 15045 77217 15048
rect 77251 15045 77263 15079
rect 77205 15039 77263 15045
rect 77294 15036 77300 15088
rect 77352 15076 77358 15088
rect 77846 15076 77852 15088
rect 77352 15048 77397 15076
rect 77807 15048 77852 15076
rect 77352 15036 77358 15048
rect 77846 15036 77852 15048
rect 77904 15036 77910 15088
rect 78674 15036 78680 15088
rect 78732 15076 78738 15088
rect 80146 15076 80152 15088
rect 78732 15048 80152 15076
rect 78732 15036 78738 15048
rect 80146 15036 80152 15048
rect 80204 15036 80210 15088
rect 68557 15011 68615 15017
rect 68557 14977 68569 15011
rect 68603 14977 68615 15011
rect 68557 14971 68615 14977
rect 69014 14968 69020 15020
rect 69072 15008 69078 15020
rect 69109 15011 69167 15017
rect 69109 15008 69121 15011
rect 69072 14980 69121 15008
rect 69072 14968 69078 14980
rect 69109 14977 69121 14980
rect 69155 14977 69167 15011
rect 69109 14971 69167 14977
rect 64874 14940 64880 14952
rect 59188 14912 61056 14940
rect 61028 14872 61056 14912
rect 61212 14912 64736 14940
rect 64835 14912 64880 14940
rect 61212 14872 61240 14912
rect 62298 14872 62304 14884
rect 61028 14844 61240 14872
rect 61488 14844 62304 14872
rect 53300 14776 55352 14804
rect 55490 14764 55496 14816
rect 55548 14804 55554 14816
rect 58161 14807 58219 14813
rect 58161 14804 58173 14807
rect 55548 14776 58173 14804
rect 55548 14764 55554 14776
rect 58161 14773 58173 14776
rect 58207 14804 58219 14807
rect 58802 14804 58808 14816
rect 58207 14776 58808 14804
rect 58207 14773 58219 14776
rect 58161 14767 58219 14773
rect 58802 14764 58808 14776
rect 58860 14764 58866 14816
rect 59446 14764 59452 14816
rect 59504 14804 59510 14816
rect 61488 14804 61516 14844
rect 62298 14832 62304 14844
rect 62356 14832 62362 14884
rect 61654 14804 61660 14816
rect 59504 14776 61516 14804
rect 61615 14776 61660 14804
rect 59504 14764 59510 14776
rect 61654 14764 61660 14776
rect 61712 14764 61718 14816
rect 63865 14807 63923 14813
rect 63865 14773 63877 14807
rect 63911 14804 63923 14807
rect 64230 14804 64236 14816
rect 63911 14776 64236 14804
rect 63911 14773 63923 14776
rect 63865 14767 63923 14773
rect 64230 14764 64236 14776
rect 64288 14764 64294 14816
rect 64708 14804 64736 14912
rect 64874 14900 64880 14912
rect 64932 14900 64938 14952
rect 65153 14943 65211 14949
rect 65153 14909 65165 14943
rect 65199 14940 65211 14943
rect 65886 14940 65892 14952
rect 65199 14912 65892 14940
rect 65199 14909 65211 14912
rect 65153 14903 65211 14909
rect 65886 14900 65892 14912
rect 65944 14900 65950 14952
rect 66438 14900 66444 14952
rect 66496 14940 66502 14952
rect 69124 14940 69152 14971
rect 71498 14968 71504 15020
rect 71556 14968 71562 15020
rect 72050 14968 72056 15020
rect 72108 15008 72114 15020
rect 72145 15011 72203 15017
rect 72145 15008 72157 15011
rect 72108 14980 72157 15008
rect 72108 14968 72114 14980
rect 72145 14977 72157 14980
rect 72191 14977 72203 15011
rect 72145 14971 72203 14977
rect 74258 14968 74264 15020
rect 74316 15008 74322 15020
rect 75822 15008 75828 15020
rect 74316 14980 75828 15008
rect 74316 14968 74322 14980
rect 75822 14968 75828 14980
rect 75880 14968 75886 15020
rect 78858 15008 78864 15020
rect 78771 14980 78864 15008
rect 78858 14968 78864 14980
rect 78916 15008 78922 15020
rect 79594 15008 79600 15020
rect 78916 14980 79600 15008
rect 78916 14968 78922 14980
rect 79594 14968 79600 14980
rect 79652 14968 79658 15020
rect 80606 15008 80612 15020
rect 80567 14980 80612 15008
rect 80606 14968 80612 14980
rect 80664 14968 80670 15020
rect 82538 15008 82544 15020
rect 82499 14980 82544 15008
rect 82538 14968 82544 14980
rect 82596 14968 82602 15020
rect 82924 15017 82952 15116
rect 84930 15104 84936 15116
rect 84988 15104 84994 15156
rect 83918 15036 83924 15088
rect 83976 15076 83982 15088
rect 84013 15079 84071 15085
rect 84013 15076 84025 15079
rect 83976 15048 84025 15076
rect 83976 15036 83982 15048
rect 84013 15045 84025 15048
rect 84059 15045 84071 15079
rect 84013 15039 84071 15045
rect 82909 15011 82967 15017
rect 82909 14977 82921 15011
rect 82955 14977 82967 15011
rect 82909 14971 82967 14977
rect 86494 14968 86500 15020
rect 86552 15008 86558 15020
rect 86865 15011 86923 15017
rect 86865 15008 86877 15011
rect 86552 14980 86877 15008
rect 86552 14968 86558 14980
rect 86865 14977 86877 14980
rect 86911 14977 86923 15011
rect 86865 14971 86923 14977
rect 69750 14940 69756 14952
rect 66496 14912 69152 14940
rect 69711 14912 69756 14940
rect 66496 14900 66502 14912
rect 69124 14872 69152 14912
rect 69750 14900 69756 14912
rect 69808 14900 69814 14952
rect 71038 14940 71044 14952
rect 69860 14912 71044 14940
rect 69860 14872 69888 14912
rect 71038 14900 71044 14912
rect 71096 14900 71102 14952
rect 73246 14900 73252 14952
rect 73304 14940 73310 14952
rect 73617 14943 73675 14949
rect 73617 14940 73629 14943
rect 73304 14912 73629 14940
rect 73304 14900 73310 14912
rect 73617 14909 73629 14912
rect 73663 14909 73675 14943
rect 80698 14940 80704 14952
rect 73617 14903 73675 14909
rect 75104 14912 80054 14940
rect 80611 14912 80704 14940
rect 66180 14844 68600 14872
rect 69124 14844 69888 14872
rect 66180 14804 66208 14844
rect 64708 14776 66208 14804
rect 66625 14807 66683 14813
rect 66625 14773 66637 14807
rect 66671 14804 66683 14807
rect 67726 14804 67732 14816
rect 66671 14776 67732 14804
rect 66671 14773 66683 14776
rect 66625 14767 66683 14773
rect 67726 14764 67732 14776
rect 67784 14764 67790 14816
rect 68462 14804 68468 14816
rect 68423 14776 68468 14804
rect 68462 14764 68468 14776
rect 68520 14764 68526 14816
rect 68572 14804 68600 14844
rect 72142 14832 72148 14884
rect 72200 14872 72206 14884
rect 72421 14875 72479 14881
rect 72421 14872 72433 14875
rect 72200 14844 72433 14872
rect 72200 14832 72206 14844
rect 72421 14841 72433 14844
rect 72467 14841 72479 14875
rect 72421 14835 72479 14841
rect 74169 14875 74227 14881
rect 74169 14841 74181 14875
rect 74215 14872 74227 14875
rect 75104 14872 75132 14912
rect 75270 14872 75276 14884
rect 74215 14844 75132 14872
rect 75231 14844 75276 14872
rect 74215 14841 74227 14844
rect 74169 14835 74227 14841
rect 75270 14832 75276 14844
rect 75328 14832 75334 14884
rect 80026 14872 80054 14912
rect 80698 14900 80704 14912
rect 80756 14940 80762 14952
rect 82814 14940 82820 14952
rect 80756 14912 82820 14940
rect 80756 14900 80762 14912
rect 82814 14900 82820 14912
rect 82872 14900 82878 14952
rect 82998 14900 83004 14952
rect 83056 14940 83062 14952
rect 83921 14943 83979 14949
rect 83921 14940 83933 14943
rect 83056 14912 83933 14940
rect 83056 14900 83062 14912
rect 83921 14909 83933 14912
rect 83967 14909 83979 14943
rect 83921 14903 83979 14909
rect 85022 14900 85028 14952
rect 85080 14940 85086 14952
rect 85669 14943 85727 14949
rect 85669 14940 85681 14943
rect 85080 14912 85681 14940
rect 85080 14900 85086 14912
rect 85669 14909 85681 14912
rect 85715 14909 85727 14943
rect 85669 14903 85727 14909
rect 86770 14900 86776 14952
rect 86828 14940 86834 14952
rect 87969 14943 88027 14949
rect 87969 14940 87981 14943
rect 86828 14912 87981 14940
rect 86828 14900 86834 14912
rect 87969 14909 87981 14912
rect 88015 14909 88027 14943
rect 87969 14903 88027 14909
rect 84473 14875 84531 14881
rect 84473 14872 84485 14875
rect 80026 14844 84485 14872
rect 84473 14841 84485 14844
rect 84519 14872 84531 14875
rect 92658 14872 92664 14884
rect 84519 14844 92664 14872
rect 84519 14841 84531 14844
rect 84473 14835 84531 14841
rect 92658 14832 92664 14844
rect 92716 14832 92722 14884
rect 74534 14804 74540 14816
rect 68572 14776 74540 14804
rect 74534 14764 74540 14776
rect 74592 14764 74598 14816
rect 74626 14764 74632 14816
rect 74684 14804 74690 14816
rect 74721 14807 74779 14813
rect 74721 14804 74733 14807
rect 74684 14776 74733 14804
rect 74684 14764 74690 14776
rect 74721 14773 74733 14776
rect 74767 14773 74779 14807
rect 74721 14767 74779 14773
rect 75914 14764 75920 14816
rect 75972 14804 75978 14816
rect 76377 14807 76435 14813
rect 76377 14804 76389 14807
rect 75972 14776 76389 14804
rect 75972 14764 75978 14776
rect 76377 14773 76389 14776
rect 76423 14773 76435 14807
rect 76377 14767 76435 14773
rect 78214 14764 78220 14816
rect 78272 14804 78278 14816
rect 78769 14807 78827 14813
rect 78769 14804 78781 14807
rect 78272 14776 78781 14804
rect 78272 14764 78278 14776
rect 78769 14773 78781 14776
rect 78815 14773 78827 14807
rect 79318 14804 79324 14816
rect 79279 14776 79324 14804
rect 78769 14767 78827 14773
rect 79318 14764 79324 14776
rect 79376 14764 79382 14816
rect 80330 14804 80336 14816
rect 80291 14776 80336 14804
rect 80330 14764 80336 14776
rect 80388 14764 80394 14816
rect 81345 14807 81403 14813
rect 81345 14773 81357 14807
rect 81391 14804 81403 14807
rect 81710 14804 81716 14816
rect 81391 14776 81716 14804
rect 81391 14773 81403 14776
rect 81345 14767 81403 14773
rect 81710 14764 81716 14776
rect 81768 14764 81774 14816
rect 85206 14804 85212 14816
rect 85167 14776 85212 14804
rect 85206 14764 85212 14776
rect 85264 14764 85270 14816
rect 86405 14807 86463 14813
rect 86405 14773 86417 14807
rect 86451 14804 86463 14807
rect 86770 14804 86776 14816
rect 86451 14776 86776 14804
rect 86451 14773 86463 14776
rect 86405 14767 86463 14773
rect 86770 14764 86776 14776
rect 86828 14764 86834 14816
rect 86954 14764 86960 14816
rect 87012 14804 87018 14816
rect 87417 14807 87475 14813
rect 87417 14804 87429 14807
rect 87012 14776 87429 14804
rect 87012 14764 87018 14776
rect 87417 14773 87429 14776
rect 87463 14773 87475 14807
rect 89070 14804 89076 14816
rect 89031 14776 89076 14804
rect 87417 14767 87475 14773
rect 89070 14764 89076 14776
rect 89128 14804 89134 14816
rect 89533 14807 89591 14813
rect 89533 14804 89545 14807
rect 89128 14776 89545 14804
rect 89128 14764 89134 14776
rect 89533 14773 89545 14776
rect 89579 14804 89591 14807
rect 90085 14807 90143 14813
rect 90085 14804 90097 14807
rect 89579 14776 90097 14804
rect 89579 14773 89591 14776
rect 89533 14767 89591 14773
rect 90085 14773 90097 14776
rect 90131 14773 90143 14807
rect 90085 14767 90143 14773
rect 90450 14764 90456 14816
rect 90508 14804 90514 14816
rect 90729 14807 90787 14813
rect 90729 14804 90741 14807
rect 90508 14776 90741 14804
rect 90508 14764 90514 14776
rect 90729 14773 90741 14776
rect 90775 14773 90787 14807
rect 90729 14767 90787 14773
rect 1104 14714 94852 14736
rect 1104 14662 12668 14714
rect 12720 14662 12732 14714
rect 12784 14662 12796 14714
rect 12848 14662 12860 14714
rect 12912 14662 12924 14714
rect 12976 14662 36105 14714
rect 36157 14662 36169 14714
rect 36221 14662 36233 14714
rect 36285 14662 36297 14714
rect 36349 14662 36361 14714
rect 36413 14662 59542 14714
rect 59594 14662 59606 14714
rect 59658 14662 59670 14714
rect 59722 14662 59734 14714
rect 59786 14662 59798 14714
rect 59850 14662 82979 14714
rect 83031 14662 83043 14714
rect 83095 14662 83107 14714
rect 83159 14662 83171 14714
rect 83223 14662 83235 14714
rect 83287 14662 94852 14714
rect 1104 14640 94852 14662
rect 24394 14600 24400 14612
rect 20916 14572 24400 14600
rect 8018 14492 8024 14544
rect 8076 14532 8082 14544
rect 11793 14535 11851 14541
rect 8076 14504 9260 14532
rect 8076 14492 8082 14504
rect 7282 14396 7288 14408
rect 7243 14368 7288 14396
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 8018 14396 8024 14408
rect 7979 14368 8024 14396
rect 8018 14356 8024 14368
rect 8076 14356 8082 14408
rect 9122 14328 9128 14340
rect 8234 14300 9128 14328
rect 9122 14288 9128 14300
rect 9180 14288 9186 14340
rect 9232 14337 9260 14504
rect 11793 14501 11805 14535
rect 11839 14532 11851 14535
rect 15378 14532 15384 14544
rect 11839 14504 15384 14532
rect 11839 14501 11851 14504
rect 11793 14495 11851 14501
rect 15378 14492 15384 14504
rect 15436 14492 15442 14544
rect 11330 14464 11336 14476
rect 11291 14436 11336 14464
rect 11330 14424 11336 14436
rect 11388 14424 11394 14476
rect 12437 14467 12495 14473
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 14550 14464 14556 14476
rect 12483 14436 14556 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 19429 14467 19487 14473
rect 19429 14464 19441 14467
rect 15252 14436 19441 14464
rect 15252 14424 15258 14436
rect 19429 14433 19441 14436
rect 19475 14433 19487 14467
rect 19429 14427 19487 14433
rect 19705 14467 19763 14473
rect 19705 14433 19717 14467
rect 19751 14464 19763 14467
rect 20916 14464 20944 14572
rect 24394 14560 24400 14572
rect 24452 14560 24458 14612
rect 24578 14600 24584 14612
rect 24539 14572 24584 14600
rect 24578 14560 24584 14572
rect 24636 14560 24642 14612
rect 25038 14560 25044 14612
rect 25096 14600 25102 14612
rect 28718 14600 28724 14612
rect 25096 14572 28724 14600
rect 25096 14560 25102 14572
rect 28718 14560 28724 14572
rect 28776 14560 28782 14612
rect 35986 14600 35992 14612
rect 28828 14572 35992 14600
rect 23750 14492 23756 14544
rect 23808 14532 23814 14544
rect 27154 14532 27160 14544
rect 23808 14504 27160 14532
rect 23808 14492 23814 14504
rect 27154 14492 27160 14504
rect 27212 14492 27218 14544
rect 28828 14532 28856 14572
rect 35986 14560 35992 14572
rect 36044 14560 36050 14612
rect 42702 14600 42708 14612
rect 38626 14572 42708 14600
rect 28552 14504 28856 14532
rect 28905 14535 28963 14541
rect 19751 14436 20944 14464
rect 21453 14467 21511 14473
rect 19751 14433 19763 14436
rect 19705 14427 19763 14433
rect 21453 14433 21465 14467
rect 21499 14464 21511 14467
rect 26878 14464 26884 14476
rect 21499 14436 26884 14464
rect 21499 14433 21511 14436
rect 21453 14427 21511 14433
rect 26878 14424 26884 14436
rect 26936 14424 26942 14476
rect 27433 14467 27491 14473
rect 27433 14433 27445 14467
rect 27479 14464 27491 14467
rect 28552 14464 28580 14504
rect 28905 14501 28917 14535
rect 28951 14532 28963 14535
rect 28951 14504 35894 14532
rect 28951 14501 28963 14504
rect 28905 14495 28963 14501
rect 27479 14436 28580 14464
rect 27479 14433 27491 14436
rect 27433 14427 27491 14433
rect 28810 14424 28816 14476
rect 28868 14464 28874 14476
rect 30650 14464 30656 14476
rect 28868 14436 30656 14464
rect 28868 14424 28874 14436
rect 30650 14424 30656 14436
rect 30708 14424 30714 14476
rect 30760 14436 31800 14464
rect 11422 14396 11428 14408
rect 11383 14368 11428 14396
rect 11422 14356 11428 14368
rect 11480 14356 11486 14408
rect 12526 14396 12532 14408
rect 12487 14368 12532 14396
rect 12526 14356 12532 14368
rect 12584 14356 12590 14408
rect 15102 14356 15108 14408
rect 15160 14396 15166 14408
rect 15657 14399 15715 14405
rect 15657 14396 15669 14399
rect 15160 14368 15669 14396
rect 15160 14356 15166 14368
rect 15657 14365 15669 14368
rect 15703 14365 15715 14399
rect 15657 14359 15715 14365
rect 20806 14356 20812 14408
rect 20864 14356 20870 14408
rect 23753 14399 23811 14405
rect 23753 14365 23765 14399
rect 23799 14396 23811 14399
rect 24486 14396 24492 14408
rect 23799 14368 24492 14396
rect 23799 14365 23811 14368
rect 23753 14359 23811 14365
rect 24486 14356 24492 14368
rect 24544 14356 24550 14408
rect 24762 14396 24768 14408
rect 24723 14368 24768 14396
rect 24762 14356 24768 14368
rect 24820 14356 24826 14408
rect 25590 14396 25596 14408
rect 24964 14368 25596 14396
rect 9217 14331 9275 14337
rect 9217 14297 9229 14331
rect 9263 14328 9275 14331
rect 12434 14328 12440 14340
rect 9263 14300 12440 14328
rect 9263 14297 9275 14300
rect 9217 14291 9275 14297
rect 12434 14288 12440 14300
rect 12492 14328 12498 14340
rect 13078 14328 13084 14340
rect 12492 14300 13084 14328
rect 12492 14288 12498 14300
rect 13078 14288 13084 14300
rect 13136 14288 13142 14340
rect 22738 14288 22744 14340
rect 22796 14288 22802 14340
rect 23477 14331 23535 14337
rect 23477 14297 23489 14331
rect 23523 14328 23535 14331
rect 24854 14328 24860 14340
rect 23523 14300 24860 14328
rect 23523 14297 23535 14300
rect 23477 14291 23535 14297
rect 24854 14288 24860 14300
rect 24912 14288 24918 14340
rect 13998 14220 14004 14272
rect 14056 14260 14062 14272
rect 14553 14263 14611 14269
rect 14553 14260 14565 14263
rect 14056 14232 14565 14260
rect 14056 14220 14062 14232
rect 14553 14229 14565 14232
rect 14599 14229 14611 14263
rect 15562 14260 15568 14272
rect 15523 14232 15568 14260
rect 14553 14223 14611 14229
rect 15562 14220 15568 14232
rect 15620 14220 15626 14272
rect 16206 14260 16212 14272
rect 16119 14232 16212 14260
rect 16206 14220 16212 14232
rect 16264 14260 16270 14272
rect 20622 14260 20628 14272
rect 16264 14232 20628 14260
rect 16264 14220 16270 14232
rect 20622 14220 20628 14232
rect 20680 14220 20686 14272
rect 22005 14263 22063 14269
rect 22005 14229 22017 14263
rect 22051 14260 22063 14263
rect 24964 14260 24992 14368
rect 25590 14356 25596 14368
rect 25648 14356 25654 14408
rect 25685 14399 25743 14405
rect 25685 14365 25697 14399
rect 25731 14396 25743 14399
rect 27154 14396 27160 14408
rect 25731 14368 27016 14396
rect 27115 14368 27160 14396
rect 25731 14365 25743 14368
rect 25685 14359 25743 14365
rect 25590 14260 25596 14272
rect 22051 14232 24992 14260
rect 25551 14232 25596 14260
rect 22051 14229 22063 14232
rect 22005 14223 22063 14229
rect 25590 14220 25596 14232
rect 25648 14220 25654 14272
rect 26234 14220 26240 14272
rect 26292 14260 26298 14272
rect 26605 14263 26663 14269
rect 26605 14260 26617 14263
rect 26292 14232 26617 14260
rect 26292 14220 26298 14232
rect 26605 14229 26617 14232
rect 26651 14229 26663 14263
rect 26988 14260 27016 14368
rect 27154 14356 27160 14368
rect 27212 14356 27218 14408
rect 28534 14356 28540 14408
rect 28592 14356 28598 14408
rect 29825 14399 29883 14405
rect 29825 14365 29837 14399
rect 29871 14365 29883 14399
rect 30466 14396 30472 14408
rect 30427 14368 30472 14396
rect 29825 14359 29883 14365
rect 27338 14288 27344 14340
rect 27396 14328 27402 14340
rect 29840 14328 29868 14359
rect 30466 14356 30472 14368
rect 30524 14356 30530 14408
rect 30760 14328 30788 14436
rect 27396 14300 27844 14328
rect 27396 14288 27402 14300
rect 27614 14260 27620 14272
rect 26988 14232 27620 14260
rect 26605 14223 26663 14229
rect 27614 14220 27620 14232
rect 27672 14220 27678 14272
rect 27816 14260 27844 14300
rect 29840 14300 30788 14328
rect 31772 14328 31800 14436
rect 31846 14424 31852 14476
rect 31904 14464 31910 14476
rect 32030 14464 32036 14476
rect 31904 14436 31949 14464
rect 31991 14436 32036 14464
rect 31904 14424 31910 14436
rect 32030 14424 32036 14436
rect 32088 14424 32094 14476
rect 32766 14424 32772 14476
rect 32824 14464 32830 14476
rect 35866 14464 35894 14504
rect 38626 14464 38654 14572
rect 42702 14560 42708 14572
rect 42760 14560 42766 14612
rect 46293 14603 46351 14609
rect 46293 14569 46305 14603
rect 46339 14600 46351 14603
rect 46658 14600 46664 14612
rect 46339 14572 46664 14600
rect 46339 14569 46351 14572
rect 46293 14563 46351 14569
rect 46658 14560 46664 14572
rect 46716 14560 46722 14612
rect 47118 14560 47124 14612
rect 47176 14600 47182 14612
rect 50706 14600 50712 14612
rect 47176 14572 50712 14600
rect 47176 14560 47182 14572
rect 50706 14560 50712 14572
rect 50764 14560 50770 14612
rect 50890 14560 50896 14612
rect 50948 14600 50954 14612
rect 51442 14600 51448 14612
rect 50948 14572 51448 14600
rect 50948 14560 50954 14572
rect 51442 14560 51448 14572
rect 51500 14560 51506 14612
rect 51534 14560 51540 14612
rect 51592 14600 51598 14612
rect 54202 14600 54208 14612
rect 51592 14572 54208 14600
rect 51592 14560 51598 14572
rect 54202 14560 54208 14572
rect 54260 14560 54266 14612
rect 56229 14603 56287 14609
rect 55784 14572 56180 14600
rect 41874 14492 41880 14544
rect 41932 14532 41938 14544
rect 49326 14532 49332 14544
rect 41932 14504 49332 14532
rect 41932 14492 41938 14504
rect 40586 14464 40592 14476
rect 32824 14436 35296 14464
rect 35866 14436 38654 14464
rect 40547 14436 40592 14464
rect 32824 14424 32830 14436
rect 34882 14356 34888 14408
rect 34940 14396 34946 14408
rect 35161 14399 35219 14405
rect 35161 14396 35173 14399
rect 34940 14368 35173 14396
rect 34940 14356 34946 14368
rect 35161 14365 35173 14368
rect 35207 14365 35219 14399
rect 35268 14396 35296 14436
rect 40586 14424 40592 14436
rect 40644 14424 40650 14476
rect 40678 14424 40684 14476
rect 40736 14464 40742 14476
rect 41322 14464 41328 14476
rect 40736 14436 41328 14464
rect 40736 14424 40742 14436
rect 41322 14424 41328 14436
rect 41380 14464 41386 14476
rect 44100 14473 44128 14504
rect 49326 14492 49332 14504
rect 49384 14492 49390 14544
rect 53098 14492 53104 14544
rect 53156 14532 53162 14544
rect 55784 14532 55812 14572
rect 53156 14504 55812 14532
rect 56152 14532 56180 14572
rect 56229 14569 56241 14603
rect 56275 14600 56287 14603
rect 64874 14600 64880 14612
rect 56275 14572 64880 14600
rect 56275 14569 56287 14572
rect 56229 14563 56287 14569
rect 64874 14560 64880 14572
rect 64932 14560 64938 14612
rect 64984 14572 72464 14600
rect 59262 14532 59268 14544
rect 56152 14504 59268 14532
rect 53156 14492 53162 14504
rect 59262 14492 59268 14504
rect 59320 14492 59326 14544
rect 59354 14492 59360 14544
rect 59412 14532 59418 14544
rect 60458 14532 60464 14544
rect 59412 14504 60464 14532
rect 59412 14492 59418 14504
rect 60458 14492 60464 14504
rect 60516 14492 60522 14544
rect 63034 14492 63040 14544
rect 63092 14532 63098 14544
rect 63221 14535 63279 14541
rect 63221 14532 63233 14535
rect 63092 14504 63233 14532
rect 63092 14492 63098 14504
rect 63221 14501 63233 14504
rect 63267 14532 63279 14535
rect 64984 14532 65012 14572
rect 63267 14504 65012 14532
rect 69860 14504 71176 14532
rect 63267 14501 63279 14504
rect 63221 14495 63279 14501
rect 44085 14467 44143 14473
rect 41380 14436 41828 14464
rect 41380 14424 41386 14436
rect 35268 14368 37044 14396
rect 35161 14359 35219 14365
rect 32950 14328 32956 14340
rect 31772 14300 32956 14328
rect 29840 14260 29868 14300
rect 32950 14288 32956 14300
rect 33008 14288 33014 14340
rect 33689 14331 33747 14337
rect 33689 14297 33701 14331
rect 33735 14328 33747 14331
rect 33962 14328 33968 14340
rect 33735 14300 33968 14328
rect 33735 14297 33747 14300
rect 33689 14291 33747 14297
rect 33962 14288 33968 14300
rect 34020 14288 34026 14340
rect 35989 14331 36047 14337
rect 35989 14328 36001 14331
rect 34256 14300 36001 14328
rect 34256 14272 34284 14300
rect 35989 14297 36001 14300
rect 36035 14297 36047 14331
rect 37016 14328 37044 14368
rect 37090 14356 37096 14408
rect 37148 14396 37154 14408
rect 37366 14396 37372 14408
rect 37148 14368 37193 14396
rect 37327 14368 37372 14396
rect 37148 14356 37154 14368
rect 37366 14356 37372 14368
rect 37424 14356 37430 14408
rect 38289 14399 38347 14405
rect 38289 14365 38301 14399
rect 38335 14365 38347 14399
rect 38838 14396 38844 14408
rect 38799 14368 38844 14396
rect 38289 14359 38347 14365
rect 38197 14331 38255 14337
rect 38197 14328 38209 14331
rect 37016 14300 38209 14328
rect 35989 14291 36047 14297
rect 38197 14297 38209 14300
rect 38243 14297 38255 14331
rect 38197 14291 38255 14297
rect 27816 14232 29868 14260
rect 29917 14263 29975 14269
rect 29917 14229 29929 14263
rect 29963 14260 29975 14263
rect 30006 14260 30012 14272
rect 29963 14232 30012 14260
rect 29963 14229 29975 14232
rect 29917 14223 29975 14229
rect 30006 14220 30012 14232
rect 30064 14220 30070 14272
rect 30190 14220 30196 14272
rect 30248 14260 30254 14272
rect 30561 14263 30619 14269
rect 30561 14260 30573 14263
rect 30248 14232 30573 14260
rect 30248 14220 30254 14232
rect 30561 14229 30573 14232
rect 30607 14229 30619 14263
rect 31386 14260 31392 14272
rect 31347 14232 31392 14260
rect 30561 14223 30619 14229
rect 31386 14220 31392 14232
rect 31444 14220 31450 14272
rect 34238 14260 34244 14272
rect 34199 14232 34244 14260
rect 34238 14220 34244 14232
rect 34296 14220 34302 14272
rect 35066 14260 35072 14272
rect 35027 14232 35072 14260
rect 35066 14220 35072 14232
rect 35124 14220 35130 14272
rect 35434 14220 35440 14272
rect 35492 14260 35498 14272
rect 36541 14263 36599 14269
rect 36541 14260 36553 14263
rect 35492 14232 36553 14260
rect 35492 14220 35498 14232
rect 36541 14229 36553 14232
rect 36587 14229 36599 14263
rect 38304 14260 38332 14359
rect 38838 14356 38844 14368
rect 38896 14356 38902 14408
rect 40126 14396 40132 14408
rect 38948 14368 40132 14396
rect 38562 14288 38568 14340
rect 38620 14328 38626 14340
rect 38948 14328 38976 14368
rect 40126 14356 40132 14368
rect 40184 14396 40190 14408
rect 40313 14399 40371 14405
rect 40313 14396 40325 14399
rect 40184 14368 40325 14396
rect 40184 14356 40190 14368
rect 40313 14365 40325 14368
rect 40359 14365 40371 14399
rect 41800 14396 41828 14436
rect 44085 14433 44097 14467
rect 44131 14433 44143 14467
rect 44085 14427 44143 14433
rect 48593 14467 48651 14473
rect 48593 14433 48605 14467
rect 48639 14464 48651 14467
rect 55766 14464 55772 14476
rect 48639 14436 55772 14464
rect 48639 14433 48651 14436
rect 48593 14427 48651 14433
rect 55766 14424 55772 14436
rect 55824 14424 55830 14476
rect 55861 14467 55919 14473
rect 55861 14433 55873 14467
rect 55907 14433 55919 14467
rect 55861 14427 55919 14433
rect 42613 14399 42671 14405
rect 42613 14396 42625 14399
rect 41800 14368 42625 14396
rect 40313 14359 40371 14365
rect 42613 14365 42625 14368
rect 42659 14365 42671 14399
rect 43806 14396 43812 14408
rect 43767 14368 43812 14396
rect 42613 14359 42671 14365
rect 43806 14356 43812 14368
rect 43864 14356 43870 14408
rect 45462 14396 45468 14408
rect 45375 14368 45468 14396
rect 45462 14356 45468 14368
rect 45520 14396 45526 14408
rect 45738 14396 45744 14408
rect 45520 14368 45744 14396
rect 45520 14356 45526 14368
rect 45738 14356 45744 14368
rect 45796 14396 45802 14408
rect 46201 14399 46259 14405
rect 46201 14396 46213 14399
rect 45796 14368 46213 14396
rect 45796 14356 45802 14368
rect 46201 14365 46213 14368
rect 46247 14396 46259 14399
rect 49234 14396 49240 14408
rect 46247 14368 49240 14396
rect 46247 14365 46259 14368
rect 46201 14359 46259 14365
rect 49234 14356 49240 14368
rect 49292 14356 49298 14408
rect 50614 14356 50620 14408
rect 50672 14396 50678 14408
rect 50985 14399 51043 14405
rect 50985 14396 50997 14399
rect 50672 14368 50997 14396
rect 50672 14356 50678 14368
rect 50985 14365 50997 14368
rect 51031 14396 51043 14399
rect 51534 14396 51540 14408
rect 51031 14368 51540 14396
rect 51031 14365 51043 14368
rect 50985 14359 51043 14365
rect 51534 14356 51540 14368
rect 51592 14356 51598 14408
rect 53742 14356 53748 14408
rect 53800 14396 53806 14408
rect 54021 14399 54079 14405
rect 54021 14396 54033 14399
rect 53800 14368 54033 14396
rect 53800 14356 53806 14368
rect 54021 14365 54033 14368
rect 54067 14365 54079 14399
rect 54021 14359 54079 14365
rect 54938 14356 54944 14408
rect 54996 14396 55002 14408
rect 55582 14396 55588 14408
rect 54996 14368 55588 14396
rect 54996 14356 55002 14368
rect 55582 14356 55588 14368
rect 55640 14356 55646 14408
rect 39114 14328 39120 14340
rect 38620 14300 38976 14328
rect 39075 14300 39120 14328
rect 38620 14288 38626 14300
rect 39114 14288 39120 14300
rect 39172 14288 39178 14340
rect 41598 14288 41604 14340
rect 41656 14288 41662 14340
rect 46842 14328 46848 14340
rect 42076 14300 45508 14328
rect 46803 14300 46848 14328
rect 41874 14260 41880 14272
rect 38304 14232 41880 14260
rect 36541 14223 36599 14229
rect 41874 14220 41880 14232
rect 41932 14220 41938 14272
rect 42076 14269 42104 14300
rect 42061 14263 42119 14269
rect 42061 14229 42073 14263
rect 42107 14229 42119 14263
rect 42702 14260 42708 14272
rect 42663 14232 42708 14260
rect 42061 14223 42119 14229
rect 42702 14220 42708 14232
rect 42760 14220 42766 14272
rect 44637 14263 44695 14269
rect 44637 14229 44649 14263
rect 44683 14260 44695 14263
rect 44910 14260 44916 14272
rect 44683 14232 44916 14260
rect 44683 14229 44695 14232
rect 44637 14223 44695 14229
rect 44910 14220 44916 14232
rect 44968 14220 44974 14272
rect 45186 14220 45192 14272
rect 45244 14260 45250 14272
rect 45373 14263 45431 14269
rect 45373 14260 45385 14263
rect 45244 14232 45385 14260
rect 45244 14220 45250 14232
rect 45373 14229 45385 14232
rect 45419 14229 45431 14263
rect 45480 14260 45508 14300
rect 46842 14288 46848 14300
rect 46900 14288 46906 14340
rect 47026 14288 47032 14340
rect 47084 14328 47090 14340
rect 51810 14328 51816 14340
rect 47084 14300 51074 14328
rect 51771 14300 51816 14328
rect 47084 14288 47090 14300
rect 47302 14260 47308 14272
rect 45480 14232 47308 14260
rect 45373 14223 45431 14229
rect 47302 14220 47308 14232
rect 47360 14220 47366 14272
rect 48314 14220 48320 14272
rect 48372 14260 48378 14272
rect 49145 14263 49203 14269
rect 49145 14260 49157 14263
rect 48372 14232 49157 14260
rect 48372 14220 48378 14232
rect 49145 14229 49157 14232
rect 49191 14229 49203 14263
rect 49694 14260 49700 14272
rect 49655 14232 49700 14260
rect 49145 14223 49203 14229
rect 49694 14220 49700 14232
rect 49752 14260 49758 14272
rect 50062 14260 50068 14272
rect 49752 14232 50068 14260
rect 49752 14220 49758 14232
rect 50062 14220 50068 14232
rect 50120 14220 50126 14272
rect 50246 14220 50252 14272
rect 50304 14260 50310 14272
rect 50341 14263 50399 14269
rect 50341 14260 50353 14263
rect 50304 14232 50353 14260
rect 50304 14220 50310 14232
rect 50341 14229 50353 14232
rect 50387 14229 50399 14263
rect 51046 14260 51074 14300
rect 51810 14288 51816 14300
rect 51868 14288 51874 14340
rect 53929 14331 53987 14337
rect 53929 14328 53941 14331
rect 53038 14300 53941 14328
rect 53929 14297 53941 14300
rect 53975 14297 53987 14331
rect 53929 14291 53987 14297
rect 54846 14288 54852 14340
rect 54904 14328 54910 14340
rect 55876 14328 55904 14427
rect 56318 14424 56324 14476
rect 56376 14464 56382 14476
rect 56376 14436 60504 14464
rect 56376 14424 56382 14436
rect 55950 14356 55956 14408
rect 56008 14396 56014 14408
rect 56008 14368 56053 14396
rect 56008 14356 56014 14368
rect 58986 14356 58992 14408
rect 59044 14396 59050 14408
rect 59906 14396 59912 14408
rect 59044 14368 59912 14396
rect 59044 14356 59050 14368
rect 59906 14356 59912 14368
rect 59964 14356 59970 14408
rect 60476 14396 60504 14436
rect 60550 14424 60556 14476
rect 60608 14464 60614 14476
rect 60645 14467 60703 14473
rect 60645 14464 60657 14467
rect 60608 14436 60657 14464
rect 60608 14424 60614 14436
rect 60645 14433 60657 14436
rect 60691 14433 60703 14467
rect 67634 14464 67640 14476
rect 60645 14427 60703 14433
rect 65260 14436 67640 14464
rect 62669 14399 62727 14405
rect 60476 14368 60688 14396
rect 56226 14328 56232 14340
rect 54904 14300 56232 14328
rect 54904 14288 54910 14300
rect 56226 14288 56232 14300
rect 56284 14288 56290 14340
rect 57238 14328 57244 14340
rect 57199 14300 57244 14328
rect 57238 14288 57244 14300
rect 57296 14288 57302 14340
rect 58250 14288 58256 14340
rect 58308 14328 58314 14340
rect 58805 14331 58863 14337
rect 58805 14328 58817 14331
rect 58308 14300 58817 14328
rect 58308 14288 58314 14300
rect 58805 14297 58817 14300
rect 58851 14297 58863 14331
rect 58805 14291 58863 14297
rect 59357 14331 59415 14337
rect 59357 14297 59369 14331
rect 59403 14328 59415 14331
rect 60550 14328 60556 14340
rect 59403 14300 60556 14328
rect 59403 14297 59415 14300
rect 59357 14291 59415 14297
rect 60550 14288 60556 14300
rect 60608 14288 60614 14340
rect 53285 14263 53343 14269
rect 53285 14260 53297 14263
rect 51046 14232 53297 14260
rect 50341 14223 50399 14229
rect 53285 14229 53297 14232
rect 53331 14229 53343 14263
rect 53285 14223 53343 14229
rect 54478 14220 54484 14272
rect 54536 14260 54542 14272
rect 54573 14263 54631 14269
rect 54573 14260 54585 14263
rect 54536 14232 54585 14260
rect 54536 14220 54542 14232
rect 54573 14229 54585 14232
rect 54619 14260 54631 14263
rect 57330 14260 57336 14272
rect 54619 14232 57336 14260
rect 54619 14229 54631 14232
rect 54573 14223 54631 14229
rect 57330 14220 57336 14232
rect 57388 14220 57394 14272
rect 59998 14260 60004 14272
rect 59959 14232 60004 14260
rect 59998 14220 60004 14232
rect 60056 14220 60062 14272
rect 60660 14260 60688 14368
rect 62669 14365 62681 14399
rect 62715 14396 62727 14399
rect 62942 14396 62948 14408
rect 62715 14368 62948 14396
rect 62715 14365 62727 14368
rect 62669 14359 62727 14365
rect 62942 14356 62948 14368
rect 63000 14356 63006 14408
rect 65260 14405 65288 14436
rect 67634 14424 67640 14436
rect 67692 14424 67698 14476
rect 68554 14424 68560 14476
rect 68612 14464 68618 14476
rect 69860 14464 69888 14504
rect 71038 14464 71044 14476
rect 68612 14436 69888 14464
rect 70999 14436 71044 14464
rect 68612 14424 68618 14436
rect 71038 14424 71044 14436
rect 71096 14424 71102 14476
rect 71148 14464 71176 14504
rect 71498 14492 71504 14544
rect 71556 14532 71562 14544
rect 72436 14532 72464 14572
rect 75822 14560 75828 14612
rect 75880 14600 75886 14612
rect 77110 14600 77116 14612
rect 75880 14572 77116 14600
rect 75880 14560 75886 14572
rect 77110 14560 77116 14572
rect 77168 14600 77174 14612
rect 77662 14600 77668 14612
rect 77168 14572 77668 14600
rect 77168 14560 77174 14572
rect 77662 14560 77668 14572
rect 77720 14560 77726 14612
rect 78490 14560 78496 14612
rect 78548 14600 78554 14612
rect 81253 14603 81311 14609
rect 81253 14600 81265 14603
rect 78548 14572 81265 14600
rect 78548 14560 78554 14572
rect 81253 14569 81265 14572
rect 81299 14569 81311 14603
rect 92658 14600 92664 14612
rect 92619 14572 92664 14600
rect 81253 14563 81311 14569
rect 92658 14560 92664 14572
rect 92716 14560 92722 14612
rect 77386 14532 77392 14544
rect 71556 14504 71601 14532
rect 72436 14504 77392 14532
rect 71556 14492 71562 14504
rect 77386 14492 77392 14504
rect 77444 14492 77450 14544
rect 83829 14535 83887 14541
rect 83829 14501 83841 14535
rect 83875 14532 83887 14535
rect 88518 14532 88524 14544
rect 83875 14504 88524 14532
rect 83875 14501 83887 14504
rect 83829 14495 83887 14501
rect 88518 14492 88524 14504
rect 88576 14492 88582 14544
rect 76929 14467 76987 14473
rect 76929 14464 76941 14467
rect 71148 14436 76941 14464
rect 76929 14433 76941 14436
rect 76975 14433 76987 14467
rect 78582 14464 78588 14476
rect 76929 14427 76987 14433
rect 77036 14436 78588 14464
rect 65245 14399 65303 14405
rect 65245 14365 65257 14399
rect 65291 14365 65303 14399
rect 65245 14359 65303 14365
rect 65426 14356 65432 14408
rect 65484 14396 65490 14408
rect 65978 14396 65984 14408
rect 65484 14368 65984 14396
rect 65484 14356 65490 14368
rect 65978 14356 65984 14368
rect 66036 14356 66042 14408
rect 66070 14356 66076 14408
rect 66128 14396 66134 14408
rect 66530 14396 66536 14408
rect 66128 14368 66536 14396
rect 66128 14356 66134 14368
rect 66530 14356 66536 14368
rect 66588 14356 66594 14408
rect 66625 14399 66683 14405
rect 66625 14365 66637 14399
rect 66671 14396 66683 14399
rect 67266 14396 67272 14408
rect 66671 14368 67272 14396
rect 66671 14365 66683 14368
rect 66625 14359 66683 14365
rect 67266 14356 67272 14368
rect 67324 14356 67330 14408
rect 67726 14396 67732 14408
rect 67687 14368 67732 14396
rect 67726 14356 67732 14368
rect 67784 14356 67790 14408
rect 68186 14396 68192 14408
rect 68147 14368 68192 14396
rect 68186 14356 68192 14368
rect 68244 14356 68250 14408
rect 70946 14356 70952 14408
rect 71004 14396 71010 14408
rect 71133 14399 71191 14405
rect 71133 14396 71145 14399
rect 71004 14368 71145 14396
rect 71004 14356 71010 14368
rect 71133 14365 71145 14368
rect 71179 14365 71191 14399
rect 71133 14359 71191 14365
rect 72145 14399 72203 14405
rect 72145 14365 72157 14399
rect 72191 14396 72203 14399
rect 73522 14396 73528 14408
rect 72191 14368 73528 14396
rect 72191 14365 72203 14368
rect 72145 14359 72203 14365
rect 73522 14356 73528 14368
rect 73580 14356 73586 14408
rect 74810 14356 74816 14408
rect 74868 14396 74874 14408
rect 77036 14396 77064 14436
rect 78582 14424 78588 14436
rect 78640 14424 78646 14476
rect 78953 14467 79011 14473
rect 78953 14433 78965 14467
rect 78999 14464 79011 14467
rect 80330 14464 80336 14476
rect 78999 14436 80336 14464
rect 78999 14433 79011 14436
rect 78953 14427 79011 14433
rect 80330 14424 80336 14436
rect 80388 14424 80394 14476
rect 80606 14424 80612 14476
rect 80664 14464 80670 14476
rect 83553 14467 83611 14473
rect 80664 14436 83504 14464
rect 80664 14424 80670 14436
rect 83476 14408 83504 14436
rect 83553 14433 83565 14467
rect 83599 14464 83611 14467
rect 84102 14464 84108 14476
rect 83599 14436 84108 14464
rect 83599 14433 83611 14436
rect 83553 14427 83611 14433
rect 84102 14424 84108 14436
rect 84160 14424 84166 14476
rect 88429 14467 88487 14473
rect 88429 14464 88441 14467
rect 86788 14436 88441 14464
rect 86788 14408 86816 14436
rect 88429 14433 88441 14436
rect 88475 14433 88487 14467
rect 88429 14427 88487 14433
rect 79594 14396 79600 14408
rect 74868 14368 77064 14396
rect 79555 14368 79600 14396
rect 74868 14356 74874 14368
rect 79594 14356 79600 14368
rect 79652 14396 79658 14408
rect 80057 14399 80115 14405
rect 80057 14396 80069 14399
rect 79652 14368 80069 14396
rect 79652 14356 79658 14368
rect 80057 14365 80069 14368
rect 80103 14365 80115 14399
rect 80057 14359 80115 14365
rect 81802 14356 81808 14408
rect 81860 14396 81866 14408
rect 82357 14399 82415 14405
rect 82357 14396 82369 14399
rect 81860 14368 82369 14396
rect 81860 14356 81866 14368
rect 82357 14365 82369 14368
rect 82403 14365 82415 14399
rect 83458 14396 83464 14408
rect 83419 14368 83464 14396
rect 82357 14359 82415 14365
rect 83458 14356 83464 14368
rect 83516 14356 83522 14408
rect 84930 14396 84936 14408
rect 84891 14368 84936 14396
rect 84930 14356 84936 14368
rect 84988 14356 84994 14408
rect 86770 14396 86776 14408
rect 86731 14368 86776 14396
rect 86770 14356 86776 14368
rect 86828 14356 86834 14408
rect 86954 14356 86960 14408
rect 87012 14396 87018 14408
rect 87049 14399 87107 14405
rect 87049 14396 87061 14399
rect 87012 14368 87061 14396
rect 87012 14356 87018 14368
rect 87049 14365 87061 14368
rect 87095 14365 87107 14399
rect 87049 14359 87107 14365
rect 88242 14356 88248 14408
rect 88300 14396 88306 14408
rect 88521 14399 88579 14405
rect 88521 14396 88533 14399
rect 88300 14368 88533 14396
rect 88300 14356 88306 14368
rect 88521 14365 88533 14368
rect 88567 14365 88579 14399
rect 89346 14396 89352 14408
rect 89307 14368 89352 14396
rect 88521 14359 88579 14365
rect 89346 14356 89352 14368
rect 89404 14356 89410 14408
rect 61654 14288 61660 14340
rect 61712 14288 61718 14340
rect 62393 14331 62451 14337
rect 62393 14297 62405 14331
rect 62439 14328 62451 14331
rect 67637 14331 67695 14337
rect 67637 14328 67649 14331
rect 62439 14300 67649 14328
rect 62439 14297 62451 14300
rect 62393 14291 62451 14297
rect 67637 14297 67649 14300
rect 67683 14297 67695 14331
rect 68462 14328 68468 14340
rect 68423 14300 68468 14328
rect 67637 14291 67695 14297
rect 68462 14288 68468 14300
rect 68520 14288 68526 14340
rect 71038 14328 71044 14340
rect 69690 14300 71044 14328
rect 71038 14288 71044 14300
rect 71096 14288 71102 14340
rect 71866 14288 71872 14340
rect 71924 14328 71930 14340
rect 72697 14331 72755 14337
rect 72697 14328 72709 14331
rect 71924 14300 72709 14328
rect 71924 14288 71930 14300
rect 72697 14297 72709 14300
rect 72743 14297 72755 14331
rect 76926 14328 76932 14340
rect 72697 14291 72755 14297
rect 73816 14300 76932 14328
rect 63218 14260 63224 14272
rect 60660 14232 63224 14260
rect 63218 14220 63224 14232
rect 63276 14220 63282 14272
rect 63678 14260 63684 14272
rect 63639 14232 63684 14260
rect 63678 14220 63684 14232
rect 63736 14220 63742 14272
rect 64230 14260 64236 14272
rect 64191 14232 64236 14260
rect 64230 14220 64236 14232
rect 64288 14220 64294 14272
rect 65150 14260 65156 14272
rect 65111 14232 65156 14260
rect 65150 14220 65156 14232
rect 65208 14220 65214 14272
rect 65886 14260 65892 14272
rect 65847 14232 65892 14260
rect 65886 14220 65892 14232
rect 65944 14220 65950 14272
rect 65978 14220 65984 14272
rect 66036 14260 66042 14272
rect 69290 14260 69296 14272
rect 66036 14232 69296 14260
rect 66036 14220 66042 14232
rect 69290 14220 69296 14232
rect 69348 14220 69354 14272
rect 69934 14260 69940 14272
rect 69895 14232 69940 14260
rect 69934 14220 69940 14232
rect 69992 14220 69998 14272
rect 72050 14260 72056 14272
rect 72011 14232 72056 14260
rect 72050 14220 72056 14232
rect 72108 14220 72114 14272
rect 72326 14220 72332 14272
rect 72384 14260 72390 14272
rect 73816 14260 73844 14300
rect 76926 14288 76932 14300
rect 76984 14288 76990 14340
rect 78214 14288 78220 14340
rect 78272 14288 78278 14340
rect 78398 14288 78404 14340
rect 78456 14328 78462 14340
rect 78677 14331 78735 14337
rect 78677 14328 78689 14331
rect 78456 14300 78689 14328
rect 78456 14288 78462 14300
rect 78677 14297 78689 14300
rect 78723 14297 78735 14331
rect 78677 14291 78735 14297
rect 79226 14288 79232 14340
rect 79284 14328 79290 14340
rect 82538 14328 82544 14340
rect 79284 14300 82544 14328
rect 79284 14288 79290 14300
rect 82538 14288 82544 14300
rect 82596 14288 82602 14340
rect 84381 14331 84439 14337
rect 84381 14297 84393 14331
rect 84427 14328 84439 14331
rect 85666 14328 85672 14340
rect 84427 14300 85672 14328
rect 84427 14297 84439 14300
rect 84381 14291 84439 14297
rect 85666 14288 85672 14300
rect 85724 14328 85730 14340
rect 89254 14328 89260 14340
rect 85724 14300 89116 14328
rect 89215 14300 89260 14328
rect 85724 14288 85730 14300
rect 73982 14260 73988 14272
rect 72384 14232 73844 14260
rect 73943 14232 73988 14260
rect 72384 14220 72390 14232
rect 73982 14220 73988 14232
rect 74040 14220 74046 14272
rect 74997 14263 75055 14269
rect 74997 14229 75009 14263
rect 75043 14260 75055 14263
rect 75086 14260 75092 14272
rect 75043 14232 75092 14260
rect 75043 14229 75055 14232
rect 74997 14223 75055 14229
rect 75086 14220 75092 14232
rect 75144 14220 75150 14272
rect 75178 14220 75184 14272
rect 75236 14260 75242 14272
rect 75549 14263 75607 14269
rect 75549 14260 75561 14263
rect 75236 14232 75561 14260
rect 75236 14220 75242 14232
rect 75549 14229 75561 14232
rect 75595 14260 75607 14263
rect 75914 14260 75920 14272
rect 75595 14232 75920 14260
rect 75595 14229 75607 14232
rect 75549 14223 75607 14229
rect 75914 14220 75920 14232
rect 75972 14220 75978 14272
rect 76190 14260 76196 14272
rect 76151 14232 76196 14260
rect 76190 14220 76196 14232
rect 76248 14220 76254 14272
rect 76944 14260 76972 14288
rect 78858 14260 78864 14272
rect 76944 14232 78864 14260
rect 78858 14220 78864 14232
rect 78916 14220 78922 14272
rect 79502 14260 79508 14272
rect 79463 14232 79508 14260
rect 79502 14220 79508 14232
rect 79560 14220 79566 14272
rect 80054 14220 80060 14272
rect 80112 14260 80118 14272
rect 80149 14263 80207 14269
rect 80149 14260 80161 14263
rect 80112 14232 80161 14260
rect 80112 14220 80118 14232
rect 80149 14229 80161 14232
rect 80195 14229 80207 14263
rect 80149 14223 80207 14229
rect 80606 14220 80612 14272
rect 80664 14260 80670 14272
rect 81342 14260 81348 14272
rect 80664 14232 81348 14260
rect 80664 14220 80670 14232
rect 81342 14220 81348 14232
rect 81400 14260 81406 14272
rect 81805 14263 81863 14269
rect 81805 14260 81817 14263
rect 81400 14232 81817 14260
rect 81400 14220 81406 14232
rect 81805 14229 81817 14232
rect 81851 14229 81863 14263
rect 85022 14260 85028 14272
rect 84983 14232 85028 14260
rect 81805 14223 81863 14229
rect 85022 14220 85028 14232
rect 85080 14220 85086 14272
rect 85577 14263 85635 14269
rect 85577 14229 85589 14263
rect 85623 14260 85635 14263
rect 85850 14260 85856 14272
rect 85623 14232 85856 14260
rect 85623 14229 85635 14232
rect 85577 14223 85635 14229
rect 85850 14220 85856 14232
rect 85908 14220 85914 14272
rect 86402 14260 86408 14272
rect 86363 14232 86408 14260
rect 86402 14220 86408 14232
rect 86460 14220 86466 14272
rect 88150 14260 88156 14272
rect 88111 14232 88156 14260
rect 88150 14220 88156 14232
rect 88208 14220 88214 14272
rect 89088 14260 89116 14300
rect 89254 14288 89260 14300
rect 89312 14288 89318 14340
rect 89530 14260 89536 14272
rect 89088 14232 89536 14260
rect 89530 14220 89536 14232
rect 89588 14260 89594 14272
rect 89993 14263 90051 14269
rect 89993 14260 90005 14263
rect 89588 14232 90005 14260
rect 89588 14220 89594 14232
rect 89993 14229 90005 14232
rect 90039 14260 90051 14263
rect 90545 14263 90603 14269
rect 90545 14260 90557 14263
rect 90039 14232 90557 14260
rect 90039 14229 90051 14232
rect 89993 14223 90051 14229
rect 90545 14229 90557 14232
rect 90591 14229 90603 14263
rect 90545 14223 90603 14229
rect 91094 14220 91100 14272
rect 91152 14260 91158 14272
rect 91557 14263 91615 14269
rect 91557 14260 91569 14263
rect 91152 14232 91569 14260
rect 91152 14220 91158 14232
rect 91557 14229 91569 14232
rect 91603 14229 91615 14263
rect 91557 14223 91615 14229
rect 92201 14263 92259 14269
rect 92201 14229 92213 14263
rect 92247 14260 92259 14263
rect 92474 14260 92480 14272
rect 92247 14232 92480 14260
rect 92247 14229 92259 14232
rect 92201 14223 92259 14229
rect 92474 14220 92480 14232
rect 92532 14220 92538 14272
rect 1104 14170 95011 14192
rect 1104 14118 24386 14170
rect 24438 14118 24450 14170
rect 24502 14118 24514 14170
rect 24566 14118 24578 14170
rect 24630 14118 24642 14170
rect 24694 14118 47823 14170
rect 47875 14118 47887 14170
rect 47939 14118 47951 14170
rect 48003 14118 48015 14170
rect 48067 14118 48079 14170
rect 48131 14118 71260 14170
rect 71312 14118 71324 14170
rect 71376 14118 71388 14170
rect 71440 14118 71452 14170
rect 71504 14118 71516 14170
rect 71568 14118 94697 14170
rect 94749 14118 94761 14170
rect 94813 14118 94825 14170
rect 94877 14118 94889 14170
rect 94941 14118 94953 14170
rect 95005 14118 95011 14170
rect 1104 14096 95011 14118
rect 9122 14016 9128 14068
rect 9180 14056 9186 14068
rect 20438 14056 20444 14068
rect 9180 14028 20444 14056
rect 9180 14016 9186 14028
rect 20438 14016 20444 14028
rect 20496 14016 20502 14068
rect 20533 14059 20591 14065
rect 20533 14025 20545 14059
rect 20579 14056 20591 14059
rect 22465 14059 22523 14065
rect 20579 14028 22094 14056
rect 20579 14025 20591 14028
rect 20533 14019 20591 14025
rect 7745 13991 7803 13997
rect 7745 13957 7757 13991
rect 7791 13988 7803 13991
rect 8018 13988 8024 14000
rect 7791 13960 8024 13988
rect 7791 13957 7803 13960
rect 7745 13951 7803 13957
rect 8018 13948 8024 13960
rect 8076 13988 8082 14000
rect 9306 13988 9312 14000
rect 8076 13960 8616 13988
rect 9219 13960 9312 13988
rect 8076 13948 8082 13960
rect 2958 13920 2964 13932
rect 2919 13892 2964 13920
rect 2958 13880 2964 13892
rect 3016 13880 3022 13932
rect 3881 13923 3939 13929
rect 3881 13889 3893 13923
rect 3927 13920 3939 13923
rect 4154 13920 4160 13932
rect 3927 13892 4160 13920
rect 3927 13889 3939 13892
rect 3881 13883 3939 13889
rect 4154 13880 4160 13892
rect 4212 13880 4218 13932
rect 7282 13880 7288 13932
rect 7340 13920 7346 13932
rect 8588 13929 8616 13960
rect 9306 13948 9312 13960
rect 9364 13988 9370 14000
rect 16206 13988 16212 14000
rect 9364 13960 16212 13988
rect 9364 13948 9370 13960
rect 8573 13923 8631 13929
rect 7340 13892 8524 13920
rect 7340 13880 7346 13892
rect 8202 13852 8208 13864
rect 8163 13824 8208 13852
rect 8202 13812 8208 13824
rect 8260 13812 8266 13864
rect 8496 13861 8524 13892
rect 8573 13889 8585 13923
rect 8619 13920 8631 13923
rect 11885 13923 11943 13929
rect 8619 13892 11192 13920
rect 8619 13889 8631 13892
rect 8573 13883 8631 13889
rect 11164 13861 11192 13892
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 12434 13920 12440 13932
rect 11931 13892 12440 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 12434 13880 12440 13892
rect 12492 13880 12498 13932
rect 13265 13923 13323 13929
rect 13265 13889 13277 13923
rect 13311 13920 13323 13923
rect 13906 13920 13912 13932
rect 13311 13892 13912 13920
rect 13311 13889 13323 13892
rect 13265 13883 13323 13889
rect 13906 13880 13912 13892
rect 13964 13880 13970 13932
rect 14936 13929 14964 13960
rect 16206 13948 16212 13960
rect 16264 13948 16270 14000
rect 16942 13988 16948 14000
rect 16903 13960 16948 13988
rect 16942 13948 16948 13960
rect 17000 13948 17006 14000
rect 20070 13948 20076 14000
rect 20128 13948 20134 14000
rect 22066 13988 22094 14028
rect 22465 14025 22477 14059
rect 22511 14056 22523 14059
rect 22646 14056 22652 14068
rect 22511 14028 22652 14056
rect 22511 14025 22523 14028
rect 22465 14019 22523 14025
rect 22646 14016 22652 14028
rect 22704 14016 22710 14068
rect 25682 14056 25688 14068
rect 23768 14028 25688 14056
rect 23658 13988 23664 14000
rect 20548 13960 21404 13988
rect 22066 13960 23664 13988
rect 14921 13923 14979 13929
rect 14921 13889 14933 13923
rect 14967 13889 14979 13923
rect 14921 13883 14979 13889
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 15933 13923 15991 13929
rect 15933 13920 15945 13923
rect 15160 13892 15945 13920
rect 15160 13880 15166 13892
rect 15933 13889 15945 13892
rect 15979 13889 15991 13923
rect 15933 13883 15991 13889
rect 8481 13855 8539 13861
rect 8481 13821 8493 13855
rect 8527 13821 8539 13855
rect 8481 13815 8539 13821
rect 11149 13855 11207 13861
rect 11149 13821 11161 13855
rect 11195 13852 11207 13855
rect 11974 13852 11980 13864
rect 11195 13824 11980 13852
rect 11195 13821 11207 13824
rect 11149 13815 11207 13821
rect 11974 13812 11980 13824
rect 12032 13812 12038 13864
rect 13998 13852 14004 13864
rect 13959 13824 14004 13852
rect 13998 13812 14004 13824
rect 14056 13812 14062 13864
rect 14458 13812 14464 13864
rect 14516 13852 14522 13864
rect 15010 13852 15016 13864
rect 14516 13824 15016 13852
rect 14516 13812 14522 13824
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 15838 13852 15844 13864
rect 15799 13824 15844 13852
rect 15838 13812 15844 13824
rect 15896 13812 15902 13864
rect 18785 13855 18843 13861
rect 18785 13852 18797 13855
rect 17052 13824 18797 13852
rect 12253 13787 12311 13793
rect 12253 13753 12265 13787
rect 12299 13784 12311 13787
rect 14277 13787 14335 13793
rect 12299 13756 13308 13784
rect 12299 13753 12311 13756
rect 12253 13747 12311 13753
rect 4798 13716 4804 13728
rect 4759 13688 4804 13716
rect 4798 13676 4804 13688
rect 4856 13676 4862 13728
rect 6641 13719 6699 13725
rect 6641 13685 6653 13719
rect 6687 13716 6699 13719
rect 6822 13716 6828 13728
rect 6687 13688 6828 13716
rect 6687 13685 6699 13688
rect 6641 13679 6699 13685
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 10134 13676 10140 13728
rect 10192 13716 10198 13728
rect 11330 13716 11336 13728
rect 10192 13688 11336 13716
rect 10192 13676 10198 13688
rect 11330 13676 11336 13688
rect 11388 13676 11394 13728
rect 13280 13716 13308 13756
rect 14277 13753 14289 13787
rect 14323 13784 14335 13787
rect 15194 13784 15200 13796
rect 14323 13756 15200 13784
rect 14323 13753 14335 13756
rect 14277 13747 14335 13753
rect 15194 13744 15200 13756
rect 15252 13744 15258 13796
rect 15289 13787 15347 13793
rect 15289 13753 15301 13787
rect 15335 13784 15347 13787
rect 17052 13784 17080 13824
rect 18785 13821 18797 13824
rect 18831 13821 18843 13855
rect 18785 13815 18843 13821
rect 19061 13855 19119 13861
rect 19061 13821 19073 13855
rect 19107 13852 19119 13855
rect 20548 13852 20576 13960
rect 21266 13920 21272 13932
rect 21227 13892 21272 13920
rect 21266 13880 21272 13892
rect 21324 13880 21330 13932
rect 21376 13920 21404 13960
rect 23658 13948 23664 13960
rect 23716 13948 23722 14000
rect 23768 13997 23796 14028
rect 25682 14016 25688 14028
rect 25740 14016 25746 14068
rect 26142 14016 26148 14068
rect 26200 14016 26206 14068
rect 27709 14059 27767 14065
rect 27709 14025 27721 14059
rect 27755 14056 27767 14059
rect 30282 14056 30288 14068
rect 27755 14028 30288 14056
rect 27755 14025 27767 14028
rect 27709 14019 27767 14025
rect 30282 14016 30288 14028
rect 30340 14016 30346 14068
rect 37366 14016 37372 14068
rect 37424 14056 37430 14068
rect 41414 14056 41420 14068
rect 37424 14028 41420 14056
rect 37424 14016 37430 14028
rect 41414 14016 41420 14028
rect 41472 14016 41478 14068
rect 47210 14056 47216 14068
rect 41524 14028 44588 14056
rect 47171 14028 47216 14056
rect 23753 13991 23811 13997
rect 23753 13957 23765 13991
rect 23799 13957 23811 13991
rect 23753 13951 23811 13957
rect 24302 13948 24308 14000
rect 24360 13988 24366 14000
rect 24581 13991 24639 13997
rect 24581 13988 24593 13991
rect 24360 13960 24593 13988
rect 24360 13948 24366 13960
rect 24581 13957 24593 13960
rect 24627 13957 24639 13991
rect 24581 13951 24639 13957
rect 25590 13948 25596 14000
rect 25648 13948 25654 14000
rect 26160 13988 26188 14016
rect 30190 13988 30196 14000
rect 26160 13960 27660 13988
rect 29394 13960 30196 13988
rect 25038 13920 25044 13932
rect 21376 13892 25044 13920
rect 25038 13880 25044 13892
rect 25096 13880 25102 13932
rect 27632 13929 27660 13960
rect 30190 13948 30196 13960
rect 30248 13948 30254 14000
rect 32398 13948 32404 14000
rect 32456 13988 32462 14000
rect 34238 13988 34244 14000
rect 32456 13960 34244 13988
rect 32456 13948 32462 13960
rect 27617 13923 27675 13929
rect 27617 13889 27629 13923
rect 27663 13920 27675 13923
rect 27890 13920 27896 13932
rect 27663 13892 27896 13920
rect 27663 13889 27675 13892
rect 27617 13883 27675 13889
rect 27890 13880 27896 13892
rect 27948 13880 27954 13932
rect 30098 13880 30104 13932
rect 30156 13920 30162 13932
rect 30837 13923 30895 13929
rect 30156 13892 30201 13920
rect 30156 13880 30162 13892
rect 30837 13889 30849 13923
rect 30883 13920 30895 13923
rect 31478 13920 31484 13932
rect 30883 13892 31484 13920
rect 30883 13889 30895 13892
rect 30837 13883 30895 13889
rect 31478 13880 31484 13892
rect 31536 13880 31542 13932
rect 31754 13920 31760 13932
rect 31715 13892 31760 13920
rect 31754 13880 31760 13892
rect 31812 13880 31818 13932
rect 32493 13923 32551 13929
rect 32493 13889 32505 13923
rect 32539 13920 32551 13923
rect 32582 13920 32588 13932
rect 32539 13892 32588 13920
rect 32539 13889 32551 13892
rect 32493 13883 32551 13889
rect 32582 13880 32588 13892
rect 32640 13880 32646 13932
rect 33152 13929 33180 13960
rect 34238 13948 34244 13960
rect 34296 13948 34302 14000
rect 35434 13988 35440 14000
rect 35395 13960 35440 13988
rect 35434 13948 35440 13960
rect 35492 13948 35498 14000
rect 35618 13948 35624 14000
rect 35676 13988 35682 14000
rect 36722 13988 36728 14000
rect 35676 13960 36728 13988
rect 35676 13948 35682 13960
rect 36722 13948 36728 13960
rect 36780 13948 36786 14000
rect 38562 13988 38568 14000
rect 37752 13960 38568 13988
rect 33137 13923 33195 13929
rect 33137 13889 33149 13923
rect 33183 13889 33195 13923
rect 33137 13883 33195 13889
rect 36357 13923 36415 13929
rect 36357 13889 36369 13923
rect 36403 13920 36415 13923
rect 37458 13920 37464 13932
rect 36403 13892 37464 13920
rect 36403 13889 36415 13892
rect 36357 13883 36415 13889
rect 37458 13880 37464 13892
rect 37516 13880 37522 13932
rect 19107 13824 20576 13852
rect 21361 13855 21419 13861
rect 19107 13821 19119 13824
rect 19061 13815 19119 13821
rect 21361 13821 21373 13855
rect 21407 13852 21419 13855
rect 22186 13852 22192 13864
rect 21407 13824 22192 13852
rect 21407 13821 21419 13824
rect 21361 13815 21419 13821
rect 22186 13812 22192 13824
rect 22244 13812 22250 13864
rect 22554 13812 22560 13864
rect 22612 13852 22618 13864
rect 25958 13852 25964 13864
rect 22612 13824 25964 13852
rect 22612 13812 22618 13824
rect 25958 13812 25964 13824
rect 26016 13812 26022 13864
rect 26329 13855 26387 13861
rect 26329 13821 26341 13855
rect 26375 13852 26387 13855
rect 26605 13855 26663 13861
rect 26375 13824 26556 13852
rect 26375 13821 26387 13824
rect 26329 13815 26387 13821
rect 15335 13756 17080 13784
rect 15335 13753 15347 13756
rect 15289 13747 15347 13753
rect 20070 13744 20076 13796
rect 20128 13784 20134 13796
rect 25314 13784 25320 13796
rect 20128 13756 25320 13784
rect 20128 13744 20134 13756
rect 25314 13744 25320 13756
rect 25372 13744 25378 13796
rect 26528 13784 26556 13824
rect 26605 13821 26617 13855
rect 26651 13852 26663 13855
rect 28258 13852 28264 13864
rect 26651 13824 28264 13852
rect 26651 13821 26663 13824
rect 26605 13815 26663 13821
rect 28258 13812 28264 13824
rect 28316 13812 28322 13864
rect 28353 13855 28411 13861
rect 28353 13821 28365 13855
rect 28399 13852 28411 13855
rect 29822 13852 29828 13864
rect 28399 13824 29828 13852
rect 28399 13821 28411 13824
rect 28353 13815 28411 13821
rect 29822 13812 29828 13824
rect 29880 13812 29886 13864
rect 30742 13852 30748 13864
rect 30392 13824 30748 13852
rect 30190 13784 30196 13796
rect 26528 13756 28856 13784
rect 15746 13716 15752 13728
rect 13280 13688 15752 13716
rect 15746 13676 15752 13688
rect 15804 13676 15810 13728
rect 17402 13716 17408 13728
rect 17363 13688 17408 13716
rect 17402 13676 17408 13688
rect 17460 13676 17466 13728
rect 17494 13676 17500 13728
rect 17552 13716 17558 13728
rect 19610 13716 19616 13728
rect 17552 13688 19616 13716
rect 17552 13676 17558 13688
rect 19610 13676 19616 13688
rect 19668 13676 19674 13728
rect 19702 13676 19708 13728
rect 19760 13716 19766 13728
rect 28534 13716 28540 13728
rect 19760 13688 28540 13716
rect 19760 13676 19766 13688
rect 28534 13676 28540 13688
rect 28592 13676 28598 13728
rect 28828 13716 28856 13756
rect 30024 13756 30196 13784
rect 29638 13716 29644 13728
rect 28828 13688 29644 13716
rect 29638 13676 29644 13688
rect 29696 13676 29702 13728
rect 29843 13719 29901 13725
rect 29843 13685 29855 13719
rect 29889 13716 29901 13719
rect 30024 13716 30052 13756
rect 30190 13744 30196 13756
rect 30248 13744 30254 13796
rect 29889 13688 30052 13716
rect 29889 13685 29901 13688
rect 29843 13679 29901 13685
rect 30098 13676 30104 13728
rect 30156 13716 30162 13728
rect 30392 13716 30420 13824
rect 30742 13812 30748 13824
rect 30800 13812 30806 13864
rect 30926 13812 30932 13864
rect 30984 13852 30990 13864
rect 32401 13855 32459 13861
rect 32401 13852 32413 13855
rect 30984 13824 32413 13852
rect 30984 13812 30990 13824
rect 32401 13821 32413 13824
rect 32447 13821 32459 13855
rect 33962 13852 33968 13864
rect 33923 13824 33968 13852
rect 32401 13815 32459 13821
rect 33962 13812 33968 13824
rect 34020 13812 34026 13864
rect 34054 13812 34060 13864
rect 34112 13852 34118 13864
rect 35066 13852 35072 13864
rect 34112 13824 35072 13852
rect 34112 13812 34118 13824
rect 35066 13812 35072 13824
rect 35124 13852 35130 13864
rect 35621 13855 35679 13861
rect 35621 13852 35633 13855
rect 35124 13824 35633 13852
rect 35124 13812 35130 13824
rect 35621 13821 35633 13824
rect 35667 13821 35679 13855
rect 35621 13815 35679 13821
rect 36909 13855 36967 13861
rect 36909 13821 36921 13855
rect 36955 13852 36967 13855
rect 37274 13852 37280 13864
rect 36955 13824 37280 13852
rect 36955 13821 36967 13824
rect 36909 13815 36967 13821
rect 37274 13812 37280 13824
rect 37332 13852 37338 13864
rect 37752 13861 37780 13960
rect 38562 13948 38568 13960
rect 38620 13988 38626 14000
rect 38620 13960 38976 13988
rect 38620 13948 38626 13960
rect 38470 13920 38476 13932
rect 38431 13892 38476 13920
rect 38470 13880 38476 13892
rect 38528 13880 38534 13932
rect 38948 13929 38976 13960
rect 39114 13948 39120 14000
rect 39172 13988 39178 14000
rect 39209 13991 39267 13997
rect 39209 13988 39221 13991
rect 39172 13960 39221 13988
rect 39172 13948 39178 13960
rect 39209 13957 39221 13960
rect 39255 13957 39267 13991
rect 39209 13951 39267 13957
rect 40218 13948 40224 14000
rect 40276 13948 40282 14000
rect 40494 13948 40500 14000
rect 40552 13988 40558 14000
rect 41524 13988 41552 14028
rect 43717 13991 43775 13997
rect 40552 13960 41552 13988
rect 41616 13960 42564 13988
rect 40552 13948 40558 13960
rect 38933 13923 38991 13929
rect 38933 13889 38945 13923
rect 38979 13889 38991 13923
rect 40954 13920 40960 13932
rect 40915 13892 40960 13920
rect 38933 13883 38991 13889
rect 40954 13880 40960 13892
rect 41012 13920 41018 13932
rect 41616 13920 41644 13960
rect 41012 13892 41644 13920
rect 41679 13923 41737 13929
rect 41012 13880 41018 13892
rect 41679 13889 41691 13923
rect 41725 13920 41737 13923
rect 41782 13920 41788 13932
rect 41725 13892 41788 13920
rect 41725 13889 41737 13892
rect 41679 13883 41737 13889
rect 41782 13880 41788 13892
rect 41840 13920 41846 13932
rect 42426 13920 42432 13932
rect 41840 13892 42432 13920
rect 41840 13880 41846 13892
rect 42426 13880 42432 13892
rect 42484 13880 42490 13932
rect 42536 13920 42564 13960
rect 43717 13957 43729 13991
rect 43763 13988 43775 13991
rect 44082 13988 44088 14000
rect 43763 13960 44088 13988
rect 43763 13957 43775 13960
rect 43717 13951 43775 13957
rect 44082 13948 44088 13960
rect 44140 13948 44146 14000
rect 42705 13923 42763 13929
rect 42705 13920 42717 13923
rect 42536 13892 42717 13920
rect 42705 13889 42717 13892
rect 42751 13889 42763 13923
rect 42705 13883 42763 13889
rect 42794 13880 42800 13932
rect 42852 13920 42858 13932
rect 44560 13929 44588 14028
rect 47210 14016 47216 14028
rect 47268 14016 47274 14068
rect 47302 14016 47308 14068
rect 47360 14056 47366 14068
rect 47360 14028 55536 14056
rect 47360 14016 47366 14028
rect 45646 13988 45652 14000
rect 45480 13960 45652 13988
rect 45480 13929 45508 13960
rect 45646 13948 45652 13960
rect 45704 13948 45710 14000
rect 46474 13948 46480 14000
rect 46532 13948 46538 14000
rect 48314 13988 48320 14000
rect 47780 13960 48320 13988
rect 47780 13929 47808 13960
rect 48314 13948 48320 13960
rect 48372 13948 48378 14000
rect 48774 13948 48780 14000
rect 48832 13948 48838 14000
rect 49510 13948 49516 14000
rect 49568 13988 49574 14000
rect 49973 13991 50031 13997
rect 49973 13988 49985 13991
rect 49568 13960 49985 13988
rect 49568 13948 49574 13960
rect 49973 13957 49985 13960
rect 50019 13957 50031 13991
rect 49973 13951 50031 13957
rect 50062 13948 50068 14000
rect 50120 13988 50126 14000
rect 51077 13991 51135 13997
rect 51077 13988 51089 13991
rect 50120 13960 51089 13988
rect 50120 13948 50126 13960
rect 51077 13957 51089 13960
rect 51123 13957 51135 13991
rect 51077 13951 51135 13957
rect 53009 13991 53067 13997
rect 53009 13957 53021 13991
rect 53055 13988 53067 13991
rect 53055 13960 55444 13988
rect 53055 13957 53067 13960
rect 53009 13951 53067 13957
rect 42889 13923 42947 13929
rect 42889 13920 42901 13923
rect 42852 13892 42901 13920
rect 42852 13880 42858 13892
rect 42889 13889 42901 13892
rect 42935 13889 42947 13923
rect 42889 13883 42947 13889
rect 44545 13923 44603 13929
rect 44545 13889 44557 13923
rect 44591 13889 44603 13923
rect 44545 13883 44603 13889
rect 45465 13923 45523 13929
rect 45465 13889 45477 13923
rect 45511 13889 45523 13923
rect 45465 13883 45523 13889
rect 47765 13923 47823 13929
rect 47765 13889 47777 13923
rect 47811 13889 47823 13923
rect 47765 13883 47823 13889
rect 49326 13880 49332 13932
rect 49384 13920 49390 13932
rect 52362 13920 52368 13932
rect 49384 13892 52368 13920
rect 49384 13880 49390 13892
rect 52362 13880 52368 13892
rect 52420 13880 52426 13932
rect 52917 13923 52975 13929
rect 52917 13889 52929 13923
rect 52963 13920 52975 13923
rect 53558 13920 53564 13932
rect 52963 13892 53564 13920
rect 52963 13889 52975 13892
rect 52917 13883 52975 13889
rect 53558 13880 53564 13892
rect 53616 13880 53622 13932
rect 53742 13920 53748 13932
rect 53703 13892 53748 13920
rect 53742 13880 53748 13892
rect 53800 13880 53806 13932
rect 54938 13920 54944 13932
rect 54036 13892 54944 13920
rect 37737 13855 37795 13861
rect 37737 13852 37749 13855
rect 37332 13824 37749 13852
rect 37332 13812 37338 13824
rect 37737 13821 37749 13824
rect 37783 13821 37795 13855
rect 37737 13815 37795 13821
rect 38194 13812 38200 13864
rect 38252 13852 38258 13864
rect 38381 13855 38439 13861
rect 38381 13852 38393 13855
rect 38252 13824 38393 13852
rect 38252 13812 38258 13824
rect 38381 13821 38393 13824
rect 38427 13821 38439 13855
rect 38381 13815 38439 13821
rect 41601 13855 41659 13861
rect 41601 13821 41613 13855
rect 41647 13821 41659 13855
rect 44818 13852 44824 13864
rect 44779 13824 44824 13852
rect 41601 13815 41659 13821
rect 30466 13744 30472 13796
rect 30524 13784 30530 13796
rect 38654 13784 38660 13796
rect 30524 13756 38660 13784
rect 30524 13744 30530 13756
rect 38654 13744 38660 13756
rect 38712 13744 38718 13796
rect 30156 13688 30420 13716
rect 30156 13676 30162 13688
rect 30650 13676 30656 13728
rect 30708 13716 30714 13728
rect 30745 13719 30803 13725
rect 30745 13716 30757 13719
rect 30708 13688 30757 13716
rect 30708 13676 30714 13688
rect 30745 13685 30757 13688
rect 30791 13685 30803 13719
rect 30745 13679 30803 13685
rect 31018 13676 31024 13728
rect 31076 13716 31082 13728
rect 33134 13716 33140 13728
rect 31076 13688 33140 13716
rect 31076 13676 31082 13688
rect 33134 13676 33140 13688
rect 33192 13676 33198 13728
rect 33229 13719 33287 13725
rect 33229 13685 33241 13719
rect 33275 13716 33287 13719
rect 33318 13716 33324 13728
rect 33275 13688 33324 13716
rect 33275 13685 33287 13688
rect 33229 13679 33287 13685
rect 33318 13676 33324 13688
rect 33376 13676 33382 13728
rect 33410 13676 33416 13728
rect 33468 13716 33474 13728
rect 35986 13716 35992 13728
rect 33468 13688 35992 13716
rect 33468 13676 33474 13688
rect 35986 13676 35992 13688
rect 36044 13676 36050 13728
rect 36446 13676 36452 13728
rect 36504 13716 36510 13728
rect 38838 13716 38844 13728
rect 36504 13688 38844 13716
rect 36504 13676 36510 13688
rect 38838 13676 38844 13688
rect 38896 13676 38902 13728
rect 41616 13716 41644 13815
rect 44818 13812 44824 13824
rect 44876 13812 44882 13864
rect 45738 13852 45744 13864
rect 45699 13824 45744 13852
rect 45738 13812 45744 13824
rect 45796 13812 45802 13864
rect 46106 13812 46112 13864
rect 46164 13852 46170 13864
rect 49513 13855 49571 13861
rect 46164 13824 49464 13852
rect 46164 13812 46170 13824
rect 41969 13787 42027 13793
rect 41969 13753 41981 13787
rect 42015 13784 42027 13787
rect 49436 13784 49464 13824
rect 49513 13821 49525 13855
rect 49559 13852 49571 13855
rect 50338 13852 50344 13864
rect 49559 13824 50344 13852
rect 49559 13821 49571 13824
rect 49513 13815 49571 13821
rect 50338 13812 50344 13824
rect 50396 13812 50402 13864
rect 51442 13812 51448 13864
rect 51500 13852 51506 13864
rect 54036 13852 54064 13892
rect 54938 13880 54944 13892
rect 54996 13880 55002 13932
rect 55033 13923 55091 13929
rect 55033 13889 55045 13923
rect 55079 13920 55091 13923
rect 55306 13920 55312 13932
rect 55079 13892 55312 13920
rect 55079 13889 55091 13892
rect 55033 13883 55091 13889
rect 55306 13880 55312 13892
rect 55364 13880 55370 13932
rect 54202 13852 54208 13864
rect 51500 13824 54064 13852
rect 54163 13824 54208 13852
rect 51500 13812 51506 13824
rect 54202 13812 54208 13824
rect 54260 13812 54266 13864
rect 49786 13784 49792 13796
rect 42015 13756 44956 13784
rect 49436 13756 49792 13784
rect 42015 13753 42027 13756
rect 41969 13747 42027 13753
rect 42242 13716 42248 13728
rect 41616 13688 42248 13716
rect 42242 13676 42248 13688
rect 42300 13676 42306 13728
rect 44928 13716 44956 13756
rect 49786 13744 49792 13756
rect 49844 13744 49850 13796
rect 52270 13744 52276 13796
rect 52328 13784 52334 13796
rect 53834 13784 53840 13796
rect 52328 13756 53840 13784
rect 52328 13744 52334 13756
rect 53834 13744 53840 13756
rect 53892 13744 53898 13796
rect 48022 13719 48080 13725
rect 48022 13716 48034 13719
rect 44928 13688 48034 13716
rect 48022 13685 48034 13688
rect 48068 13685 48080 13719
rect 48022 13679 48080 13685
rect 48774 13676 48780 13728
rect 48832 13716 48838 13728
rect 49694 13716 49700 13728
rect 48832 13688 49700 13716
rect 48832 13676 48838 13688
rect 49694 13676 49700 13688
rect 49752 13676 49758 13728
rect 50430 13676 50436 13728
rect 50488 13716 50494 13728
rect 50525 13719 50583 13725
rect 50525 13716 50537 13719
rect 50488 13688 50537 13716
rect 50488 13676 50494 13688
rect 50525 13685 50537 13688
rect 50571 13685 50583 13719
rect 51626 13716 51632 13728
rect 51587 13688 51632 13716
rect 50525 13679 50583 13685
rect 51626 13676 51632 13688
rect 51684 13676 51690 13728
rect 52178 13716 52184 13728
rect 52139 13688 52184 13716
rect 52178 13676 52184 13688
rect 52236 13676 52242 13728
rect 53650 13716 53656 13728
rect 53611 13688 53656 13716
rect 53650 13676 53656 13688
rect 53708 13676 53714 13728
rect 55416 13716 55444 13960
rect 55508 13852 55536 14028
rect 55766 14016 55772 14068
rect 55824 14056 55830 14068
rect 58250 14056 58256 14068
rect 55824 14028 58112 14056
rect 58211 14028 58256 14056
rect 55824 14016 55830 14028
rect 56042 13948 56048 14000
rect 56100 13948 56106 14000
rect 56686 13948 56692 14000
rect 56744 13988 56750 14000
rect 57974 13988 57980 14000
rect 56744 13960 57980 13988
rect 56744 13948 56750 13960
rect 57974 13948 57980 13960
rect 58032 13948 58038 14000
rect 57057 13924 57115 13929
rect 57057 13923 57192 13924
rect 57057 13889 57069 13923
rect 57103 13920 57192 13923
rect 57330 13920 57336 13932
rect 57103 13896 57336 13920
rect 57103 13889 57115 13896
rect 57164 13892 57336 13896
rect 57057 13883 57115 13889
rect 57330 13880 57336 13892
rect 57388 13880 57394 13932
rect 58084 13929 58112 14028
rect 58250 14016 58256 14028
rect 58308 14016 58314 14068
rect 58342 14016 58348 14068
rect 58400 14056 58406 14068
rect 58400 14028 61240 14056
rect 58400 14016 58406 14028
rect 59262 13988 59268 14000
rect 59223 13960 59268 13988
rect 59262 13948 59268 13960
rect 59320 13948 59326 14000
rect 59998 13948 60004 14000
rect 60056 13948 60062 14000
rect 61013 13991 61071 13997
rect 61013 13957 61025 13991
rect 61059 13988 61071 13991
rect 61102 13988 61108 14000
rect 61059 13960 61108 13988
rect 61059 13957 61071 13960
rect 61013 13951 61071 13957
rect 61102 13948 61108 13960
rect 61160 13948 61166 14000
rect 61212 13988 61240 14028
rect 61654 14016 61660 14068
rect 61712 14056 61718 14068
rect 62206 14056 62212 14068
rect 61712 14028 62212 14056
rect 61712 14016 61718 14028
rect 62206 14016 62212 14028
rect 62264 14056 62270 14068
rect 67450 14056 67456 14068
rect 62264 14028 65840 14056
rect 67411 14028 67456 14056
rect 62264 14016 62270 14028
rect 62393 13991 62451 13997
rect 62393 13988 62405 13991
rect 61212 13960 62405 13988
rect 62393 13957 62405 13960
rect 62439 13988 62451 13991
rect 63862 13988 63868 14000
rect 62439 13960 63868 13988
rect 62439 13957 62451 13960
rect 62393 13951 62451 13957
rect 63862 13948 63868 13960
rect 63920 13948 63926 14000
rect 65150 13948 65156 14000
rect 65208 13948 65214 14000
rect 65812 13988 65840 14028
rect 67450 14016 67456 14028
rect 67508 14016 67514 14068
rect 74810 14056 74816 14068
rect 67606 14028 70394 14056
rect 74771 14028 74816 14056
rect 67606 13988 67634 14028
rect 65812 13960 67634 13988
rect 67726 13948 67732 14000
rect 67784 13988 67790 14000
rect 67784 13960 69336 13988
rect 67784 13948 67790 13960
rect 58069 13923 58127 13929
rect 58069 13889 58081 13923
rect 58115 13920 58127 13923
rect 59446 13920 59452 13932
rect 58115 13892 59452 13920
rect 58115 13889 58127 13892
rect 58069 13883 58127 13889
rect 59446 13880 59452 13892
rect 59504 13880 59510 13932
rect 61289 13923 61347 13929
rect 61289 13889 61301 13923
rect 61335 13920 61347 13923
rect 61470 13920 61476 13932
rect 61335 13892 61476 13920
rect 61335 13889 61347 13892
rect 61289 13883 61347 13889
rect 61470 13880 61476 13892
rect 61528 13920 61534 13932
rect 63589 13923 63647 13929
rect 61528 13892 62896 13920
rect 61528 13880 61534 13892
rect 56686 13852 56692 13864
rect 55508 13824 56692 13852
rect 56686 13812 56692 13824
rect 56744 13812 56750 13864
rect 57146 13812 57152 13864
rect 57204 13852 57210 13864
rect 57204 13824 57974 13852
rect 57204 13812 57210 13824
rect 57946 13784 57974 13824
rect 60458 13812 60464 13864
rect 60516 13852 60522 13864
rect 61562 13852 61568 13864
rect 60516 13824 61240 13852
rect 60516 13812 60522 13824
rect 58805 13787 58863 13793
rect 58805 13784 58817 13787
rect 57946 13756 58817 13784
rect 58805 13753 58817 13756
rect 58851 13784 58863 13787
rect 59998 13784 60004 13796
rect 58851 13756 60004 13784
rect 58851 13753 58863 13756
rect 58805 13747 58863 13753
rect 59998 13744 60004 13756
rect 60056 13744 60062 13796
rect 61212 13784 61240 13824
rect 61396 13824 61568 13852
rect 61396 13784 61424 13824
rect 61562 13812 61568 13824
rect 61620 13852 61626 13864
rect 61749 13855 61807 13861
rect 61749 13852 61761 13855
rect 61620 13824 61761 13852
rect 61620 13812 61626 13824
rect 61749 13821 61761 13824
rect 61795 13821 61807 13855
rect 62868 13852 62896 13892
rect 63589 13889 63601 13923
rect 63635 13920 63647 13923
rect 64598 13920 64604 13932
rect 63635 13892 64604 13920
rect 63635 13889 63647 13892
rect 63589 13883 63647 13889
rect 64598 13880 64604 13892
rect 64656 13880 64662 13932
rect 66530 13880 66536 13932
rect 66588 13920 66594 13932
rect 69308 13929 69336 13960
rect 68925 13923 68983 13929
rect 68925 13920 68937 13923
rect 66588 13892 68937 13920
rect 66588 13880 66594 13892
rect 68925 13889 68937 13892
rect 68971 13889 68983 13923
rect 68925 13883 68983 13889
rect 69293 13923 69351 13929
rect 69293 13889 69305 13923
rect 69339 13889 69351 13923
rect 69293 13883 69351 13889
rect 64049 13855 64107 13861
rect 64049 13852 64061 13855
rect 62868 13824 64061 13852
rect 61749 13815 61807 13821
rect 64049 13821 64061 13824
rect 64095 13852 64107 13855
rect 64230 13852 64236 13864
rect 64095 13824 64236 13852
rect 64095 13821 64107 13824
rect 64049 13815 64107 13821
rect 64230 13812 64236 13824
rect 64288 13812 64294 13864
rect 66441 13855 66499 13861
rect 66441 13852 66453 13855
rect 65168 13824 66453 13852
rect 65168 13784 65196 13824
rect 66441 13821 66453 13824
rect 66487 13821 66499 13855
rect 66441 13815 66499 13821
rect 66622 13812 66628 13864
rect 66680 13852 66686 13864
rect 66901 13855 66959 13861
rect 66901 13852 66913 13855
rect 66680 13824 66913 13852
rect 66680 13812 66686 13824
rect 66901 13821 66913 13824
rect 66947 13821 66959 13855
rect 70366 13852 70394 14028
rect 74810 14016 74816 14028
rect 74868 14016 74874 14068
rect 76193 14059 76251 14065
rect 76193 14025 76205 14059
rect 76239 14056 76251 14059
rect 78398 14056 78404 14068
rect 76239 14028 78404 14056
rect 76239 14025 76251 14028
rect 76193 14019 76251 14025
rect 78398 14016 78404 14028
rect 78456 14016 78462 14068
rect 78582 14016 78588 14068
rect 78640 14056 78646 14068
rect 80977 14059 81035 14065
rect 80977 14056 80989 14059
rect 78640 14028 80989 14056
rect 78640 14016 78646 14028
rect 80977 14025 80989 14028
rect 81023 14025 81035 14059
rect 80977 14019 81035 14025
rect 81342 14016 81348 14068
rect 81400 14056 81406 14068
rect 82633 14059 82691 14065
rect 82633 14056 82645 14059
rect 81400 14028 82645 14056
rect 81400 14016 81406 14028
rect 82633 14025 82645 14028
rect 82679 14025 82691 14059
rect 82633 14019 82691 14025
rect 83458 14016 83464 14068
rect 83516 14056 83522 14068
rect 83516 14028 86264 14056
rect 83516 14016 83522 14028
rect 71590 13948 71596 14000
rect 71648 13948 71654 14000
rect 73706 13948 73712 14000
rect 73764 13988 73770 14000
rect 75549 13991 75607 13997
rect 75549 13988 75561 13991
rect 73764 13960 75561 13988
rect 73764 13948 73770 13960
rect 75549 13957 75561 13960
rect 75595 13957 75607 13991
rect 78953 13991 79011 13997
rect 75549 13951 75607 13957
rect 75656 13960 78352 13988
rect 72602 13880 72608 13932
rect 72660 13920 72666 13932
rect 73522 13920 73528 13932
rect 72660 13892 72705 13920
rect 73483 13892 73528 13920
rect 72660 13880 72666 13892
rect 73522 13880 73528 13892
rect 73580 13880 73586 13932
rect 73798 13880 73804 13932
rect 73856 13920 73862 13932
rect 74350 13920 74356 13932
rect 73856 13892 74356 13920
rect 73856 13880 73862 13892
rect 74350 13880 74356 13892
rect 74408 13920 74414 13932
rect 75178 13920 75184 13932
rect 74408 13892 75184 13920
rect 74408 13880 74414 13892
rect 75178 13880 75184 13892
rect 75236 13880 75242 13932
rect 75656 13929 75684 13960
rect 75641 13923 75699 13929
rect 75641 13889 75653 13923
rect 75687 13889 75699 13923
rect 75641 13883 75699 13889
rect 76101 13923 76159 13929
rect 76101 13889 76113 13923
rect 76147 13889 76159 13923
rect 76926 13920 76932 13932
rect 76887 13892 76932 13920
rect 76101 13883 76159 13889
rect 70857 13855 70915 13861
rect 70857 13852 70869 13855
rect 70366 13824 70869 13852
rect 66901 13815 66959 13821
rect 70857 13821 70869 13824
rect 70903 13821 70915 13855
rect 70857 13815 70915 13821
rect 70964 13824 72556 13852
rect 61212 13756 61424 13784
rect 61672 13756 65196 13784
rect 56793 13719 56851 13725
rect 56793 13716 56805 13719
rect 55416 13688 56805 13716
rect 56793 13685 56805 13688
rect 56839 13685 56851 13719
rect 56793 13679 56851 13685
rect 56962 13676 56968 13728
rect 57020 13716 57026 13728
rect 61672 13716 61700 13756
rect 68646 13744 68652 13796
rect 68704 13784 68710 13796
rect 70670 13784 70676 13796
rect 68704 13756 70676 13784
rect 68704 13744 68710 13756
rect 70670 13744 70676 13756
rect 70728 13744 70734 13796
rect 70762 13744 70768 13796
rect 70820 13784 70826 13796
rect 70964 13784 70992 13824
rect 70820 13756 70992 13784
rect 72528 13784 72556 13824
rect 72970 13812 72976 13864
rect 73028 13852 73034 13864
rect 73617 13855 73675 13861
rect 73617 13852 73629 13855
rect 73028 13824 73629 13852
rect 73028 13812 73034 13824
rect 73617 13821 73629 13824
rect 73663 13821 73675 13855
rect 73617 13815 73675 13821
rect 73890 13812 73896 13864
rect 73948 13852 73954 13864
rect 76116 13852 76144 13883
rect 76926 13880 76932 13892
rect 76984 13880 76990 13932
rect 77389 13923 77447 13929
rect 77389 13889 77401 13923
rect 77435 13889 77447 13923
rect 77389 13883 77447 13889
rect 77481 13923 77539 13929
rect 77481 13889 77493 13923
rect 77527 13920 77539 13923
rect 78214 13920 78220 13932
rect 77527 13892 78220 13920
rect 77527 13889 77539 13892
rect 77481 13883 77539 13889
rect 73948 13824 76144 13852
rect 73948 13812 73954 13824
rect 73706 13784 73712 13796
rect 72528 13756 73712 13784
rect 70820 13744 70826 13756
rect 73706 13744 73712 13756
rect 73764 13744 73770 13796
rect 74258 13784 74264 13796
rect 74219 13756 74264 13784
rect 74258 13744 74264 13756
rect 74316 13744 74322 13796
rect 77404 13784 77432 13883
rect 78214 13880 78220 13892
rect 78272 13880 78278 13932
rect 78122 13852 78128 13864
rect 78083 13824 78128 13852
rect 78122 13812 78128 13824
rect 78180 13812 78186 13864
rect 78324 13852 78352 13960
rect 78953 13957 78965 13991
rect 78999 13988 79011 13991
rect 79042 13988 79048 14000
rect 78999 13960 79048 13988
rect 78999 13957 79011 13960
rect 78953 13951 79011 13957
rect 79042 13948 79048 13960
rect 79100 13948 79106 14000
rect 78674 13920 78680 13932
rect 78635 13892 78680 13920
rect 78674 13880 78680 13892
rect 78732 13880 78738 13932
rect 80054 13880 80060 13932
rect 80112 13880 80118 13932
rect 81342 13880 81348 13932
rect 81400 13920 81406 13932
rect 83185 13923 83243 13929
rect 83185 13920 83197 13923
rect 81400 13892 83197 13920
rect 81400 13880 81406 13892
rect 83185 13889 83197 13892
rect 83231 13889 83243 13923
rect 83185 13883 83243 13889
rect 84102 13880 84108 13932
rect 84160 13920 84166 13932
rect 86236 13929 86264 14028
rect 86954 14016 86960 14068
rect 87012 14056 87018 14068
rect 88242 14056 88248 14068
rect 87012 14028 88248 14056
rect 87012 14016 87018 14028
rect 88242 14016 88248 14028
rect 88300 14016 88306 14068
rect 92753 14059 92811 14065
rect 92753 14025 92765 14059
rect 92799 14056 92811 14059
rect 94038 14056 94044 14068
rect 92799 14028 94044 14056
rect 92799 14025 92811 14028
rect 92753 14019 92811 14025
rect 94038 14016 94044 14028
rect 94096 14016 94102 14068
rect 89254 13988 89260 14000
rect 89215 13960 89260 13988
rect 89254 13948 89260 13960
rect 89312 13948 89318 14000
rect 89806 13948 89812 14000
rect 89864 13948 89870 14000
rect 85301 13923 85359 13929
rect 85301 13920 85313 13923
rect 84160 13892 85313 13920
rect 84160 13880 84166 13892
rect 85301 13889 85313 13892
rect 85347 13889 85359 13923
rect 85301 13883 85359 13889
rect 86221 13923 86279 13929
rect 86221 13889 86233 13923
rect 86267 13920 86279 13923
rect 87141 13923 87199 13929
rect 87141 13920 87153 13923
rect 86267 13892 87153 13920
rect 86267 13889 86279 13892
rect 86221 13883 86279 13889
rect 87141 13889 87153 13892
rect 87187 13889 87199 13923
rect 87141 13883 87199 13889
rect 90726 13880 90732 13932
rect 90784 13920 90790 13932
rect 91833 13923 91891 13929
rect 91833 13920 91845 13923
rect 90784 13892 91845 13920
rect 90784 13880 90790 13892
rect 91833 13889 91845 13892
rect 91879 13889 91891 13923
rect 91833 13883 91891 13889
rect 92569 13923 92627 13929
rect 92569 13889 92581 13923
rect 92615 13920 92627 13923
rect 92658 13920 92664 13932
rect 92615 13892 92664 13920
rect 92615 13889 92627 13892
rect 92569 13883 92627 13889
rect 92658 13880 92664 13892
rect 92716 13880 92722 13932
rect 78324 13824 80054 13852
rect 76668 13756 77432 13784
rect 80026 13784 80054 13824
rect 83550 13812 83556 13864
rect 83608 13852 83614 13864
rect 83829 13855 83887 13861
rect 83829 13852 83841 13855
rect 83608 13824 83841 13852
rect 83608 13812 83614 13824
rect 83829 13821 83841 13824
rect 83875 13821 83887 13855
rect 83829 13815 83887 13821
rect 84654 13812 84660 13864
rect 84712 13852 84718 13864
rect 84930 13852 84936 13864
rect 84712 13824 84936 13852
rect 84712 13812 84718 13824
rect 84930 13812 84936 13824
rect 84988 13812 84994 13864
rect 87693 13855 87751 13861
rect 87693 13852 87705 13855
rect 86604 13824 87705 13852
rect 80026 13756 80468 13784
rect 63494 13716 63500 13728
rect 57020 13688 61700 13716
rect 63455 13688 63500 13716
rect 57020 13676 57026 13688
rect 63494 13676 63500 13688
rect 63552 13676 63558 13728
rect 64690 13716 64696 13728
rect 64651 13688 64696 13716
rect 64690 13676 64696 13688
rect 64748 13676 64754 13728
rect 66183 13719 66241 13725
rect 66183 13685 66195 13719
rect 66229 13716 66241 13719
rect 66530 13716 66536 13728
rect 66229 13688 66536 13716
rect 66229 13685 66241 13688
rect 66183 13679 66241 13685
rect 66530 13676 66536 13688
rect 66588 13676 66594 13728
rect 68002 13676 68008 13728
rect 68060 13716 68066 13728
rect 68373 13719 68431 13725
rect 68373 13716 68385 13719
rect 68060 13688 68385 13716
rect 68060 13676 68066 13688
rect 68373 13685 68385 13688
rect 68419 13685 68431 13719
rect 68373 13679 68431 13685
rect 70854 13676 70860 13728
rect 70912 13716 70918 13728
rect 72341 13719 72399 13725
rect 72341 13716 72353 13719
rect 70912 13688 72353 13716
rect 70912 13676 70918 13688
rect 72341 13685 72353 13688
rect 72387 13685 72399 13719
rect 72341 13679 72399 13685
rect 73062 13676 73068 13728
rect 73120 13716 73126 13728
rect 76668 13716 76696 13756
rect 76834 13716 76840 13728
rect 73120 13688 76696 13716
rect 76795 13688 76840 13716
rect 73120 13676 73126 13688
rect 76834 13676 76840 13688
rect 76892 13676 76898 13728
rect 77202 13676 77208 13728
rect 77260 13716 77266 13728
rect 79686 13716 79692 13728
rect 77260 13688 79692 13716
rect 77260 13676 77266 13688
rect 79686 13676 79692 13688
rect 79744 13676 79750 13728
rect 80440 13725 80468 13756
rect 80790 13744 80796 13796
rect 80848 13784 80854 13796
rect 81529 13787 81587 13793
rect 81529 13784 81541 13787
rect 80848 13756 81541 13784
rect 80848 13744 80854 13756
rect 81529 13753 81541 13756
rect 81575 13753 81587 13787
rect 81529 13747 81587 13753
rect 85022 13744 85028 13796
rect 85080 13784 85086 13796
rect 86604 13784 86632 13824
rect 87693 13821 87705 13824
rect 87739 13852 87751 13855
rect 87966 13852 87972 13864
rect 87739 13824 87972 13852
rect 87739 13821 87751 13824
rect 87693 13815 87751 13821
rect 87966 13812 87972 13824
rect 88024 13812 88030 13864
rect 88978 13852 88984 13864
rect 88939 13824 88984 13852
rect 88978 13812 88984 13824
rect 89036 13852 89042 13864
rect 91281 13855 91339 13861
rect 91281 13852 91293 13855
rect 89036 13824 91293 13852
rect 89036 13812 89042 13824
rect 91281 13821 91293 13824
rect 91327 13821 91339 13855
rect 91281 13815 91339 13821
rect 85080 13756 86632 13784
rect 85080 13744 85086 13756
rect 80425 13719 80483 13725
rect 80425 13685 80437 13719
rect 80471 13716 80483 13719
rect 80514 13716 80520 13728
rect 80471 13688 80520 13716
rect 80471 13685 80483 13688
rect 80425 13679 80483 13685
rect 80514 13676 80520 13688
rect 80572 13676 80578 13728
rect 81066 13676 81072 13728
rect 81124 13716 81130 13728
rect 82081 13719 82139 13725
rect 82081 13716 82093 13719
rect 81124 13688 82093 13716
rect 81124 13676 81130 13688
rect 82081 13685 82093 13688
rect 82127 13716 82139 13719
rect 85850 13716 85856 13728
rect 82127 13688 85856 13716
rect 82127 13685 82139 13688
rect 82081 13679 82139 13685
rect 85850 13676 85856 13688
rect 85908 13676 85914 13728
rect 90542 13676 90548 13728
rect 90600 13716 90606 13728
rect 90729 13719 90787 13725
rect 90729 13716 90741 13719
rect 90600 13688 90741 13716
rect 90600 13676 90606 13688
rect 90729 13685 90741 13688
rect 90775 13685 90787 13719
rect 90729 13679 90787 13685
rect 92658 13676 92664 13728
rect 92716 13716 92722 13728
rect 93213 13719 93271 13725
rect 93213 13716 93225 13719
rect 92716 13688 93225 13716
rect 92716 13676 92722 13688
rect 93213 13685 93225 13688
rect 93259 13685 93271 13719
rect 94130 13716 94136 13728
rect 94091 13688 94136 13716
rect 93213 13679 93271 13685
rect 94130 13676 94136 13688
rect 94188 13676 94194 13728
rect 1104 13626 94852 13648
rect 1104 13574 12668 13626
rect 12720 13574 12732 13626
rect 12784 13574 12796 13626
rect 12848 13574 12860 13626
rect 12912 13574 12924 13626
rect 12976 13574 36105 13626
rect 36157 13574 36169 13626
rect 36221 13574 36233 13626
rect 36285 13574 36297 13626
rect 36349 13574 36361 13626
rect 36413 13574 59542 13626
rect 59594 13574 59606 13626
rect 59658 13574 59670 13626
rect 59722 13574 59734 13626
rect 59786 13574 59798 13626
rect 59850 13574 82979 13626
rect 83031 13574 83043 13626
rect 83095 13574 83107 13626
rect 83159 13574 83171 13626
rect 83223 13574 83235 13626
rect 83287 13574 94852 13626
rect 1104 13552 94852 13574
rect 5074 13512 5080 13524
rect 5035 13484 5080 13512
rect 5074 13472 5080 13484
rect 5132 13472 5138 13524
rect 6822 13472 6828 13524
rect 6880 13512 6886 13524
rect 6880 13484 7512 13512
rect 6880 13472 6886 13484
rect 5721 13447 5779 13453
rect 5721 13413 5733 13447
rect 5767 13444 5779 13447
rect 7282 13444 7288 13456
rect 5767 13416 7288 13444
rect 5767 13413 5779 13416
rect 5721 13407 5779 13413
rect 7282 13404 7288 13416
rect 7340 13404 7346 13456
rect 7484 13453 7512 13484
rect 8110 13472 8116 13524
rect 8168 13512 8174 13524
rect 19426 13512 19432 13524
rect 8168 13484 19432 13512
rect 8168 13472 8174 13484
rect 19426 13472 19432 13484
rect 19484 13472 19490 13524
rect 21082 13512 21088 13524
rect 19536 13484 21088 13512
rect 7469 13447 7527 13453
rect 7469 13413 7481 13447
rect 7515 13444 7527 13447
rect 11238 13444 11244 13456
rect 7515 13416 11244 13444
rect 7515 13413 7527 13416
rect 7469 13407 7527 13413
rect 11238 13404 11244 13416
rect 11296 13404 11302 13456
rect 13354 13404 13360 13456
rect 13412 13444 13418 13456
rect 13449 13447 13507 13453
rect 13449 13444 13461 13447
rect 13412 13416 13461 13444
rect 13412 13404 13418 13416
rect 13449 13413 13461 13416
rect 13495 13444 13507 13447
rect 13998 13444 14004 13456
rect 13495 13416 14004 13444
rect 13495 13413 13507 13416
rect 13449 13407 13507 13413
rect 13998 13404 14004 13416
rect 14056 13404 14062 13456
rect 19536 13444 19564 13484
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 21177 13515 21235 13521
rect 21177 13481 21189 13515
rect 21223 13512 21235 13515
rect 21910 13512 21916 13524
rect 21223 13484 21916 13512
rect 21223 13481 21235 13484
rect 21177 13475 21235 13481
rect 21910 13472 21916 13484
rect 21968 13472 21974 13524
rect 22002 13472 22008 13524
rect 22060 13512 22066 13524
rect 22094 13512 22100 13524
rect 22060 13484 22100 13512
rect 22060 13472 22066 13484
rect 22094 13472 22100 13484
rect 22152 13472 22158 13524
rect 22296 13484 24072 13512
rect 16316 13416 19564 13444
rect 2958 13376 2964 13388
rect 2919 13348 2964 13376
rect 2958 13336 2964 13348
rect 3016 13336 3022 13388
rect 4062 13376 4068 13388
rect 4023 13348 4068 13376
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 7374 13336 7380 13388
rect 7432 13376 7438 13388
rect 8113 13379 8171 13385
rect 8113 13376 8125 13379
rect 7432 13348 8125 13376
rect 7432 13336 7438 13348
rect 8113 13345 8125 13348
rect 8159 13345 8171 13379
rect 8113 13339 8171 13345
rect 8478 13336 8484 13388
rect 8536 13376 8542 13388
rect 9766 13376 9772 13388
rect 8536 13348 9444 13376
rect 9727 13348 9772 13376
rect 8536 13336 8542 13348
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13308 3111 13311
rect 4154 13308 4160 13320
rect 3099 13280 4160 13308
rect 3099 13277 3111 13280
rect 3053 13271 3111 13277
rect 4154 13268 4160 13280
rect 4212 13268 4218 13320
rect 5810 13308 5816 13320
rect 5771 13280 5816 13308
rect 5810 13268 5816 13280
rect 5868 13268 5874 13320
rect 5997 13311 6055 13317
rect 5997 13277 6009 13311
rect 6043 13308 6055 13311
rect 6822 13308 6828 13320
rect 6043 13280 6828 13308
rect 6043 13277 6055 13280
rect 5997 13271 6055 13277
rect 6822 13268 6828 13280
rect 6880 13268 6886 13320
rect 8205 13311 8263 13317
rect 8205 13277 8217 13311
rect 8251 13308 8263 13311
rect 9306 13308 9312 13320
rect 8251 13280 9312 13308
rect 8251 13277 8263 13280
rect 8205 13271 8263 13277
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 9416 13308 9444 13348
rect 9766 13336 9772 13348
rect 9824 13336 9830 13388
rect 11422 13336 11428 13388
rect 11480 13376 11486 13388
rect 12069 13379 12127 13385
rect 12069 13376 12081 13379
rect 11480 13348 12081 13376
rect 11480 13336 11486 13348
rect 12069 13345 12081 13348
rect 12115 13345 12127 13379
rect 14550 13376 14556 13388
rect 12069 13339 12127 13345
rect 12406 13348 14136 13376
rect 14511 13348 14556 13376
rect 10134 13308 10140 13320
rect 9416 13280 10140 13308
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 10502 13308 10508 13320
rect 10463 13280 10508 13308
rect 10502 13268 10508 13280
rect 10560 13268 10566 13320
rect 12406 13308 12434 13348
rect 10612 13280 12434 13308
rect 12621 13311 12679 13317
rect 4430 13200 4436 13252
rect 4488 13240 4494 13252
rect 10612 13240 10640 13280
rect 12621 13277 12633 13311
rect 12667 13308 12679 13311
rect 13998 13308 14004 13320
rect 12667 13280 14004 13308
rect 12667 13277 12679 13280
rect 12621 13271 12679 13277
rect 13998 13268 14004 13280
rect 14056 13268 14062 13320
rect 4488 13212 10640 13240
rect 4488 13200 4494 13212
rect 10686 13200 10692 13252
rect 10744 13240 10750 13252
rect 11422 13240 11428 13252
rect 10744 13212 11428 13240
rect 10744 13200 10750 13212
rect 11422 13200 11428 13212
rect 11480 13200 11486 13252
rect 3418 13172 3424 13184
rect 3379 13144 3424 13172
rect 3418 13132 3424 13144
rect 3476 13132 3482 13184
rect 4522 13172 4528 13184
rect 4483 13144 4528 13172
rect 4522 13132 4528 13144
rect 4580 13132 4586 13184
rect 6917 13175 6975 13181
rect 6917 13141 6929 13175
rect 6963 13172 6975 13175
rect 7006 13172 7012 13184
rect 6963 13144 7012 13172
rect 6963 13141 6975 13144
rect 6917 13135 6975 13141
rect 7006 13132 7012 13144
rect 7064 13132 7070 13184
rect 7650 13132 7656 13184
rect 7708 13172 7714 13184
rect 8478 13172 8484 13184
rect 7708 13144 8484 13172
rect 7708 13132 7714 13144
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 8573 13175 8631 13181
rect 8573 13141 8585 13175
rect 8619 13172 8631 13175
rect 13262 13172 13268 13184
rect 8619 13144 13268 13172
rect 8619 13141 8631 13144
rect 8573 13135 8631 13141
rect 13262 13132 13268 13144
rect 13320 13132 13326 13184
rect 14108 13172 14136 13348
rect 14550 13336 14556 13348
rect 14608 13336 14614 13388
rect 15010 13336 15016 13388
rect 15068 13376 15074 13388
rect 16114 13376 16120 13388
rect 15068 13348 16120 13376
rect 15068 13336 15074 13348
rect 16114 13336 16120 13348
rect 16172 13336 16178 13388
rect 16316 13385 16344 13416
rect 20714 13404 20720 13456
rect 20772 13444 20778 13456
rect 22296 13444 22324 13484
rect 20772 13416 22324 13444
rect 20772 13404 20778 13416
rect 16301 13379 16359 13385
rect 16301 13345 16313 13379
rect 16347 13345 16359 13379
rect 21266 13376 21272 13388
rect 16301 13339 16359 13345
rect 18248 13348 21272 13376
rect 14274 13308 14280 13320
rect 14235 13280 14280 13308
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 16758 13268 16764 13320
rect 16816 13308 16822 13320
rect 17037 13311 17095 13317
rect 17037 13308 17049 13311
rect 16816 13280 17049 13308
rect 16816 13268 16822 13280
rect 17037 13277 17049 13280
rect 17083 13308 17095 13311
rect 17402 13308 17408 13320
rect 17083 13280 17408 13308
rect 17083 13277 17095 13280
rect 17037 13271 17095 13277
rect 17402 13268 17408 13280
rect 17460 13268 17466 13320
rect 18248 13317 18276 13348
rect 21266 13336 21272 13348
rect 21324 13336 21330 13388
rect 22094 13336 22100 13388
rect 22152 13376 22158 13388
rect 23937 13379 23995 13385
rect 22152 13348 23888 13376
rect 22152 13336 22158 13348
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13277 18291 13311
rect 18233 13271 18291 13277
rect 18877 13311 18935 13317
rect 18877 13277 18889 13311
rect 18923 13308 18935 13311
rect 19242 13308 19248 13320
rect 18923 13280 19248 13308
rect 18923 13277 18935 13280
rect 18877 13271 18935 13277
rect 19242 13268 19248 13280
rect 19300 13268 19306 13320
rect 19426 13308 19432 13320
rect 19387 13280 19432 13308
rect 19426 13268 19432 13280
rect 19484 13268 19490 13320
rect 22186 13308 22192 13320
rect 22147 13280 22192 13308
rect 22186 13268 22192 13280
rect 22244 13268 22250 13320
rect 15562 13200 15568 13252
rect 15620 13200 15626 13252
rect 17494 13240 17500 13252
rect 15856 13212 17500 13240
rect 15856 13172 15884 13212
rect 17494 13200 17500 13212
rect 17552 13200 17558 13252
rect 18141 13243 18199 13249
rect 18141 13209 18153 13243
rect 18187 13240 18199 13243
rect 19334 13240 19340 13252
rect 18187 13212 19340 13240
rect 18187 13209 18199 13212
rect 18141 13203 18199 13209
rect 19334 13200 19340 13212
rect 19392 13200 19398 13252
rect 19702 13240 19708 13252
rect 19663 13212 19708 13240
rect 19702 13200 19708 13212
rect 19760 13200 19766 13252
rect 19812 13212 20194 13240
rect 16850 13172 16856 13184
rect 14108 13144 15884 13172
rect 16811 13144 16856 13172
rect 16850 13132 16856 13144
rect 16908 13132 16914 13184
rect 17589 13175 17647 13181
rect 17589 13141 17601 13175
rect 17635 13172 17647 13175
rect 17954 13172 17960 13184
rect 17635 13144 17960 13172
rect 17635 13141 17647 13144
rect 17589 13135 17647 13141
rect 17954 13132 17960 13144
rect 18012 13132 18018 13184
rect 18785 13175 18843 13181
rect 18785 13141 18797 13175
rect 18831 13172 18843 13175
rect 19812 13172 19840 13212
rect 21450 13200 21456 13252
rect 21508 13240 21514 13252
rect 22465 13243 22523 13249
rect 22465 13240 22477 13243
rect 21508 13212 22477 13240
rect 21508 13200 21514 13212
rect 22465 13209 22477 13212
rect 22511 13209 22523 13243
rect 22465 13203 22523 13209
rect 23198 13200 23204 13252
rect 23256 13200 23262 13252
rect 23860 13240 23888 13348
rect 23937 13345 23949 13379
rect 23983 13345 23995 13379
rect 24044 13376 24072 13484
rect 25314 13472 25320 13524
rect 25372 13512 25378 13524
rect 27430 13512 27436 13524
rect 25372 13484 27436 13512
rect 25372 13472 25378 13484
rect 27430 13472 27436 13484
rect 27488 13472 27494 13524
rect 27525 13515 27583 13521
rect 27525 13481 27537 13515
rect 27571 13512 27583 13515
rect 27614 13512 27620 13524
rect 27571 13484 27620 13512
rect 27571 13481 27583 13484
rect 27525 13475 27583 13481
rect 27614 13472 27620 13484
rect 27672 13472 27678 13524
rect 28442 13512 28448 13524
rect 28403 13484 28448 13512
rect 28442 13472 28448 13484
rect 28500 13472 28506 13524
rect 28534 13472 28540 13524
rect 28592 13512 28598 13524
rect 29454 13512 29460 13524
rect 28592 13484 29460 13512
rect 28592 13472 28598 13484
rect 29454 13472 29460 13484
rect 29512 13472 29518 13524
rect 30190 13472 30196 13524
rect 30248 13512 30254 13524
rect 31018 13512 31024 13524
rect 30248 13484 31024 13512
rect 30248 13472 30254 13484
rect 31018 13472 31024 13484
rect 31076 13472 31082 13524
rect 31478 13512 31484 13524
rect 31439 13484 31484 13512
rect 31478 13472 31484 13484
rect 31536 13472 31542 13524
rect 31754 13472 31760 13524
rect 31812 13512 31818 13524
rect 32766 13512 32772 13524
rect 31812 13484 32772 13512
rect 31812 13472 31818 13484
rect 32766 13472 32772 13484
rect 32824 13472 32830 13524
rect 32858 13472 32864 13524
rect 32916 13512 32922 13524
rect 33410 13512 33416 13524
rect 32916 13484 33416 13512
rect 32916 13472 32922 13484
rect 33410 13472 33416 13484
rect 33468 13472 33474 13524
rect 35894 13472 35900 13524
rect 35952 13512 35958 13524
rect 35989 13515 36047 13521
rect 35989 13512 36001 13515
rect 35952 13484 36001 13512
rect 35952 13472 35958 13484
rect 35989 13481 36001 13484
rect 36035 13481 36047 13515
rect 37274 13512 37280 13524
rect 37235 13484 37280 13512
rect 35989 13475 36047 13481
rect 37274 13472 37280 13484
rect 37332 13472 37338 13524
rect 38197 13515 38255 13521
rect 38197 13481 38209 13515
rect 38243 13512 38255 13515
rect 38470 13512 38476 13524
rect 38243 13484 38476 13512
rect 38243 13481 38255 13484
rect 38197 13475 38255 13481
rect 38470 13472 38476 13484
rect 38528 13472 38534 13524
rect 42426 13472 42432 13524
rect 42484 13512 42490 13524
rect 44361 13515 44419 13521
rect 44361 13512 44373 13515
rect 42484 13484 44373 13512
rect 42484 13472 42490 13484
rect 44361 13481 44373 13484
rect 44407 13512 44419 13515
rect 46842 13512 46848 13524
rect 44407 13484 46848 13512
rect 44407 13481 44419 13484
rect 44361 13475 44419 13481
rect 46842 13472 46848 13484
rect 46900 13472 46906 13524
rect 49326 13512 49332 13524
rect 46952 13484 49332 13512
rect 26786 13404 26792 13456
rect 26844 13444 26850 13456
rect 29546 13444 29552 13456
rect 26844 13416 29552 13444
rect 26844 13404 26850 13416
rect 29546 13404 29552 13416
rect 29604 13404 29610 13456
rect 36446 13444 36452 13456
rect 31312 13416 36452 13444
rect 25409 13379 25467 13385
rect 25409 13376 25421 13379
rect 24044 13348 25421 13376
rect 23937 13339 23995 13345
rect 25409 13345 25421 13348
rect 25455 13376 25467 13379
rect 30558 13376 30564 13388
rect 25455 13348 30564 13376
rect 25455 13345 25467 13348
rect 25409 13339 25467 13345
rect 23952 13308 23980 13339
rect 30558 13336 30564 13348
rect 30616 13336 30622 13388
rect 25133 13311 25191 13317
rect 25133 13308 25145 13311
rect 23952 13280 25145 13308
rect 25133 13277 25145 13280
rect 25179 13277 25191 13311
rect 25133 13271 25191 13277
rect 25958 13268 25964 13320
rect 26016 13308 26022 13320
rect 26053 13311 26111 13317
rect 26053 13308 26065 13311
rect 26016 13280 26065 13308
rect 26016 13268 26022 13280
rect 26053 13277 26065 13280
rect 26099 13277 26111 13311
rect 26053 13271 26111 13277
rect 27706 13268 27712 13320
rect 27764 13308 27770 13320
rect 28261 13311 28319 13317
rect 28261 13308 28273 13311
rect 27764 13280 28273 13308
rect 27764 13268 27770 13280
rect 28261 13277 28273 13280
rect 28307 13277 28319 13311
rect 29730 13308 29736 13320
rect 29691 13280 29736 13308
rect 28261 13271 28319 13277
rect 29730 13268 29736 13280
rect 29788 13268 29794 13320
rect 24581 13243 24639 13249
rect 24581 13240 24593 13243
rect 23860 13212 24593 13240
rect 24581 13209 24593 13212
rect 24627 13240 24639 13243
rect 26326 13240 26332 13252
rect 24627 13212 26332 13240
rect 24627 13209 24639 13212
rect 24581 13203 24639 13209
rect 26326 13200 26332 13212
rect 26384 13200 26390 13252
rect 30006 13240 30012 13252
rect 26896 13212 29886 13240
rect 29967 13212 30012 13240
rect 18831 13144 19840 13172
rect 18831 13141 18843 13144
rect 18785 13135 18843 13141
rect 21082 13132 21088 13184
rect 21140 13172 21146 13184
rect 26896 13172 26924 13212
rect 21140 13144 26924 13172
rect 21140 13132 21146 13144
rect 27430 13132 27436 13184
rect 27488 13172 27494 13184
rect 29086 13172 29092 13184
rect 27488 13144 29092 13172
rect 27488 13132 27494 13144
rect 29086 13132 29092 13144
rect 29144 13132 29150 13184
rect 29181 13175 29239 13181
rect 29181 13141 29193 13175
rect 29227 13172 29239 13175
rect 29638 13172 29644 13184
rect 29227 13144 29644 13172
rect 29227 13141 29239 13144
rect 29181 13135 29239 13141
rect 29638 13132 29644 13144
rect 29696 13132 29702 13184
rect 29858 13172 29886 13212
rect 30006 13200 30012 13212
rect 30064 13200 30070 13252
rect 30466 13200 30472 13252
rect 30524 13200 30530 13252
rect 31312 13172 31340 13416
rect 36446 13404 36452 13416
rect 36504 13404 36510 13456
rect 36630 13404 36636 13456
rect 36688 13444 36694 13456
rect 41141 13447 41199 13453
rect 41141 13444 41153 13447
rect 36688 13416 41153 13444
rect 36688 13404 36694 13416
rect 41141 13413 41153 13416
rect 41187 13444 41199 13447
rect 42518 13444 42524 13456
rect 41187 13416 42524 13444
rect 41187 13413 41199 13416
rect 41141 13407 41199 13413
rect 42518 13404 42524 13416
rect 42576 13404 42582 13456
rect 44284 13416 45324 13444
rect 32674 13376 32680 13388
rect 32635 13348 32680 13376
rect 32674 13336 32680 13348
rect 32732 13336 32738 13388
rect 32766 13336 32772 13388
rect 32824 13376 32830 13388
rect 32824 13348 35894 13376
rect 32824 13336 32830 13348
rect 32490 13308 32496 13320
rect 32451 13280 32496 13308
rect 32490 13268 32496 13280
rect 32548 13268 32554 13320
rect 35434 13308 35440 13320
rect 35395 13280 35440 13308
rect 35434 13268 35440 13280
rect 35492 13268 35498 13320
rect 31478 13200 31484 13252
rect 31536 13240 31542 13252
rect 33962 13240 33968 13252
rect 31536 13212 33968 13240
rect 31536 13200 31542 13212
rect 33962 13200 33968 13212
rect 34020 13240 34026 13252
rect 34333 13243 34391 13249
rect 34333 13240 34345 13243
rect 34020 13212 34345 13240
rect 34020 13200 34026 13212
rect 34333 13209 34345 13212
rect 34379 13240 34391 13243
rect 35710 13240 35716 13252
rect 34379 13212 35716 13240
rect 34379 13209 34391 13212
rect 34333 13203 34391 13209
rect 35710 13200 35716 13212
rect 35768 13200 35774 13252
rect 35866 13240 35894 13348
rect 35986 13336 35992 13388
rect 36044 13376 36050 13388
rect 44284 13376 44312 13416
rect 45186 13376 45192 13388
rect 36044 13348 44312 13376
rect 45147 13348 45192 13376
rect 36044 13336 36050 13348
rect 45186 13336 45192 13348
rect 45244 13336 45250 13388
rect 45296 13376 45324 13416
rect 46952 13376 46980 13484
rect 49326 13472 49332 13484
rect 49384 13472 49390 13524
rect 52362 13472 52368 13524
rect 52420 13512 52426 13524
rect 52825 13515 52883 13521
rect 52825 13512 52837 13515
rect 52420 13484 52837 13512
rect 52420 13472 52426 13484
rect 52825 13481 52837 13484
rect 52871 13481 52883 13515
rect 52825 13475 52883 13481
rect 52932 13484 54708 13512
rect 49602 13404 49608 13456
rect 49660 13444 49666 13456
rect 49660 13416 50476 13444
rect 49660 13404 49666 13416
rect 50448 13385 50476 13416
rect 51718 13404 51724 13456
rect 51776 13444 51782 13456
rect 52932 13444 52960 13484
rect 51776 13416 52960 13444
rect 51776 13404 51782 13416
rect 45296 13348 46980 13376
rect 47397 13379 47455 13385
rect 47397 13345 47409 13379
rect 47443 13376 47455 13379
rect 49697 13379 49755 13385
rect 49697 13376 49709 13379
rect 47443 13348 49709 13376
rect 47443 13345 47455 13348
rect 47397 13339 47455 13345
rect 49697 13345 49709 13348
rect 49743 13345 49755 13379
rect 49697 13339 49755 13345
rect 50433 13379 50491 13385
rect 50433 13345 50445 13379
rect 50479 13376 50491 13379
rect 51534 13376 51540 13388
rect 50479 13348 51540 13376
rect 50479 13345 50491 13348
rect 50433 13339 50491 13345
rect 51534 13336 51540 13348
rect 51592 13336 51598 13388
rect 54297 13379 54355 13385
rect 54297 13376 54309 13379
rect 52012 13348 54309 13376
rect 36081 13311 36139 13317
rect 36081 13277 36093 13311
rect 36127 13308 36139 13311
rect 36446 13308 36452 13320
rect 36127 13280 36452 13308
rect 36127 13277 36139 13280
rect 36081 13271 36139 13277
rect 36446 13268 36452 13280
rect 36504 13268 36510 13320
rect 36725 13311 36783 13317
rect 36725 13277 36737 13311
rect 36771 13308 36783 13311
rect 38286 13308 38292 13320
rect 36771 13280 38292 13308
rect 36771 13277 36783 13280
rect 36725 13271 36783 13277
rect 38286 13268 38292 13280
rect 38344 13268 38350 13320
rect 38470 13268 38476 13320
rect 38528 13308 38534 13320
rect 40221 13311 40279 13317
rect 40221 13308 40233 13311
rect 38528 13280 40233 13308
rect 38528 13268 38534 13280
rect 40221 13277 40233 13280
rect 40267 13308 40279 13311
rect 40310 13308 40316 13320
rect 40267 13280 40316 13308
rect 40267 13277 40279 13280
rect 40221 13271 40279 13277
rect 40310 13268 40316 13280
rect 40368 13268 40374 13320
rect 42426 13308 42432 13320
rect 42387 13280 42432 13308
rect 42426 13268 42432 13280
rect 42484 13268 42490 13320
rect 48774 13268 48780 13320
rect 48832 13268 48838 13320
rect 49234 13268 49240 13320
rect 49292 13308 49298 13320
rect 49605 13311 49663 13317
rect 49605 13308 49617 13311
rect 49292 13280 49617 13308
rect 49292 13268 49298 13280
rect 49605 13277 49617 13280
rect 49651 13277 49663 13311
rect 49605 13271 49663 13277
rect 50338 13268 50344 13320
rect 50396 13308 50402 13320
rect 51813 13311 51871 13317
rect 51813 13308 51825 13311
rect 50396 13280 51825 13308
rect 50396 13268 50402 13280
rect 51813 13277 51825 13280
rect 51859 13277 51871 13311
rect 51813 13271 51871 13277
rect 39390 13240 39396 13252
rect 35866 13212 39396 13240
rect 39390 13200 39396 13212
rect 39448 13200 39454 13252
rect 39485 13243 39543 13249
rect 39485 13209 39497 13243
rect 39531 13240 39543 13243
rect 42886 13240 42892 13252
rect 39531 13212 40724 13240
rect 42847 13212 42892 13240
rect 39531 13209 39543 13212
rect 39485 13203 39543 13209
rect 29858 13144 31340 13172
rect 32033 13175 32091 13181
rect 32033 13141 32045 13175
rect 32079 13172 32091 13175
rect 32214 13172 32220 13184
rect 32079 13144 32220 13172
rect 32079 13141 32091 13144
rect 32033 13135 32091 13141
rect 32214 13132 32220 13144
rect 32272 13132 32278 13184
rect 32858 13132 32864 13184
rect 32916 13172 32922 13184
rect 35345 13175 35403 13181
rect 35345 13172 35357 13175
rect 32916 13144 35357 13172
rect 32916 13132 32922 13144
rect 35345 13141 35357 13144
rect 35391 13141 35403 13175
rect 35345 13135 35403 13141
rect 35618 13132 35624 13184
rect 35676 13172 35682 13184
rect 39942 13172 39948 13184
rect 35676 13144 39948 13172
rect 35676 13132 35682 13144
rect 39942 13132 39948 13144
rect 40000 13132 40006 13184
rect 40126 13172 40132 13184
rect 40087 13144 40132 13172
rect 40126 13132 40132 13144
rect 40184 13132 40190 13184
rect 40696 13172 40724 13212
rect 42886 13200 42892 13212
rect 42944 13200 42950 13252
rect 43162 13200 43168 13252
rect 43220 13240 43226 13252
rect 45465 13243 45523 13249
rect 45465 13240 45477 13243
rect 43220 13212 45477 13240
rect 43220 13200 43226 13212
rect 45465 13209 45477 13212
rect 45511 13209 45523 13243
rect 45465 13203 45523 13209
rect 46474 13200 46480 13252
rect 46532 13200 46538 13252
rect 47670 13240 47676 13252
rect 47631 13212 47676 13240
rect 47670 13200 47676 13212
rect 47728 13200 47734 13252
rect 49050 13200 49056 13252
rect 49108 13240 49114 13252
rect 52012 13240 52040 13348
rect 54297 13345 54309 13348
rect 54343 13345 54355 13379
rect 54297 13339 54355 13345
rect 54573 13311 54631 13317
rect 54573 13277 54585 13311
rect 54619 13277 54631 13311
rect 54573 13271 54631 13277
rect 49108 13212 52040 13240
rect 49108 13200 49114 13212
rect 52086 13200 52092 13252
rect 52144 13240 52150 13252
rect 52144 13212 52189 13240
rect 52144 13200 52150 13212
rect 53650 13200 53656 13252
rect 53708 13200 53714 13252
rect 44726 13172 44732 13184
rect 40696 13144 44732 13172
rect 44726 13132 44732 13144
rect 44784 13132 44790 13184
rect 46750 13132 46756 13184
rect 46808 13172 46814 13184
rect 46937 13175 46995 13181
rect 46937 13172 46949 13175
rect 46808 13144 46949 13172
rect 46808 13132 46814 13144
rect 46937 13141 46949 13144
rect 46983 13141 46995 13175
rect 46937 13135 46995 13141
rect 48958 13132 48964 13184
rect 49016 13172 49022 13184
rect 49145 13175 49203 13181
rect 49145 13172 49157 13175
rect 49016 13144 49157 13172
rect 49016 13132 49022 13144
rect 49145 13141 49157 13144
rect 49191 13141 49203 13175
rect 49145 13135 49203 13141
rect 50985 13175 51043 13181
rect 50985 13141 50997 13175
rect 51031 13172 51043 13175
rect 51258 13172 51264 13184
rect 51031 13144 51264 13172
rect 51031 13141 51043 13144
rect 50985 13135 51043 13141
rect 51258 13132 51264 13144
rect 51316 13172 51322 13184
rect 52178 13172 52184 13184
rect 51316 13144 52184 13172
rect 51316 13132 51322 13144
rect 52178 13132 52184 13144
rect 52236 13132 52242 13184
rect 54588 13172 54616 13271
rect 54680 13240 54708 13484
rect 56594 13472 56600 13524
rect 56652 13512 56658 13524
rect 57238 13512 57244 13524
rect 56652 13484 57244 13512
rect 56652 13472 56658 13484
rect 57238 13472 57244 13484
rect 57296 13472 57302 13524
rect 57882 13472 57888 13524
rect 57940 13512 57946 13524
rect 60458 13512 60464 13524
rect 57940 13484 60464 13512
rect 57940 13472 57946 13484
rect 60458 13472 60464 13484
rect 60516 13472 60522 13524
rect 60752 13484 60964 13512
rect 60752 13444 60780 13484
rect 56152 13416 60780 13444
rect 60936 13444 60964 13484
rect 61010 13472 61016 13524
rect 61068 13512 61074 13524
rect 65153 13515 65211 13521
rect 65153 13512 65165 13515
rect 61068 13484 65165 13512
rect 61068 13472 61074 13484
rect 65153 13481 65165 13484
rect 65199 13481 65211 13515
rect 69014 13512 69020 13524
rect 65153 13475 65211 13481
rect 65260 13484 69020 13512
rect 62114 13444 62120 13456
rect 60936 13416 62120 13444
rect 56152 13317 56180 13416
rect 62114 13404 62120 13416
rect 62172 13404 62178 13456
rect 64230 13404 64236 13456
rect 64288 13444 64294 13456
rect 65260 13444 65288 13484
rect 69014 13472 69020 13484
rect 69072 13472 69078 13524
rect 69937 13515 69995 13521
rect 69937 13481 69949 13515
rect 69983 13512 69995 13515
rect 70854 13512 70860 13524
rect 69983 13484 70860 13512
rect 69983 13481 69995 13484
rect 69937 13475 69995 13481
rect 70854 13472 70860 13484
rect 70912 13472 70918 13524
rect 71038 13512 71044 13524
rect 70999 13484 71044 13512
rect 71038 13472 71044 13484
rect 71096 13472 71102 13524
rect 71866 13512 71872 13524
rect 71516 13484 71872 13512
rect 64288 13416 65288 13444
rect 66625 13447 66683 13453
rect 64288 13404 64294 13416
rect 66625 13413 66637 13447
rect 66671 13444 66683 13447
rect 71516 13444 71544 13484
rect 71866 13472 71872 13484
rect 71924 13472 71930 13524
rect 72510 13472 72516 13524
rect 72568 13512 72574 13524
rect 76098 13512 76104 13524
rect 72568 13484 75960 13512
rect 76059 13484 76104 13512
rect 72568 13472 72574 13484
rect 66671 13416 71544 13444
rect 66671 13413 66683 13416
rect 66625 13407 66683 13413
rect 73062 13404 73068 13456
rect 73120 13444 73126 13456
rect 73341 13447 73399 13453
rect 73341 13444 73353 13447
rect 73120 13416 73353 13444
rect 73120 13404 73126 13416
rect 73341 13413 73353 13416
rect 73387 13413 73399 13447
rect 75932 13444 75960 13484
rect 76098 13472 76104 13484
rect 76156 13472 76162 13524
rect 78950 13512 78956 13524
rect 77128 13484 78956 13512
rect 77128 13444 77156 13484
rect 78950 13472 78956 13484
rect 79008 13472 79014 13524
rect 79042 13472 79048 13524
rect 79100 13512 79106 13524
rect 79413 13515 79471 13521
rect 79413 13512 79425 13515
rect 79100 13484 79425 13512
rect 79100 13472 79106 13484
rect 79413 13481 79425 13484
rect 79459 13481 79471 13515
rect 79413 13475 79471 13481
rect 79686 13472 79692 13524
rect 79744 13512 79750 13524
rect 81805 13515 81863 13521
rect 81805 13512 81817 13515
rect 79744 13484 81817 13512
rect 79744 13472 79750 13484
rect 81805 13481 81817 13484
rect 81851 13481 81863 13515
rect 81805 13475 81863 13481
rect 84194 13472 84200 13524
rect 84252 13512 84258 13524
rect 85206 13512 85212 13524
rect 84252 13484 85212 13512
rect 84252 13472 84258 13484
rect 85206 13472 85212 13484
rect 85264 13472 85270 13524
rect 88978 13512 88984 13524
rect 86696 13484 88984 13512
rect 75932 13416 77156 13444
rect 73341 13407 73399 13413
rect 78306 13404 78312 13456
rect 78364 13444 78370 13456
rect 78769 13447 78827 13453
rect 78769 13444 78781 13447
rect 78364 13416 78781 13444
rect 78364 13404 78370 13416
rect 78769 13413 78781 13416
rect 78815 13413 78827 13447
rect 78769 13407 78827 13413
rect 79962 13404 79968 13456
rect 80020 13444 80026 13456
rect 81158 13444 81164 13456
rect 80020 13416 81164 13444
rect 80020 13404 80026 13416
rect 81158 13404 81164 13416
rect 81216 13404 81222 13456
rect 86696 13453 86724 13484
rect 88978 13472 88984 13484
rect 89036 13472 89042 13524
rect 89165 13515 89223 13521
rect 89165 13481 89177 13515
rect 89211 13512 89223 13515
rect 89346 13512 89352 13524
rect 89211 13484 89352 13512
rect 89211 13481 89223 13484
rect 89165 13475 89223 13481
rect 89346 13472 89352 13484
rect 89404 13472 89410 13524
rect 89806 13512 89812 13524
rect 89767 13484 89812 13512
rect 89806 13472 89812 13484
rect 89864 13472 89870 13524
rect 85669 13447 85727 13453
rect 85669 13444 85681 13447
rect 84212 13416 85681 13444
rect 56226 13336 56232 13388
rect 56284 13376 56290 13388
rect 58434 13376 58440 13388
rect 56284 13348 58440 13376
rect 56284 13336 56290 13348
rect 58434 13336 58440 13348
rect 58492 13336 58498 13388
rect 58986 13376 58992 13388
rect 58947 13348 58992 13376
rect 58986 13336 58992 13348
rect 59044 13336 59050 13388
rect 62482 13376 62488 13388
rect 59188 13348 59400 13376
rect 56137 13311 56195 13317
rect 56137 13277 56149 13311
rect 56183 13277 56195 13311
rect 56137 13271 56195 13277
rect 56413 13311 56471 13317
rect 56413 13277 56425 13311
rect 56459 13308 56471 13311
rect 59188 13308 59216 13348
rect 56459 13280 59216 13308
rect 56459 13277 56471 13280
rect 56413 13271 56471 13277
rect 57238 13240 57244 13252
rect 54680 13212 57100 13240
rect 57199 13212 57244 13240
rect 55858 13172 55864 13184
rect 54588 13144 55864 13172
rect 55858 13132 55864 13144
rect 55916 13132 55922 13184
rect 56781 13175 56839 13181
rect 56781 13141 56793 13175
rect 56827 13172 56839 13175
rect 56962 13172 56968 13184
rect 56827 13144 56968 13172
rect 56827 13141 56839 13144
rect 56781 13135 56839 13141
rect 56962 13132 56968 13144
rect 57020 13132 57026 13184
rect 57072 13172 57100 13212
rect 57238 13200 57244 13212
rect 57296 13200 57302 13252
rect 59170 13240 59176 13252
rect 57348 13212 59176 13240
rect 57348 13172 57376 13212
rect 59170 13200 59176 13212
rect 59228 13200 59234 13252
rect 59372 13240 59400 13348
rect 62224 13348 62488 13376
rect 59446 13268 59452 13320
rect 59504 13308 59510 13320
rect 59633 13311 59691 13317
rect 59633 13308 59645 13311
rect 59504 13280 59645 13308
rect 59504 13268 59510 13280
rect 59633 13277 59645 13280
rect 59679 13277 59691 13311
rect 60642 13308 60648 13320
rect 60603 13280 60648 13308
rect 59633 13271 59691 13277
rect 60642 13268 60648 13280
rect 60700 13268 60706 13320
rect 61565 13311 61623 13317
rect 61565 13277 61577 13311
rect 61611 13308 61623 13311
rect 61654 13308 61660 13320
rect 61611 13280 61660 13308
rect 61611 13277 61623 13280
rect 61565 13271 61623 13277
rect 61654 13268 61660 13280
rect 61712 13268 61718 13320
rect 62224 13317 62252 13348
rect 62482 13336 62488 13348
rect 62540 13336 62546 13388
rect 62942 13336 62948 13388
rect 63000 13376 63006 13388
rect 73982 13376 73988 13388
rect 63000 13348 67220 13376
rect 63000 13336 63006 13348
rect 62209 13311 62267 13317
rect 62209 13277 62221 13311
rect 62255 13277 62267 13311
rect 62209 13271 62267 13277
rect 64598 13268 64604 13320
rect 64656 13308 64662 13320
rect 64693 13311 64751 13317
rect 64693 13308 64705 13311
rect 64656 13280 64705 13308
rect 64656 13268 64662 13280
rect 64693 13277 64705 13280
rect 64739 13308 64751 13311
rect 65978 13308 65984 13320
rect 64739 13280 65984 13308
rect 64739 13277 64751 13280
rect 64693 13271 64751 13277
rect 65978 13268 65984 13280
rect 66036 13268 66042 13320
rect 66162 13268 66168 13320
rect 66220 13308 66226 13320
rect 66441 13311 66499 13317
rect 66441 13308 66453 13311
rect 66220 13280 66453 13308
rect 66220 13268 66226 13280
rect 66441 13277 66453 13280
rect 66487 13277 66499 13311
rect 66441 13271 66499 13277
rect 60660 13240 60688 13268
rect 59372 13212 60688 13240
rect 61746 13200 61752 13252
rect 61804 13240 61810 13252
rect 62485 13243 62543 13249
rect 62485 13240 62497 13243
rect 61804 13212 62497 13240
rect 61804 13200 61810 13212
rect 62485 13209 62497 13212
rect 62531 13209 62543 13243
rect 62485 13203 62543 13209
rect 63494 13200 63500 13252
rect 63552 13200 63558 13252
rect 66622 13240 66628 13252
rect 63972 13212 66628 13240
rect 57072 13144 57376 13172
rect 59078 13132 59084 13184
rect 59136 13172 59142 13184
rect 59541 13175 59599 13181
rect 59541 13172 59553 13175
rect 59136 13144 59553 13172
rect 59136 13132 59142 13144
rect 59541 13141 59553 13144
rect 59587 13141 59599 13175
rect 59541 13135 59599 13141
rect 60734 13132 60740 13184
rect 60792 13172 60798 13184
rect 61657 13175 61715 13181
rect 60792 13144 60837 13172
rect 60792 13132 60798 13144
rect 61657 13141 61669 13175
rect 61703 13172 61715 13175
rect 63310 13172 63316 13184
rect 61703 13144 63316 13172
rect 61703 13141 61715 13144
rect 61657 13135 61715 13141
rect 63310 13132 63316 13144
rect 63368 13132 63374 13184
rect 63402 13132 63408 13184
rect 63460 13172 63466 13184
rect 63972 13181 64000 13212
rect 66622 13200 66628 13212
rect 66680 13200 66686 13252
rect 63957 13175 64015 13181
rect 63957 13172 63969 13175
rect 63460 13144 63969 13172
rect 63460 13132 63466 13144
rect 63957 13141 63969 13144
rect 64003 13141 64015 13175
rect 63957 13135 64015 13141
rect 64601 13175 64659 13181
rect 64601 13141 64613 13175
rect 64647 13172 64659 13175
rect 64690 13172 64696 13184
rect 64647 13144 64696 13172
rect 64647 13141 64659 13144
rect 64601 13135 64659 13141
rect 64690 13132 64696 13144
rect 64748 13132 64754 13184
rect 65886 13172 65892 13184
rect 65847 13144 65892 13172
rect 65886 13132 65892 13144
rect 65944 13132 65950 13184
rect 67082 13172 67088 13184
rect 67043 13144 67088 13172
rect 67082 13132 67088 13144
rect 67140 13132 67146 13184
rect 67192 13172 67220 13348
rect 69400 13348 73988 13376
rect 69400 13317 69428 13348
rect 69385 13311 69443 13317
rect 69385 13277 69397 13311
rect 69431 13277 69443 13311
rect 69842 13308 69848 13320
rect 69803 13280 69848 13308
rect 69385 13271 69443 13277
rect 69842 13268 69848 13280
rect 69900 13268 69906 13320
rect 70302 13268 70308 13320
rect 70360 13308 70366 13320
rect 71133 13311 71191 13317
rect 71133 13308 71145 13311
rect 70360 13280 71145 13308
rect 70360 13268 70366 13280
rect 71133 13277 71145 13280
rect 71179 13277 71191 13311
rect 71133 13271 71191 13277
rect 71593 13311 71651 13317
rect 71593 13277 71605 13311
rect 71639 13277 71651 13311
rect 71593 13271 71651 13277
rect 67821 13243 67879 13249
rect 67821 13209 67833 13243
rect 67867 13240 67879 13243
rect 70320 13240 70348 13268
rect 67867 13212 70348 13240
rect 71608 13240 71636 13271
rect 72970 13268 72976 13320
rect 73028 13268 73034 13320
rect 73816 13317 73844 13348
rect 73982 13336 73988 13348
rect 74040 13336 74046 13388
rect 75549 13379 75607 13385
rect 75549 13345 75561 13379
rect 75595 13376 75607 13379
rect 79594 13376 79600 13388
rect 75595 13348 79600 13376
rect 75595 13345 75607 13348
rect 75549 13339 75607 13345
rect 79594 13336 79600 13348
rect 79652 13336 79658 13388
rect 80057 13379 80115 13385
rect 80057 13345 80069 13379
rect 80103 13376 80115 13379
rect 80103 13348 80284 13376
rect 80103 13345 80115 13348
rect 80057 13339 80115 13345
rect 73801 13311 73859 13317
rect 73801 13277 73813 13311
rect 73847 13277 73859 13311
rect 73801 13271 73859 13277
rect 76285 13311 76343 13317
rect 76285 13277 76297 13311
rect 76331 13308 76343 13311
rect 76558 13308 76564 13320
rect 76331 13280 76564 13308
rect 76331 13277 76343 13280
rect 76285 13271 76343 13277
rect 76558 13268 76564 13280
rect 76616 13268 76622 13320
rect 77018 13308 77024 13320
rect 76979 13280 77024 13308
rect 77018 13268 77024 13280
rect 77076 13268 77082 13320
rect 78950 13268 78956 13320
rect 79008 13308 79014 13320
rect 79410 13308 79416 13320
rect 79008 13280 79416 13308
rect 79008 13268 79014 13280
rect 79410 13268 79416 13280
rect 79468 13308 79474 13320
rect 79505 13311 79563 13317
rect 79505 13308 79517 13311
rect 79468 13280 79517 13308
rect 79468 13268 79474 13280
rect 79505 13277 79517 13280
rect 79551 13277 79563 13311
rect 79612 13308 79640 13336
rect 79957 13311 80015 13317
rect 79957 13308 79969 13311
rect 79612 13280 79969 13308
rect 79505 13271 79563 13277
rect 79957 13277 79969 13280
rect 80003 13277 80015 13311
rect 79957 13271 80015 13277
rect 71774 13240 71780 13252
rect 71608 13212 71780 13240
rect 67867 13209 67879 13212
rect 67821 13203 67879 13209
rect 71774 13200 71780 13212
rect 71832 13200 71838 13252
rect 71869 13243 71927 13249
rect 71869 13209 71881 13243
rect 71915 13209 71927 13243
rect 76834 13240 76840 13252
rect 71869 13203 71927 13209
rect 73172 13212 76840 13240
rect 71682 13172 71688 13184
rect 67192 13144 71688 13172
rect 71682 13132 71688 13144
rect 71740 13132 71746 13184
rect 71884 13172 71912 13203
rect 73172 13172 73200 13212
rect 76834 13200 76840 13212
rect 76892 13200 76898 13252
rect 76926 13200 76932 13252
rect 76984 13240 76990 13252
rect 77297 13243 77355 13249
rect 77297 13240 77309 13243
rect 76984 13212 77309 13240
rect 76984 13200 76990 13212
rect 77297 13209 77309 13212
rect 77343 13209 77355 13243
rect 80256 13240 80284 13348
rect 80330 13336 80336 13388
rect 80388 13376 80394 13388
rect 82909 13379 82967 13385
rect 82909 13376 82921 13379
rect 80388 13348 82921 13376
rect 80388 13336 80394 13348
rect 82909 13345 82921 13348
rect 82955 13376 82967 13379
rect 84212 13376 84240 13416
rect 85669 13413 85681 13416
rect 85715 13413 85727 13447
rect 86681 13447 86739 13453
rect 86681 13444 86693 13447
rect 85669 13407 85727 13413
rect 86328 13416 86693 13444
rect 82955 13348 84240 13376
rect 84657 13379 84715 13385
rect 82955 13345 82967 13348
rect 82909 13339 82967 13345
rect 84657 13345 84669 13379
rect 84703 13376 84715 13379
rect 86218 13376 86224 13388
rect 84703 13348 86224 13376
rect 84703 13345 84715 13348
rect 84657 13339 84715 13345
rect 86218 13336 86224 13348
rect 86276 13336 86282 13388
rect 84470 13268 84476 13320
rect 84528 13308 84534 13320
rect 86328 13308 86356 13416
rect 86681 13413 86693 13416
rect 86727 13413 86739 13447
rect 86681 13407 86739 13413
rect 87693 13379 87751 13385
rect 87693 13345 87705 13379
rect 87739 13376 87751 13379
rect 90453 13379 90511 13385
rect 90453 13376 90465 13379
rect 87739 13348 90465 13376
rect 87739 13345 87751 13348
rect 87693 13339 87751 13345
rect 90453 13345 90465 13348
rect 90499 13345 90511 13379
rect 90453 13339 90511 13345
rect 92566 13336 92572 13388
rect 92624 13376 92630 13388
rect 93581 13379 93639 13385
rect 93581 13376 93593 13379
rect 92624 13348 93593 13376
rect 92624 13336 92630 13348
rect 93581 13345 93593 13348
rect 93627 13345 93639 13379
rect 93581 13339 93639 13345
rect 84528 13280 86356 13308
rect 84528 13268 84534 13280
rect 86402 13268 86408 13320
rect 86460 13308 86466 13320
rect 86678 13308 86684 13320
rect 86460 13280 86684 13308
rect 86460 13268 86466 13280
rect 86678 13268 86684 13280
rect 86736 13308 86742 13320
rect 87417 13311 87475 13317
rect 87417 13308 87429 13311
rect 86736 13280 87429 13308
rect 86736 13268 86742 13280
rect 87417 13277 87429 13280
rect 87463 13277 87475 13311
rect 87417 13271 87475 13277
rect 89070 13268 89076 13320
rect 89128 13308 89134 13320
rect 89717 13311 89775 13317
rect 89717 13308 89729 13311
rect 89128 13280 89729 13308
rect 89128 13268 89134 13280
rect 89717 13277 89729 13280
rect 89763 13277 89775 13311
rect 90542 13308 90548 13320
rect 90503 13280 90548 13308
rect 89717 13271 89775 13277
rect 90542 13268 90548 13280
rect 90600 13268 90606 13320
rect 82357 13243 82415 13249
rect 82357 13240 82369 13243
rect 78522 13212 80284 13240
rect 80532 13212 82369 13240
rect 77297 13203 77355 13209
rect 71884 13144 73200 13172
rect 73246 13132 73252 13184
rect 73304 13172 73310 13184
rect 79870 13172 79876 13184
rect 73304 13144 79876 13172
rect 73304 13132 73310 13144
rect 79870 13132 79876 13144
rect 79928 13132 79934 13184
rect 79962 13132 79968 13184
rect 80020 13172 80026 13184
rect 80532 13172 80560 13212
rect 82357 13209 82369 13212
rect 82403 13209 82415 13243
rect 83182 13240 83188 13252
rect 83143 13212 83188 13240
rect 82357 13203 82415 13209
rect 83182 13200 83188 13212
rect 83240 13200 83246 13252
rect 84562 13240 84568 13252
rect 84410 13212 84568 13240
rect 84562 13200 84568 13212
rect 84620 13200 84626 13252
rect 87782 13200 87788 13252
rect 87840 13240 87846 13252
rect 87840 13212 88182 13240
rect 87840 13200 87846 13212
rect 89438 13200 89444 13252
rect 89496 13240 89502 13252
rect 93302 13240 93308 13252
rect 89496 13212 92138 13240
rect 93263 13212 93308 13240
rect 89496 13200 89502 13212
rect 80020 13144 80560 13172
rect 80020 13132 80026 13144
rect 80606 13132 80612 13184
rect 80664 13172 80670 13184
rect 80664 13144 80709 13172
rect 80664 13132 80670 13144
rect 81158 13132 81164 13184
rect 81216 13172 81222 13184
rect 81345 13175 81403 13181
rect 81345 13172 81357 13175
rect 81216 13144 81357 13172
rect 81216 13132 81222 13144
rect 81345 13141 81357 13144
rect 81391 13172 81403 13175
rect 86494 13172 86500 13184
rect 81391 13144 86500 13172
rect 81391 13141 81403 13144
rect 81345 13135 81403 13141
rect 86494 13132 86500 13144
rect 86552 13132 86558 13184
rect 91830 13172 91836 13184
rect 91791 13144 91836 13172
rect 91830 13132 91836 13144
rect 91888 13132 91894 13184
rect 92032 13172 92060 13212
rect 93302 13200 93308 13212
rect 93360 13200 93366 13252
rect 92566 13172 92572 13184
rect 92032 13144 92572 13172
rect 92566 13132 92572 13144
rect 92624 13172 92630 13184
rect 94041 13175 94099 13181
rect 94041 13172 94053 13175
rect 92624 13144 94053 13172
rect 92624 13132 92630 13144
rect 94041 13141 94053 13144
rect 94087 13141 94099 13175
rect 94041 13135 94099 13141
rect 1104 13082 95011 13104
rect 1104 13030 24386 13082
rect 24438 13030 24450 13082
rect 24502 13030 24514 13082
rect 24566 13030 24578 13082
rect 24630 13030 24642 13082
rect 24694 13030 47823 13082
rect 47875 13030 47887 13082
rect 47939 13030 47951 13082
rect 48003 13030 48015 13082
rect 48067 13030 48079 13082
rect 48131 13030 71260 13082
rect 71312 13030 71324 13082
rect 71376 13030 71388 13082
rect 71440 13030 71452 13082
rect 71504 13030 71516 13082
rect 71568 13030 94697 13082
rect 94749 13030 94761 13082
rect 94813 13030 94825 13082
rect 94877 13030 94889 13082
rect 94941 13030 94953 13082
rect 95005 13030 95011 13082
rect 1104 13008 95011 13030
rect 4430 12968 4436 12980
rect 4391 12940 4436 12968
rect 4430 12928 4436 12940
rect 4488 12928 4494 12980
rect 6546 12968 6552 12980
rect 6507 12940 6552 12968
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 9582 12968 9588 12980
rect 6656 12940 9588 12968
rect 4154 12900 4160 12912
rect 3804 12872 4160 12900
rect 3804 12841 3832 12872
rect 4154 12860 4160 12872
rect 4212 12900 4218 12912
rect 6656 12900 6684 12940
rect 9582 12928 9588 12940
rect 9640 12928 9646 12980
rect 9953 12971 10011 12977
rect 9953 12937 9965 12971
rect 9999 12937 10011 12971
rect 11882 12968 11888 12980
rect 11843 12940 11888 12968
rect 9953 12931 10011 12937
rect 7650 12900 7656 12912
rect 4212 12872 6684 12900
rect 6748 12872 7656 12900
rect 4212 12860 4218 12872
rect 3789 12835 3847 12841
rect 3789 12801 3801 12835
rect 3835 12801 3847 12835
rect 3789 12795 3847 12801
rect 4985 12835 5043 12841
rect 4985 12801 4997 12835
rect 5031 12832 5043 12835
rect 5074 12832 5080 12844
rect 5031 12804 5080 12832
rect 5031 12801 5043 12804
rect 4985 12795 5043 12801
rect 5074 12792 5080 12804
rect 5132 12792 5138 12844
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12764 3939 12767
rect 5166 12764 5172 12776
rect 3927 12736 5172 12764
rect 3927 12733 3939 12736
rect 3881 12727 3939 12733
rect 5166 12724 5172 12736
rect 5224 12764 5230 12776
rect 6748 12764 6776 12872
rect 7650 12860 7656 12872
rect 7708 12860 7714 12912
rect 8938 12860 8944 12912
rect 8996 12900 9002 12912
rect 9968 12900 9996 12931
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 13262 12928 13268 12980
rect 13320 12968 13326 12980
rect 21450 12968 21456 12980
rect 13320 12940 21456 12968
rect 13320 12928 13326 12940
rect 21450 12928 21456 12940
rect 21508 12928 21514 12980
rect 22572 12940 25268 12968
rect 14274 12900 14280 12912
rect 8996 12872 9812 12900
rect 9968 12872 14280 12900
rect 8996 12860 9002 12872
rect 6822 12792 6828 12844
rect 6880 12832 6886 12844
rect 6917 12835 6975 12841
rect 6917 12832 6929 12835
rect 6880 12804 6929 12832
rect 6880 12792 6886 12804
rect 6917 12801 6929 12804
rect 6963 12801 6975 12835
rect 6917 12795 6975 12801
rect 7745 12835 7803 12841
rect 7745 12801 7757 12835
rect 7791 12832 7803 12835
rect 8573 12835 8631 12841
rect 8573 12832 8585 12835
rect 7791 12804 8585 12832
rect 7791 12801 7803 12804
rect 7745 12795 7803 12801
rect 8573 12801 8585 12804
rect 8619 12832 8631 12835
rect 8662 12832 8668 12844
rect 8619 12804 8668 12832
rect 8619 12801 8631 12804
rect 8573 12795 8631 12801
rect 8662 12792 8668 12804
rect 8720 12792 8726 12844
rect 9582 12832 9588 12844
rect 9495 12804 9588 12832
rect 9582 12792 9588 12804
rect 9640 12792 9646 12844
rect 9784 12832 9812 12872
rect 14274 12860 14280 12872
rect 14332 12860 14338 12912
rect 14737 12903 14795 12909
rect 14737 12869 14749 12903
rect 14783 12900 14795 12903
rect 15010 12900 15016 12912
rect 14783 12872 15016 12900
rect 14783 12869 14795 12872
rect 14737 12863 14795 12869
rect 15010 12860 15016 12872
rect 15068 12860 15074 12912
rect 16850 12860 16856 12912
rect 16908 12900 16914 12912
rect 16945 12903 17003 12909
rect 16945 12900 16957 12903
rect 16908 12872 16957 12900
rect 16908 12860 16914 12872
rect 16945 12869 16957 12872
rect 16991 12900 17003 12903
rect 21085 12903 21143 12909
rect 16991 12872 20576 12900
rect 16991 12869 17003 12872
rect 16945 12863 17003 12869
rect 11701 12835 11759 12841
rect 11701 12832 11713 12835
rect 9784 12804 11713 12832
rect 11701 12801 11713 12804
rect 11747 12801 11759 12835
rect 13906 12832 13912 12844
rect 13867 12804 13912 12832
rect 11701 12795 11759 12801
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 15838 12792 15844 12844
rect 15896 12792 15902 12844
rect 17957 12835 18015 12841
rect 17957 12801 17969 12835
rect 18003 12832 18015 12835
rect 18509 12835 18567 12841
rect 18509 12832 18521 12835
rect 18003 12804 18521 12832
rect 18003 12801 18015 12804
rect 17957 12795 18015 12801
rect 18509 12801 18521 12804
rect 18555 12801 18567 12835
rect 20438 12832 20444 12844
rect 18509 12795 18567 12801
rect 19076 12804 20444 12832
rect 7006 12764 7012 12776
rect 5224 12736 6776 12764
rect 6967 12736 7012 12764
rect 5224 12724 5230 12736
rect 7006 12724 7012 12736
rect 7064 12724 7070 12776
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12764 7895 12767
rect 7926 12764 7932 12776
rect 7883 12736 7932 12764
rect 7883 12733 7895 12736
rect 7837 12727 7895 12733
rect 7926 12724 7932 12736
rect 7984 12724 7990 12776
rect 8110 12764 8116 12776
rect 8071 12736 8116 12764
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 8478 12724 8484 12776
rect 8536 12764 8542 12776
rect 9493 12767 9551 12773
rect 9493 12764 9505 12767
rect 8536 12736 9505 12764
rect 8536 12724 8542 12736
rect 9493 12733 9505 12736
rect 9539 12733 9551 12767
rect 9600 12764 9628 12792
rect 10502 12764 10508 12776
rect 9600 12736 10508 12764
rect 9493 12727 9551 12733
rect 10502 12724 10508 12736
rect 10560 12724 10566 12776
rect 14461 12767 14519 12773
rect 14461 12764 14473 12767
rect 12406 12736 14473 12764
rect 3418 12656 3424 12708
rect 3476 12696 3482 12708
rect 12406 12696 12434 12736
rect 14461 12733 14473 12736
rect 14507 12733 14519 12767
rect 14461 12727 14519 12733
rect 15102 12724 15108 12776
rect 15160 12764 15166 12776
rect 17972 12764 18000 12795
rect 15160 12736 18000 12764
rect 15160 12724 15166 12736
rect 19076 12696 19104 12804
rect 20438 12792 20444 12804
rect 20496 12792 20502 12844
rect 20548 12764 20576 12872
rect 21085 12869 21097 12903
rect 21131 12900 21143 12903
rect 22370 12900 22376 12912
rect 21131 12872 22376 12900
rect 21131 12869 21143 12872
rect 21085 12863 21143 12869
rect 22370 12860 22376 12872
rect 22428 12860 22434 12912
rect 21266 12792 21272 12844
rect 21324 12832 21330 12844
rect 22572 12841 22600 12940
rect 23198 12860 23204 12912
rect 23256 12900 23262 12912
rect 24489 12903 24547 12909
rect 23256 12872 23322 12900
rect 23256 12860 23262 12872
rect 24489 12869 24501 12903
rect 24535 12900 24547 12903
rect 25130 12900 25136 12912
rect 24535 12872 25136 12900
rect 24535 12869 24547 12872
rect 24489 12863 24547 12869
rect 25130 12860 25136 12872
rect 25188 12860 25194 12912
rect 25240 12847 25268 12940
rect 26142 12928 26148 12980
rect 26200 12968 26206 12980
rect 30466 12968 30472 12980
rect 26200 12940 29316 12968
rect 30427 12940 30472 12968
rect 26200 12928 26206 12940
rect 25314 12860 25320 12912
rect 25372 12900 25378 12912
rect 29288 12909 29316 12940
rect 30466 12928 30472 12940
rect 30524 12928 30530 12980
rect 30558 12928 30564 12980
rect 30616 12968 30622 12980
rect 45462 12968 45468 12980
rect 30616 12940 45324 12968
rect 45423 12940 45468 12968
rect 30616 12928 30622 12940
rect 29273 12903 29331 12909
rect 25372 12872 29224 12900
rect 25372 12860 25378 12872
rect 25225 12841 25283 12847
rect 22557 12835 22615 12841
rect 22557 12832 22569 12835
rect 21324 12804 22569 12832
rect 21324 12792 21330 12804
rect 22557 12801 22569 12804
rect 22603 12801 22615 12835
rect 25225 12807 25237 12841
rect 25271 12807 25283 12841
rect 26234 12832 26240 12844
rect 25225 12801 25283 12807
rect 26195 12804 26240 12832
rect 22557 12795 22615 12801
rect 26234 12792 26240 12804
rect 26292 12792 26298 12844
rect 27338 12832 27344 12844
rect 26344 12804 27344 12832
rect 26344 12776 26372 12804
rect 27338 12792 27344 12804
rect 27396 12792 27402 12844
rect 22186 12764 22192 12776
rect 20548 12736 22192 12764
rect 22186 12724 22192 12736
rect 22244 12724 22250 12776
rect 24765 12767 24823 12773
rect 23492 12736 24716 12764
rect 3476 12668 12434 12696
rect 16132 12668 19104 12696
rect 3476 12656 3482 12668
rect 5261 12631 5319 12637
rect 5261 12597 5273 12631
rect 5307 12628 5319 12631
rect 5626 12628 5632 12640
rect 5307 12600 5632 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 5626 12588 5632 12600
rect 5684 12588 5690 12640
rect 5810 12588 5816 12640
rect 5868 12628 5874 12640
rect 5997 12631 6055 12637
rect 5997 12628 6009 12631
rect 5868 12600 6009 12628
rect 5868 12588 5874 12600
rect 5997 12597 6009 12600
rect 6043 12628 6055 12631
rect 11146 12628 11152 12640
rect 6043 12600 11152 12628
rect 6043 12597 6055 12600
rect 5997 12591 6055 12597
rect 11146 12588 11152 12600
rect 11204 12588 11210 12640
rect 12526 12588 12532 12640
rect 12584 12628 12590 12640
rect 13173 12631 13231 12637
rect 13173 12628 13185 12631
rect 12584 12600 13185 12628
rect 12584 12588 12590 12600
rect 13173 12597 13185 12600
rect 13219 12597 13231 12631
rect 13814 12628 13820 12640
rect 13775 12600 13820 12628
rect 13173 12591 13231 12597
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 13998 12588 14004 12640
rect 14056 12628 14062 12640
rect 16132 12628 16160 12668
rect 19150 12656 19156 12708
rect 19208 12696 19214 12708
rect 23492 12696 23520 12736
rect 19208 12668 23520 12696
rect 24688 12696 24716 12736
rect 24765 12733 24777 12767
rect 24811 12764 24823 12767
rect 25317 12767 25375 12773
rect 25317 12764 25329 12767
rect 24811 12736 25329 12764
rect 24811 12733 24823 12736
rect 24765 12727 24823 12733
rect 25317 12733 25329 12736
rect 25363 12733 25375 12767
rect 26326 12764 26332 12776
rect 26287 12736 26332 12764
rect 25317 12727 25375 12733
rect 26326 12724 26332 12736
rect 26384 12724 26390 12776
rect 26605 12767 26663 12773
rect 26605 12733 26617 12767
rect 26651 12764 26663 12767
rect 27154 12764 27160 12776
rect 26651 12736 27160 12764
rect 26651 12733 26663 12736
rect 26605 12727 26663 12733
rect 27154 12724 27160 12736
rect 27212 12724 27218 12776
rect 27433 12767 27491 12773
rect 27433 12733 27445 12767
rect 27479 12733 27491 12767
rect 27433 12727 27491 12733
rect 27617 12767 27675 12773
rect 27617 12733 27629 12767
rect 27663 12764 27675 12767
rect 27663 12736 29040 12764
rect 27663 12733 27675 12736
rect 27617 12727 27675 12733
rect 27448 12696 27476 12727
rect 24688 12668 27660 12696
rect 19208 12656 19214 12668
rect 27632 12640 27660 12668
rect 14056 12600 16160 12628
rect 16209 12631 16267 12637
rect 14056 12588 14062 12600
rect 16209 12597 16221 12631
rect 16255 12628 16267 12631
rect 16298 12628 16304 12640
rect 16255 12600 16304 12628
rect 16255 12597 16267 12600
rect 16209 12591 16267 12597
rect 16298 12588 16304 12600
rect 16356 12588 16362 12640
rect 16850 12588 16856 12640
rect 16908 12628 16914 12640
rect 17037 12631 17095 12637
rect 17037 12628 17049 12631
rect 16908 12600 17049 12628
rect 16908 12588 16914 12600
rect 17037 12597 17049 12600
rect 17083 12597 17095 12631
rect 17037 12591 17095 12597
rect 17494 12588 17500 12640
rect 17552 12628 17558 12640
rect 17865 12631 17923 12637
rect 17865 12628 17877 12631
rect 17552 12600 17877 12628
rect 17552 12588 17558 12600
rect 17865 12597 17877 12600
rect 17911 12597 17923 12631
rect 18598 12628 18604 12640
rect 18559 12600 18604 12628
rect 17865 12591 17923 12597
rect 18598 12588 18604 12600
rect 18656 12588 18662 12640
rect 19610 12628 19616 12640
rect 19571 12600 19616 12628
rect 19610 12588 19616 12600
rect 19668 12588 19674 12640
rect 22278 12588 22284 12640
rect 22336 12628 22342 12640
rect 22465 12631 22523 12637
rect 22465 12628 22477 12631
rect 22336 12600 22477 12628
rect 22336 12588 22342 12600
rect 22465 12597 22477 12600
rect 22511 12597 22523 12631
rect 22465 12591 22523 12597
rect 23017 12631 23075 12637
rect 23017 12597 23029 12631
rect 23063 12628 23075 12631
rect 27246 12628 27252 12640
rect 23063 12600 27252 12628
rect 23063 12597 23075 12600
rect 23017 12591 23075 12597
rect 27246 12588 27252 12600
rect 27304 12588 27310 12640
rect 27614 12588 27620 12640
rect 27672 12588 27678 12640
rect 29012 12628 29040 12736
rect 29196 12696 29224 12872
rect 29273 12869 29285 12903
rect 29319 12900 29331 12903
rect 32398 12900 32404 12912
rect 29319 12872 30328 12900
rect 29319 12869 29331 12872
rect 29273 12863 29331 12869
rect 29546 12792 29552 12844
rect 29604 12832 29610 12844
rect 30098 12832 30104 12844
rect 29604 12804 30104 12832
rect 29604 12792 29610 12804
rect 30098 12792 30104 12804
rect 30156 12792 30162 12844
rect 29270 12724 29276 12776
rect 29328 12764 29334 12776
rect 29822 12764 29828 12776
rect 29328 12736 29828 12764
rect 29328 12724 29334 12736
rect 29822 12724 29828 12736
rect 29880 12724 29886 12776
rect 30300 12764 30328 12872
rect 30392 12872 32404 12900
rect 30392 12841 30420 12872
rect 32398 12860 32404 12872
rect 32456 12860 32462 12912
rect 32858 12900 32864 12912
rect 32819 12872 32864 12900
rect 32858 12860 32864 12872
rect 32916 12860 32922 12912
rect 33318 12860 33324 12912
rect 33376 12860 33382 12912
rect 38654 12900 38660 12912
rect 38615 12872 38660 12900
rect 38654 12860 38660 12872
rect 38712 12860 38718 12912
rect 40126 12900 40132 12912
rect 39882 12872 40132 12900
rect 40126 12860 40132 12872
rect 40184 12860 40190 12912
rect 44177 12903 44235 12909
rect 41708 12872 44128 12900
rect 41708 12844 41736 12872
rect 30377 12835 30435 12841
rect 30377 12801 30389 12835
rect 30423 12801 30435 12835
rect 30377 12795 30435 12801
rect 30466 12792 30472 12844
rect 30524 12832 30530 12844
rect 31294 12832 31300 12844
rect 30524 12804 31300 12832
rect 30524 12792 30530 12804
rect 31294 12792 31300 12804
rect 31352 12792 31358 12844
rect 31386 12792 31392 12844
rect 31444 12832 31450 12844
rect 31573 12835 31631 12841
rect 31573 12832 31585 12835
rect 31444 12804 31585 12832
rect 31444 12792 31450 12804
rect 31573 12801 31585 12804
rect 31619 12832 31631 12835
rect 32582 12832 32588 12844
rect 31619 12804 32444 12832
rect 32543 12804 32588 12832
rect 31619 12801 31631 12804
rect 31573 12795 31631 12801
rect 31478 12764 31484 12776
rect 30300 12736 31484 12764
rect 31478 12724 31484 12736
rect 31536 12724 31542 12776
rect 31662 12764 31668 12776
rect 31623 12736 31668 12764
rect 31662 12724 31668 12736
rect 31720 12724 31726 12776
rect 32416 12764 32444 12804
rect 32582 12792 32588 12804
rect 32640 12792 32646 12844
rect 34974 12832 34980 12844
rect 34935 12804 34980 12832
rect 34974 12792 34980 12804
rect 35032 12792 35038 12844
rect 35161 12835 35219 12841
rect 35161 12801 35173 12835
rect 35207 12832 35219 12835
rect 35526 12832 35532 12844
rect 35207 12804 35532 12832
rect 35207 12801 35219 12804
rect 35161 12795 35219 12801
rect 35526 12792 35532 12804
rect 35584 12792 35590 12844
rect 35897 12835 35955 12841
rect 35897 12801 35909 12835
rect 35943 12801 35955 12835
rect 37734 12832 37740 12844
rect 37695 12804 37740 12832
rect 35897 12795 35955 12801
rect 35618 12764 35624 12776
rect 32416 12736 35624 12764
rect 35618 12724 35624 12736
rect 35676 12724 35682 12776
rect 31386 12696 31392 12708
rect 29196 12668 31392 12696
rect 31386 12656 31392 12668
rect 31444 12656 31450 12708
rect 35161 12699 35219 12705
rect 35161 12696 35173 12699
rect 33888 12668 35173 12696
rect 30834 12628 30840 12640
rect 29012 12600 30840 12628
rect 30834 12588 30840 12600
rect 30892 12588 30898 12640
rect 31294 12628 31300 12640
rect 31255 12600 31300 12628
rect 31294 12588 31300 12600
rect 31352 12588 31358 12640
rect 33594 12588 33600 12640
rect 33652 12628 33658 12640
rect 33888 12628 33916 12668
rect 35161 12665 35173 12668
rect 35207 12665 35219 12699
rect 35161 12659 35219 12665
rect 33652 12600 33916 12628
rect 33652 12588 33658 12600
rect 33962 12588 33968 12640
rect 34020 12628 34026 12640
rect 34333 12631 34391 12637
rect 34333 12628 34345 12631
rect 34020 12600 34345 12628
rect 34020 12588 34026 12600
rect 34333 12597 34345 12600
rect 34379 12628 34391 12631
rect 35912 12628 35940 12795
rect 37734 12792 37740 12804
rect 37792 12792 37798 12844
rect 39942 12792 39948 12844
rect 40000 12832 40006 12844
rect 41690 12832 41696 12844
rect 40000 12804 41696 12832
rect 40000 12792 40006 12804
rect 41690 12792 41696 12804
rect 41748 12792 41754 12844
rect 42797 12835 42855 12841
rect 42797 12801 42809 12835
rect 42843 12832 42855 12835
rect 43070 12832 43076 12844
rect 42843 12804 43076 12832
rect 42843 12801 42855 12804
rect 42797 12795 42855 12801
rect 43070 12792 43076 12804
rect 43128 12832 43134 12844
rect 43990 12832 43996 12844
rect 43128 12804 43996 12832
rect 43128 12792 43134 12804
rect 43990 12792 43996 12804
rect 44048 12792 44054 12844
rect 44100 12832 44128 12872
rect 44177 12869 44189 12903
rect 44223 12900 44235 12903
rect 44726 12900 44732 12912
rect 44223 12872 44732 12900
rect 44223 12869 44235 12872
rect 44177 12863 44235 12869
rect 44726 12860 44732 12872
rect 44784 12860 44790 12912
rect 45296 12900 45324 12940
rect 45462 12928 45468 12940
rect 45520 12928 45526 12980
rect 45922 12928 45928 12980
rect 45980 12968 45986 12980
rect 46474 12968 46480 12980
rect 45980 12940 46480 12968
rect 45980 12928 45986 12940
rect 46474 12928 46480 12940
rect 46532 12928 46538 12980
rect 46934 12928 46940 12980
rect 46992 12968 46998 12980
rect 47765 12971 47823 12977
rect 47765 12968 47777 12971
rect 46992 12940 47777 12968
rect 46992 12928 46998 12940
rect 47765 12937 47777 12940
rect 47811 12937 47823 12971
rect 47765 12931 47823 12937
rect 50338 12928 50344 12980
rect 50396 12968 50402 12980
rect 51994 12968 52000 12980
rect 50396 12940 52000 12968
rect 50396 12928 50402 12940
rect 51994 12928 52000 12940
rect 52052 12928 52058 12980
rect 53377 12971 53435 12977
rect 53377 12937 53389 12971
rect 53423 12968 53435 12971
rect 53742 12968 53748 12980
rect 53423 12940 53748 12968
rect 53423 12937 53435 12940
rect 53377 12931 53435 12937
rect 53742 12928 53748 12940
rect 53800 12928 53806 12980
rect 55030 12968 55036 12980
rect 54588 12940 55036 12968
rect 54588 12900 54616 12940
rect 55030 12928 55036 12940
rect 55088 12968 55094 12980
rect 55950 12968 55956 12980
rect 55088 12940 55956 12968
rect 55088 12928 55094 12940
rect 55950 12928 55956 12940
rect 56008 12968 56014 12980
rect 56781 12971 56839 12977
rect 56008 12940 56732 12968
rect 56008 12928 56014 12940
rect 45296 12872 54616 12900
rect 54665 12903 54723 12909
rect 54665 12869 54677 12903
rect 54711 12900 54723 12903
rect 56594 12900 56600 12912
rect 54711 12872 56600 12900
rect 54711 12869 54723 12872
rect 54665 12863 54723 12869
rect 56594 12860 56600 12872
rect 56652 12860 56658 12912
rect 56704 12900 56732 12940
rect 56781 12937 56793 12971
rect 56827 12968 56839 12971
rect 57146 12968 57152 12980
rect 56827 12940 57152 12968
rect 56827 12937 56839 12940
rect 56781 12931 56839 12937
rect 57146 12928 57152 12940
rect 57204 12968 57210 12980
rect 60366 12968 60372 12980
rect 57204 12940 60372 12968
rect 57204 12928 57210 12940
rect 60366 12928 60372 12940
rect 60424 12928 60430 12980
rect 60642 12928 60648 12980
rect 60700 12968 60706 12980
rect 61286 12968 61292 12980
rect 60700 12940 61292 12968
rect 60700 12928 60706 12940
rect 61286 12928 61292 12940
rect 61344 12928 61350 12980
rect 61562 12968 61568 12980
rect 61523 12940 61568 12968
rect 61562 12928 61568 12940
rect 61620 12928 61626 12980
rect 62114 12928 62120 12980
rect 62172 12968 62178 12980
rect 64969 12971 65027 12977
rect 64969 12968 64981 12971
rect 62172 12940 64981 12968
rect 62172 12928 62178 12940
rect 64969 12937 64981 12940
rect 65015 12968 65027 12971
rect 66530 12968 66536 12980
rect 65015 12940 66300 12968
rect 66491 12940 66536 12968
rect 65015 12937 65027 12940
rect 64969 12931 65027 12937
rect 59354 12900 59360 12912
rect 56704 12872 59360 12900
rect 59354 12860 59360 12872
rect 59412 12860 59418 12912
rect 60734 12860 60740 12912
rect 60792 12900 60798 12912
rect 63497 12903 63555 12909
rect 63497 12900 63509 12903
rect 60792 12872 63509 12900
rect 60792 12860 60798 12872
rect 63497 12869 63509 12872
rect 63543 12869 63555 12903
rect 65886 12900 65892 12912
rect 64722 12872 65892 12900
rect 63497 12863 63555 12869
rect 65886 12860 65892 12872
rect 65944 12860 65950 12912
rect 44266 12832 44272 12844
rect 44100 12804 44272 12832
rect 44266 12792 44272 12804
rect 44324 12832 44330 12844
rect 44818 12832 44824 12844
rect 44324 12804 44824 12832
rect 44324 12792 44330 12804
rect 44818 12792 44824 12804
rect 44876 12792 44882 12844
rect 46750 12832 46756 12844
rect 46711 12804 46756 12832
rect 46750 12792 46756 12804
rect 46808 12792 46814 12844
rect 48130 12832 48136 12844
rect 46860 12804 47164 12832
rect 48091 12804 48136 12832
rect 36173 12767 36231 12773
rect 36173 12733 36185 12767
rect 36219 12764 36231 12767
rect 36998 12764 37004 12776
rect 36219 12736 37004 12764
rect 36219 12733 36231 12736
rect 36173 12727 36231 12733
rect 36998 12724 37004 12736
rect 37056 12724 37062 12776
rect 37274 12724 37280 12776
rect 37332 12764 37338 12776
rect 38381 12767 38439 12773
rect 38381 12764 38393 12767
rect 37332 12736 38393 12764
rect 37332 12724 37338 12736
rect 38381 12733 38393 12736
rect 38427 12764 38439 12767
rect 39298 12764 39304 12776
rect 38427 12736 39304 12764
rect 38427 12733 38439 12736
rect 38381 12727 38439 12733
rect 39298 12724 39304 12736
rect 39356 12724 39362 12776
rect 39390 12724 39396 12776
rect 39448 12764 39454 12776
rect 40129 12767 40187 12773
rect 40129 12764 40141 12767
rect 39448 12736 40141 12764
rect 39448 12724 39454 12736
rect 40129 12733 40141 12736
rect 40175 12733 40187 12767
rect 40129 12727 40187 12733
rect 41598 12724 41604 12776
rect 41656 12764 41662 12776
rect 41785 12767 41843 12773
rect 41785 12764 41797 12767
rect 41656 12736 41797 12764
rect 41656 12724 41662 12736
rect 41785 12733 41797 12736
rect 41831 12764 41843 12767
rect 42334 12764 42340 12776
rect 41831 12736 42340 12764
rect 41831 12733 41843 12736
rect 41785 12727 41843 12733
rect 42334 12724 42340 12736
rect 42392 12724 42398 12776
rect 42886 12764 42892 12776
rect 42847 12736 42892 12764
rect 42886 12724 42892 12736
rect 42944 12724 42950 12776
rect 46860 12764 46888 12804
rect 47026 12764 47032 12776
rect 42996 12736 46888 12764
rect 46987 12736 47032 12764
rect 40034 12656 40040 12708
rect 40092 12696 40098 12708
rect 42996 12696 43024 12736
rect 47026 12724 47032 12736
rect 47084 12724 47090 12776
rect 47136 12764 47164 12804
rect 48130 12792 48136 12804
rect 48188 12792 48194 12844
rect 48958 12832 48964 12844
rect 48919 12804 48964 12832
rect 48958 12792 48964 12804
rect 49016 12792 49022 12844
rect 49326 12832 49332 12844
rect 49287 12804 49332 12832
rect 49326 12792 49332 12804
rect 49384 12792 49390 12844
rect 50893 12835 50951 12841
rect 50893 12801 50905 12835
rect 50939 12832 50951 12835
rect 51718 12832 51724 12844
rect 50939 12804 51724 12832
rect 50939 12801 50951 12804
rect 50893 12795 50951 12801
rect 51718 12792 51724 12804
rect 51776 12792 51782 12844
rect 51813 12835 51871 12841
rect 51813 12801 51825 12835
rect 51859 12832 51871 12835
rect 51994 12832 52000 12844
rect 51859 12804 52000 12832
rect 51859 12801 51871 12804
rect 51813 12795 51871 12801
rect 51994 12792 52000 12804
rect 52052 12792 52058 12844
rect 55030 12792 55036 12844
rect 55088 12832 55094 12844
rect 55401 12835 55459 12841
rect 55401 12832 55413 12835
rect 55088 12804 55413 12832
rect 55088 12792 55094 12804
rect 55401 12801 55413 12804
rect 55447 12801 55459 12835
rect 55401 12795 55459 12801
rect 58069 12835 58127 12841
rect 58069 12801 58081 12835
rect 58115 12832 58127 12835
rect 58710 12832 58716 12844
rect 58115 12804 58716 12832
rect 58115 12801 58127 12804
rect 58069 12795 58127 12801
rect 58710 12792 58716 12804
rect 58768 12792 58774 12844
rect 59078 12832 59084 12844
rect 59039 12804 59084 12832
rect 59078 12792 59084 12804
rect 59136 12792 59142 12844
rect 61010 12832 61016 12844
rect 60490 12804 61016 12832
rect 61010 12792 61016 12804
rect 61068 12792 61074 12844
rect 61105 12835 61163 12841
rect 61105 12801 61117 12835
rect 61151 12832 61163 12835
rect 62022 12832 62028 12844
rect 61151 12804 62028 12832
rect 61151 12801 61163 12804
rect 61105 12795 61163 12801
rect 62022 12792 62028 12804
rect 62080 12792 62086 12844
rect 63218 12832 63224 12844
rect 63179 12804 63224 12832
rect 63218 12792 63224 12804
rect 63276 12792 63282 12844
rect 65521 12835 65579 12841
rect 65521 12801 65533 12835
rect 65567 12832 65579 12835
rect 66162 12832 66168 12844
rect 65567 12804 66168 12832
rect 65567 12801 65579 12804
rect 65521 12795 65579 12801
rect 66162 12792 66168 12804
rect 66220 12792 66226 12844
rect 66272 12832 66300 12940
rect 66530 12928 66536 12940
rect 66588 12928 66594 12980
rect 66622 12928 66628 12980
rect 66680 12968 66686 12980
rect 76926 12968 76932 12980
rect 66680 12940 76788 12968
rect 76887 12940 76932 12968
rect 66680 12928 66686 12940
rect 66714 12860 66720 12912
rect 66772 12900 66778 12912
rect 66772 12872 68692 12900
rect 66772 12860 66778 12872
rect 66441 12835 66499 12841
rect 66441 12832 66453 12835
rect 66272 12804 66453 12832
rect 66441 12801 66453 12804
rect 66487 12801 66499 12835
rect 66441 12795 66499 12801
rect 66898 12792 66904 12844
rect 66956 12832 66962 12844
rect 67545 12835 67603 12841
rect 67545 12832 67557 12835
rect 66956 12804 67557 12832
rect 66956 12792 66962 12804
rect 67545 12801 67557 12804
rect 67591 12801 67603 12835
rect 67545 12795 67603 12801
rect 67637 12835 67695 12841
rect 67637 12801 67649 12835
rect 67683 12832 67695 12835
rect 67818 12832 67824 12844
rect 67683 12804 67824 12832
rect 67683 12801 67695 12804
rect 67637 12795 67695 12801
rect 67818 12792 67824 12804
rect 67876 12792 67882 12844
rect 67910 12792 67916 12844
rect 67968 12832 67974 12844
rect 68373 12835 68431 12841
rect 68373 12832 68385 12835
rect 67968 12804 68385 12832
rect 67968 12792 67974 12804
rect 68373 12801 68385 12804
rect 68419 12832 68431 12835
rect 68462 12832 68468 12844
rect 68419 12804 68468 12832
rect 68419 12801 68431 12804
rect 68373 12795 68431 12801
rect 68462 12792 68468 12804
rect 68520 12792 68526 12844
rect 68664 12841 68692 12872
rect 69014 12860 69020 12912
rect 69072 12900 69078 12912
rect 70762 12900 70768 12912
rect 69072 12872 70394 12900
rect 70723 12872 70768 12900
rect 69072 12860 69078 12872
rect 68649 12835 68707 12841
rect 68649 12801 68661 12835
rect 68695 12832 68707 12835
rect 68695 12804 68784 12832
rect 68695 12801 68707 12804
rect 68649 12795 68707 12801
rect 48041 12767 48099 12773
rect 48041 12764 48053 12767
rect 47136 12736 48053 12764
rect 48041 12733 48053 12736
rect 48087 12764 48099 12767
rect 49694 12764 49700 12776
rect 48087 12736 49700 12764
rect 48087 12733 48099 12736
rect 48041 12727 48099 12733
rect 49694 12724 49700 12736
rect 49752 12724 49758 12776
rect 49970 12724 49976 12776
rect 50028 12764 50034 12776
rect 50065 12767 50123 12773
rect 50065 12764 50077 12767
rect 50028 12736 50077 12764
rect 50028 12724 50034 12736
rect 50065 12733 50077 12736
rect 50111 12733 50123 12767
rect 50065 12727 50123 12733
rect 50985 12767 51043 12773
rect 50985 12733 50997 12767
rect 51031 12764 51043 12767
rect 51166 12764 51172 12776
rect 51031 12736 51172 12764
rect 51031 12733 51043 12736
rect 50985 12727 51043 12733
rect 51166 12724 51172 12736
rect 51224 12764 51230 12776
rect 51626 12764 51632 12776
rect 51224 12736 51632 12764
rect 51224 12724 51230 12736
rect 51626 12724 51632 12736
rect 51684 12724 51690 12776
rect 51905 12767 51963 12773
rect 51905 12733 51917 12767
rect 51951 12764 51963 12767
rect 52178 12764 52184 12776
rect 51951 12736 52184 12764
rect 51951 12733 51963 12736
rect 51905 12727 51963 12733
rect 52178 12724 52184 12736
rect 52236 12724 52242 12776
rect 54846 12724 54852 12776
rect 54904 12764 54910 12776
rect 55309 12767 55367 12773
rect 55309 12764 55321 12767
rect 54904 12736 55321 12764
rect 54904 12724 54910 12736
rect 55309 12733 55321 12736
rect 55355 12733 55367 12767
rect 56226 12764 56232 12776
rect 56187 12736 56232 12764
rect 55309 12727 55367 12733
rect 56226 12724 56232 12736
rect 56284 12724 56290 12776
rect 56870 12764 56876 12776
rect 56336 12736 56876 12764
rect 43162 12696 43168 12708
rect 40092 12668 43024 12696
rect 43123 12668 43168 12696
rect 40092 12656 40098 12668
rect 43162 12656 43168 12668
rect 43220 12656 43226 12708
rect 43254 12656 43260 12708
rect 43312 12696 43318 12708
rect 55398 12696 55404 12708
rect 43312 12668 55404 12696
rect 43312 12656 43318 12668
rect 55398 12656 55404 12668
rect 55456 12656 55462 12708
rect 55508 12668 56180 12696
rect 36906 12628 36912 12640
rect 34379 12600 35940 12628
rect 36867 12600 36912 12628
rect 34379 12597 34391 12600
rect 34333 12591 34391 12597
rect 36906 12588 36912 12600
rect 36964 12588 36970 12640
rect 37829 12631 37887 12637
rect 37829 12597 37841 12631
rect 37875 12628 37887 12631
rect 39206 12628 39212 12640
rect 37875 12600 39212 12628
rect 37875 12597 37887 12600
rect 37829 12591 37887 12597
rect 39206 12588 39212 12600
rect 39264 12588 39270 12640
rect 41049 12631 41107 12637
rect 41049 12597 41061 12631
rect 41095 12628 41107 12631
rect 41690 12628 41696 12640
rect 41095 12600 41696 12628
rect 41095 12597 41107 12600
rect 41049 12591 41107 12597
rect 41690 12588 41696 12600
rect 41748 12588 41754 12640
rect 41782 12588 41788 12640
rect 41840 12628 41846 12640
rect 41969 12631 42027 12637
rect 41969 12628 41981 12631
rect 41840 12600 41981 12628
rect 41840 12588 41846 12600
rect 41969 12597 41981 12600
rect 42015 12597 42027 12631
rect 41969 12591 42027 12597
rect 43717 12631 43775 12637
rect 43717 12597 43729 12631
rect 43763 12628 43775 12631
rect 43898 12628 43904 12640
rect 43763 12600 43904 12628
rect 43763 12597 43775 12600
rect 43717 12591 43775 12597
rect 43898 12588 43904 12600
rect 43956 12588 43962 12640
rect 43990 12588 43996 12640
rect 44048 12628 44054 12640
rect 47026 12628 47032 12640
rect 44048 12600 47032 12628
rect 44048 12588 44054 12600
rect 47026 12588 47032 12600
rect 47084 12628 47090 12640
rect 50338 12628 50344 12640
rect 47084 12600 50344 12628
rect 47084 12588 47090 12600
rect 50338 12588 50344 12600
rect 50396 12588 50402 12640
rect 52181 12631 52239 12637
rect 52181 12597 52193 12631
rect 52227 12628 52239 12631
rect 55508 12628 55536 12668
rect 52227 12600 55536 12628
rect 56152 12628 56180 12668
rect 56336 12628 56364 12736
rect 56870 12724 56876 12736
rect 56928 12724 56934 12776
rect 58161 12767 58219 12773
rect 58161 12733 58173 12767
rect 58207 12764 58219 12767
rect 59357 12767 59415 12773
rect 59357 12764 59369 12767
rect 58207 12736 59369 12764
rect 58207 12733 58219 12736
rect 58161 12727 58219 12733
rect 59357 12733 59369 12736
rect 59403 12733 59415 12767
rect 59357 12727 59415 12733
rect 61654 12724 61660 12776
rect 61712 12764 61718 12776
rect 62117 12767 62175 12773
rect 62117 12764 62129 12767
rect 61712 12736 62129 12764
rect 61712 12724 61718 12736
rect 62117 12733 62129 12736
rect 62163 12733 62175 12767
rect 62117 12727 62175 12733
rect 67082 12724 67088 12776
rect 67140 12764 67146 12776
rect 68278 12764 68284 12776
rect 67140 12736 68284 12764
rect 67140 12724 67146 12736
rect 68278 12724 68284 12736
rect 68336 12724 68342 12776
rect 56410 12656 56416 12708
rect 56468 12696 56474 12708
rect 56468 12668 57376 12696
rect 56468 12656 56474 12668
rect 57348 12637 57376 12668
rect 57698 12656 57704 12708
rect 57756 12696 57762 12708
rect 57756 12668 58388 12696
rect 57756 12656 57762 12668
rect 56152 12600 56364 12628
rect 57333 12631 57391 12637
rect 52227 12597 52239 12600
rect 52181 12591 52239 12597
rect 57333 12597 57345 12631
rect 57379 12628 57391 12631
rect 58250 12628 58256 12640
rect 57379 12600 58256 12628
rect 57379 12597 57391 12600
rect 57333 12591 57391 12597
rect 58250 12588 58256 12600
rect 58308 12588 58314 12640
rect 58360 12628 58388 12668
rect 58434 12656 58440 12708
rect 58492 12696 58498 12708
rect 59078 12696 59084 12708
rect 58492 12668 59084 12696
rect 58492 12656 58498 12668
rect 59078 12656 59084 12668
rect 59136 12656 59142 12708
rect 60458 12656 60464 12708
rect 60516 12696 60522 12708
rect 65705 12699 65763 12705
rect 60516 12668 62804 12696
rect 60516 12656 60522 12668
rect 60642 12628 60648 12640
rect 58360 12600 60648 12628
rect 60642 12588 60648 12600
rect 60700 12588 60706 12640
rect 61010 12588 61016 12640
rect 61068 12628 61074 12640
rect 61930 12628 61936 12640
rect 61068 12600 61936 12628
rect 61068 12588 61074 12600
rect 61930 12588 61936 12600
rect 61988 12628 61994 12640
rect 62206 12628 62212 12640
rect 61988 12600 62212 12628
rect 61988 12588 61994 12600
rect 62206 12588 62212 12600
rect 62264 12588 62270 12640
rect 62776 12628 62804 12668
rect 65705 12665 65717 12699
rect 65751 12696 65763 12699
rect 68370 12696 68376 12708
rect 65751 12668 68376 12696
rect 65751 12665 65763 12668
rect 65705 12659 65763 12665
rect 68370 12656 68376 12668
rect 68428 12656 68434 12708
rect 68646 12696 68652 12708
rect 68559 12668 68652 12696
rect 68646 12656 68652 12668
rect 68704 12656 68710 12708
rect 68756 12696 68784 12804
rect 68830 12792 68836 12844
rect 68888 12832 68894 12844
rect 69753 12835 69811 12841
rect 69753 12832 69765 12835
rect 68888 12804 69765 12832
rect 68888 12792 68894 12804
rect 69753 12801 69765 12804
rect 69799 12801 69811 12835
rect 70366 12832 70394 12872
rect 70762 12860 70768 12872
rect 70820 12860 70826 12912
rect 72050 12900 72056 12912
rect 71990 12872 72056 12900
rect 72050 12860 72056 12872
rect 72108 12860 72114 12912
rect 72418 12860 72424 12912
rect 72476 12900 72482 12912
rect 72476 12872 75684 12900
rect 72476 12860 72482 12872
rect 70486 12832 70492 12844
rect 70366 12804 70492 12832
rect 69753 12795 69811 12801
rect 70486 12792 70492 12804
rect 70544 12792 70550 12844
rect 73522 12792 73528 12844
rect 73580 12832 73586 12844
rect 73617 12835 73675 12841
rect 73617 12832 73629 12835
rect 73580 12804 73629 12832
rect 73580 12792 73586 12804
rect 73617 12801 73629 12804
rect 73663 12801 73675 12835
rect 73617 12795 73675 12801
rect 75181 12835 75239 12841
rect 75181 12801 75193 12835
rect 75227 12832 75239 12835
rect 75270 12832 75276 12844
rect 75227 12804 75276 12832
rect 75227 12801 75239 12804
rect 75181 12795 75239 12801
rect 75270 12792 75276 12804
rect 75328 12792 75334 12844
rect 75656 12841 75684 12872
rect 75730 12860 75736 12912
rect 75788 12900 75794 12912
rect 75788 12872 75833 12900
rect 75788 12860 75794 12872
rect 76760 12841 76788 12940
rect 76926 12928 76932 12940
rect 76984 12928 76990 12980
rect 77018 12928 77024 12980
rect 77076 12968 77082 12980
rect 77076 12940 79824 12968
rect 77076 12928 77082 12940
rect 77202 12860 77208 12912
rect 77260 12900 77266 12912
rect 77757 12903 77815 12909
rect 77757 12900 77769 12903
rect 77260 12872 77769 12900
rect 77260 12860 77266 12872
rect 77757 12869 77769 12872
rect 77803 12869 77815 12903
rect 77757 12863 77815 12869
rect 79502 12860 79508 12912
rect 79560 12860 79566 12912
rect 79796 12900 79824 12940
rect 79870 12928 79876 12980
rect 79928 12968 79934 12980
rect 79928 12940 83136 12968
rect 79928 12928 79934 12940
rect 83108 12900 83136 12940
rect 83182 12928 83188 12980
rect 83240 12968 83246 12980
rect 83921 12971 83979 12977
rect 83921 12968 83933 12971
rect 83240 12940 83933 12968
rect 83240 12928 83246 12940
rect 83921 12937 83933 12940
rect 83967 12937 83979 12971
rect 83921 12931 83979 12937
rect 84562 12928 84568 12980
rect 84620 12968 84626 12980
rect 84657 12971 84715 12977
rect 84657 12968 84669 12971
rect 84620 12940 84669 12968
rect 84620 12928 84626 12940
rect 84657 12937 84669 12940
rect 84703 12937 84715 12971
rect 87782 12968 87788 12980
rect 87743 12940 87788 12968
rect 84657 12931 84715 12937
rect 87782 12928 87788 12940
rect 87840 12928 87846 12980
rect 93302 12968 93308 12980
rect 93263 12940 93308 12968
rect 93302 12928 93308 12940
rect 93360 12928 93366 12980
rect 85022 12900 85028 12912
rect 79796 12872 83044 12900
rect 83108 12872 85028 12900
rect 75641 12835 75699 12841
rect 75641 12801 75653 12835
rect 75687 12801 75699 12835
rect 75641 12795 75699 12801
rect 76745 12835 76803 12841
rect 76745 12801 76757 12835
rect 76791 12801 76803 12835
rect 76745 12795 76803 12801
rect 77110 12792 77116 12844
rect 77168 12832 77174 12844
rect 77481 12835 77539 12841
rect 77481 12832 77493 12835
rect 77168 12804 77493 12832
rect 77168 12792 77174 12804
rect 77481 12801 77493 12804
rect 77527 12832 77539 12835
rect 78674 12832 78680 12844
rect 77527 12804 78680 12832
rect 77527 12801 77539 12804
rect 77481 12795 77539 12801
rect 78674 12792 78680 12804
rect 78732 12792 78738 12844
rect 80514 12792 80520 12844
rect 80572 12832 80578 12844
rect 81897 12835 81955 12841
rect 81897 12832 81909 12835
rect 80572 12804 81909 12832
rect 80572 12792 80578 12804
rect 81897 12801 81909 12804
rect 81943 12801 81955 12835
rect 82262 12832 82268 12844
rect 82223 12804 82268 12832
rect 81897 12795 81955 12801
rect 82262 12792 82268 12804
rect 82320 12792 82326 12844
rect 83016 12832 83044 12872
rect 85022 12860 85028 12872
rect 85080 12860 85086 12912
rect 85500 12872 87736 12900
rect 84102 12832 84108 12844
rect 83016 12804 83964 12832
rect 84063 12804 84108 12832
rect 69290 12764 69296 12776
rect 69203 12736 69296 12764
rect 69290 12724 69296 12736
rect 69348 12764 69354 12776
rect 71958 12764 71964 12776
rect 69348 12736 71964 12764
rect 69348 12724 69354 12736
rect 71958 12724 71964 12736
rect 72016 12724 72022 12776
rect 72510 12764 72516 12776
rect 72471 12736 72516 12764
rect 72510 12724 72516 12736
rect 72568 12724 72574 12776
rect 78214 12724 78220 12776
rect 78272 12764 78278 12776
rect 80149 12767 80207 12773
rect 80149 12764 80161 12767
rect 78272 12736 80161 12764
rect 78272 12724 78278 12736
rect 80149 12733 80161 12736
rect 80195 12733 80207 12767
rect 80149 12727 80207 12733
rect 80425 12767 80483 12773
rect 80425 12733 80437 12767
rect 80471 12733 80483 12767
rect 80425 12727 80483 12733
rect 73890 12696 73896 12708
rect 68756 12668 70256 12696
rect 68664 12628 68692 12656
rect 62776 12600 68692 12628
rect 69937 12631 69995 12637
rect 69937 12597 69949 12631
rect 69983 12628 69995 12631
rect 70118 12628 70124 12640
rect 69983 12600 70124 12628
rect 69983 12597 69995 12600
rect 69937 12591 69995 12597
rect 70118 12588 70124 12600
rect 70176 12588 70182 12640
rect 70228 12628 70256 12668
rect 72712 12668 73896 12696
rect 70946 12628 70952 12640
rect 70228 12600 70952 12628
rect 70946 12588 70952 12600
rect 71004 12588 71010 12640
rect 71222 12588 71228 12640
rect 71280 12628 71286 12640
rect 72712 12628 72740 12668
rect 73890 12656 73896 12668
rect 73948 12656 73954 12708
rect 75822 12656 75828 12708
rect 75880 12696 75886 12708
rect 80440 12696 80468 12727
rect 83826 12696 83832 12708
rect 75880 12668 78812 12696
rect 80440 12668 83832 12696
rect 75880 12656 75886 12668
rect 71280 12600 72740 12628
rect 71280 12588 71286 12600
rect 73522 12588 73528 12640
rect 73580 12628 73586 12640
rect 73709 12631 73767 12637
rect 73709 12628 73721 12631
rect 73580 12600 73721 12628
rect 73580 12588 73586 12600
rect 73709 12597 73721 12600
rect 73755 12597 73767 12631
rect 73709 12591 73767 12597
rect 73982 12588 73988 12640
rect 74040 12628 74046 12640
rect 74261 12631 74319 12637
rect 74261 12628 74273 12631
rect 74040 12600 74273 12628
rect 74040 12588 74046 12600
rect 74261 12597 74273 12600
rect 74307 12597 74319 12631
rect 74994 12628 75000 12640
rect 74955 12600 75000 12628
rect 74261 12591 74319 12597
rect 74994 12588 75000 12600
rect 75052 12588 75058 12640
rect 75178 12588 75184 12640
rect 75236 12628 75242 12640
rect 78306 12628 78312 12640
rect 75236 12600 78312 12628
rect 75236 12588 75242 12600
rect 78306 12588 78312 12600
rect 78364 12588 78370 12640
rect 78582 12588 78588 12640
rect 78640 12628 78646 12640
rect 78677 12631 78735 12637
rect 78677 12628 78689 12631
rect 78640 12600 78689 12628
rect 78640 12588 78646 12600
rect 78677 12597 78689 12600
rect 78723 12597 78735 12631
rect 78784 12628 78812 12668
rect 83826 12656 83832 12668
rect 83884 12656 83890 12708
rect 83936 12696 83964 12804
rect 84102 12792 84108 12804
rect 84160 12792 84166 12844
rect 84749 12835 84807 12841
rect 84749 12801 84761 12835
rect 84795 12801 84807 12835
rect 84749 12795 84807 12801
rect 84470 12696 84476 12708
rect 83936 12668 84476 12696
rect 84470 12656 84476 12668
rect 84528 12656 84534 12708
rect 84764 12696 84792 12795
rect 85206 12792 85212 12844
rect 85264 12832 85270 12844
rect 85500 12841 85528 12872
rect 85485 12835 85543 12841
rect 85485 12832 85497 12835
rect 85264 12804 85497 12832
rect 85264 12792 85270 12804
rect 85485 12801 85497 12804
rect 85531 12801 85543 12835
rect 86218 12832 86224 12844
rect 86179 12804 86224 12832
rect 85485 12795 85543 12801
rect 86218 12792 86224 12804
rect 86276 12792 86282 12844
rect 86862 12832 86868 12844
rect 86823 12804 86868 12832
rect 86862 12792 86868 12804
rect 86920 12792 86926 12844
rect 87708 12841 87736 12872
rect 89346 12860 89352 12912
rect 89404 12900 89410 12912
rect 89404 12872 91140 12900
rect 89404 12860 89410 12872
rect 87693 12835 87751 12841
rect 87693 12801 87705 12835
rect 87739 12832 87751 12835
rect 87782 12832 87788 12844
rect 87739 12804 87788 12832
rect 87739 12801 87751 12804
rect 87693 12795 87751 12801
rect 87782 12792 87788 12804
rect 87840 12792 87846 12844
rect 89438 12832 89444 12844
rect 89399 12804 89444 12832
rect 89438 12792 89444 12804
rect 89496 12792 89502 12844
rect 89530 12792 89536 12844
rect 89588 12832 89594 12844
rect 89588 12804 89633 12832
rect 89588 12792 89594 12804
rect 90542 12792 90548 12844
rect 90600 12832 90606 12844
rect 91112 12841 91140 12872
rect 92474 12860 92480 12912
rect 92532 12900 92538 12912
rect 94225 12903 94283 12909
rect 94225 12900 94237 12903
rect 92532 12872 94237 12900
rect 92532 12860 92538 12872
rect 90729 12835 90787 12841
rect 90729 12832 90741 12835
rect 90600 12804 90741 12832
rect 90600 12792 90606 12804
rect 90729 12801 90741 12804
rect 90775 12801 90787 12835
rect 90729 12795 90787 12801
rect 91097 12835 91155 12841
rect 91097 12801 91109 12835
rect 91143 12801 91155 12835
rect 92566 12832 92572 12844
rect 92527 12804 92572 12832
rect 91097 12795 91155 12801
rect 92566 12792 92572 12804
rect 92624 12792 92630 12844
rect 92768 12841 92796 12872
rect 94225 12869 94237 12872
rect 94271 12869 94283 12903
rect 94225 12863 94283 12869
rect 92753 12835 92811 12841
rect 92753 12801 92765 12835
rect 92799 12801 92811 12835
rect 92753 12795 92811 12801
rect 93213 12835 93271 12841
rect 93213 12801 93225 12835
rect 93259 12801 93271 12835
rect 93213 12795 93271 12801
rect 86770 12764 86776 12776
rect 86731 12736 86776 12764
rect 86770 12724 86776 12736
rect 86828 12724 86834 12776
rect 88337 12767 88395 12773
rect 88337 12764 88349 12767
rect 87156 12736 88349 12764
rect 87156 12696 87184 12736
rect 88337 12733 88349 12736
rect 88383 12764 88395 12767
rect 89070 12764 89076 12776
rect 88383 12736 89076 12764
rect 88383 12733 88395 12736
rect 88337 12727 88395 12733
rect 89070 12724 89076 12736
rect 89128 12724 89134 12776
rect 92106 12724 92112 12776
rect 92164 12764 92170 12776
rect 93228 12764 93256 12795
rect 93302 12792 93308 12844
rect 93360 12832 93366 12844
rect 94133 12835 94191 12841
rect 94133 12832 94145 12835
rect 93360 12804 94145 12832
rect 93360 12792 93366 12804
rect 94133 12801 94145 12804
rect 94179 12801 94191 12835
rect 94133 12795 94191 12801
rect 92164 12736 93256 12764
rect 92164 12724 92170 12736
rect 84764 12668 87184 12696
rect 87233 12699 87291 12705
rect 87233 12665 87245 12699
rect 87279 12696 87291 12699
rect 89622 12696 89628 12708
rect 87279 12668 89628 12696
rect 87279 12665 87291 12668
rect 87233 12659 87291 12665
rect 89622 12656 89628 12668
rect 89680 12656 89686 12708
rect 80146 12628 80152 12640
rect 78784 12600 80152 12628
rect 78677 12591 78735 12597
rect 80146 12588 80152 12600
rect 80204 12588 80210 12640
rect 81526 12628 81532 12640
rect 81487 12600 81532 12628
rect 81526 12588 81532 12600
rect 81584 12588 81590 12640
rect 85114 12588 85120 12640
rect 85172 12628 85178 12640
rect 85393 12631 85451 12637
rect 85393 12628 85405 12631
rect 85172 12600 85405 12628
rect 85172 12588 85178 12600
rect 85393 12597 85405 12600
rect 85439 12597 85451 12631
rect 85393 12591 85451 12597
rect 85574 12588 85580 12640
rect 85632 12628 85638 12640
rect 86129 12631 86187 12637
rect 86129 12628 86141 12631
rect 85632 12600 86141 12628
rect 85632 12588 85638 12600
rect 86129 12597 86141 12600
rect 86175 12597 86187 12631
rect 90174 12628 90180 12640
rect 90135 12600 90180 12628
rect 86129 12591 86187 12597
rect 90174 12588 90180 12600
rect 90232 12588 90238 12640
rect 92753 12631 92811 12637
rect 92753 12597 92765 12631
rect 92799 12628 92811 12631
rect 92934 12628 92940 12640
rect 92799 12600 92940 12628
rect 92799 12597 92811 12600
rect 92753 12591 92811 12597
rect 92934 12588 92940 12600
rect 92992 12588 92998 12640
rect 1104 12538 94852 12560
rect 1104 12486 12668 12538
rect 12720 12486 12732 12538
rect 12784 12486 12796 12538
rect 12848 12486 12860 12538
rect 12912 12486 12924 12538
rect 12976 12486 36105 12538
rect 36157 12486 36169 12538
rect 36221 12486 36233 12538
rect 36285 12486 36297 12538
rect 36349 12486 36361 12538
rect 36413 12486 59542 12538
rect 59594 12486 59606 12538
rect 59658 12486 59670 12538
rect 59722 12486 59734 12538
rect 59786 12486 59798 12538
rect 59850 12486 82979 12538
rect 83031 12486 83043 12538
rect 83095 12486 83107 12538
rect 83159 12486 83171 12538
rect 83223 12486 83235 12538
rect 83287 12486 94852 12538
rect 1104 12464 94852 12486
rect 4522 12384 4528 12436
rect 4580 12424 4586 12436
rect 4580 12396 13860 12424
rect 4580 12384 4586 12396
rect 13832 12356 13860 12396
rect 13906 12384 13912 12436
rect 13964 12424 13970 12436
rect 15102 12424 15108 12436
rect 13964 12396 15108 12424
rect 13964 12384 13970 12396
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 15746 12384 15752 12436
rect 15804 12424 15810 12436
rect 15804 12396 19564 12424
rect 15804 12384 15810 12396
rect 13832 12328 13952 12356
rect 3329 12291 3387 12297
rect 3329 12257 3341 12291
rect 3375 12288 3387 12291
rect 4062 12288 4068 12300
rect 3375 12260 4068 12288
rect 3375 12257 3387 12260
rect 3329 12251 3387 12257
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 8018 12288 8024 12300
rect 7979 12260 8024 12288
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 13725 12291 13783 12297
rect 13725 12257 13737 12291
rect 13771 12288 13783 12291
rect 13814 12288 13820 12300
rect 13771 12260 13820 12288
rect 13771 12257 13783 12260
rect 13725 12251 13783 12257
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 13924 12288 13952 12328
rect 16114 12316 16120 12368
rect 16172 12356 16178 12368
rect 19242 12356 19248 12368
rect 16172 12328 17080 12356
rect 16172 12316 16178 12328
rect 15746 12288 15752 12300
rect 13924 12260 15752 12288
rect 15746 12248 15752 12260
rect 15804 12248 15810 12300
rect 15841 12291 15899 12297
rect 15841 12257 15853 12291
rect 15887 12288 15899 12291
rect 16942 12288 16948 12300
rect 15887 12260 16948 12288
rect 15887 12257 15899 12260
rect 15841 12251 15899 12257
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 17052 12288 17080 12328
rect 18432 12328 19248 12356
rect 18432 12288 18460 12328
rect 19242 12316 19248 12328
rect 19300 12316 19306 12368
rect 17052 12260 18460 12288
rect 18509 12291 18567 12297
rect 18509 12257 18521 12291
rect 18555 12288 18567 12291
rect 18598 12288 18604 12300
rect 18555 12260 18604 12288
rect 18555 12257 18567 12260
rect 18509 12251 18567 12257
rect 18598 12248 18604 12260
rect 18656 12248 18662 12300
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 19429 12291 19487 12297
rect 19429 12288 19441 12291
rect 19392 12260 19441 12288
rect 19392 12248 19398 12260
rect 19429 12257 19441 12260
rect 19475 12257 19487 12291
rect 19536 12288 19564 12396
rect 20438 12384 20444 12436
rect 20496 12424 20502 12436
rect 21177 12427 21235 12433
rect 21177 12424 21189 12427
rect 20496 12396 21189 12424
rect 20496 12384 20502 12396
rect 21177 12393 21189 12396
rect 21223 12393 21235 12427
rect 21177 12387 21235 12393
rect 21821 12427 21879 12433
rect 21821 12393 21833 12427
rect 21867 12424 21879 12427
rect 22094 12424 22100 12436
rect 21867 12396 22100 12424
rect 21867 12393 21879 12396
rect 21821 12387 21879 12393
rect 22094 12384 22100 12396
rect 22152 12384 22158 12436
rect 22186 12384 22192 12436
rect 22244 12424 22250 12436
rect 22738 12424 22744 12436
rect 22244 12396 22744 12424
rect 22244 12384 22250 12396
rect 22738 12384 22744 12396
rect 22796 12384 22802 12436
rect 24857 12427 24915 12433
rect 24857 12393 24869 12427
rect 24903 12424 24915 12427
rect 26418 12424 26424 12436
rect 24903 12396 26424 12424
rect 24903 12393 24915 12396
rect 24857 12387 24915 12393
rect 26418 12384 26424 12396
rect 26476 12424 26482 12436
rect 29914 12424 29920 12436
rect 26476 12396 27384 12424
rect 29875 12396 29920 12424
rect 26476 12384 26482 12396
rect 24026 12356 24032 12368
rect 23987 12328 24032 12356
rect 24026 12316 24032 12328
rect 24084 12316 24090 12368
rect 26234 12316 26240 12368
rect 26292 12356 26298 12368
rect 27154 12356 27160 12368
rect 26292 12328 27160 12356
rect 26292 12316 26298 12328
rect 27154 12316 27160 12328
rect 27212 12316 27218 12368
rect 19705 12291 19763 12297
rect 19705 12288 19717 12291
rect 19536 12260 19717 12288
rect 19429 12251 19487 12257
rect 19705 12257 19717 12260
rect 19751 12257 19763 12291
rect 22278 12288 22284 12300
rect 22239 12260 22284 12288
rect 19705 12251 19763 12257
rect 22278 12248 22284 12260
rect 22336 12248 22342 12300
rect 22557 12291 22615 12297
rect 22557 12257 22569 12291
rect 22603 12288 22615 12291
rect 26329 12291 26387 12297
rect 22603 12260 26188 12288
rect 22603 12257 22615 12260
rect 22557 12251 22615 12257
rect 2958 12180 2964 12232
rect 3016 12220 3022 12232
rect 3237 12223 3295 12229
rect 3237 12220 3249 12223
rect 3016 12192 3249 12220
rect 3016 12180 3022 12192
rect 3237 12189 3249 12192
rect 3283 12220 3295 12223
rect 5077 12223 5135 12229
rect 5077 12220 5089 12223
rect 3283 12192 5089 12220
rect 3283 12189 3295 12192
rect 3237 12183 3295 12189
rect 5077 12189 5089 12192
rect 5123 12220 5135 12223
rect 5166 12220 5172 12232
rect 5123 12192 5172 12220
rect 5123 12189 5135 12192
rect 5077 12183 5135 12189
rect 5166 12180 5172 12192
rect 5224 12180 5230 12232
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12220 8539 12223
rect 9674 12220 9680 12232
rect 8527 12192 9680 12220
rect 8527 12189 8539 12192
rect 8481 12183 8539 12189
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 16114 12180 16120 12232
rect 16172 12220 16178 12232
rect 21634 12220 21640 12232
rect 16172 12192 16217 12220
rect 21595 12192 21640 12220
rect 16172 12180 16178 12192
rect 21634 12180 21640 12192
rect 21692 12180 21698 12232
rect 4341 12155 4399 12161
rect 4341 12121 4353 12155
rect 4387 12152 4399 12155
rect 4522 12152 4528 12164
rect 4387 12124 4528 12152
rect 4387 12121 4399 12124
rect 4341 12115 4399 12121
rect 4522 12112 4528 12124
rect 4580 12112 4586 12164
rect 5534 12112 5540 12164
rect 5592 12152 5598 12164
rect 6089 12155 6147 12161
rect 6089 12152 6101 12155
rect 5592 12124 6101 12152
rect 5592 12112 5598 12124
rect 6089 12121 6101 12124
rect 6135 12121 6147 12155
rect 6089 12115 6147 12121
rect 12986 12112 12992 12164
rect 13044 12112 13050 12164
rect 13446 12152 13452 12164
rect 13407 12124 13452 12152
rect 13446 12112 13452 12124
rect 13504 12112 13510 12164
rect 13998 12112 14004 12164
rect 14056 12152 14062 12164
rect 14056 12124 14674 12152
rect 14056 12112 14062 12124
rect 15562 12112 15568 12164
rect 15620 12152 15626 12164
rect 16850 12152 16856 12164
rect 15620 12124 16856 12152
rect 15620 12112 15626 12124
rect 16850 12112 16856 12124
rect 16908 12152 16914 12164
rect 18230 12152 18236 12164
rect 16908 12124 17066 12152
rect 18191 12124 18236 12152
rect 16908 12112 16914 12124
rect 2869 12087 2927 12093
rect 2869 12053 2881 12087
rect 2915 12084 2927 12087
rect 3050 12084 3056 12096
rect 2915 12056 3056 12084
rect 2915 12053 2927 12056
rect 2869 12047 2927 12053
rect 3050 12044 3056 12056
rect 3108 12044 3114 12096
rect 5994 12084 6000 12096
rect 5955 12056 6000 12084
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6822 12084 6828 12096
rect 6783 12056 6828 12084
rect 6822 12044 6828 12056
rect 6880 12044 6886 12096
rect 7282 12084 7288 12096
rect 7243 12056 7288 12084
rect 7282 12044 7288 12056
rect 7340 12084 7346 12096
rect 7926 12084 7932 12096
rect 7340 12056 7932 12084
rect 7340 12044 7346 12056
rect 7926 12044 7932 12056
rect 7984 12044 7990 12096
rect 11974 12084 11980 12096
rect 11935 12056 11980 12084
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 14366 12084 14372 12096
rect 14327 12056 14372 12084
rect 14366 12044 14372 12056
rect 14424 12044 14430 12096
rect 15470 12044 15476 12096
rect 15528 12084 15534 12096
rect 16761 12087 16819 12093
rect 16761 12084 16773 12087
rect 15528 12056 16773 12084
rect 15528 12044 15534 12056
rect 16761 12053 16773 12056
rect 16807 12053 16819 12087
rect 16960 12084 16988 12124
rect 18230 12112 18236 12124
rect 18288 12112 18294 12164
rect 26160 12152 26188 12260
rect 26329 12257 26341 12291
rect 26375 12288 26387 12291
rect 27356 12288 27384 12396
rect 29914 12384 29920 12396
rect 29972 12384 29978 12436
rect 30742 12384 30748 12436
rect 30800 12424 30806 12436
rect 30837 12427 30895 12433
rect 30837 12424 30849 12427
rect 30800 12396 30849 12424
rect 30800 12384 30806 12396
rect 30837 12393 30849 12396
rect 30883 12393 30895 12427
rect 34974 12424 34980 12436
rect 34935 12396 34980 12424
rect 30837 12387 30895 12393
rect 34974 12384 34980 12396
rect 35032 12384 35038 12436
rect 36446 12384 36452 12436
rect 36504 12424 36510 12436
rect 37737 12427 37795 12433
rect 37737 12424 37749 12427
rect 36504 12396 37749 12424
rect 36504 12384 36510 12396
rect 37737 12393 37749 12396
rect 37783 12393 37795 12427
rect 37737 12387 37795 12393
rect 37826 12384 37832 12436
rect 37884 12424 37890 12436
rect 40313 12427 40371 12433
rect 37884 12396 39436 12424
rect 37884 12384 37890 12396
rect 29181 12359 29239 12365
rect 29181 12325 29193 12359
rect 29227 12356 29239 12359
rect 30650 12356 30656 12368
rect 29227 12328 30656 12356
rect 29227 12325 29239 12328
rect 29181 12319 29239 12325
rect 30650 12316 30656 12328
rect 30708 12316 30714 12368
rect 31036 12328 31340 12356
rect 28169 12291 28227 12297
rect 28169 12288 28181 12291
rect 26375 12260 27016 12288
rect 27356 12260 28181 12288
rect 26375 12257 26387 12260
rect 26329 12251 26387 12257
rect 26237 12223 26295 12229
rect 26237 12189 26249 12223
rect 26283 12220 26295 12223
rect 26418 12220 26424 12232
rect 26283 12192 26424 12220
rect 26283 12189 26295 12192
rect 26237 12183 26295 12189
rect 26418 12180 26424 12192
rect 26476 12180 26482 12232
rect 26878 12152 26884 12164
rect 19306 12124 20194 12152
rect 22756 12124 23046 12152
rect 26160 12124 26884 12152
rect 18414 12084 18420 12096
rect 16960 12056 18420 12084
rect 16761 12047 16819 12053
rect 18414 12044 18420 12056
rect 18472 12084 18478 12096
rect 19306 12084 19334 12124
rect 18472 12056 19334 12084
rect 20088 12084 20116 12124
rect 22756 12096 22784 12124
rect 26878 12112 26884 12124
rect 26936 12112 26942 12164
rect 22738 12084 22744 12096
rect 20088 12056 22744 12084
rect 18472 12044 18478 12056
rect 22738 12044 22744 12056
rect 22796 12084 22802 12096
rect 23198 12084 23204 12096
rect 22796 12056 23204 12084
rect 22796 12044 22802 12056
rect 23198 12044 23204 12056
rect 23256 12044 23262 12096
rect 25406 12084 25412 12096
rect 25367 12056 25412 12084
rect 25406 12044 25412 12056
rect 25464 12044 25470 12096
rect 25866 12084 25872 12096
rect 25827 12056 25872 12084
rect 25866 12044 25872 12056
rect 25924 12044 25930 12096
rect 26988 12084 27016 12260
rect 28169 12257 28181 12260
rect 28215 12257 28227 12291
rect 30282 12288 30288 12300
rect 30195 12260 30288 12288
rect 28169 12251 28227 12257
rect 27062 12180 27068 12232
rect 27120 12220 27126 12232
rect 27120 12192 27165 12220
rect 27120 12180 27126 12192
rect 27246 12180 27252 12232
rect 27304 12220 27310 12232
rect 27985 12223 28043 12229
rect 27985 12220 27997 12223
rect 27304 12192 27997 12220
rect 27304 12180 27310 12192
rect 27985 12189 27997 12192
rect 28031 12189 28043 12223
rect 28184 12220 28212 12251
rect 30282 12248 30288 12260
rect 30340 12288 30346 12300
rect 31036 12288 31064 12328
rect 30340 12260 31064 12288
rect 30340 12248 30346 12260
rect 31110 12248 31116 12300
rect 31168 12288 31174 12300
rect 31312 12288 31340 12328
rect 31386 12316 31392 12368
rect 31444 12356 31450 12368
rect 33413 12359 33471 12365
rect 33413 12356 33425 12359
rect 31444 12328 33425 12356
rect 31444 12316 31450 12328
rect 33413 12325 33425 12328
rect 33459 12325 33471 12359
rect 39408 12356 39436 12396
rect 40313 12393 40325 12427
rect 40359 12424 40371 12427
rect 40494 12424 40500 12436
rect 40359 12396 40500 12424
rect 40359 12393 40371 12396
rect 40313 12387 40371 12393
rect 40494 12384 40500 12396
rect 40552 12384 40558 12436
rect 42610 12424 42616 12436
rect 40604 12396 42616 12424
rect 40604 12356 40632 12396
rect 42610 12384 42616 12396
rect 42668 12384 42674 12436
rect 42705 12427 42763 12433
rect 42705 12393 42717 12427
rect 42751 12424 42763 12427
rect 43438 12424 43444 12436
rect 42751 12396 43444 12424
rect 42751 12393 42763 12396
rect 42705 12387 42763 12393
rect 43438 12384 43444 12396
rect 43496 12384 43502 12436
rect 47578 12424 47584 12436
rect 45480 12396 47584 12424
rect 45278 12356 45284 12368
rect 33413 12319 33471 12325
rect 33704 12328 34008 12356
rect 39408 12328 40632 12356
rect 41984 12328 45284 12356
rect 31168 12260 31213 12288
rect 31312 12260 32260 12288
rect 31168 12248 31174 12260
rect 32232 12232 32260 12260
rect 32398 12248 32404 12300
rect 32456 12288 32462 12300
rect 33704 12297 33732 12328
rect 33689 12291 33747 12297
rect 33689 12288 33701 12291
rect 32456 12260 33701 12288
rect 32456 12248 32462 12260
rect 33689 12257 33701 12260
rect 33735 12257 33747 12291
rect 33689 12251 33747 12257
rect 28350 12220 28356 12232
rect 28184 12192 28356 12220
rect 27985 12183 28043 12189
rect 28350 12180 28356 12192
rect 28408 12220 28414 12232
rect 30190 12220 30196 12232
rect 28408 12192 30196 12220
rect 28408 12180 28414 12192
rect 30190 12180 30196 12192
rect 30248 12180 30254 12232
rect 31205 12223 31263 12229
rect 31205 12189 31217 12223
rect 31251 12220 31263 12223
rect 31294 12220 31300 12232
rect 31251 12192 31300 12220
rect 31251 12189 31263 12192
rect 31205 12183 31263 12189
rect 31294 12180 31300 12192
rect 31352 12180 31358 12232
rect 31754 12180 31760 12232
rect 31812 12220 31818 12232
rect 31941 12223 31999 12229
rect 31941 12220 31953 12223
rect 31812 12192 31953 12220
rect 31812 12180 31818 12192
rect 31941 12189 31953 12192
rect 31987 12189 31999 12223
rect 32122 12220 32128 12232
rect 32083 12192 32128 12220
rect 31941 12183 31999 12189
rect 32122 12180 32128 12192
rect 32180 12180 32186 12232
rect 32214 12180 32220 12232
rect 32272 12220 32278 12232
rect 33778 12220 33784 12232
rect 32272 12192 33784 12220
rect 32272 12180 32278 12192
rect 33778 12180 33784 12192
rect 33836 12180 33842 12232
rect 27154 12112 27160 12164
rect 27212 12152 27218 12164
rect 27341 12155 27399 12161
rect 27341 12152 27353 12155
rect 27212 12124 27353 12152
rect 27212 12112 27218 12124
rect 27341 12121 27353 12124
rect 27387 12121 27399 12155
rect 32398 12152 32404 12164
rect 27341 12115 27399 12121
rect 27448 12124 32404 12152
rect 27448 12084 27476 12124
rect 32398 12112 32404 12124
rect 32456 12112 32462 12164
rect 33042 12152 33048 12164
rect 32508 12124 33048 12152
rect 26988 12056 27476 12084
rect 27890 12044 27896 12096
rect 27948 12084 27954 12096
rect 32508 12084 32536 12124
rect 33042 12112 33048 12124
rect 33100 12112 33106 12164
rect 33980 12152 34008 12328
rect 36630 12288 36636 12300
rect 35820 12260 36636 12288
rect 34238 12180 34244 12232
rect 34296 12220 34302 12232
rect 35069 12223 35127 12229
rect 35069 12220 35081 12223
rect 34296 12192 35081 12220
rect 34296 12180 34302 12192
rect 35069 12189 35081 12192
rect 35115 12220 35127 12223
rect 35820 12220 35848 12260
rect 36630 12248 36636 12260
rect 36688 12248 36694 12300
rect 36998 12288 37004 12300
rect 36959 12260 37004 12288
rect 36998 12248 37004 12260
rect 37056 12248 37062 12300
rect 39206 12288 39212 12300
rect 39167 12260 39212 12288
rect 39206 12248 39212 12260
rect 39264 12248 39270 12300
rect 39482 12288 39488 12300
rect 39395 12260 39488 12288
rect 39482 12248 39488 12260
rect 39540 12288 39546 12300
rect 41984 12288 42012 12328
rect 45278 12316 45284 12328
rect 45336 12316 45342 12368
rect 39540 12260 42012 12288
rect 42061 12291 42119 12297
rect 39540 12248 39546 12260
rect 42061 12257 42073 12291
rect 42107 12288 42119 12291
rect 42702 12288 42708 12300
rect 42107 12260 42708 12288
rect 42107 12257 42119 12260
rect 42061 12251 42119 12257
rect 42702 12248 42708 12260
rect 42760 12248 42766 12300
rect 45480 12288 45508 12396
rect 47578 12384 47584 12396
rect 47636 12384 47642 12436
rect 49602 12424 49608 12436
rect 49563 12396 49608 12424
rect 49602 12384 49608 12396
rect 49660 12384 49666 12436
rect 49694 12384 49700 12436
rect 49752 12424 49758 12436
rect 53377 12427 53435 12433
rect 53377 12424 53389 12427
rect 49752 12396 53389 12424
rect 49752 12384 49758 12396
rect 53377 12393 53389 12396
rect 53423 12393 53435 12427
rect 59354 12424 59360 12436
rect 53377 12387 53435 12393
rect 56520 12396 58756 12424
rect 59315 12396 59360 12424
rect 45554 12316 45560 12368
rect 45612 12356 45618 12368
rect 51534 12356 51540 12368
rect 45612 12328 46520 12356
rect 45612 12316 45618 12328
rect 43640 12260 45508 12288
rect 46201 12291 46259 12297
rect 35115 12192 35848 12220
rect 35115 12189 35127 12192
rect 35069 12183 35127 12189
rect 37274 12180 37280 12232
rect 37332 12220 37338 12232
rect 42518 12220 42524 12232
rect 37332 12192 37377 12220
rect 42479 12192 42524 12220
rect 37332 12180 37338 12192
rect 42518 12180 42524 12192
rect 42576 12180 42582 12232
rect 42610 12180 42616 12232
rect 42668 12220 42674 12232
rect 43640 12220 43668 12260
rect 46201 12257 46213 12291
rect 46247 12288 46259 12291
rect 46290 12288 46296 12300
rect 46247 12260 46296 12288
rect 46247 12257 46259 12260
rect 46201 12251 46259 12257
rect 46290 12248 46296 12260
rect 46348 12248 46354 12300
rect 46492 12297 46520 12328
rect 49436 12328 51540 12356
rect 46477 12291 46535 12297
rect 46477 12257 46489 12291
rect 46523 12257 46535 12291
rect 46477 12251 46535 12257
rect 46750 12248 46756 12300
rect 46808 12288 46814 12300
rect 48130 12288 48136 12300
rect 46808 12260 48136 12288
rect 46808 12248 46814 12260
rect 48130 12248 48136 12260
rect 48188 12248 48194 12300
rect 43806 12220 43812 12232
rect 42668 12192 43668 12220
rect 43767 12192 43812 12220
rect 42668 12180 42674 12192
rect 43806 12180 43812 12192
rect 43864 12180 43870 12232
rect 43990 12220 43996 12232
rect 43951 12192 43996 12220
rect 43990 12180 43996 12192
rect 44048 12180 44054 12232
rect 45365 12223 45423 12229
rect 45365 12220 45377 12223
rect 45296 12192 45377 12220
rect 33980 12124 35664 12152
rect 27948 12056 32536 12084
rect 27948 12044 27954 12056
rect 32858 12044 32864 12096
rect 32916 12084 32922 12096
rect 32953 12087 33011 12093
rect 32953 12084 32965 12087
rect 32916 12056 32965 12084
rect 32916 12044 32922 12056
rect 32953 12053 32965 12056
rect 32999 12053 33011 12087
rect 32953 12047 33011 12053
rect 34974 12044 34980 12096
rect 35032 12084 35038 12096
rect 35434 12084 35440 12096
rect 35032 12056 35440 12084
rect 35032 12044 35038 12056
rect 35434 12044 35440 12056
rect 35492 12084 35498 12096
rect 35529 12087 35587 12093
rect 35529 12084 35541 12087
rect 35492 12056 35541 12084
rect 35492 12044 35498 12056
rect 35529 12053 35541 12056
rect 35575 12053 35587 12087
rect 35636 12084 35664 12124
rect 36538 12112 36544 12164
rect 36596 12112 36602 12164
rect 38194 12112 38200 12164
rect 38252 12112 38258 12164
rect 38930 12112 38936 12164
rect 38988 12152 38994 12164
rect 41782 12152 41788 12164
rect 38988 12124 40618 12152
rect 41743 12124 41788 12152
rect 38988 12112 38994 12124
rect 41782 12112 41788 12124
rect 41840 12112 41846 12164
rect 44542 12152 44548 12164
rect 44503 12124 44548 12152
rect 44542 12112 44548 12124
rect 44600 12112 44606 12164
rect 45296 12152 45324 12192
rect 45365 12189 45377 12192
rect 45411 12189 45423 12223
rect 46014 12220 46020 12232
rect 45975 12192 46020 12220
rect 45365 12183 45423 12189
rect 46014 12180 46020 12192
rect 46072 12180 46078 12232
rect 48498 12220 48504 12232
rect 48459 12192 48504 12220
rect 48498 12180 48504 12192
rect 48556 12180 48562 12232
rect 49436 12229 49464 12328
rect 51534 12316 51540 12328
rect 51592 12316 51598 12368
rect 51718 12316 51724 12368
rect 51776 12356 51782 12368
rect 54665 12359 54723 12365
rect 54665 12356 54677 12359
rect 51776 12328 54677 12356
rect 51776 12316 51782 12328
rect 54665 12325 54677 12328
rect 54711 12356 54723 12359
rect 56134 12356 56140 12368
rect 54711 12328 56140 12356
rect 54711 12325 54723 12328
rect 54665 12319 54723 12325
rect 56134 12316 56140 12328
rect 56192 12316 56198 12368
rect 56410 12316 56416 12368
rect 56468 12316 56474 12368
rect 49712 12260 50752 12288
rect 49421 12223 49479 12229
rect 49421 12189 49433 12223
rect 49467 12189 49479 12223
rect 49421 12183 49479 12189
rect 49510 12180 49516 12232
rect 49568 12220 49574 12232
rect 49568 12192 49661 12220
rect 49568 12180 49574 12192
rect 47118 12152 47124 12164
rect 45296 12124 47124 12152
rect 36722 12084 36728 12096
rect 35636 12056 36728 12084
rect 35529 12047 35587 12053
rect 36722 12044 36728 12056
rect 36780 12044 36786 12096
rect 36998 12044 37004 12096
rect 37056 12084 37062 12096
rect 43714 12084 43720 12096
rect 37056 12056 43720 12084
rect 37056 12044 37062 12056
rect 43714 12044 43720 12056
rect 43772 12084 43778 12096
rect 45296 12084 45324 12124
rect 47118 12112 47124 12124
rect 47176 12112 47182 12164
rect 48774 12152 48780 12164
rect 48735 12124 48780 12152
rect 48774 12112 48780 12124
rect 48832 12112 48838 12164
rect 49234 12112 49240 12164
rect 49292 12152 49298 12164
rect 49528 12152 49556 12180
rect 49292 12124 49556 12152
rect 49292 12112 49298 12124
rect 45462 12084 45468 12096
rect 43772 12056 45324 12084
rect 45423 12056 45468 12084
rect 43772 12044 43778 12056
rect 45462 12044 45468 12056
rect 45520 12044 45526 12096
rect 45646 12044 45652 12096
rect 45704 12084 45710 12096
rect 49712 12084 49740 12260
rect 50338 12180 50344 12232
rect 50396 12220 50402 12232
rect 50617 12223 50675 12229
rect 50617 12220 50629 12223
rect 50396 12192 50629 12220
rect 50396 12180 50402 12192
rect 50617 12189 50629 12192
rect 50663 12189 50675 12223
rect 50724 12220 50752 12260
rect 52178 12248 52184 12300
rect 52236 12288 52242 12300
rect 54021 12291 54079 12297
rect 54021 12288 54033 12291
rect 52236 12260 54033 12288
rect 52236 12248 52242 12260
rect 54021 12257 54033 12260
rect 54067 12288 54079 12291
rect 55950 12288 55956 12300
rect 54067 12260 55956 12288
rect 54067 12257 54079 12260
rect 54021 12251 54079 12257
rect 55950 12248 55956 12260
rect 56008 12248 56014 12300
rect 56428 12288 56456 12316
rect 56520 12297 56548 12396
rect 58066 12356 58072 12368
rect 57164 12328 58072 12356
rect 56060 12260 56456 12288
rect 56505 12291 56563 12297
rect 51169 12223 51227 12229
rect 51169 12220 51181 12223
rect 50724 12192 51181 12220
rect 50617 12183 50675 12189
rect 51169 12189 51181 12192
rect 51215 12220 51227 12223
rect 51258 12220 51264 12232
rect 51215 12192 51264 12220
rect 51215 12189 51227 12192
rect 51169 12183 51227 12189
rect 51258 12180 51264 12192
rect 51316 12180 51322 12232
rect 51626 12180 51632 12232
rect 51684 12220 51690 12232
rect 52822 12220 52828 12232
rect 51684 12192 52828 12220
rect 51684 12180 51690 12192
rect 52822 12180 52828 12192
rect 52880 12180 52886 12232
rect 52914 12180 52920 12232
rect 52972 12220 52978 12232
rect 53282 12220 53288 12232
rect 52972 12192 53288 12220
rect 52972 12180 52978 12192
rect 53282 12180 53288 12192
rect 53340 12220 53346 12232
rect 56060 12220 56088 12260
rect 56505 12257 56517 12291
rect 56551 12257 56563 12291
rect 56505 12251 56563 12257
rect 53340 12192 56088 12220
rect 56413 12223 56471 12229
rect 53340 12180 53346 12192
rect 56413 12189 56425 12223
rect 56459 12220 56471 12223
rect 57054 12220 57060 12232
rect 56459 12192 57060 12220
rect 56459 12189 56471 12192
rect 56413 12183 56471 12189
rect 57054 12180 57060 12192
rect 57112 12180 57118 12232
rect 57164 12229 57192 12328
rect 58066 12316 58072 12328
rect 58124 12316 58130 12368
rect 58728 12288 58756 12396
rect 59354 12384 59360 12396
rect 59412 12384 59418 12436
rect 60826 12384 60832 12436
rect 60884 12424 60890 12436
rect 61565 12427 61623 12433
rect 61565 12424 61577 12427
rect 60884 12396 61577 12424
rect 60884 12384 60890 12396
rect 61565 12393 61577 12396
rect 61611 12393 61623 12427
rect 67082 12424 67088 12436
rect 61565 12387 61623 12393
rect 62684 12396 67088 12424
rect 58805 12359 58863 12365
rect 58805 12325 58817 12359
rect 58851 12356 58863 12359
rect 61746 12356 61752 12368
rect 58851 12328 61752 12356
rect 58851 12325 58863 12328
rect 58805 12319 58863 12325
rect 61746 12316 61752 12328
rect 61804 12316 61810 12368
rect 62574 12356 62580 12368
rect 62040 12328 62580 12356
rect 62040 12288 62068 12328
rect 62574 12316 62580 12328
rect 62632 12316 62638 12368
rect 58728 12260 62068 12288
rect 62114 12248 62120 12300
rect 62172 12288 62178 12300
rect 62684 12297 62712 12396
rect 67082 12384 67088 12396
rect 67140 12384 67146 12436
rect 67634 12384 67640 12436
rect 67692 12424 67698 12436
rect 67692 12396 69244 12424
rect 67692 12384 67698 12396
rect 69216 12368 69244 12396
rect 69934 12384 69940 12436
rect 69992 12424 69998 12436
rect 69992 12396 74948 12424
rect 69992 12384 69998 12396
rect 66533 12359 66591 12365
rect 66533 12356 66545 12359
rect 63972 12328 66545 12356
rect 62669 12291 62727 12297
rect 62669 12288 62681 12291
rect 62172 12260 62681 12288
rect 62172 12248 62178 12260
rect 62669 12257 62681 12260
rect 62715 12257 62727 12291
rect 62669 12251 62727 12257
rect 62945 12291 63003 12297
rect 62945 12257 62957 12291
rect 62991 12288 63003 12291
rect 63972 12288 64000 12328
rect 66533 12325 66545 12328
rect 66579 12325 66591 12359
rect 66533 12319 66591 12325
rect 69198 12316 69204 12368
rect 69256 12356 69262 12368
rect 71222 12356 71228 12368
rect 69256 12328 71228 12356
rect 69256 12316 69262 12328
rect 71222 12316 71228 12328
rect 71280 12316 71286 12368
rect 73356 12328 73660 12356
rect 64690 12288 64696 12300
rect 62991 12260 64000 12288
rect 64064 12260 64696 12288
rect 62991 12257 63003 12260
rect 62945 12251 63003 12257
rect 57149 12223 57207 12229
rect 57149 12189 57161 12223
rect 57195 12189 57207 12223
rect 57149 12183 57207 12189
rect 57333 12223 57391 12229
rect 57333 12189 57345 12223
rect 57379 12220 57391 12223
rect 57698 12220 57704 12232
rect 57379 12192 57704 12220
rect 57379 12189 57391 12192
rect 57333 12183 57391 12189
rect 50154 12112 50160 12164
rect 50212 12152 50218 12164
rect 50890 12152 50896 12164
rect 50212 12124 50896 12152
rect 50212 12112 50218 12124
rect 50890 12112 50896 12124
rect 50948 12112 50954 12164
rect 53745 12155 53803 12161
rect 51460 12124 51566 12152
rect 45704 12056 49740 12084
rect 49789 12087 49847 12093
rect 45704 12044 45710 12056
rect 49789 12053 49801 12087
rect 49835 12084 49847 12087
rect 50062 12084 50068 12096
rect 49835 12056 50068 12084
rect 49835 12053 49847 12056
rect 49789 12047 49847 12053
rect 50062 12044 50068 12056
rect 50120 12044 50126 12096
rect 50338 12044 50344 12096
rect 50396 12084 50402 12096
rect 51460 12084 51488 12124
rect 53745 12121 53757 12155
rect 53791 12152 53803 12155
rect 54202 12152 54208 12164
rect 53791 12124 54208 12152
rect 53791 12121 53803 12124
rect 53745 12115 53803 12121
rect 54202 12112 54208 12124
rect 54260 12112 54266 12164
rect 54294 12112 54300 12164
rect 54352 12152 54358 12164
rect 54352 12124 55720 12152
rect 54352 12112 54358 12124
rect 51994 12084 52000 12096
rect 50396 12056 52000 12084
rect 50396 12044 50402 12056
rect 51994 12044 52000 12056
rect 52052 12044 52058 12096
rect 52362 12044 52368 12096
rect 52420 12084 52426 12096
rect 53837 12087 53895 12093
rect 53837 12084 53849 12087
rect 52420 12056 53849 12084
rect 52420 12044 52426 12056
rect 53837 12053 53849 12056
rect 53883 12084 53895 12087
rect 54478 12084 54484 12096
rect 53883 12056 54484 12084
rect 53883 12053 53895 12056
rect 53837 12047 53895 12053
rect 54478 12044 54484 12056
rect 54536 12044 54542 12096
rect 55214 12044 55220 12096
rect 55272 12084 55278 12096
rect 55585 12087 55643 12093
rect 55585 12084 55597 12087
rect 55272 12056 55597 12084
rect 55272 12044 55278 12056
rect 55585 12053 55597 12056
rect 55631 12053 55643 12087
rect 55692 12084 55720 12124
rect 55766 12112 55772 12164
rect 55824 12152 55830 12164
rect 57164 12152 57192 12183
rect 57698 12180 57704 12192
rect 57756 12180 57762 12232
rect 57793 12223 57851 12229
rect 57793 12189 57805 12223
rect 57839 12189 57851 12223
rect 57793 12183 57851 12189
rect 55824 12124 57192 12152
rect 57241 12155 57299 12161
rect 55824 12112 55830 12124
rect 57241 12121 57253 12155
rect 57287 12152 57299 12155
rect 57514 12152 57520 12164
rect 57287 12124 57520 12152
rect 57287 12121 57299 12124
rect 57241 12115 57299 12121
rect 57514 12112 57520 12124
rect 57572 12152 57578 12164
rect 57808 12152 57836 12183
rect 57974 12180 57980 12232
rect 58032 12220 58038 12232
rect 58032 12192 58077 12220
rect 58032 12180 58038 12192
rect 58342 12180 58348 12232
rect 58400 12220 58406 12232
rect 58710 12220 58716 12232
rect 58400 12192 58716 12220
rect 58400 12180 58406 12192
rect 58710 12180 58716 12192
rect 58768 12180 58774 12232
rect 58894 12220 58900 12232
rect 58855 12192 58900 12220
rect 58894 12180 58900 12192
rect 58952 12180 58958 12232
rect 59998 12180 60004 12232
rect 60056 12220 60062 12232
rect 60642 12220 60648 12232
rect 60056 12192 60648 12220
rect 60056 12180 60062 12192
rect 60642 12180 60648 12192
rect 60700 12180 60706 12232
rect 61654 12180 61660 12232
rect 61712 12220 61718 12232
rect 61712 12192 62068 12220
rect 64064 12206 64092 12260
rect 64690 12248 64696 12260
rect 64748 12248 64754 12300
rect 66226 12260 67312 12288
rect 65978 12220 65984 12232
rect 65939 12192 65984 12220
rect 61712 12180 61718 12192
rect 57572 12124 57836 12152
rect 57885 12155 57943 12161
rect 57572 12112 57578 12124
rect 57885 12121 57897 12155
rect 57931 12152 57943 12155
rect 58526 12152 58532 12164
rect 57931 12124 58532 12152
rect 57931 12121 57943 12124
rect 57885 12115 57943 12121
rect 58526 12112 58532 12124
rect 58584 12152 58590 12164
rect 62040 12161 62068 12192
rect 65978 12180 65984 12192
rect 66036 12220 66042 12232
rect 66226 12220 66254 12260
rect 66622 12220 66628 12232
rect 66036 12192 66254 12220
rect 66583 12192 66628 12220
rect 66036 12180 66042 12192
rect 66622 12180 66628 12192
rect 66680 12180 66686 12232
rect 67284 12229 67312 12260
rect 67542 12248 67548 12300
rect 67600 12288 67606 12300
rect 71038 12288 71044 12300
rect 67600 12260 71044 12288
rect 67600 12248 67606 12260
rect 71038 12248 71044 12260
rect 71096 12248 71102 12300
rect 72234 12248 72240 12300
rect 72292 12288 72298 12300
rect 73356 12288 73384 12328
rect 73522 12288 73528 12300
rect 72292 12260 73384 12288
rect 73483 12260 73528 12288
rect 72292 12248 72298 12260
rect 73522 12248 73528 12260
rect 73580 12248 73586 12300
rect 73632 12288 73660 12328
rect 74810 12288 74816 12300
rect 73632 12260 74816 12288
rect 74810 12248 74816 12260
rect 74868 12248 74874 12300
rect 74920 12288 74948 12396
rect 74994 12384 75000 12436
rect 75052 12424 75058 12436
rect 78582 12424 78588 12436
rect 75052 12396 78588 12424
rect 75052 12384 75058 12396
rect 78582 12384 78588 12396
rect 78640 12384 78646 12436
rect 78674 12384 78680 12436
rect 78732 12424 78738 12436
rect 79962 12424 79968 12436
rect 78732 12396 79968 12424
rect 78732 12384 78738 12396
rect 79962 12384 79968 12396
rect 80020 12384 80026 12436
rect 80238 12424 80244 12436
rect 80151 12396 80244 12424
rect 80238 12384 80244 12396
rect 80296 12424 80302 12436
rect 80790 12424 80796 12436
rect 80296 12396 80796 12424
rect 80296 12384 80302 12396
rect 80790 12384 80796 12396
rect 80848 12384 80854 12436
rect 84102 12424 84108 12436
rect 84015 12396 84108 12424
rect 84102 12384 84108 12396
rect 84160 12424 84166 12436
rect 84160 12396 85988 12424
rect 84160 12384 84166 12396
rect 77938 12356 77944 12368
rect 77404 12328 77944 12356
rect 74920 12260 75040 12288
rect 67269 12223 67327 12229
rect 67269 12189 67281 12223
rect 67315 12189 67327 12223
rect 67269 12183 67327 12189
rect 67361 12223 67419 12229
rect 67361 12189 67373 12223
rect 67407 12220 67419 12223
rect 67913 12223 67971 12229
rect 67913 12220 67925 12223
rect 67407 12192 67925 12220
rect 67407 12189 67419 12192
rect 67361 12183 67419 12189
rect 67913 12189 67925 12192
rect 67959 12189 67971 12223
rect 67913 12183 67971 12189
rect 70397 12223 70455 12229
rect 70397 12189 70409 12223
rect 70443 12220 70455 12223
rect 71498 12220 71504 12232
rect 70443 12192 71504 12220
rect 70443 12189 70455 12192
rect 70397 12183 70455 12189
rect 71498 12180 71504 12192
rect 71556 12180 71562 12232
rect 73065 12223 73123 12229
rect 73065 12189 73077 12223
rect 73111 12189 73123 12223
rect 75012 12220 75040 12260
rect 75362 12248 75368 12300
rect 75420 12288 75426 12300
rect 75549 12291 75607 12297
rect 75549 12288 75561 12291
rect 75420 12260 75561 12288
rect 75420 12248 75426 12260
rect 75549 12257 75561 12260
rect 75595 12257 75607 12291
rect 75549 12251 75607 12257
rect 75638 12248 75644 12300
rect 75696 12288 75702 12300
rect 77110 12288 77116 12300
rect 75696 12260 77116 12288
rect 75696 12248 75702 12260
rect 77110 12248 77116 12260
rect 77168 12248 77174 12300
rect 76285 12223 76343 12229
rect 76285 12220 76297 12223
rect 75012 12192 76297 12220
rect 73065 12183 73123 12189
rect 76285 12189 76297 12192
rect 76331 12189 76343 12223
rect 76285 12183 76343 12189
rect 61841 12155 61899 12161
rect 61841 12152 61853 12155
rect 58584 12124 61853 12152
rect 58584 12112 58590 12124
rect 61841 12121 61853 12124
rect 61887 12121 61899 12155
rect 61841 12115 61899 12121
rect 62025 12155 62083 12161
rect 62025 12121 62037 12155
rect 62071 12121 62083 12155
rect 62025 12115 62083 12121
rect 62117 12155 62175 12161
rect 62117 12121 62129 12155
rect 62163 12121 62175 12155
rect 62117 12115 62175 12121
rect 64693 12155 64751 12161
rect 64693 12121 64705 12155
rect 64739 12152 64751 12155
rect 64739 12124 66208 12152
rect 64739 12121 64751 12124
rect 64693 12115 64751 12121
rect 56594 12084 56600 12096
rect 55692 12056 56600 12084
rect 55585 12047 55643 12053
rect 56594 12044 56600 12056
rect 56652 12044 56658 12096
rect 59446 12044 59452 12096
rect 59504 12084 59510 12096
rect 59909 12087 59967 12093
rect 59909 12084 59921 12087
rect 59504 12056 59921 12084
rect 59504 12044 59510 12056
rect 59909 12053 59921 12056
rect 59955 12084 59967 12087
rect 60642 12084 60648 12096
rect 59955 12056 60648 12084
rect 59955 12053 59967 12056
rect 59909 12047 59967 12053
rect 60642 12044 60648 12056
rect 60700 12044 60706 12096
rect 60737 12087 60795 12093
rect 60737 12053 60749 12087
rect 60783 12084 60795 12087
rect 61746 12084 61752 12096
rect 60783 12056 61752 12084
rect 60783 12053 60795 12056
rect 60737 12047 60795 12053
rect 61746 12044 61752 12056
rect 61804 12044 61810 12096
rect 61930 12044 61936 12096
rect 61988 12084 61994 12096
rect 62132 12084 62160 12115
rect 63678 12084 63684 12096
rect 61988 12056 63684 12084
rect 61988 12044 61994 12056
rect 63678 12044 63684 12056
rect 63736 12044 63742 12096
rect 64782 12044 64788 12096
rect 64840 12084 64846 12096
rect 65153 12087 65211 12093
rect 65153 12084 65165 12087
rect 64840 12056 65165 12084
rect 64840 12044 64846 12056
rect 65153 12053 65165 12056
rect 65199 12053 65211 12087
rect 65886 12084 65892 12096
rect 65847 12056 65892 12084
rect 65153 12047 65211 12053
rect 65886 12044 65892 12056
rect 65944 12044 65950 12096
rect 66180 12084 66208 12124
rect 66530 12112 66536 12164
rect 66588 12152 66594 12164
rect 68189 12155 68247 12161
rect 68189 12152 68201 12155
rect 66588 12124 68201 12152
rect 66588 12112 66594 12124
rect 68189 12121 68201 12124
rect 68235 12121 68247 12155
rect 68189 12115 68247 12121
rect 68738 12112 68744 12164
rect 68796 12112 68802 12164
rect 70762 12112 70768 12164
rect 70820 12152 70826 12164
rect 72510 12152 72516 12164
rect 70820 12124 71544 12152
rect 72358 12124 72516 12152
rect 70820 12112 70826 12124
rect 67634 12084 67640 12096
rect 66180 12056 67640 12084
rect 67634 12044 67640 12056
rect 67692 12044 67698 12096
rect 67726 12044 67732 12096
rect 67784 12084 67790 12096
rect 69661 12087 69719 12093
rect 69661 12084 69673 12087
rect 67784 12056 69673 12084
rect 67784 12044 67790 12056
rect 69661 12053 69673 12056
rect 69707 12053 69719 12087
rect 70302 12084 70308 12096
rect 70263 12056 70308 12084
rect 69661 12047 69719 12053
rect 70302 12044 70308 12056
rect 70360 12044 70366 12096
rect 71130 12044 71136 12096
rect 71188 12084 71194 12096
rect 71314 12084 71320 12096
rect 71188 12056 71320 12084
rect 71188 12044 71194 12056
rect 71314 12044 71320 12056
rect 71372 12044 71378 12096
rect 71516 12084 71544 12124
rect 72510 12112 72516 12124
rect 72568 12112 72574 12164
rect 72694 12112 72700 12164
rect 72752 12152 72758 12164
rect 72789 12155 72847 12161
rect 72789 12152 72801 12155
rect 72752 12124 72801 12152
rect 72752 12112 72758 12124
rect 72789 12121 72801 12124
rect 72835 12121 72847 12155
rect 72789 12115 72847 12121
rect 73080 12084 73108 12183
rect 76374 12180 76380 12232
rect 76432 12220 76438 12232
rect 76432 12192 76477 12220
rect 76432 12180 76438 12192
rect 76650 12180 76656 12232
rect 76708 12220 76714 12232
rect 77018 12220 77024 12232
rect 76708 12192 77024 12220
rect 76708 12180 76714 12192
rect 77018 12180 77024 12192
rect 77076 12180 77082 12232
rect 77205 12223 77263 12229
rect 77205 12189 77217 12223
rect 77251 12189 77263 12223
rect 77205 12183 77263 12189
rect 77297 12223 77355 12229
rect 77297 12189 77309 12223
rect 77343 12220 77355 12223
rect 77404 12220 77432 12328
rect 77938 12316 77944 12328
rect 77996 12316 78002 12368
rect 78033 12359 78091 12365
rect 78033 12325 78045 12359
rect 78079 12356 78091 12359
rect 78079 12328 78904 12356
rect 78079 12325 78091 12328
rect 78033 12319 78091 12325
rect 77570 12248 77576 12300
rect 77628 12288 77634 12300
rect 78490 12288 78496 12300
rect 77628 12260 78352 12288
rect 78451 12260 78496 12288
rect 77628 12248 77634 12260
rect 77343 12192 77432 12220
rect 77343 12189 77355 12192
rect 77297 12183 77355 12189
rect 73801 12155 73859 12161
rect 73801 12121 73813 12155
rect 73847 12152 73859 12155
rect 73890 12152 73896 12164
rect 73847 12124 73896 12152
rect 73847 12121 73859 12124
rect 73801 12115 73859 12121
rect 73890 12112 73896 12124
rect 73948 12112 73954 12164
rect 74534 12112 74540 12164
rect 74592 12112 74598 12164
rect 75546 12112 75552 12164
rect 75604 12152 75610 12164
rect 75604 12124 75776 12152
rect 75604 12112 75610 12124
rect 75086 12084 75092 12096
rect 71516 12056 75092 12084
rect 75086 12044 75092 12056
rect 75144 12084 75150 12096
rect 75638 12084 75644 12096
rect 75144 12056 75644 12084
rect 75144 12044 75150 12056
rect 75638 12044 75644 12056
rect 75696 12044 75702 12096
rect 75748 12084 75776 12124
rect 75914 12112 75920 12164
rect 75972 12152 75978 12164
rect 77220 12152 77248 12183
rect 77478 12180 77484 12232
rect 77536 12220 77542 12232
rect 78324 12229 78352 12260
rect 78490 12248 78496 12260
rect 78548 12248 78554 12300
rect 78876 12288 78904 12328
rect 78950 12316 78956 12368
rect 79008 12356 79014 12368
rect 79594 12356 79600 12368
rect 79008 12328 79600 12356
rect 79008 12316 79014 12328
rect 79594 12316 79600 12328
rect 79652 12316 79658 12368
rect 79870 12316 79876 12368
rect 79928 12356 79934 12368
rect 81066 12356 81072 12368
rect 79928 12328 81072 12356
rect 79928 12316 79934 12328
rect 81066 12316 81072 12328
rect 81124 12316 81130 12368
rect 81250 12356 81256 12368
rect 81211 12328 81256 12356
rect 81250 12316 81256 12328
rect 81308 12316 81314 12368
rect 84010 12356 84016 12368
rect 81544 12328 84016 12356
rect 79226 12288 79232 12300
rect 78876 12260 79232 12288
rect 79226 12248 79232 12260
rect 79284 12248 79290 12300
rect 79778 12248 79784 12300
rect 79836 12288 79842 12300
rect 80330 12288 80336 12300
rect 79836 12260 80336 12288
rect 79836 12248 79842 12260
rect 80330 12248 80336 12260
rect 80388 12248 80394 12300
rect 77941 12223 77999 12229
rect 77941 12220 77953 12223
rect 77536 12192 77953 12220
rect 77536 12180 77542 12192
rect 77941 12189 77953 12192
rect 77987 12189 77999 12223
rect 77941 12183 77999 12189
rect 78309 12223 78367 12229
rect 78309 12189 78321 12223
rect 78355 12220 78367 12223
rect 78398 12220 78404 12232
rect 78355 12192 78404 12220
rect 78355 12189 78367 12192
rect 78309 12183 78367 12189
rect 78398 12180 78404 12192
rect 78456 12180 78462 12232
rect 78953 12223 79011 12229
rect 78953 12189 78965 12223
rect 78999 12220 79011 12223
rect 79870 12220 79876 12232
rect 78999 12192 79876 12220
rect 78999 12189 79011 12192
rect 78953 12183 79011 12189
rect 78968 12152 78996 12183
rect 79870 12180 79876 12192
rect 79928 12180 79934 12232
rect 81544 12220 81572 12328
rect 84010 12316 84016 12328
rect 84068 12356 84074 12368
rect 84562 12356 84568 12368
rect 84068 12328 84568 12356
rect 84068 12316 84074 12328
rect 84562 12316 84568 12328
rect 84620 12316 84626 12368
rect 81710 12288 81716 12300
rect 81671 12260 81716 12288
rect 81710 12248 81716 12260
rect 81768 12248 81774 12300
rect 85206 12288 85212 12300
rect 81912 12260 85212 12288
rect 80026 12192 81572 12220
rect 81621 12223 81679 12229
rect 75972 12124 77248 12152
rect 77404 12124 78996 12152
rect 75972 12112 75978 12124
rect 76190 12084 76196 12096
rect 75748 12056 76196 12084
rect 76190 12044 76196 12056
rect 76248 12084 76254 12096
rect 77404 12084 77432 12124
rect 79042 12112 79048 12164
rect 79100 12152 79106 12164
rect 79778 12152 79784 12164
rect 79100 12124 79784 12152
rect 79100 12112 79106 12124
rect 79778 12112 79784 12124
rect 79836 12112 79842 12164
rect 76248 12056 77432 12084
rect 77481 12087 77539 12093
rect 76248 12044 76254 12056
rect 77481 12053 77493 12087
rect 77527 12084 77539 12087
rect 77846 12084 77852 12096
rect 77527 12056 77852 12084
rect 77527 12053 77539 12056
rect 77481 12047 77539 12053
rect 77846 12044 77852 12056
rect 77904 12044 77910 12096
rect 77938 12044 77944 12096
rect 77996 12084 78002 12096
rect 78674 12084 78680 12096
rect 77996 12056 78680 12084
rect 77996 12044 78002 12056
rect 78674 12044 78680 12056
rect 78732 12044 78738 12096
rect 79594 12044 79600 12096
rect 79652 12084 79658 12096
rect 80026 12084 80054 12192
rect 81621 12189 81633 12223
rect 81667 12220 81679 12223
rect 81802 12220 81808 12232
rect 81667 12192 81808 12220
rect 81667 12189 81679 12192
rect 81621 12183 81679 12189
rect 81802 12180 81808 12192
rect 81860 12180 81866 12232
rect 81158 12112 81164 12164
rect 81216 12152 81222 12164
rect 81912 12152 81940 12260
rect 85206 12248 85212 12260
rect 85264 12248 85270 12300
rect 85574 12288 85580 12300
rect 85535 12260 85580 12288
rect 85574 12248 85580 12260
rect 85632 12248 85638 12300
rect 85850 12288 85856 12300
rect 85811 12260 85856 12288
rect 85850 12248 85856 12260
rect 85908 12248 85914 12300
rect 85960 12288 85988 12396
rect 87782 12384 87788 12436
rect 87840 12424 87846 12436
rect 89717 12427 89775 12433
rect 89717 12424 89729 12427
rect 87840 12396 89729 12424
rect 87840 12384 87846 12396
rect 89717 12393 89729 12396
rect 89763 12393 89775 12427
rect 93302 12424 93308 12436
rect 93263 12396 93308 12424
rect 89717 12387 89775 12393
rect 93302 12384 93308 12396
rect 93360 12384 93366 12436
rect 94222 12424 94228 12436
rect 94183 12396 94228 12424
rect 94222 12384 94228 12396
rect 94280 12384 94286 12436
rect 86218 12316 86224 12368
rect 86276 12356 86282 12368
rect 86276 12328 87736 12356
rect 86276 12316 86282 12328
rect 87601 12291 87659 12297
rect 87601 12288 87613 12291
rect 85960 12260 87613 12288
rect 87601 12257 87613 12260
rect 87647 12257 87659 12291
rect 87601 12251 87659 12257
rect 82265 12223 82323 12229
rect 82265 12189 82277 12223
rect 82311 12189 82323 12223
rect 82265 12183 82323 12189
rect 83001 12223 83059 12229
rect 83001 12189 83013 12223
rect 83047 12220 83059 12223
rect 84102 12220 84108 12232
rect 83047 12192 84108 12220
rect 83047 12189 83059 12192
rect 83001 12183 83059 12189
rect 81216 12124 81940 12152
rect 82280 12152 82308 12183
rect 84102 12180 84108 12192
rect 84160 12180 84166 12232
rect 84194 12180 84200 12232
rect 84252 12180 84258 12232
rect 86218 12180 86224 12232
rect 86276 12220 86282 12232
rect 87708 12229 87736 12328
rect 91833 12291 91891 12297
rect 91833 12257 91845 12291
rect 91879 12288 91891 12291
rect 92474 12288 92480 12300
rect 91879 12260 92480 12288
rect 91879 12257 91891 12260
rect 91833 12251 91891 12257
rect 92474 12248 92480 12260
rect 92532 12248 92538 12300
rect 86589 12223 86647 12229
rect 86589 12220 86601 12223
rect 86276 12192 86601 12220
rect 86276 12180 86282 12192
rect 86589 12189 86601 12192
rect 86635 12189 86647 12223
rect 86589 12183 86647 12189
rect 87693 12223 87751 12229
rect 87693 12189 87705 12223
rect 87739 12189 87751 12223
rect 87693 12183 87751 12189
rect 89530 12180 89536 12232
rect 89588 12220 89594 12232
rect 90361 12223 90419 12229
rect 90361 12220 90373 12223
rect 89588 12192 90373 12220
rect 89588 12180 89594 12192
rect 90361 12189 90373 12192
rect 90407 12189 90419 12223
rect 90361 12183 90419 12189
rect 90637 12223 90695 12229
rect 90637 12189 90649 12223
rect 90683 12220 90695 12223
rect 91557 12223 91615 12229
rect 91557 12220 91569 12223
rect 90683 12192 91569 12220
rect 90683 12189 90695 12192
rect 90637 12183 90695 12189
rect 91557 12189 91569 12192
rect 91603 12189 91615 12223
rect 94038 12220 94044 12232
rect 93999 12192 94044 12220
rect 91557 12183 91615 12189
rect 94038 12180 94044 12192
rect 94096 12180 94102 12232
rect 83553 12155 83611 12161
rect 83553 12152 83565 12155
rect 82280 12124 83565 12152
rect 81216 12112 81222 12124
rect 83553 12121 83565 12124
rect 83599 12152 83611 12155
rect 83642 12152 83648 12164
rect 83599 12124 83648 12152
rect 83599 12121 83611 12124
rect 83553 12115 83611 12121
rect 83642 12112 83648 12124
rect 83700 12152 83706 12164
rect 84212 12152 84240 12180
rect 83700 12124 84240 12152
rect 83700 12112 83706 12124
rect 85114 12112 85120 12164
rect 85172 12112 85178 12164
rect 85574 12112 85580 12164
rect 85632 12152 85638 12164
rect 87049 12155 87107 12161
rect 87049 12152 87061 12155
rect 85632 12124 87061 12152
rect 85632 12112 85638 12124
rect 87049 12121 87061 12124
rect 87095 12121 87107 12155
rect 87049 12115 87107 12121
rect 91094 12112 91100 12164
rect 91152 12152 91158 12164
rect 91152 12124 92322 12152
rect 91152 12112 91158 12124
rect 82354 12084 82360 12096
rect 79652 12056 80054 12084
rect 82315 12056 82360 12084
rect 79652 12044 79658 12056
rect 82354 12044 82360 12056
rect 82412 12044 82418 12096
rect 84194 12044 84200 12096
rect 84252 12084 84258 12096
rect 86497 12087 86555 12093
rect 86497 12084 86509 12087
rect 84252 12056 86509 12084
rect 84252 12044 84258 12056
rect 86497 12053 86509 12056
rect 86543 12053 86555 12087
rect 86497 12047 86555 12053
rect 86954 12044 86960 12096
rect 87012 12084 87018 12096
rect 88613 12087 88671 12093
rect 88613 12084 88625 12087
rect 87012 12056 88625 12084
rect 87012 12044 87018 12056
rect 88613 12053 88625 12056
rect 88659 12053 88671 12087
rect 89162 12084 89168 12096
rect 89123 12056 89168 12084
rect 88613 12047 88671 12053
rect 89162 12044 89168 12056
rect 89220 12044 89226 12096
rect 1104 11994 95011 12016
rect 1104 11942 24386 11994
rect 24438 11942 24450 11994
rect 24502 11942 24514 11994
rect 24566 11942 24578 11994
rect 24630 11942 24642 11994
rect 24694 11942 47823 11994
rect 47875 11942 47887 11994
rect 47939 11942 47951 11994
rect 48003 11942 48015 11994
rect 48067 11942 48079 11994
rect 48131 11942 71260 11994
rect 71312 11942 71324 11994
rect 71376 11942 71388 11994
rect 71440 11942 71452 11994
rect 71504 11942 71516 11994
rect 71568 11942 94697 11994
rect 94749 11942 94761 11994
rect 94813 11942 94825 11994
rect 94877 11942 94889 11994
rect 94941 11942 94953 11994
rect 95005 11942 95011 11994
rect 1104 11920 95011 11942
rect 3970 11840 3976 11892
rect 4028 11880 4034 11892
rect 4522 11880 4528 11892
rect 4028 11852 4384 11880
rect 4483 11852 4528 11880
rect 4028 11840 4034 11852
rect 3050 11812 3056 11824
rect 3011 11784 3056 11812
rect 3050 11772 3056 11784
rect 3108 11772 3114 11824
rect 4356 11812 4384 11852
rect 4522 11840 4528 11852
rect 4580 11840 4586 11892
rect 9674 11880 9680 11892
rect 9635 11852 9680 11880
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 13998 11880 14004 11892
rect 13959 11852 14004 11880
rect 13998 11840 14004 11852
rect 14056 11840 14062 11892
rect 16301 11883 16359 11889
rect 16301 11849 16313 11883
rect 16347 11880 16359 11883
rect 16347 11852 20208 11880
rect 16347 11849 16359 11852
rect 16301 11843 16359 11849
rect 5994 11812 6000 11824
rect 4278 11784 6000 11812
rect 5994 11772 6000 11784
rect 6052 11772 6058 11824
rect 8202 11812 8208 11824
rect 8163 11784 8208 11812
rect 8202 11772 8208 11784
rect 8260 11772 8266 11824
rect 8846 11772 8852 11824
rect 8904 11772 8910 11824
rect 15378 11772 15384 11824
rect 15436 11772 15442 11824
rect 18046 11812 18052 11824
rect 17144 11784 18052 11812
rect 17144 11756 17172 11784
rect 18046 11772 18052 11784
rect 18104 11772 18110 11824
rect 18414 11772 18420 11824
rect 18472 11772 18478 11824
rect 6733 11747 6791 11753
rect 6733 11713 6745 11747
rect 6779 11744 6791 11747
rect 6822 11744 6828 11756
rect 6779 11716 6828 11744
rect 6779 11713 6791 11716
rect 6733 11707 6791 11713
rect 6822 11704 6828 11716
rect 6880 11744 6886 11756
rect 10134 11744 10140 11756
rect 6880 11716 7788 11744
rect 10095 11716 10140 11744
rect 6880 11704 6886 11716
rect 2314 11636 2320 11688
rect 2372 11676 2378 11688
rect 2777 11679 2835 11685
rect 2777 11676 2789 11679
rect 2372 11648 2789 11676
rect 2372 11636 2378 11648
rect 2777 11645 2789 11648
rect 2823 11645 2835 11679
rect 2777 11639 2835 11645
rect 6641 11679 6699 11685
rect 6641 11645 6653 11679
rect 6687 11676 6699 11679
rect 6914 11676 6920 11688
rect 6687 11648 6920 11676
rect 6687 11645 6699 11648
rect 6641 11639 6699 11645
rect 6914 11636 6920 11648
rect 6972 11636 6978 11688
rect 7098 11608 7104 11620
rect 7059 11580 7104 11608
rect 7098 11568 7104 11580
rect 7156 11568 7162 11620
rect 7760 11608 7788 11716
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11744 13139 11747
rect 13354 11744 13360 11756
rect 13127 11716 13360 11744
rect 13127 11713 13139 11716
rect 13081 11707 13139 11713
rect 13354 11704 13360 11716
rect 13412 11704 13418 11756
rect 13906 11744 13912 11756
rect 13867 11716 13912 11744
rect 13906 11704 13912 11716
rect 13964 11704 13970 11756
rect 17126 11744 17132 11756
rect 17039 11716 17132 11744
rect 17126 11704 17132 11716
rect 17184 11704 17190 11756
rect 17494 11704 17500 11756
rect 17552 11744 17558 11756
rect 17681 11747 17739 11753
rect 17681 11744 17693 11747
rect 17552 11716 17693 11744
rect 17552 11704 17558 11716
rect 17681 11713 17693 11716
rect 17727 11713 17739 11747
rect 17681 11707 17739 11713
rect 19242 11704 19248 11756
rect 19300 11744 19306 11756
rect 20180 11753 20208 11852
rect 20364 11852 26924 11880
rect 20165 11747 20223 11753
rect 19300 11716 20116 11744
rect 19300 11704 19306 11716
rect 7926 11676 7932 11688
rect 7887 11648 7932 11676
rect 7926 11636 7932 11648
rect 7984 11636 7990 11688
rect 10413 11679 10471 11685
rect 10413 11676 10425 11679
rect 8036 11648 10425 11676
rect 8036 11608 8064 11648
rect 10413 11645 10425 11648
rect 10459 11645 10471 11679
rect 10413 11639 10471 11645
rect 12253 11679 12311 11685
rect 12253 11645 12265 11679
rect 12299 11676 12311 11679
rect 13170 11676 13176 11688
rect 12299 11648 13176 11676
rect 12299 11645 12311 11648
rect 12253 11639 12311 11645
rect 7760 11580 8064 11608
rect 10428 11608 10456 11639
rect 13170 11636 13176 11648
rect 13228 11636 13234 11688
rect 13538 11636 13544 11688
rect 13596 11676 13602 11688
rect 14553 11679 14611 11685
rect 14553 11676 14565 11679
rect 13596 11648 14565 11676
rect 13596 11636 13602 11648
rect 14553 11645 14565 11648
rect 14599 11645 14611 11679
rect 14826 11676 14832 11688
rect 14787 11648 14832 11676
rect 14553 11639 14611 11645
rect 14458 11608 14464 11620
rect 10428 11580 14464 11608
rect 14458 11568 14464 11580
rect 14516 11568 14522 11620
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 5074 11540 5080 11552
rect 5035 11512 5080 11540
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 5534 11540 5540 11552
rect 5495 11512 5540 11540
rect 5534 11500 5540 11512
rect 5592 11540 5598 11552
rect 11882 11540 11888 11552
rect 5592 11512 11888 11540
rect 5592 11500 5598 11512
rect 11882 11500 11888 11512
rect 11940 11500 11946 11552
rect 12805 11543 12863 11549
rect 12805 11509 12817 11543
rect 12851 11540 12863 11543
rect 12986 11540 12992 11552
rect 12851 11512 12992 11540
rect 12851 11509 12863 11512
rect 12805 11503 12863 11509
rect 12986 11500 12992 11512
rect 13044 11500 13050 11552
rect 14568 11540 14596 11639
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 15194 11636 15200 11688
rect 15252 11676 15258 11688
rect 16114 11676 16120 11688
rect 15252 11648 16120 11676
rect 15252 11636 15258 11648
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 17221 11679 17279 11685
rect 17221 11645 17233 11679
rect 17267 11676 17279 11679
rect 17957 11679 18015 11685
rect 17957 11676 17969 11679
rect 17267 11648 17969 11676
rect 17267 11645 17279 11648
rect 17221 11639 17279 11645
rect 17957 11645 17969 11648
rect 18003 11645 18015 11679
rect 17957 11639 18015 11645
rect 18046 11636 18052 11688
rect 18104 11676 18110 11688
rect 19705 11679 19763 11685
rect 19705 11676 19717 11679
rect 18104 11648 19717 11676
rect 18104 11636 18110 11648
rect 19705 11645 19717 11648
rect 19751 11645 19763 11679
rect 20088 11676 20116 11716
rect 20165 11713 20177 11747
rect 20211 11713 20223 11747
rect 20165 11707 20223 11713
rect 20364 11676 20392 11852
rect 21453 11815 21511 11821
rect 21453 11781 21465 11815
rect 21499 11812 21511 11815
rect 22281 11815 22339 11821
rect 22281 11812 22293 11815
rect 21499 11784 22293 11812
rect 21499 11781 21511 11784
rect 21453 11775 21511 11781
rect 22281 11781 22293 11784
rect 22327 11812 22339 11815
rect 22554 11812 22560 11824
rect 22327 11784 22560 11812
rect 22327 11781 22339 11784
rect 22281 11775 22339 11781
rect 22554 11772 22560 11784
rect 22612 11772 22618 11824
rect 22830 11772 22836 11824
rect 22888 11772 22894 11824
rect 24305 11815 24363 11821
rect 24305 11781 24317 11815
rect 24351 11812 24363 11815
rect 26234 11812 26240 11824
rect 24351 11784 26240 11812
rect 24351 11781 24363 11784
rect 24305 11775 24363 11781
rect 26234 11772 26240 11784
rect 26292 11772 26298 11824
rect 26421 11815 26479 11821
rect 26421 11781 26433 11815
rect 26467 11812 26479 11815
rect 26896 11812 26924 11852
rect 26970 11840 26976 11892
rect 27028 11880 27034 11892
rect 29089 11883 29147 11889
rect 29089 11880 29101 11883
rect 27028 11852 29101 11880
rect 27028 11840 27034 11852
rect 29089 11849 29101 11852
rect 29135 11849 29147 11883
rect 29089 11843 29147 11849
rect 32490 11840 32496 11892
rect 32548 11880 32554 11892
rect 36354 11880 36360 11892
rect 32548 11852 36360 11880
rect 32548 11840 32554 11852
rect 36354 11840 36360 11852
rect 36412 11840 36418 11892
rect 36538 11880 36544 11892
rect 36499 11852 36544 11880
rect 36538 11840 36544 11852
rect 36596 11840 36602 11892
rect 36722 11840 36728 11892
rect 36780 11880 36786 11892
rect 41049 11883 41107 11889
rect 41049 11880 41061 11883
rect 36780 11852 41061 11880
rect 36780 11840 36786 11852
rect 41049 11849 41061 11852
rect 41095 11849 41107 11883
rect 41049 11843 41107 11849
rect 41417 11883 41475 11889
rect 41417 11849 41429 11883
rect 41463 11880 41475 11883
rect 41966 11880 41972 11892
rect 41463 11852 41972 11880
rect 41463 11849 41475 11852
rect 41417 11843 41475 11849
rect 41966 11840 41972 11852
rect 42024 11840 42030 11892
rect 42610 11880 42616 11892
rect 42571 11852 42616 11880
rect 42610 11840 42616 11852
rect 42668 11840 42674 11892
rect 43714 11840 43720 11892
rect 43772 11880 43778 11892
rect 43809 11883 43867 11889
rect 43809 11880 43821 11883
rect 43772 11852 43821 11880
rect 43772 11840 43778 11852
rect 43809 11849 43821 11852
rect 43855 11849 43867 11883
rect 44358 11880 44364 11892
rect 43809 11843 43867 11849
rect 44008 11852 44364 11880
rect 28810 11812 28816 11824
rect 26467 11784 26832 11812
rect 26896 11784 28816 11812
rect 26467 11781 26479 11784
rect 26421 11775 26479 11781
rect 20441 11747 20499 11753
rect 20441 11713 20453 11747
rect 20487 11744 20499 11747
rect 21910 11744 21916 11756
rect 20487 11716 21916 11744
rect 20487 11713 20499 11716
rect 20441 11707 20499 11713
rect 21910 11704 21916 11716
rect 21968 11704 21974 11756
rect 21634 11676 21640 11688
rect 20088 11648 20392 11676
rect 20456 11648 21640 11676
rect 19705 11639 19763 11645
rect 20456 11608 20484 11648
rect 21634 11636 21640 11648
rect 21692 11676 21698 11688
rect 22005 11679 22063 11685
rect 22005 11676 22017 11679
rect 21692 11648 22017 11676
rect 21692 11636 21698 11648
rect 22005 11645 22017 11648
rect 22051 11645 22063 11679
rect 25038 11676 25044 11688
rect 24999 11648 25044 11676
rect 22005 11639 22063 11645
rect 25038 11636 25044 11648
rect 25096 11676 25102 11688
rect 26050 11676 26056 11688
rect 25096 11648 26056 11676
rect 25096 11636 25102 11648
rect 26050 11636 26056 11648
rect 26108 11636 26114 11688
rect 26602 11676 26608 11688
rect 26563 11648 26608 11676
rect 26602 11636 26608 11648
rect 26660 11636 26666 11688
rect 26804 11676 26832 11784
rect 28810 11772 28816 11784
rect 28868 11772 28874 11824
rect 30650 11812 30656 11824
rect 30563 11784 30656 11812
rect 30650 11772 30656 11784
rect 30708 11812 30714 11824
rect 31110 11812 31116 11824
rect 30708 11784 31116 11812
rect 30708 11772 30714 11784
rect 31110 11772 31116 11784
rect 31168 11772 31174 11824
rect 33778 11772 33784 11824
rect 33836 11812 33842 11824
rect 37182 11812 37188 11824
rect 33836 11784 37188 11812
rect 33836 11772 33842 11784
rect 37182 11772 37188 11784
rect 37240 11772 37246 11824
rect 37458 11772 37464 11824
rect 37516 11812 37522 11824
rect 38838 11812 38844 11824
rect 37516 11784 38844 11812
rect 37516 11772 37522 11784
rect 27154 11704 27160 11756
rect 27212 11744 27218 11756
rect 27525 11747 27583 11753
rect 27525 11744 27537 11747
rect 27212 11716 27537 11744
rect 27212 11704 27218 11716
rect 27525 11713 27537 11716
rect 27571 11744 27583 11747
rect 28994 11744 29000 11756
rect 27571 11716 29000 11744
rect 27571 11713 27583 11716
rect 27525 11707 27583 11713
rect 28994 11704 29000 11716
rect 29052 11704 29058 11756
rect 29454 11744 29460 11756
rect 29415 11716 29460 11744
rect 29454 11704 29460 11716
rect 29512 11704 29518 11756
rect 30387 11747 30445 11753
rect 30387 11713 30399 11747
rect 30433 11713 30445 11747
rect 30387 11707 30445 11713
rect 26804 11648 27384 11676
rect 27157 11611 27215 11617
rect 27157 11608 27169 11611
rect 16224 11580 17816 11608
rect 16224 11540 16252 11580
rect 14568 11512 16252 11540
rect 17788 11540 17816 11580
rect 19996 11580 20484 11608
rect 23308 11580 27169 11608
rect 19996 11552 20024 11580
rect 19978 11540 19984 11552
rect 17788 11512 19984 11540
rect 19978 11500 19984 11512
rect 20036 11500 20042 11552
rect 20162 11500 20168 11552
rect 20220 11540 20226 11552
rect 23308 11540 23336 11580
rect 27157 11577 27169 11580
rect 27203 11577 27215 11611
rect 27356 11608 27384 11648
rect 27430 11636 27436 11688
rect 27488 11676 27494 11688
rect 27488 11648 27533 11676
rect 27488 11636 27494 11648
rect 27798 11636 27804 11688
rect 27856 11676 27862 11688
rect 28537 11679 28595 11685
rect 28537 11676 28549 11679
rect 27856 11648 28549 11676
rect 27856 11636 27862 11648
rect 28537 11645 28549 11648
rect 28583 11676 28595 11679
rect 28810 11676 28816 11688
rect 28583 11648 28816 11676
rect 28583 11645 28595 11648
rect 28537 11639 28595 11645
rect 28810 11636 28816 11648
rect 28868 11636 28874 11688
rect 28902 11636 28908 11688
rect 28960 11676 28966 11688
rect 29178 11676 29184 11688
rect 28960 11648 29184 11676
rect 28960 11636 28966 11648
rect 29178 11636 29184 11648
rect 29236 11636 29242 11688
rect 29362 11636 29368 11688
rect 29420 11676 29426 11688
rect 30392 11676 30420 11707
rect 31570 11704 31576 11756
rect 31628 11744 31634 11756
rect 33962 11744 33968 11756
rect 31628 11716 33824 11744
rect 33923 11716 33968 11744
rect 31628 11704 31634 11716
rect 29420 11648 29465 11676
rect 30300 11648 30420 11676
rect 33229 11679 33287 11685
rect 29420 11636 29426 11648
rect 27890 11608 27896 11620
rect 27356 11580 27896 11608
rect 27157 11571 27215 11577
rect 27890 11568 27896 11580
rect 27948 11568 27954 11620
rect 30300 11608 30328 11648
rect 33229 11645 33241 11679
rect 33275 11676 33287 11679
rect 33502 11676 33508 11688
rect 33275 11648 33508 11676
rect 33275 11645 33287 11648
rect 33229 11639 33287 11645
rect 33502 11636 33508 11648
rect 33560 11636 33566 11688
rect 33796 11676 33824 11716
rect 33962 11704 33968 11716
rect 34020 11704 34026 11756
rect 34149 11747 34207 11753
rect 34149 11713 34161 11747
rect 34195 11744 34207 11747
rect 34974 11744 34980 11756
rect 34195 11716 34980 11744
rect 34195 11713 34207 11716
rect 34149 11707 34207 11713
rect 34974 11704 34980 11716
rect 35032 11704 35038 11756
rect 35253 11747 35311 11753
rect 35253 11713 35265 11747
rect 35299 11744 35311 11747
rect 35529 11747 35587 11753
rect 35299 11716 35388 11744
rect 35299 11713 35311 11716
rect 35253 11707 35311 11713
rect 35360 11676 35388 11716
rect 35529 11713 35541 11747
rect 35575 11744 35587 11747
rect 36446 11744 36452 11756
rect 35575 11716 36452 11744
rect 35575 11713 35587 11716
rect 35529 11707 35587 11713
rect 36446 11704 36452 11716
rect 36504 11704 36510 11756
rect 36630 11744 36636 11756
rect 36591 11716 36636 11744
rect 36630 11704 36636 11716
rect 36688 11704 36694 11756
rect 38013 11747 38071 11753
rect 38013 11713 38025 11747
rect 38059 11713 38071 11747
rect 38580 11730 38608 11784
rect 38838 11772 38844 11784
rect 38896 11772 38902 11824
rect 39022 11812 39028 11824
rect 38983 11784 39028 11812
rect 39022 11772 39028 11784
rect 39080 11772 39086 11824
rect 40586 11772 40592 11824
rect 40644 11812 40650 11824
rect 41509 11815 41567 11821
rect 40644 11784 40689 11812
rect 40644 11772 40650 11784
rect 41509 11781 41521 11815
rect 41555 11812 41567 11815
rect 44008 11812 44036 11852
rect 44358 11840 44364 11852
rect 44416 11840 44422 11892
rect 51997 11883 52055 11889
rect 51997 11880 52009 11883
rect 44468 11852 52009 11880
rect 41555 11784 44036 11812
rect 41555 11781 41567 11784
rect 41509 11775 41567 11781
rect 44082 11772 44088 11824
rect 44140 11812 44146 11824
rect 44468 11812 44496 11852
rect 51997 11849 52009 11852
rect 52043 11849 52055 11883
rect 51997 11843 52055 11849
rect 52822 11840 52828 11892
rect 52880 11880 52886 11892
rect 53009 11883 53067 11889
rect 53009 11880 53021 11883
rect 52880 11852 53021 11880
rect 52880 11840 52886 11852
rect 53009 11849 53021 11852
rect 53055 11880 53067 11883
rect 53742 11880 53748 11892
rect 53055 11852 53748 11880
rect 53055 11849 53067 11852
rect 53009 11843 53067 11849
rect 53742 11840 53748 11852
rect 53800 11840 53806 11892
rect 58802 11880 58808 11892
rect 56152 11852 58808 11880
rect 45646 11812 45652 11824
rect 44140 11784 44496 11812
rect 44560 11784 45652 11812
rect 44140 11772 44146 11784
rect 40224 11756 40276 11762
rect 38013 11707 38071 11713
rect 33796 11648 35388 11676
rect 28552 11580 30328 11608
rect 20220 11512 23336 11540
rect 23753 11543 23811 11549
rect 20220 11500 20226 11512
rect 23753 11509 23765 11543
rect 23799 11540 23811 11543
rect 28552 11540 28580 11580
rect 31478 11568 31484 11620
rect 31536 11608 31542 11620
rect 35360 11608 35388 11648
rect 35434 11636 35440 11688
rect 35492 11676 35498 11688
rect 35805 11679 35863 11685
rect 35805 11676 35817 11679
rect 35492 11648 35817 11676
rect 35492 11636 35498 11648
rect 35805 11645 35817 11648
rect 35851 11645 35863 11679
rect 35805 11639 35863 11645
rect 36354 11636 36360 11688
rect 36412 11676 36418 11688
rect 38028 11676 38056 11707
rect 41414 11704 41420 11756
rect 41472 11744 41478 11756
rect 42981 11747 43039 11753
rect 42981 11744 42993 11747
rect 41472 11716 42993 11744
rect 41472 11704 41478 11716
rect 42981 11713 42993 11716
rect 43027 11744 43039 11747
rect 44560 11744 44588 11784
rect 45646 11772 45652 11784
rect 45704 11772 45710 11824
rect 46566 11812 46572 11824
rect 46527 11784 46572 11812
rect 46566 11772 46572 11784
rect 46624 11772 46630 11824
rect 50246 11812 50252 11824
rect 48424 11784 50252 11812
rect 43027 11716 44588 11744
rect 44836 11716 45416 11744
rect 43027 11713 43039 11716
rect 42981 11707 43039 11713
rect 40224 11698 40276 11704
rect 36412 11648 38056 11676
rect 36412 11636 36418 11648
rect 37734 11608 37740 11620
rect 31536 11580 32260 11608
rect 35360 11580 37740 11608
rect 31536 11568 31542 11580
rect 23799 11512 28580 11540
rect 23799 11509 23811 11512
rect 23753 11503 23811 11509
rect 28626 11500 28632 11552
rect 28684 11540 28690 11552
rect 31570 11540 31576 11552
rect 28684 11512 31576 11540
rect 28684 11500 28690 11512
rect 31570 11500 31576 11512
rect 31628 11540 31634 11552
rect 31757 11543 31815 11549
rect 31757 11540 31769 11543
rect 31628 11512 31769 11540
rect 31628 11500 31634 11512
rect 31757 11509 31769 11512
rect 31803 11509 31815 11543
rect 32232 11540 32260 11580
rect 37734 11568 37740 11580
rect 37792 11568 37798 11620
rect 38028 11608 38056 11648
rect 38378 11636 38384 11688
rect 38436 11676 38442 11688
rect 39574 11676 39580 11688
rect 38436 11648 39580 11676
rect 38436 11636 38442 11648
rect 39574 11636 39580 11648
rect 39632 11636 39638 11688
rect 39758 11676 39764 11688
rect 39719 11648 39764 11676
rect 39758 11636 39764 11648
rect 39816 11636 39822 11688
rect 41598 11636 41604 11688
rect 41656 11676 41662 11688
rect 41656 11648 41701 11676
rect 41656 11636 41662 11648
rect 42886 11636 42892 11688
rect 42944 11676 42950 11688
rect 43073 11679 43131 11685
rect 43073 11676 43085 11679
rect 42944 11648 43085 11676
rect 42944 11636 42950 11648
rect 43073 11645 43085 11648
rect 43119 11676 43131 11679
rect 44082 11676 44088 11688
rect 43119 11648 44088 11676
rect 43119 11645 43131 11648
rect 43073 11639 43131 11645
rect 44082 11636 44088 11648
rect 44140 11636 44146 11688
rect 44358 11676 44364 11688
rect 44319 11648 44364 11676
rect 44358 11636 44364 11648
rect 44416 11676 44422 11688
rect 44836 11676 44864 11716
rect 44416 11648 44864 11676
rect 44913 11679 44971 11685
rect 44416 11636 44422 11648
rect 44913 11645 44925 11679
rect 44959 11645 44971 11679
rect 45388 11676 45416 11716
rect 46842 11704 46848 11756
rect 46900 11744 46906 11756
rect 48424 11744 48452 11784
rect 50246 11772 50252 11784
rect 50304 11812 50310 11824
rect 51261 11815 51319 11821
rect 50304 11784 51074 11812
rect 50304 11772 50310 11784
rect 50154 11744 50160 11756
rect 46900 11730 48452 11744
rect 46900 11716 48438 11730
rect 49068 11716 50160 11744
rect 46900 11704 46906 11716
rect 46014 11676 46020 11688
rect 45388 11648 46020 11676
rect 44913 11639 44971 11645
rect 38194 11608 38200 11620
rect 38028 11580 38200 11608
rect 38194 11568 38200 11580
rect 38252 11568 38258 11620
rect 38286 11568 38292 11620
rect 38344 11608 38350 11620
rect 44928 11608 44956 11639
rect 46014 11636 46020 11648
rect 46072 11636 46078 11688
rect 46290 11636 46296 11688
rect 46348 11676 46354 11688
rect 46753 11679 46811 11685
rect 46753 11676 46765 11679
rect 46348 11648 46765 11676
rect 46348 11636 46354 11648
rect 46753 11645 46765 11648
rect 46799 11645 46811 11679
rect 46753 11639 46811 11645
rect 47578 11636 47584 11688
rect 47636 11676 47642 11688
rect 48501 11679 48559 11685
rect 48501 11676 48513 11679
rect 47636 11648 48513 11676
rect 47636 11636 47642 11648
rect 48501 11645 48513 11648
rect 48547 11676 48559 11679
rect 49068 11676 49096 11716
rect 50154 11704 50160 11716
rect 50212 11744 50218 11756
rect 50212 11716 50292 11744
rect 50356 11730 50384 11784
rect 51046 11744 51074 11784
rect 51261 11781 51273 11815
rect 51307 11812 51319 11815
rect 52270 11812 52276 11824
rect 51307 11784 52276 11812
rect 51307 11781 51319 11784
rect 51261 11775 51319 11781
rect 52270 11772 52276 11784
rect 52328 11772 52334 11824
rect 54294 11812 54300 11824
rect 53760 11784 54300 11812
rect 51902 11744 51908 11756
rect 51046 11716 51908 11744
rect 50212 11704 50218 11716
rect 49326 11676 49332 11688
rect 48547 11648 49096 11676
rect 49287 11648 49332 11676
rect 48547 11645 48559 11648
rect 48501 11639 48559 11645
rect 49326 11636 49332 11648
rect 49384 11636 49390 11688
rect 50264 11676 50292 11716
rect 51902 11704 51908 11716
rect 51960 11704 51966 11756
rect 52178 11744 52184 11756
rect 52139 11716 52184 11744
rect 52178 11704 52184 11716
rect 52236 11704 52242 11756
rect 52362 11744 52368 11756
rect 52323 11716 52368 11744
rect 52362 11704 52368 11716
rect 52420 11704 52426 11756
rect 52914 11744 52920 11756
rect 52875 11716 52920 11744
rect 52914 11704 52920 11716
rect 52972 11704 52978 11756
rect 53006 11704 53012 11756
rect 53064 11744 53070 11756
rect 53101 11747 53159 11753
rect 53101 11744 53113 11747
rect 53064 11716 53113 11744
rect 53064 11704 53070 11716
rect 53101 11713 53113 11716
rect 53147 11713 53159 11747
rect 53101 11707 53159 11713
rect 50433 11679 50491 11685
rect 50433 11676 50445 11679
rect 50264 11648 50445 11676
rect 50433 11645 50445 11648
rect 50479 11645 50491 11679
rect 50433 11639 50491 11645
rect 50522 11636 50528 11688
rect 50580 11676 50586 11688
rect 50580 11648 51212 11676
rect 50580 11636 50586 11648
rect 45186 11608 45192 11620
rect 38344 11580 45192 11608
rect 38344 11568 38350 11580
rect 45186 11568 45192 11580
rect 45244 11608 45250 11620
rect 45554 11608 45560 11620
rect 45244 11580 45560 11608
rect 45244 11568 45250 11580
rect 45554 11568 45560 11580
rect 45612 11568 45618 11620
rect 49602 11608 49608 11620
rect 45664 11580 49608 11608
rect 32585 11543 32643 11549
rect 32585 11540 32597 11543
rect 32232 11512 32597 11540
rect 31757 11503 31815 11509
rect 32585 11509 32597 11512
rect 32631 11540 32643 11543
rect 33410 11540 33416 11552
rect 32631 11512 33416 11540
rect 32631 11509 32643 11512
rect 32585 11503 32643 11509
rect 33410 11500 33416 11512
rect 33468 11500 33474 11552
rect 35710 11500 35716 11552
rect 35768 11540 35774 11552
rect 37458 11540 37464 11552
rect 35768 11512 37464 11540
rect 35768 11500 35774 11512
rect 37458 11500 37464 11512
rect 37516 11500 37522 11552
rect 41966 11500 41972 11552
rect 42024 11540 42030 11552
rect 45664 11540 45692 11580
rect 49602 11568 49608 11580
rect 49660 11568 49666 11620
rect 51184 11608 51212 11648
rect 51258 11636 51264 11688
rect 51316 11676 51322 11688
rect 52196 11676 52224 11704
rect 51316 11648 52224 11676
rect 51316 11636 51322 11648
rect 52270 11636 52276 11688
rect 52328 11676 52334 11688
rect 53760 11685 53788 11784
rect 54294 11772 54300 11784
rect 54352 11772 54358 11824
rect 54389 11747 54447 11753
rect 54389 11713 54401 11747
rect 54435 11744 54447 11747
rect 54846 11744 54852 11756
rect 54435 11716 54852 11744
rect 54435 11713 54447 11716
rect 54389 11707 54447 11713
rect 54846 11704 54852 11716
rect 54904 11704 54910 11756
rect 55030 11744 55036 11756
rect 54991 11716 55036 11744
rect 55030 11704 55036 11716
rect 55088 11704 55094 11756
rect 56152 11753 56180 11852
rect 58802 11840 58808 11852
rect 58860 11880 58866 11892
rect 61565 11883 61623 11889
rect 58860 11852 58940 11880
rect 58860 11840 58866 11852
rect 57514 11812 57520 11824
rect 57475 11784 57520 11812
rect 57514 11772 57520 11784
rect 57572 11772 57578 11824
rect 58912 11812 58940 11852
rect 61565 11849 61577 11883
rect 61611 11880 61623 11883
rect 62298 11880 62304 11892
rect 61611 11852 62304 11880
rect 61611 11849 61623 11852
rect 61565 11843 61623 11849
rect 62298 11840 62304 11852
rect 62356 11840 62362 11892
rect 63310 11840 63316 11892
rect 63368 11840 63374 11892
rect 63678 11840 63684 11892
rect 63736 11880 63742 11892
rect 65613 11883 65671 11889
rect 65613 11880 65625 11883
rect 63736 11852 65625 11880
rect 63736 11840 63742 11852
rect 65613 11849 65625 11852
rect 65659 11849 65671 11883
rect 69842 11880 69848 11892
rect 65613 11843 65671 11849
rect 65996 11852 69848 11880
rect 62114 11812 62120 11824
rect 58912 11784 62120 11812
rect 62114 11772 62120 11784
rect 62172 11772 62178 11824
rect 63218 11812 63224 11824
rect 62408 11784 63224 11812
rect 56137 11747 56195 11753
rect 56137 11713 56149 11747
rect 56183 11713 56195 11747
rect 56686 11744 56692 11756
rect 56647 11716 56692 11744
rect 56137 11707 56195 11713
rect 56686 11704 56692 11716
rect 56744 11704 56750 11756
rect 57333 11747 57391 11753
rect 57333 11713 57345 11747
rect 57379 11744 57391 11747
rect 57790 11744 57796 11756
rect 57379 11716 57796 11744
rect 57379 11713 57391 11716
rect 57333 11707 57391 11713
rect 57790 11704 57796 11716
rect 57848 11704 57854 11756
rect 58250 11744 58256 11756
rect 58211 11716 58256 11744
rect 58250 11704 58256 11716
rect 58308 11704 58314 11756
rect 58416 11747 58474 11753
rect 58416 11744 58428 11747
rect 58360 11716 58428 11744
rect 53745 11679 53803 11685
rect 53745 11676 53757 11679
rect 52328 11648 53757 11676
rect 52328 11636 52334 11648
rect 53745 11645 53757 11648
rect 53791 11645 53803 11679
rect 53745 11639 53803 11645
rect 56318 11636 56324 11688
rect 56376 11676 56382 11688
rect 57149 11679 57207 11685
rect 57149 11676 57161 11679
rect 56376 11648 57161 11676
rect 56376 11636 56382 11648
rect 57149 11645 57161 11648
rect 57195 11676 57207 11679
rect 58360 11676 58388 11716
rect 58416 11713 58428 11716
rect 58462 11713 58474 11747
rect 58416 11707 58474 11713
rect 58526 11704 58532 11756
rect 58584 11744 58590 11756
rect 58710 11753 58716 11756
rect 58667 11747 58716 11753
rect 58584 11716 58629 11744
rect 58584 11704 58590 11716
rect 58667 11713 58679 11747
rect 58713 11713 58716 11747
rect 58667 11707 58716 11713
rect 58710 11704 58716 11707
rect 58768 11704 58774 11756
rect 58894 11704 58900 11756
rect 58952 11744 58958 11756
rect 62408 11753 62436 11784
rect 63218 11772 63224 11784
rect 63276 11772 63282 11824
rect 63328 11812 63356 11840
rect 63589 11815 63647 11821
rect 63589 11812 63601 11815
rect 63328 11784 63601 11812
rect 63589 11781 63601 11784
rect 63635 11781 63647 11815
rect 65886 11812 65892 11824
rect 64814 11784 65892 11812
rect 63589 11775 63647 11781
rect 65886 11772 65892 11784
rect 65944 11772 65950 11824
rect 61933 11747 61991 11753
rect 61933 11744 61945 11747
rect 58952 11716 61945 11744
rect 58952 11704 58958 11716
rect 61933 11713 61945 11716
rect 61979 11713 61991 11747
rect 61933 11707 61991 11713
rect 62393 11747 62451 11753
rect 62393 11713 62405 11747
rect 62439 11713 62451 11747
rect 62393 11707 62451 11713
rect 57195 11648 58388 11676
rect 61948 11676 61976 11707
rect 63126 11704 63132 11756
rect 63184 11744 63190 11756
rect 63313 11747 63371 11753
rect 63313 11744 63325 11747
rect 63184 11716 63325 11744
rect 63184 11704 63190 11716
rect 63313 11713 63325 11716
rect 63359 11713 63371 11747
rect 63313 11707 63371 11713
rect 63586 11676 63592 11688
rect 61948 11648 63592 11676
rect 57195 11645 57207 11648
rect 57149 11639 57207 11645
rect 63586 11636 63592 11648
rect 63644 11676 63650 11688
rect 64782 11676 64788 11688
rect 63644 11648 64788 11676
rect 63644 11636 63650 11648
rect 64782 11636 64788 11648
rect 64840 11636 64846 11688
rect 65058 11676 65064 11688
rect 64971 11648 65064 11676
rect 65058 11636 65064 11648
rect 65116 11676 65122 11688
rect 65996 11676 66024 11852
rect 69842 11840 69848 11852
rect 69900 11840 69906 11892
rect 71774 11840 71780 11892
rect 71832 11880 71838 11892
rect 72602 11880 72608 11892
rect 71832 11852 72608 11880
rect 71832 11840 71838 11852
rect 72602 11840 72608 11852
rect 72660 11840 72666 11892
rect 73614 11880 73620 11892
rect 73575 11852 73620 11880
rect 73614 11840 73620 11852
rect 73672 11840 73678 11892
rect 75362 11880 75368 11892
rect 74000 11852 75368 11880
rect 74000 11824 74028 11852
rect 75362 11840 75368 11852
rect 75420 11840 75426 11892
rect 77110 11840 77116 11892
rect 77168 11880 77174 11892
rect 78674 11880 78680 11892
rect 77168 11852 78680 11880
rect 77168 11840 77174 11852
rect 78674 11840 78680 11852
rect 78732 11880 78738 11892
rect 78769 11883 78827 11889
rect 78769 11880 78781 11883
rect 78732 11852 78781 11880
rect 78732 11840 78738 11852
rect 78769 11849 78781 11852
rect 78815 11880 78827 11883
rect 79318 11880 79324 11892
rect 78815 11852 79324 11880
rect 78815 11849 78827 11852
rect 78769 11843 78827 11849
rect 79318 11840 79324 11852
rect 79376 11840 79382 11892
rect 80606 11880 80612 11892
rect 79612 11852 80612 11880
rect 79612 11824 79640 11852
rect 80606 11840 80612 11852
rect 80664 11840 80670 11892
rect 84194 11880 84200 11892
rect 81820 11852 84200 11880
rect 66070 11772 66076 11824
rect 66128 11812 66134 11824
rect 67726 11812 67732 11824
rect 66128 11784 67732 11812
rect 66128 11772 66134 11784
rect 67726 11772 67732 11784
rect 67784 11772 67790 11824
rect 68370 11812 68376 11824
rect 68331 11784 68376 11812
rect 68370 11772 68376 11784
rect 68428 11772 68434 11824
rect 69934 11772 69940 11824
rect 69992 11812 69998 11824
rect 73982 11812 73988 11824
rect 69992 11784 71268 11812
rect 69992 11772 69998 11784
rect 67358 11744 67364 11756
rect 67319 11716 67364 11744
rect 67358 11704 67364 11716
rect 67416 11704 67422 11756
rect 67545 11747 67603 11753
rect 67545 11713 67557 11747
rect 67591 11744 67603 11747
rect 67818 11744 67824 11756
rect 67591 11716 67824 11744
rect 67591 11713 67603 11716
rect 67545 11707 67603 11713
rect 67818 11704 67824 11716
rect 67876 11704 67882 11756
rect 68002 11704 68008 11756
rect 68060 11744 68066 11756
rect 71130 11744 71136 11756
rect 68060 11716 70164 11744
rect 71091 11716 71136 11744
rect 68060 11704 68066 11716
rect 65116 11648 66024 11676
rect 65116 11636 65122 11648
rect 66162 11636 66168 11688
rect 66220 11676 66226 11688
rect 66533 11679 66591 11685
rect 66533 11676 66545 11679
rect 66220 11648 66545 11676
rect 66220 11636 66226 11648
rect 66533 11645 66545 11648
rect 66579 11645 66591 11679
rect 67266 11676 67272 11688
rect 66533 11639 66591 11645
rect 66640 11648 67272 11676
rect 52914 11608 52920 11620
rect 51184 11580 52920 11608
rect 52914 11568 52920 11580
rect 52972 11568 52978 11620
rect 56502 11568 56508 11620
rect 56560 11608 56566 11620
rect 56597 11611 56655 11617
rect 56597 11608 56609 11611
rect 56560 11580 56609 11608
rect 56560 11568 56566 11580
rect 56597 11577 56609 11580
rect 56643 11577 56655 11611
rect 59909 11611 59967 11617
rect 59909 11608 59921 11611
rect 56597 11571 56655 11577
rect 59004 11580 59921 11608
rect 59004 11552 59032 11580
rect 59909 11577 59921 11580
rect 59955 11608 59967 11611
rect 60090 11608 60096 11620
rect 59955 11580 60096 11608
rect 59955 11577 59967 11580
rect 59909 11571 59967 11577
rect 60090 11568 60096 11580
rect 60148 11568 60154 11620
rect 61013 11611 61071 11617
rect 61013 11608 61025 11611
rect 60292 11580 61025 11608
rect 42024 11512 45692 11540
rect 42024 11500 42030 11512
rect 45738 11500 45744 11552
rect 45796 11540 45802 11552
rect 46842 11540 46848 11552
rect 45796 11512 46848 11540
rect 45796 11500 45802 11512
rect 46842 11500 46848 11512
rect 46900 11500 46906 11552
rect 50430 11500 50436 11552
rect 50488 11540 50494 11552
rect 51166 11540 51172 11552
rect 50488 11512 51172 11540
rect 50488 11500 50494 11512
rect 51166 11500 51172 11512
rect 51224 11500 51230 11552
rect 51258 11500 51264 11552
rect 51316 11540 51322 11552
rect 52270 11540 52276 11552
rect 51316 11512 52276 11540
rect 51316 11500 51322 11512
rect 52270 11500 52276 11512
rect 52328 11500 52334 11552
rect 52365 11543 52423 11549
rect 52365 11509 52377 11543
rect 52411 11540 52423 11543
rect 53006 11540 53012 11552
rect 52411 11512 53012 11540
rect 52411 11509 52423 11512
rect 52365 11503 52423 11509
rect 53006 11500 53012 11512
rect 53064 11500 53070 11552
rect 53650 11500 53656 11552
rect 53708 11540 53714 11552
rect 56134 11540 56140 11552
rect 53708 11512 56140 11540
rect 53708 11500 53714 11512
rect 56134 11500 56140 11512
rect 56192 11540 56198 11552
rect 57882 11540 57888 11552
rect 56192 11512 57888 11540
rect 56192 11500 56198 11512
rect 57882 11500 57888 11512
rect 57940 11500 57946 11552
rect 57974 11500 57980 11552
rect 58032 11540 58038 11552
rect 58618 11540 58624 11552
rect 58032 11512 58624 11540
rect 58032 11500 58038 11512
rect 58618 11500 58624 11512
rect 58676 11500 58682 11552
rect 58894 11540 58900 11552
rect 58855 11512 58900 11540
rect 58894 11500 58900 11512
rect 58952 11500 58958 11552
rect 58986 11500 58992 11552
rect 59044 11500 59050 11552
rect 59354 11540 59360 11552
rect 59315 11512 59360 11540
rect 59354 11500 59360 11512
rect 59412 11500 59418 11552
rect 59998 11500 60004 11552
rect 60056 11540 60062 11552
rect 60292 11540 60320 11580
rect 61013 11577 61025 11580
rect 61059 11577 61071 11611
rect 61013 11571 61071 11577
rect 64966 11568 64972 11620
rect 65024 11608 65030 11620
rect 65886 11608 65892 11620
rect 65024 11580 65892 11608
rect 65024 11568 65030 11580
rect 65886 11568 65892 11580
rect 65944 11608 65950 11620
rect 66640 11608 66668 11648
rect 67266 11636 67272 11648
rect 67324 11636 67330 11688
rect 70136 11676 70164 11716
rect 71130 11704 71136 11716
rect 71188 11704 71194 11756
rect 71240 11753 71268 11784
rect 71976 11784 73988 11812
rect 71225 11747 71283 11753
rect 71225 11713 71237 11747
rect 71271 11713 71283 11747
rect 71225 11707 71283 11713
rect 70581 11679 70639 11685
rect 70581 11676 70593 11679
rect 70136 11648 70593 11676
rect 70581 11645 70593 11648
rect 70627 11645 70639 11679
rect 70581 11639 70639 11645
rect 70670 11636 70676 11688
rect 70728 11676 70734 11688
rect 71976 11676 72004 11784
rect 73982 11772 73988 11784
rect 74040 11772 74046 11824
rect 74166 11812 74172 11824
rect 74127 11784 74172 11812
rect 74166 11772 74172 11784
rect 74224 11772 74230 11824
rect 75457 11815 75515 11821
rect 75457 11781 75469 11815
rect 75503 11812 75515 11815
rect 75730 11812 75736 11824
rect 75503 11784 75736 11812
rect 75503 11781 75515 11784
rect 75457 11775 75515 11781
rect 75730 11772 75736 11784
rect 75788 11772 75794 11824
rect 79594 11812 79600 11824
rect 76116 11784 79600 11812
rect 72050 11704 72056 11756
rect 72108 11744 72114 11756
rect 72145 11747 72203 11753
rect 72145 11744 72157 11747
rect 72108 11716 72157 11744
rect 72108 11704 72114 11716
rect 72145 11713 72157 11716
rect 72191 11713 72203 11747
rect 72145 11707 72203 11713
rect 72234 11704 72240 11756
rect 72292 11744 72298 11756
rect 72329 11747 72387 11753
rect 72329 11744 72341 11747
rect 72292 11716 72341 11744
rect 72292 11704 72298 11716
rect 72329 11713 72341 11716
rect 72375 11713 72387 11747
rect 72329 11707 72387 11713
rect 72421 11747 72479 11753
rect 72421 11713 72433 11747
rect 72467 11744 72479 11747
rect 72602 11744 72608 11756
rect 72467 11716 72608 11744
rect 72467 11713 72479 11716
rect 72421 11707 72479 11713
rect 72602 11704 72608 11716
rect 72660 11704 72666 11756
rect 72697 11747 72755 11753
rect 72697 11713 72709 11747
rect 72743 11744 72755 11747
rect 72786 11744 72792 11756
rect 72743 11716 72792 11744
rect 72743 11713 72755 11716
rect 72697 11707 72755 11713
rect 72786 11704 72792 11716
rect 72844 11704 72850 11756
rect 73522 11744 73528 11756
rect 73483 11716 73528 11744
rect 73522 11704 73528 11716
rect 73580 11704 73586 11756
rect 75362 11744 75368 11756
rect 75323 11716 75368 11744
rect 75362 11704 75368 11716
rect 75420 11704 75426 11756
rect 75546 11744 75552 11756
rect 75507 11716 75552 11744
rect 75546 11704 75552 11716
rect 75604 11704 75610 11756
rect 75914 11704 75920 11756
rect 75972 11744 75978 11756
rect 76009 11747 76067 11753
rect 76009 11744 76021 11747
rect 75972 11716 76021 11744
rect 75972 11704 75978 11716
rect 76009 11713 76021 11716
rect 76055 11713 76067 11747
rect 76009 11707 76067 11713
rect 70728 11648 72004 11676
rect 72513 11679 72571 11685
rect 70728 11636 70734 11648
rect 72513 11645 72525 11679
rect 72559 11676 72571 11679
rect 74074 11676 74080 11688
rect 72559 11648 74080 11676
rect 72559 11645 72571 11648
rect 72513 11639 72571 11645
rect 74074 11636 74080 11648
rect 74132 11636 74138 11688
rect 74718 11676 74724 11688
rect 74679 11648 74724 11676
rect 74718 11636 74724 11648
rect 74776 11676 74782 11688
rect 75822 11676 75828 11688
rect 74776 11648 75828 11676
rect 74776 11636 74782 11648
rect 75822 11636 75828 11648
rect 75880 11636 75886 11688
rect 65944 11580 66668 11608
rect 65944 11568 65950 11580
rect 66898 11568 66904 11620
rect 66956 11568 66962 11620
rect 67082 11568 67088 11620
rect 67140 11608 67146 11620
rect 76116 11608 76144 11784
rect 76742 11744 76748 11756
rect 76703 11716 76748 11744
rect 76742 11704 76748 11716
rect 76800 11704 76806 11756
rect 76929 11747 76987 11753
rect 76929 11713 76941 11747
rect 76975 11744 76987 11747
rect 77110 11744 77116 11756
rect 76975 11716 77116 11744
rect 76975 11713 76987 11716
rect 76929 11707 76987 11713
rect 77110 11704 77116 11716
rect 77168 11704 77174 11756
rect 77220 11753 77248 11784
rect 79594 11772 79600 11784
rect 79652 11772 79658 11824
rect 80146 11812 80152 11824
rect 80107 11784 80152 11812
rect 80146 11772 80152 11784
rect 80204 11772 80210 11824
rect 80517 11815 80575 11821
rect 80517 11781 80529 11815
rect 80563 11812 80575 11815
rect 81250 11812 81256 11824
rect 80563 11784 81256 11812
rect 80563 11781 80575 11784
rect 80517 11775 80575 11781
rect 81250 11772 81256 11784
rect 81308 11772 81314 11824
rect 81820 11821 81848 11852
rect 84194 11840 84200 11852
rect 84252 11840 84258 11892
rect 84286 11840 84292 11892
rect 84344 11880 84350 11892
rect 85209 11883 85267 11889
rect 85209 11880 85221 11883
rect 84344 11852 85221 11880
rect 84344 11840 84350 11852
rect 85209 11849 85221 11852
rect 85255 11880 85267 11883
rect 85666 11880 85672 11892
rect 85255 11852 85672 11880
rect 85255 11849 85267 11852
rect 85209 11843 85267 11849
rect 85666 11840 85672 11852
rect 85724 11880 85730 11892
rect 86126 11880 86132 11892
rect 85724 11852 86132 11880
rect 85724 11840 85730 11852
rect 86126 11840 86132 11852
rect 86184 11840 86190 11892
rect 89162 11880 89168 11892
rect 86420 11852 89168 11880
rect 81805 11815 81863 11821
rect 81805 11781 81817 11815
rect 81851 11781 81863 11815
rect 81805 11775 81863 11781
rect 82354 11772 82360 11824
rect 82412 11772 82418 11824
rect 85942 11812 85948 11824
rect 84212 11784 85948 11812
rect 77205 11747 77263 11753
rect 77205 11713 77217 11747
rect 77251 11713 77263 11747
rect 77205 11707 77263 11713
rect 77389 11747 77447 11753
rect 77389 11713 77401 11747
rect 77435 11744 77447 11747
rect 77478 11744 77484 11756
rect 77435 11716 77484 11744
rect 77435 11713 77447 11716
rect 77389 11707 77447 11713
rect 77478 11704 77484 11716
rect 77536 11704 77542 11756
rect 77849 11747 77907 11753
rect 77849 11713 77861 11747
rect 77895 11744 77907 11747
rect 77938 11744 77944 11756
rect 77895 11716 77944 11744
rect 77895 11713 77907 11716
rect 77849 11707 77907 11713
rect 77938 11704 77944 11716
rect 77996 11704 78002 11756
rect 78033 11747 78091 11753
rect 78033 11713 78045 11747
rect 78079 11744 78091 11747
rect 79042 11744 79048 11756
rect 78079 11716 78168 11744
rect 79003 11716 79048 11744
rect 78079 11713 78091 11716
rect 78033 11707 78091 11713
rect 76190 11636 76196 11688
rect 76248 11676 76254 11688
rect 78140 11676 78168 11716
rect 79042 11704 79048 11716
rect 79100 11704 79106 11756
rect 79502 11704 79508 11756
rect 79560 11744 79566 11756
rect 80609 11747 80667 11753
rect 80609 11744 80621 11747
rect 79560 11716 80621 11744
rect 79560 11704 79566 11716
rect 80609 11713 80621 11716
rect 80655 11713 80667 11747
rect 80609 11707 80667 11713
rect 80238 11676 80244 11688
rect 76248 11648 80244 11676
rect 76248 11636 76254 11648
rect 80238 11636 80244 11648
rect 80296 11636 80302 11688
rect 67140 11580 73108 11608
rect 67140 11568 67146 11580
rect 60056 11512 60320 11540
rect 60056 11500 60062 11512
rect 60366 11500 60372 11552
rect 60424 11540 60430 11552
rect 60553 11543 60611 11549
rect 60553 11540 60565 11543
rect 60424 11512 60565 11540
rect 60424 11500 60430 11512
rect 60553 11509 60565 11512
rect 60599 11509 60611 11543
rect 60553 11503 60611 11509
rect 62574 11500 62580 11552
rect 62632 11540 62638 11552
rect 63586 11540 63592 11552
rect 62632 11512 63592 11540
rect 62632 11500 62638 11512
rect 63586 11500 63592 11512
rect 63644 11540 63650 11552
rect 66916 11540 66944 11568
rect 63644 11512 66944 11540
rect 63644 11500 63650 11512
rect 67266 11500 67272 11552
rect 67324 11540 67330 11552
rect 69474 11540 69480 11552
rect 67324 11512 69480 11540
rect 67324 11500 67330 11512
rect 69474 11500 69480 11512
rect 69532 11500 69538 11552
rect 69658 11540 69664 11552
rect 69619 11512 69664 11540
rect 69658 11500 69664 11512
rect 69716 11500 69722 11552
rect 71590 11500 71596 11552
rect 71648 11540 71654 11552
rect 72694 11540 72700 11552
rect 71648 11512 72700 11540
rect 71648 11500 71654 11512
rect 72694 11500 72700 11512
rect 72752 11500 72758 11552
rect 72878 11540 72884 11552
rect 72839 11512 72884 11540
rect 72878 11500 72884 11512
rect 72936 11500 72942 11552
rect 73080 11540 73108 11580
rect 75288 11580 76144 11608
rect 73982 11540 73988 11552
rect 73080 11512 73988 11540
rect 73982 11500 73988 11512
rect 74040 11540 74046 11552
rect 75288 11540 75316 11580
rect 76926 11568 76932 11620
rect 76984 11608 76990 11620
rect 77021 11611 77079 11617
rect 77021 11608 77033 11611
rect 76984 11580 77033 11608
rect 76984 11568 76990 11580
rect 77021 11577 77033 11580
rect 77067 11577 77079 11611
rect 77021 11571 77079 11577
rect 77113 11611 77171 11617
rect 77113 11577 77125 11611
rect 77159 11608 77171 11611
rect 78858 11608 78864 11620
rect 77159 11580 78864 11608
rect 77159 11577 77171 11580
rect 77113 11571 77171 11577
rect 78858 11568 78864 11580
rect 78916 11568 78922 11620
rect 76190 11540 76196 11552
rect 74040 11512 75316 11540
rect 76151 11512 76196 11540
rect 74040 11500 74046 11512
rect 76190 11500 76196 11512
rect 76248 11500 76254 11552
rect 77202 11500 77208 11552
rect 77260 11540 77266 11552
rect 78033 11543 78091 11549
rect 78033 11540 78045 11543
rect 77260 11512 78045 11540
rect 77260 11500 77266 11512
rect 78033 11509 78045 11512
rect 78079 11509 78091 11543
rect 80624 11540 80652 11707
rect 80698 11704 80704 11756
rect 80756 11744 80762 11756
rect 80756 11716 80801 11744
rect 80756 11704 80762 11716
rect 83734 11704 83740 11756
rect 83792 11744 83798 11756
rect 84212 11753 84240 11784
rect 85942 11772 85948 11784
rect 86000 11772 86006 11824
rect 84197 11747 84255 11753
rect 84197 11744 84209 11747
rect 83792 11716 84209 11744
rect 83792 11704 83798 11716
rect 84197 11713 84209 11716
rect 84243 11713 84255 11747
rect 84197 11707 84255 11713
rect 84378 11704 84384 11756
rect 84436 11744 84442 11756
rect 84933 11747 84991 11753
rect 84933 11744 84945 11747
rect 84436 11716 84945 11744
rect 84436 11704 84442 11716
rect 84933 11713 84945 11716
rect 84979 11744 84991 11747
rect 86420 11744 86448 11852
rect 89162 11840 89168 11852
rect 89220 11840 89226 11892
rect 94225 11883 94283 11889
rect 94225 11880 94237 11883
rect 90100 11852 94237 11880
rect 90100 11821 90128 11852
rect 94225 11849 94237 11852
rect 94271 11849 94283 11883
rect 94225 11843 94283 11849
rect 89073 11815 89131 11821
rect 89073 11812 89085 11815
rect 87262 11784 89085 11812
rect 89073 11781 89085 11784
rect 89119 11781 89131 11815
rect 89073 11775 89131 11781
rect 90085 11815 90143 11821
rect 90085 11781 90097 11815
rect 90131 11781 90143 11815
rect 90085 11775 90143 11781
rect 90542 11772 90548 11824
rect 90600 11772 90606 11824
rect 89162 11744 89168 11756
rect 84979 11716 86448 11744
rect 89123 11716 89168 11744
rect 84979 11713 84991 11716
rect 84933 11707 84991 11713
rect 89162 11704 89168 11716
rect 89220 11704 89226 11756
rect 92106 11744 92112 11756
rect 92067 11716 92112 11744
rect 92106 11704 92112 11716
rect 92164 11704 92170 11756
rect 92290 11744 92296 11756
rect 92251 11716 92296 11744
rect 92290 11704 92296 11716
rect 92348 11704 92354 11756
rect 93302 11704 93308 11756
rect 93360 11744 93366 11756
rect 94133 11747 94191 11753
rect 94133 11744 94145 11747
rect 93360 11716 94145 11744
rect 93360 11704 93366 11716
rect 94133 11713 94145 11716
rect 94179 11713 94191 11747
rect 94133 11707 94191 11713
rect 80885 11679 80943 11685
rect 80885 11645 80897 11679
rect 80931 11676 80943 11679
rect 81529 11679 81587 11685
rect 81529 11676 81541 11679
rect 80931 11648 81541 11676
rect 80931 11645 80943 11648
rect 80885 11639 80943 11645
rect 81529 11645 81541 11648
rect 81575 11676 81587 11679
rect 81575 11648 82860 11676
rect 81575 11645 81587 11648
rect 81529 11639 81587 11645
rect 82832 11608 82860 11648
rect 82998 11636 83004 11688
rect 83056 11676 83062 11688
rect 83550 11676 83556 11688
rect 83056 11648 83556 11676
rect 83056 11636 83062 11648
rect 83550 11636 83556 11648
rect 83608 11636 83614 11688
rect 83826 11676 83832 11688
rect 83787 11648 83832 11676
rect 83826 11636 83832 11648
rect 83884 11636 83890 11688
rect 84286 11676 84292 11688
rect 84199 11648 84292 11676
rect 84286 11636 84292 11648
rect 84344 11676 84350 11688
rect 86954 11676 86960 11688
rect 84344 11648 86960 11676
rect 84344 11636 84350 11648
rect 86954 11636 86960 11648
rect 87012 11636 87018 11688
rect 87690 11676 87696 11688
rect 87651 11648 87696 11676
rect 87690 11636 87696 11648
rect 87748 11636 87754 11688
rect 87966 11676 87972 11688
rect 87879 11648 87972 11676
rect 87966 11636 87972 11648
rect 88024 11636 88030 11688
rect 88978 11636 88984 11688
rect 89036 11676 89042 11688
rect 89809 11679 89867 11685
rect 89809 11676 89821 11679
rect 89036 11648 89821 11676
rect 89036 11636 89042 11648
rect 89809 11645 89821 11648
rect 89855 11645 89867 11679
rect 89809 11639 89867 11645
rect 91557 11679 91615 11685
rect 91557 11645 91569 11679
rect 91603 11676 91615 11679
rect 92474 11676 92480 11688
rect 91603 11648 92480 11676
rect 91603 11645 91615 11648
rect 91557 11639 91615 11645
rect 92474 11636 92480 11648
rect 92532 11636 92538 11688
rect 93121 11679 93179 11685
rect 93121 11645 93133 11679
rect 93167 11676 93179 11679
rect 93394 11676 93400 11688
rect 93167 11648 93400 11676
rect 93167 11645 93179 11648
rect 93121 11639 93179 11645
rect 93394 11636 93400 11648
rect 93452 11636 93458 11688
rect 84654 11608 84660 11620
rect 82832 11580 84660 11608
rect 84654 11568 84660 11580
rect 84712 11568 84718 11620
rect 84746 11568 84752 11620
rect 84804 11608 84810 11620
rect 87984 11608 88012 11636
rect 89714 11608 89720 11620
rect 84804 11580 86356 11608
rect 87984 11580 89720 11608
rect 84804 11568 84810 11580
rect 82998 11540 83004 11552
rect 80624 11512 83004 11540
rect 78033 11503 78091 11509
rect 82998 11500 83004 11512
rect 83056 11500 83062 11552
rect 83277 11543 83335 11549
rect 83277 11509 83289 11543
rect 83323 11540 83335 11543
rect 86034 11540 86040 11552
rect 83323 11512 86040 11540
rect 83323 11509 83335 11512
rect 83277 11503 83335 11509
rect 86034 11500 86040 11512
rect 86092 11500 86098 11552
rect 86218 11540 86224 11552
rect 86179 11512 86224 11540
rect 86218 11500 86224 11512
rect 86276 11500 86282 11552
rect 86328 11540 86356 11580
rect 89714 11568 89720 11580
rect 89772 11568 89778 11620
rect 91094 11540 91100 11552
rect 86328 11512 91100 11540
rect 91094 11500 91100 11512
rect 91152 11500 91158 11552
rect 1104 11450 94852 11472
rect 1104 11398 12668 11450
rect 12720 11398 12732 11450
rect 12784 11398 12796 11450
rect 12848 11398 12860 11450
rect 12912 11398 12924 11450
rect 12976 11398 36105 11450
rect 36157 11398 36169 11450
rect 36221 11398 36233 11450
rect 36285 11398 36297 11450
rect 36349 11398 36361 11450
rect 36413 11398 59542 11450
rect 59594 11398 59606 11450
rect 59658 11398 59670 11450
rect 59722 11398 59734 11450
rect 59786 11398 59798 11450
rect 59850 11398 82979 11450
rect 83031 11398 83043 11450
rect 83095 11398 83107 11450
rect 83159 11398 83171 11450
rect 83223 11398 83235 11450
rect 83287 11398 94852 11450
rect 1104 11376 94852 11398
rect 1762 11336 1768 11348
rect 1675 11308 1768 11336
rect 1762 11296 1768 11308
rect 1820 11336 1826 11348
rect 2498 11336 2504 11348
rect 1820 11308 2504 11336
rect 1820 11296 1826 11308
rect 2498 11296 2504 11308
rect 2556 11336 2562 11348
rect 2556 11308 4844 11336
rect 2556 11296 2562 11308
rect 4816 11268 4844 11308
rect 5074 11296 5080 11348
rect 5132 11336 5138 11348
rect 5132 11308 5580 11336
rect 5132 11296 5138 11308
rect 5442 11268 5448 11280
rect 4816 11240 5448 11268
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11132 2283 11135
rect 2498 11132 2504 11144
rect 2271 11104 2360 11132
rect 2459 11104 2504 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 2332 11076 2360 11104
rect 2498 11092 2504 11104
rect 2556 11092 2562 11144
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11132 3295 11135
rect 3878 11132 3884 11144
rect 3283 11104 3884 11132
rect 3283 11101 3295 11104
rect 3237 11095 3295 11101
rect 3878 11092 3884 11104
rect 3936 11092 3942 11144
rect 3973 11135 4031 11141
rect 3973 11101 3985 11135
rect 4019 11132 4031 11135
rect 4249 11135 4307 11141
rect 4019 11104 4108 11132
rect 4019 11101 4031 11104
rect 3973 11095 4031 11101
rect 2314 11024 2320 11076
rect 2372 11024 2378 11076
rect 3418 10996 3424 11008
rect 3379 10968 3424 10996
rect 3418 10956 3424 10968
rect 3476 10956 3482 11008
rect 4080 10996 4108 11104
rect 4249 11101 4261 11135
rect 4295 11132 4307 11135
rect 4816 11132 4844 11240
rect 5442 11228 5448 11240
rect 5500 11228 5506 11280
rect 5552 11268 5580 11308
rect 6914 11296 6920 11348
rect 6972 11336 6978 11348
rect 7374 11336 7380 11348
rect 6972 11308 7380 11336
rect 6972 11296 6978 11308
rect 7374 11296 7380 11308
rect 7432 11336 7438 11348
rect 9125 11339 9183 11345
rect 9125 11336 9137 11339
rect 7432 11308 9137 11336
rect 7432 11296 7438 11308
rect 9125 11305 9137 11308
rect 9171 11305 9183 11339
rect 9125 11299 9183 11305
rect 9490 11296 9496 11348
rect 9548 11336 9554 11348
rect 9585 11339 9643 11345
rect 9585 11336 9597 11339
rect 9548 11308 9597 11336
rect 9548 11296 9554 11308
rect 9585 11305 9597 11308
rect 9631 11336 9643 11339
rect 11241 11339 11299 11345
rect 11241 11336 11253 11339
rect 9631 11308 11253 11336
rect 9631 11305 9643 11308
rect 9585 11299 9643 11305
rect 11241 11305 11253 11308
rect 11287 11305 11299 11339
rect 11241 11299 11299 11305
rect 11882 11296 11888 11348
rect 11940 11336 11946 11348
rect 11977 11339 12035 11345
rect 11977 11336 11989 11339
rect 11940 11308 11989 11336
rect 11940 11296 11946 11308
rect 11977 11305 11989 11308
rect 12023 11336 12035 11339
rect 12023 11308 13400 11336
rect 12023 11305 12035 11308
rect 11977 11299 12035 11305
rect 12526 11268 12532 11280
rect 5552 11240 8616 11268
rect 5169 11203 5227 11209
rect 5169 11169 5181 11203
rect 5215 11200 5227 11203
rect 6914 11200 6920 11212
rect 5215 11172 6920 11200
rect 5215 11169 5227 11172
rect 5169 11163 5227 11169
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 7561 11203 7619 11209
rect 7561 11169 7573 11203
rect 7607 11200 7619 11203
rect 8478 11200 8484 11212
rect 7607 11172 8484 11200
rect 7607 11169 7619 11172
rect 7561 11163 7619 11169
rect 8478 11160 8484 11172
rect 8536 11160 8542 11212
rect 4295 11104 4844 11132
rect 4893 11135 4951 11141
rect 4295 11101 4307 11104
rect 4249 11095 4307 11101
rect 4893 11101 4905 11135
rect 4939 11101 4951 11135
rect 4893 11095 4951 11101
rect 4908 11064 4936 11095
rect 4982 11092 4988 11144
rect 5040 11132 5046 11144
rect 6365 11135 6423 11141
rect 6365 11132 6377 11135
rect 5040 11104 6377 11132
rect 5040 11092 5046 11104
rect 6365 11101 6377 11104
rect 6411 11101 6423 11135
rect 6365 11095 6423 11101
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11101 8447 11135
rect 8588 11132 8616 11240
rect 10704 11240 12532 11268
rect 9401 11203 9459 11209
rect 9401 11169 9413 11203
rect 9447 11200 9459 11203
rect 9766 11200 9772 11212
rect 9447 11172 9772 11200
rect 9447 11169 9459 11172
rect 9401 11163 9459 11169
rect 9766 11160 9772 11172
rect 9824 11200 9830 11212
rect 10704 11209 10732 11240
rect 12526 11228 12532 11240
rect 12584 11228 12590 11280
rect 13372 11268 13400 11308
rect 13446 11296 13452 11348
rect 13504 11336 13510 11348
rect 13541 11339 13599 11345
rect 13541 11336 13553 11339
rect 13504 11308 13553 11336
rect 13504 11296 13510 11308
rect 13541 11305 13553 11308
rect 13587 11305 13599 11339
rect 13541 11299 13599 11305
rect 14826 11296 14832 11348
rect 14884 11336 14890 11348
rect 20162 11336 20168 11348
rect 14884 11308 20168 11336
rect 14884 11296 14890 11308
rect 20162 11296 20168 11308
rect 20220 11296 20226 11348
rect 20257 11339 20315 11345
rect 20257 11305 20269 11339
rect 20303 11336 20315 11339
rect 20530 11336 20536 11348
rect 20303 11308 20536 11336
rect 20303 11305 20315 11308
rect 20257 11299 20315 11305
rect 20530 11296 20536 11308
rect 20588 11296 20594 11348
rect 27614 11296 27620 11348
rect 27672 11336 27678 11348
rect 27709 11339 27767 11345
rect 27709 11336 27721 11339
rect 27672 11308 27721 11336
rect 27672 11296 27678 11308
rect 27709 11305 27721 11308
rect 27755 11305 27767 11339
rect 27709 11299 27767 11305
rect 28350 11296 28356 11348
rect 28408 11336 28414 11348
rect 28537 11339 28595 11345
rect 28537 11336 28549 11339
rect 28408 11308 28549 11336
rect 28408 11296 28414 11308
rect 28537 11305 28549 11308
rect 28583 11305 28595 11339
rect 30006 11336 30012 11348
rect 29967 11308 30012 11336
rect 28537 11299 28595 11305
rect 30006 11296 30012 11308
rect 30064 11296 30070 11348
rect 31478 11336 31484 11348
rect 31439 11308 31484 11336
rect 31478 11296 31484 11308
rect 31536 11296 31542 11348
rect 34514 11296 34520 11348
rect 34572 11336 34578 11348
rect 37090 11336 37096 11348
rect 34572 11308 37096 11336
rect 34572 11296 34578 11308
rect 37090 11296 37096 11308
rect 37148 11296 37154 11348
rect 37182 11296 37188 11348
rect 37240 11336 37246 11348
rect 39114 11336 39120 11348
rect 37240 11308 39120 11336
rect 37240 11296 37246 11308
rect 39114 11296 39120 11308
rect 39172 11336 39178 11348
rect 39485 11339 39543 11345
rect 39485 11336 39497 11339
rect 39172 11308 39497 11336
rect 39172 11296 39178 11308
rect 39485 11305 39497 11308
rect 39531 11336 39543 11339
rect 41690 11336 41696 11348
rect 39531 11308 41696 11336
rect 39531 11305 39543 11308
rect 39485 11299 39543 11305
rect 41690 11296 41696 11308
rect 41748 11296 41754 11348
rect 41966 11336 41972 11348
rect 41927 11308 41972 11336
rect 41966 11296 41972 11308
rect 42024 11296 42030 11348
rect 42886 11296 42892 11348
rect 42944 11336 42950 11348
rect 43073 11339 43131 11345
rect 43073 11336 43085 11339
rect 42944 11308 43085 11336
rect 42944 11296 42950 11308
rect 43073 11305 43085 11308
rect 43119 11336 43131 11339
rect 43898 11336 43904 11348
rect 43119 11308 43904 11336
rect 43119 11305 43131 11308
rect 43073 11299 43131 11305
rect 43898 11296 43904 11308
rect 43956 11296 43962 11348
rect 45462 11296 45468 11348
rect 45520 11336 45526 11348
rect 51810 11336 51816 11348
rect 45520 11308 51816 11336
rect 45520 11296 45526 11308
rect 51810 11296 51816 11308
rect 51868 11296 51874 11348
rect 51994 11296 52000 11348
rect 52052 11336 52058 11348
rect 54481 11339 54539 11345
rect 54481 11336 54493 11339
rect 52052 11308 54493 11336
rect 52052 11296 52058 11308
rect 54481 11305 54493 11308
rect 54527 11305 54539 11339
rect 54481 11299 54539 11305
rect 56321 11339 56379 11345
rect 56321 11305 56333 11339
rect 56367 11336 56379 11339
rect 57330 11336 57336 11348
rect 56367 11308 57336 11336
rect 56367 11305 56379 11308
rect 56321 11299 56379 11305
rect 14090 11268 14096 11280
rect 13372 11240 14096 11268
rect 14090 11228 14096 11240
rect 14148 11228 14154 11280
rect 14366 11228 14372 11280
rect 14424 11268 14430 11280
rect 19334 11268 19340 11280
rect 14424 11240 19340 11268
rect 14424 11228 14430 11240
rect 19334 11228 19340 11240
rect 19392 11228 19398 11280
rect 19426 11228 19432 11280
rect 19484 11228 19490 11280
rect 19521 11271 19579 11277
rect 19521 11237 19533 11271
rect 19567 11237 19579 11271
rect 25866 11268 25872 11280
rect 19521 11231 19579 11237
rect 23032 11240 25872 11268
rect 10689 11203 10747 11209
rect 10689 11200 10701 11203
rect 9824 11172 10701 11200
rect 9824 11160 9830 11172
rect 10689 11169 10701 11172
rect 10735 11169 10747 11203
rect 10689 11163 10747 11169
rect 12250 11160 12256 11212
rect 12308 11200 12314 11212
rect 13173 11203 13231 11209
rect 13173 11200 13185 11203
rect 12308 11172 13185 11200
rect 12308 11160 12314 11172
rect 13173 11169 13185 11172
rect 13219 11169 13231 11203
rect 13173 11163 13231 11169
rect 13354 11160 13360 11212
rect 13412 11200 13418 11212
rect 15930 11200 15936 11212
rect 13412 11172 15936 11200
rect 13412 11160 13418 11172
rect 15930 11160 15936 11172
rect 15988 11160 15994 11212
rect 19444 11200 19472 11228
rect 18800 11172 19472 11200
rect 19536 11200 19564 11231
rect 20806 11200 20812 11212
rect 19536 11172 20812 11200
rect 9677 11135 9735 11141
rect 9677 11132 9689 11135
rect 8588 11104 9689 11132
rect 8389 11095 8447 11101
rect 9677 11101 9689 11104
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 5994 11064 6000 11076
rect 4908 11036 6000 11064
rect 5994 11024 6000 11036
rect 6052 11024 6058 11076
rect 6917 11067 6975 11073
rect 6917 11064 6929 11067
rect 6104 11036 6929 11064
rect 4614 10996 4620 11008
rect 4080 10968 4620 10996
rect 4614 10956 4620 10968
rect 4672 10956 4678 11008
rect 5813 10999 5871 11005
rect 5813 10965 5825 10999
rect 5859 10996 5871 10999
rect 6104 10996 6132 11036
rect 6917 11033 6929 11036
rect 6963 11064 6975 11067
rect 7282 11064 7288 11076
rect 6963 11036 7288 11064
rect 6963 11033 6975 11036
rect 6917 11027 6975 11033
rect 7282 11024 7288 11036
rect 7340 11064 7346 11076
rect 8404 11064 8432 11095
rect 8478 11064 8484 11076
rect 7340 11036 8484 11064
rect 7340 11024 7346 11036
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 9692 11064 9720 11095
rect 11790 11092 11796 11144
rect 11848 11132 11854 11144
rect 13265 11135 13323 11141
rect 13265 11132 13277 11135
rect 11848 11104 13277 11132
rect 11848 11092 11854 11104
rect 13265 11101 13277 11104
rect 13311 11101 13323 11135
rect 15194 11132 15200 11144
rect 13265 11095 13323 11101
rect 14476 11104 15200 11132
rect 10229 11067 10287 11073
rect 10229 11064 10241 11067
rect 9692 11036 10241 11064
rect 10229 11033 10241 11036
rect 10275 11064 10287 11067
rect 10275 11036 12434 11064
rect 10275 11033 10287 11036
rect 10229 11027 10287 11033
rect 8018 10996 8024 11008
rect 5859 10968 6132 10996
rect 7979 10968 8024 10996
rect 5859 10965 5871 10968
rect 5813 10959 5871 10965
rect 8018 10956 8024 10968
rect 8076 10956 8082 11008
rect 12406 10996 12434 11036
rect 12526 11024 12532 11076
rect 12584 11064 12590 11076
rect 12621 11067 12679 11073
rect 12621 11064 12633 11067
rect 12584 11036 12633 11064
rect 12584 11024 12590 11036
rect 12621 11033 12633 11036
rect 12667 11064 12679 11067
rect 14476 11064 14504 11104
rect 15194 11092 15200 11104
rect 15252 11092 15258 11144
rect 15381 11135 15439 11141
rect 15381 11101 15393 11135
rect 15427 11132 15439 11135
rect 15470 11132 15476 11144
rect 15427 11104 15476 11132
rect 15427 11101 15439 11104
rect 15381 11095 15439 11101
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 15562 11092 15568 11144
rect 15620 11132 15626 11144
rect 16577 11135 16635 11141
rect 16577 11132 16589 11135
rect 15620 11104 16589 11132
rect 15620 11092 15626 11104
rect 16577 11101 16589 11104
rect 16623 11101 16635 11135
rect 17126 11132 17132 11144
rect 17087 11104 17132 11132
rect 16577 11095 16635 11101
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 18322 11132 18328 11144
rect 17512 11104 18328 11132
rect 12667 11036 14504 11064
rect 14553 11067 14611 11073
rect 12667 11033 12679 11036
rect 12621 11027 12679 11033
rect 14553 11033 14565 11067
rect 14599 11064 14611 11067
rect 16482 11064 16488 11076
rect 14599 11036 16488 11064
rect 14599 11033 14611 11036
rect 14553 11027 14611 11033
rect 16482 11024 16488 11036
rect 16540 11024 16546 11076
rect 17512 11050 17540 11104
rect 18322 11092 18328 11104
rect 18380 11092 18386 11144
rect 18414 11092 18420 11144
rect 18472 11132 18478 11144
rect 18800 11141 18828 11172
rect 20806 11160 20812 11172
rect 20864 11160 20870 11212
rect 21637 11203 21695 11209
rect 21637 11169 21649 11203
rect 21683 11200 21695 11203
rect 23032 11200 23060 11240
rect 25866 11228 25872 11240
rect 25924 11228 25930 11280
rect 28810 11228 28816 11280
rect 28868 11268 28874 11280
rect 30466 11268 30472 11280
rect 28868 11240 30472 11268
rect 28868 11228 28874 11240
rect 30466 11228 30472 11240
rect 30524 11228 30530 11280
rect 30653 11271 30711 11277
rect 30653 11237 30665 11271
rect 30699 11268 30711 11271
rect 31294 11268 31300 11280
rect 30699 11240 31300 11268
rect 30699 11237 30711 11240
rect 30653 11231 30711 11237
rect 31294 11228 31300 11240
rect 31352 11268 31358 11280
rect 32490 11268 32496 11280
rect 31352 11240 32496 11268
rect 31352 11228 31358 11240
rect 32490 11228 32496 11240
rect 32548 11228 32554 11280
rect 33796 11240 41460 11268
rect 21683 11172 23060 11200
rect 23109 11203 23167 11209
rect 21683 11169 21695 11172
rect 21637 11163 21695 11169
rect 23109 11169 23121 11203
rect 23155 11200 23167 11203
rect 26237 11203 26295 11209
rect 26237 11200 26249 11203
rect 23155 11172 24992 11200
rect 23155 11169 23167 11172
rect 23109 11163 23167 11169
rect 18785 11135 18843 11141
rect 18785 11132 18797 11135
rect 18472 11104 18797 11132
rect 18472 11092 18478 11104
rect 18785 11101 18797 11104
rect 18831 11101 18843 11135
rect 19334 11132 19340 11144
rect 18785 11095 18843 11101
rect 19306 11092 19340 11132
rect 19392 11092 19398 11144
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11101 19487 11135
rect 19429 11095 19487 11101
rect 17862 11024 17868 11076
rect 17920 11064 17926 11076
rect 19306 11064 19334 11092
rect 17920 11036 19334 11064
rect 17920 11024 17926 11036
rect 19444 11008 19472 11095
rect 19610 11092 19616 11144
rect 19668 11132 19674 11144
rect 19668 11104 19713 11132
rect 19668 11092 19674 11104
rect 19978 11092 19984 11144
rect 20036 11132 20042 11144
rect 20073 11135 20131 11141
rect 20073 11132 20085 11135
rect 20036 11104 20085 11132
rect 20036 11092 20042 11104
rect 20073 11101 20085 11104
rect 20119 11132 20131 11135
rect 21361 11135 21419 11141
rect 21361 11132 21373 11135
rect 20119 11104 21373 11132
rect 20119 11101 20131 11104
rect 20073 11095 20131 11101
rect 21361 11101 21373 11104
rect 21407 11101 21419 11135
rect 21361 11095 21419 11101
rect 22738 11092 22744 11144
rect 22796 11092 22802 11144
rect 24964 11141 24992 11172
rect 25056 11172 26249 11200
rect 24949 11135 25007 11141
rect 24949 11101 24961 11135
rect 24995 11101 25007 11135
rect 24949 11095 25007 11101
rect 22922 11024 22928 11076
rect 22980 11064 22986 11076
rect 25056 11064 25084 11172
rect 26237 11169 26249 11172
rect 26283 11169 26295 11203
rect 26237 11163 26295 11169
rect 27430 11160 27436 11212
rect 27488 11200 27494 11212
rect 29362 11200 29368 11212
rect 27488 11172 29368 11200
rect 27488 11160 27494 11172
rect 29362 11160 29368 11172
rect 29420 11160 29426 11212
rect 33796 11200 33824 11240
rect 32324 11172 33824 11200
rect 34241 11203 34299 11209
rect 25866 11092 25872 11144
rect 25924 11132 25930 11144
rect 25961 11135 26019 11141
rect 25961 11132 25973 11135
rect 25924 11104 25973 11132
rect 25924 11092 25930 11104
rect 25961 11101 25973 11104
rect 26007 11101 26019 11135
rect 25961 11095 26019 11101
rect 27522 11092 27528 11144
rect 27580 11132 27586 11144
rect 29454 11132 29460 11144
rect 27580 11104 29460 11132
rect 27580 11092 27586 11104
rect 29454 11092 29460 11104
rect 29512 11132 29518 11144
rect 32324 11132 32352 11172
rect 34241 11169 34253 11203
rect 34287 11200 34299 11203
rect 36538 11200 36544 11212
rect 34287 11172 36544 11200
rect 34287 11169 34299 11172
rect 34241 11163 34299 11169
rect 36538 11160 36544 11172
rect 36596 11160 36602 11212
rect 36814 11160 36820 11212
rect 36872 11200 36878 11212
rect 37550 11200 37556 11212
rect 36872 11172 37556 11200
rect 36872 11160 36878 11172
rect 37550 11160 37556 11172
rect 37608 11160 37614 11212
rect 38010 11200 38016 11212
rect 37971 11172 38016 11200
rect 38010 11160 38016 11172
rect 38068 11160 38074 11212
rect 38286 11160 38292 11212
rect 38344 11200 38350 11212
rect 38344 11172 38389 11200
rect 38344 11160 38350 11172
rect 38654 11160 38660 11212
rect 38712 11200 38718 11212
rect 41432 11200 41460 11240
rect 44450 11228 44456 11280
rect 44508 11268 44514 11280
rect 52362 11268 52368 11280
rect 44508 11240 52368 11268
rect 44508 11228 44514 11240
rect 52362 11228 52368 11240
rect 52420 11228 52426 11280
rect 53466 11228 53472 11280
rect 53524 11268 53530 11280
rect 53650 11268 53656 11280
rect 53524 11240 53656 11268
rect 53524 11228 53530 11240
rect 53650 11228 53656 11240
rect 53708 11228 53714 11280
rect 38712 11172 40172 11200
rect 41432 11172 43944 11200
rect 38712 11160 38718 11172
rect 32490 11132 32496 11144
rect 29512 11104 32352 11132
rect 32451 11104 32496 11132
rect 29512 11092 29518 11104
rect 32490 11092 32496 11104
rect 32548 11092 32554 11144
rect 35250 11092 35256 11144
rect 35308 11132 35314 11144
rect 35345 11135 35403 11141
rect 35345 11132 35357 11135
rect 35308 11104 35357 11132
rect 35308 11092 35314 11104
rect 35345 11101 35357 11104
rect 35391 11101 35403 11135
rect 35345 11095 35403 11101
rect 38381 11135 38439 11141
rect 38381 11101 38393 11135
rect 38427 11132 38439 11135
rect 38838 11132 38844 11144
rect 38427 11104 38844 11132
rect 38427 11101 38439 11104
rect 38381 11095 38439 11101
rect 38838 11092 38844 11104
rect 38896 11132 38902 11144
rect 39758 11132 39764 11144
rect 38896 11104 39764 11132
rect 38896 11092 38902 11104
rect 39758 11092 39764 11104
rect 39816 11092 39822 11144
rect 40144 11132 40172 11172
rect 40494 11132 40500 11144
rect 40144 11104 40500 11132
rect 40494 11092 40500 11104
rect 40552 11092 40558 11144
rect 41417 11135 41475 11141
rect 41417 11101 41429 11135
rect 41463 11132 41475 11135
rect 41782 11132 41788 11144
rect 41463 11104 41788 11132
rect 41463 11101 41475 11104
rect 41417 11095 41475 11101
rect 41782 11092 41788 11104
rect 41840 11092 41846 11144
rect 42150 11092 42156 11144
rect 42208 11132 42214 11144
rect 42429 11135 42487 11141
rect 42429 11132 42441 11135
rect 42208 11104 42441 11132
rect 42208 11092 42214 11104
rect 42429 11101 42441 11104
rect 42475 11132 42487 11135
rect 43806 11132 43812 11144
rect 42475 11104 43812 11132
rect 42475 11101 42487 11104
rect 42429 11095 42487 11101
rect 43806 11092 43812 11104
rect 43864 11092 43870 11144
rect 43916 11132 43944 11172
rect 43990 11160 43996 11212
rect 44048 11200 44054 11212
rect 44634 11200 44640 11212
rect 44048 11172 44093 11200
rect 44595 11172 44640 11200
rect 44048 11160 44054 11172
rect 44634 11160 44640 11172
rect 44692 11160 44698 11212
rect 48958 11200 48964 11212
rect 48919 11172 48964 11200
rect 48958 11160 48964 11172
rect 49016 11160 49022 11212
rect 50430 11200 50436 11212
rect 49436 11172 50436 11200
rect 45557 11135 45615 11141
rect 45557 11132 45569 11135
rect 43916 11104 45569 11132
rect 45557 11101 45569 11104
rect 45603 11132 45615 11135
rect 45738 11132 45744 11144
rect 45603 11104 45744 11132
rect 45603 11101 45615 11104
rect 45557 11095 45615 11101
rect 45738 11092 45744 11104
rect 45796 11092 45802 11144
rect 46750 11132 46756 11144
rect 46711 11104 46756 11132
rect 46750 11092 46756 11104
rect 46808 11092 46814 11144
rect 47489 11135 47547 11141
rect 47489 11132 47501 11135
rect 46860 11104 47501 11132
rect 22980 11036 25084 11064
rect 25225 11067 25283 11073
rect 22980 11024 22986 11036
rect 25225 11033 25237 11067
rect 25271 11064 25283 11067
rect 25271 11036 26648 11064
rect 25271 11033 25283 11036
rect 25225 11027 25283 11033
rect 13630 10996 13636 11008
rect 12406 10968 13636 10996
rect 13630 10956 13636 10968
rect 13688 10956 13694 11008
rect 15010 10956 15016 11008
rect 15068 10996 15074 11008
rect 15289 10999 15347 11005
rect 15289 10996 15301 10999
rect 15068 10968 15301 10996
rect 15068 10956 15074 10968
rect 15289 10965 15301 10968
rect 15335 10996 15347 10999
rect 19058 10996 19064 11008
rect 15335 10968 19064 10996
rect 15335 10965 15347 10968
rect 15289 10959 15347 10965
rect 19058 10956 19064 10968
rect 19116 10996 19122 11008
rect 19288 10996 19294 11008
rect 19116 10968 19294 10996
rect 19116 10956 19122 10968
rect 19288 10956 19294 10968
rect 19346 10956 19352 11008
rect 19426 10956 19432 11008
rect 19484 10956 19490 11008
rect 19794 10956 19800 11008
rect 19852 10996 19858 11008
rect 20809 10999 20867 11005
rect 20809 10996 20821 10999
rect 19852 10968 20821 10996
rect 19852 10956 19858 10968
rect 20809 10965 20821 10968
rect 20855 10965 20867 10999
rect 20809 10959 20867 10965
rect 20990 10956 20996 11008
rect 21048 10996 21054 11008
rect 23934 10996 23940 11008
rect 21048 10968 23940 10996
rect 21048 10956 21054 10968
rect 23934 10956 23940 10968
rect 23992 10956 23998 11008
rect 24029 10999 24087 11005
rect 24029 10965 24041 10999
rect 24075 10996 24087 10999
rect 24762 10996 24768 11008
rect 24075 10968 24768 10996
rect 24075 10965 24087 10968
rect 24029 10959 24087 10965
rect 24762 10956 24768 10968
rect 24820 10996 24826 11008
rect 26234 10996 26240 11008
rect 24820 10968 26240 10996
rect 24820 10956 24826 10968
rect 26234 10956 26240 10968
rect 26292 10956 26298 11008
rect 26620 10996 26648 11036
rect 26694 11024 26700 11076
rect 26752 11024 26758 11076
rect 29086 11064 29092 11076
rect 27540 11036 29092 11064
rect 27540 10996 27568 11036
rect 29086 11024 29092 11036
rect 29144 11064 29150 11076
rect 30282 11064 30288 11076
rect 29144 11036 30288 11064
rect 29144 11024 29150 11036
rect 30282 11024 30288 11036
rect 30340 11024 30346 11076
rect 30374 11024 30380 11076
rect 30432 11064 30438 11076
rect 31205 11067 31263 11073
rect 31205 11064 31217 11067
rect 30432 11036 31217 11064
rect 30432 11024 30438 11036
rect 31205 11033 31217 11036
rect 31251 11033 31263 11067
rect 31205 11027 31263 11033
rect 32769 11067 32827 11073
rect 32769 11033 32781 11067
rect 32815 11064 32827 11067
rect 33042 11064 33048 11076
rect 32815 11036 33048 11064
rect 32815 11033 32827 11036
rect 32769 11027 32827 11033
rect 33042 11024 33048 11036
rect 33100 11024 33106 11076
rect 34330 11064 34336 11076
rect 33994 11036 34336 11064
rect 34330 11024 34336 11036
rect 34388 11024 34394 11076
rect 34790 11024 34796 11076
rect 34848 11064 34854 11076
rect 35529 11067 35587 11073
rect 35529 11064 35541 11067
rect 34848 11036 35541 11064
rect 34848 11024 34854 11036
rect 35529 11033 35541 11036
rect 35575 11033 35587 11067
rect 35529 11027 35587 11033
rect 35618 11024 35624 11076
rect 35676 11064 35682 11076
rect 37185 11067 37243 11073
rect 37185 11064 37197 11067
rect 35676 11036 37197 11064
rect 35676 11024 35682 11036
rect 37185 11033 37197 11036
rect 37231 11064 37243 11067
rect 38194 11064 38200 11076
rect 37231 11036 38200 11064
rect 37231 11033 37243 11036
rect 37185 11027 37243 11033
rect 38194 11024 38200 11036
rect 38252 11024 38258 11076
rect 41966 11064 41972 11076
rect 38396 11036 41972 11064
rect 38396 11008 38424 11036
rect 41966 11024 41972 11036
rect 42024 11024 42030 11076
rect 42794 11064 42800 11076
rect 42076 11036 42800 11064
rect 26620 10968 27568 10996
rect 28994 10956 29000 11008
rect 29052 10996 29058 11008
rect 29181 10999 29239 11005
rect 29181 10996 29193 10999
rect 29052 10968 29193 10996
rect 29052 10956 29058 10968
rect 29181 10965 29193 10968
rect 29227 10965 29239 10999
rect 29181 10959 29239 10965
rect 30006 10956 30012 11008
rect 30064 10996 30070 11008
rect 31754 10996 31760 11008
rect 30064 10968 31760 10996
rect 30064 10956 30070 10968
rect 31754 10956 31760 10968
rect 31812 10956 31818 11008
rect 31846 10956 31852 11008
rect 31904 10996 31910 11008
rect 37366 10996 37372 11008
rect 31904 10968 37372 10996
rect 31904 10956 31910 10968
rect 37366 10956 37372 10968
rect 37424 10956 37430 11008
rect 37458 10956 37464 11008
rect 37516 10996 37522 11008
rect 38286 10996 38292 11008
rect 37516 10968 38292 10996
rect 37516 10956 37522 10968
rect 38286 10956 38292 10968
rect 38344 10956 38350 11008
rect 38378 10956 38384 11008
rect 38436 10956 38442 11008
rect 39758 10956 39764 11008
rect 39816 10996 39822 11008
rect 42076 10996 42104 11036
rect 42794 11024 42800 11036
rect 42852 11064 42858 11076
rect 46860 11064 46888 11104
rect 47489 11101 47501 11104
rect 47535 11132 47547 11135
rect 48774 11132 48780 11144
rect 47535 11104 48780 11132
rect 47535 11101 47547 11104
rect 47489 11095 47547 11101
rect 48774 11092 48780 11104
rect 48832 11092 48838 11144
rect 49436 11141 49464 11172
rect 50430 11160 50436 11172
rect 50488 11160 50494 11212
rect 51902 11160 51908 11212
rect 51960 11200 51966 11212
rect 51960 11172 52132 11200
rect 51960 11160 51966 11172
rect 49421 11135 49479 11141
rect 49421 11101 49433 11135
rect 49467 11101 49479 11135
rect 49602 11132 49608 11144
rect 49563 11104 49608 11132
rect 49421 11095 49479 11101
rect 49602 11092 49608 11104
rect 49660 11092 49666 11144
rect 49694 11092 49700 11144
rect 49752 11132 49758 11144
rect 49752 11104 49797 11132
rect 49752 11092 49758 11104
rect 50062 11092 50068 11144
rect 50120 11132 50126 11144
rect 50341 11135 50399 11141
rect 50341 11132 50353 11135
rect 50120 11104 50353 11132
rect 50120 11092 50126 11104
rect 50341 11101 50353 11104
rect 50387 11101 50399 11135
rect 50614 11132 50620 11144
rect 50575 11104 50620 11132
rect 50341 11095 50399 11101
rect 50614 11092 50620 11104
rect 50672 11092 50678 11144
rect 50706 11092 50712 11144
rect 50764 11132 50770 11144
rect 51258 11132 51264 11144
rect 50764 11104 51264 11132
rect 50764 11092 50770 11104
rect 51258 11092 51264 11104
rect 51316 11092 51322 11144
rect 51445 11135 51503 11141
rect 51445 11101 51457 11135
rect 51491 11132 51503 11135
rect 51718 11132 51724 11144
rect 51491 11104 51724 11132
rect 51491 11101 51503 11104
rect 51445 11095 51503 11101
rect 51718 11092 51724 11104
rect 51776 11092 51782 11144
rect 51997 11135 52055 11141
rect 51997 11101 52009 11135
rect 52043 11101 52055 11135
rect 52104 11132 52132 11172
rect 53558 11160 53564 11212
rect 53616 11200 53622 11212
rect 54386 11200 54392 11212
rect 53616 11172 54392 11200
rect 53616 11160 53622 11172
rect 54386 11160 54392 11172
rect 54444 11160 54450 11212
rect 54496 11200 54524 11299
rect 57330 11296 57336 11308
rect 57388 11296 57394 11348
rect 57606 11296 57612 11348
rect 57664 11336 57670 11348
rect 59630 11336 59636 11348
rect 57664 11308 59636 11336
rect 57664 11296 57670 11308
rect 59630 11296 59636 11308
rect 59688 11296 59694 11348
rect 62482 11296 62488 11348
rect 62540 11336 62546 11348
rect 63586 11336 63592 11348
rect 62540 11308 63264 11336
rect 63547 11308 63592 11336
rect 62540 11296 62546 11308
rect 63236 11280 63264 11308
rect 63586 11296 63592 11308
rect 63644 11296 63650 11348
rect 64414 11296 64420 11348
rect 64472 11336 64478 11348
rect 64877 11339 64935 11345
rect 64877 11336 64889 11339
rect 64472 11308 64889 11336
rect 64472 11296 64478 11308
rect 64877 11305 64889 11308
rect 64923 11336 64935 11339
rect 64966 11336 64972 11348
rect 64923 11308 64972 11336
rect 64923 11305 64935 11308
rect 64877 11299 64935 11305
rect 64966 11296 64972 11308
rect 65024 11296 65030 11348
rect 66530 11336 66536 11348
rect 66364 11308 66536 11336
rect 54662 11268 54668 11280
rect 54623 11240 54668 11268
rect 54662 11228 54668 11240
rect 54720 11228 54726 11280
rect 54754 11228 54760 11280
rect 54812 11268 54818 11280
rect 55861 11271 55919 11277
rect 55861 11268 55873 11271
rect 54812 11240 55873 11268
rect 54812 11228 54818 11240
rect 55861 11237 55873 11240
rect 55907 11237 55919 11271
rect 55861 11231 55919 11237
rect 55950 11228 55956 11280
rect 56008 11268 56014 11280
rect 56965 11271 57023 11277
rect 56965 11268 56977 11271
rect 56008 11240 56977 11268
rect 56008 11228 56014 11240
rect 56965 11237 56977 11240
rect 57011 11237 57023 11271
rect 56965 11231 57023 11237
rect 57422 11228 57428 11280
rect 57480 11268 57486 11280
rect 58713 11271 58771 11277
rect 58713 11268 58725 11271
rect 57480 11240 58725 11268
rect 57480 11228 57486 11240
rect 58713 11237 58725 11240
rect 58759 11268 58771 11271
rect 59170 11268 59176 11280
rect 58759 11240 59176 11268
rect 58759 11237 58771 11240
rect 58713 11231 58771 11237
rect 59170 11228 59176 11240
rect 59228 11228 59234 11280
rect 61654 11268 61660 11280
rect 59464 11240 61660 11268
rect 58158 11200 58164 11212
rect 54496 11172 58164 11200
rect 58158 11160 58164 11172
rect 58216 11200 58222 11212
rect 58434 11200 58440 11212
rect 58216 11172 58440 11200
rect 58216 11160 58222 11172
rect 58434 11160 58440 11172
rect 58492 11160 58498 11212
rect 58618 11200 58624 11212
rect 58579 11172 58624 11200
rect 58618 11160 58624 11172
rect 58676 11160 58682 11212
rect 58842 11203 58900 11209
rect 58842 11169 58854 11203
rect 58888 11200 58900 11203
rect 59078 11200 59084 11212
rect 58888 11172 59084 11200
rect 58888 11169 58900 11172
rect 58842 11163 58900 11169
rect 59078 11160 59084 11172
rect 59136 11160 59142 11212
rect 52825 11135 52883 11141
rect 52825 11132 52837 11135
rect 52104 11104 52837 11132
rect 51997 11095 52055 11101
rect 52825 11101 52837 11104
rect 52871 11132 52883 11135
rect 52871 11104 54524 11132
rect 52871 11101 52883 11104
rect 52825 11095 52883 11101
rect 50522 11064 50528 11076
rect 42852 11036 46888 11064
rect 47702 11036 50528 11064
rect 42852 11024 42858 11036
rect 50522 11024 50528 11036
rect 50580 11024 50586 11076
rect 50890 11024 50896 11076
rect 50948 11064 50954 11076
rect 51350 11064 51356 11076
rect 50948 11036 51074 11064
rect 51311 11036 51356 11064
rect 50948 11024 50954 11036
rect 39816 10968 42104 10996
rect 39816 10956 39822 10968
rect 42702 10956 42708 11008
rect 42760 10996 42766 11008
rect 49234 10996 49240 11008
rect 42760 10968 49240 10996
rect 42760 10956 42766 10968
rect 49234 10956 49240 10968
rect 49292 10956 49298 11008
rect 49694 10956 49700 11008
rect 49752 10996 49758 11008
rect 50433 10999 50491 11005
rect 50433 10996 50445 10999
rect 49752 10968 50445 10996
rect 49752 10956 49758 10968
rect 50433 10965 50445 10968
rect 50479 10965 50491 10999
rect 50798 10996 50804 11008
rect 50759 10968 50804 10996
rect 50433 10959 50491 10965
rect 50798 10956 50804 10968
rect 50856 10956 50862 11008
rect 51046 10996 51074 11036
rect 51350 11024 51356 11036
rect 51408 11024 51414 11076
rect 52012 11064 52040 11095
rect 52730 11064 52736 11076
rect 51460 11036 52736 11064
rect 51460 10996 51488 11036
rect 52730 11024 52736 11036
rect 52788 11024 52794 11076
rect 53006 11024 53012 11076
rect 53064 11024 53070 11076
rect 54297 11067 54355 11073
rect 54297 11033 54309 11067
rect 54343 11064 54355 11067
rect 54386 11064 54392 11076
rect 54343 11036 54392 11064
rect 54343 11033 54355 11036
rect 54297 11027 54355 11033
rect 54386 11024 54392 11036
rect 54444 11024 54450 11076
rect 54496 11064 54524 11104
rect 54662 11092 54668 11144
rect 54720 11132 54726 11144
rect 55122 11132 55128 11144
rect 54720 11104 55128 11132
rect 54720 11092 54726 11104
rect 55122 11092 55128 11104
rect 55180 11132 55186 11144
rect 56042 11132 56048 11144
rect 55180 11104 56048 11132
rect 55180 11092 55186 11104
rect 56042 11092 56048 11104
rect 56100 11092 56106 11144
rect 56134 11092 56140 11144
rect 56192 11132 56198 11144
rect 56192 11104 56237 11132
rect 56192 11092 56198 11104
rect 56318 11092 56324 11144
rect 56376 11132 56382 11144
rect 57330 11132 57336 11144
rect 56376 11104 56421 11132
rect 57291 11104 57336 11132
rect 56376 11092 56382 11104
rect 57330 11092 57336 11104
rect 57388 11092 57394 11144
rect 57698 11092 57704 11144
rect 57756 11132 57762 11144
rect 59464 11141 59492 11240
rect 61654 11228 61660 11240
rect 61712 11228 61718 11280
rect 61746 11228 61752 11280
rect 61804 11268 61810 11280
rect 61804 11240 61976 11268
rect 61804 11228 61810 11240
rect 60734 11160 60740 11212
rect 60792 11200 60798 11212
rect 60792 11172 60837 11200
rect 60792 11160 60798 11172
rect 60918 11160 60924 11212
rect 60976 11200 60982 11212
rect 61838 11200 61844 11212
rect 60976 11172 61021 11200
rect 61799 11172 61844 11200
rect 60976 11160 60982 11172
rect 61838 11160 61844 11172
rect 61896 11160 61902 11212
rect 61948 11200 61976 11240
rect 63218 11228 63224 11280
rect 63276 11268 63282 11280
rect 64432 11268 64460 11296
rect 66364 11277 66392 11308
rect 66530 11296 66536 11308
rect 66588 11296 66594 11348
rect 67266 11296 67272 11348
rect 67324 11336 67330 11348
rect 67450 11336 67456 11348
rect 67324 11308 67456 11336
rect 67324 11296 67330 11308
rect 67450 11296 67456 11308
rect 67508 11296 67514 11348
rect 67606 11308 69980 11336
rect 63276 11240 64460 11268
rect 66349 11271 66407 11277
rect 63276 11228 63282 11240
rect 66349 11237 66361 11271
rect 66395 11237 66407 11271
rect 66349 11231 66407 11237
rect 66438 11228 66444 11280
rect 66496 11268 66502 11280
rect 67606 11268 67634 11308
rect 66496 11240 67634 11268
rect 66496 11228 66502 11240
rect 62117 11203 62175 11209
rect 62117 11200 62129 11203
rect 61948 11172 62129 11200
rect 62117 11169 62129 11172
rect 62163 11169 62175 11203
rect 62117 11163 62175 11169
rect 62482 11160 62488 11212
rect 62540 11200 62546 11212
rect 65889 11203 65947 11209
rect 65889 11200 65901 11203
rect 62540 11172 65901 11200
rect 62540 11160 62546 11172
rect 65889 11169 65901 11172
rect 65935 11169 65947 11203
rect 65889 11163 65947 11169
rect 66622 11160 66628 11212
rect 66680 11200 66686 11212
rect 69750 11200 69756 11212
rect 66680 11172 67634 11200
rect 69711 11172 69756 11200
rect 66680 11160 66686 11172
rect 59449 11135 59507 11141
rect 59449 11132 59461 11135
rect 57756 11104 59461 11132
rect 57756 11092 57762 11104
rect 59449 11101 59461 11104
rect 59495 11101 59507 11135
rect 59630 11132 59636 11144
rect 59591 11104 59636 11132
rect 59449 11095 59507 11101
rect 59630 11092 59636 11104
rect 59688 11092 59694 11144
rect 61013 11135 61071 11141
rect 61013 11132 61025 11135
rect 60706 11104 61025 11132
rect 56502 11064 56508 11076
rect 54496 11036 56508 11064
rect 56502 11024 56508 11036
rect 56560 11024 56566 11076
rect 57149 11067 57207 11073
rect 57149 11033 57161 11067
rect 57195 11064 57207 11067
rect 57974 11064 57980 11076
rect 57195 11036 57980 11064
rect 57195 11033 57207 11036
rect 57149 11027 57207 11033
rect 57974 11024 57980 11036
rect 58032 11024 58038 11076
rect 58250 11064 58256 11076
rect 58211 11036 58256 11064
rect 58250 11024 58256 11036
rect 58308 11024 58314 11076
rect 58434 11024 58440 11076
rect 58492 11064 58498 11076
rect 58986 11064 58992 11076
rect 58492 11036 58992 11064
rect 58492 11024 58498 11036
rect 58986 11024 58992 11036
rect 59044 11024 59050 11076
rect 59078 11024 59084 11076
rect 59136 11064 59142 11076
rect 59541 11067 59599 11073
rect 59541 11064 59553 11067
rect 59136 11036 59553 11064
rect 59136 11024 59142 11036
rect 59541 11033 59553 11036
rect 59587 11033 59599 11067
rect 59541 11027 59599 11033
rect 51046 10968 51488 10996
rect 51810 10956 51816 11008
rect 51868 10996 51874 11008
rect 53558 10996 53564 11008
rect 51868 10968 53564 10996
rect 51868 10956 51874 10968
rect 53558 10956 53564 10968
rect 53616 10956 53622 11008
rect 54202 10956 54208 11008
rect 54260 10996 54266 11008
rect 54497 10999 54555 11005
rect 54497 10996 54509 10999
rect 54260 10968 54509 10996
rect 54260 10956 54266 10968
rect 54497 10965 54509 10968
rect 54543 10965 54555 10999
rect 54497 10959 54555 10965
rect 54938 10956 54944 11008
rect 54996 10996 55002 11008
rect 59446 10996 59452 11008
rect 54996 10968 59452 10996
rect 54996 10956 55002 10968
rect 59446 10956 59452 10968
rect 59504 10956 59510 11008
rect 60550 10956 60556 11008
rect 60608 10996 60614 11008
rect 60706 10996 60734 11104
rect 61013 11101 61025 11104
rect 61059 11132 61071 11135
rect 61470 11132 61476 11144
rect 61059 11104 61476 11132
rect 61059 11101 61071 11104
rect 61013 11095 61071 11101
rect 61470 11092 61476 11104
rect 61528 11092 61534 11144
rect 64325 11135 64383 11141
rect 64325 11101 64337 11135
rect 64371 11132 64383 11135
rect 64598 11132 64604 11144
rect 64371 11104 64604 11132
rect 64371 11101 64383 11104
rect 64325 11095 64383 11101
rect 64598 11092 64604 11104
rect 64656 11132 64662 11144
rect 65426 11132 65432 11144
rect 64656 11104 65432 11132
rect 64656 11092 64662 11104
rect 65426 11092 65432 11104
rect 65484 11092 65490 11144
rect 65978 11132 65984 11144
rect 65939 11104 65984 11132
rect 65978 11092 65984 11104
rect 66036 11092 66042 11144
rect 62114 11064 62120 11076
rect 61396 11036 62120 11064
rect 61396 11005 61424 11036
rect 62114 11024 62120 11036
rect 62172 11064 62178 11076
rect 62390 11064 62396 11076
rect 62172 11036 62396 11064
rect 62172 11024 62178 11036
rect 62390 11024 62396 11036
rect 62448 11024 62454 11076
rect 64233 11067 64291 11073
rect 64233 11064 64245 11067
rect 63342 11036 64245 11064
rect 64233 11033 64245 11036
rect 64279 11033 64291 11067
rect 67082 11064 67088 11076
rect 67043 11036 67088 11064
rect 64233 11027 64291 11033
rect 67082 11024 67088 11036
rect 67140 11024 67146 11076
rect 67606 11064 67634 11172
rect 69750 11160 69756 11172
rect 69808 11160 69814 11212
rect 69952 11200 69980 11308
rect 72694 11296 72700 11348
rect 72752 11336 72758 11348
rect 74074 11336 74080 11348
rect 72752 11308 73936 11336
rect 74035 11308 74080 11336
rect 72752 11296 72758 11308
rect 70029 11271 70087 11277
rect 70029 11237 70041 11271
rect 70075 11268 70087 11271
rect 73798 11268 73804 11280
rect 70075 11240 73804 11268
rect 70075 11237 70087 11240
rect 70029 11231 70087 11237
rect 73798 11228 73804 11240
rect 73856 11228 73862 11280
rect 73908 11268 73936 11308
rect 74074 11296 74080 11308
rect 74132 11296 74138 11348
rect 74442 11296 74448 11348
rect 74500 11336 74506 11348
rect 75270 11336 75276 11348
rect 74500 11308 75276 11336
rect 74500 11296 74506 11308
rect 75270 11296 75276 11308
rect 75328 11336 75334 11348
rect 76650 11336 76656 11348
rect 75328 11308 76656 11336
rect 75328 11296 75334 11308
rect 76650 11296 76656 11308
rect 76708 11296 76714 11348
rect 76926 11336 76932 11348
rect 76887 11308 76932 11336
rect 76926 11296 76932 11308
rect 76984 11296 76990 11348
rect 77110 11296 77116 11348
rect 77168 11336 77174 11348
rect 77389 11339 77447 11345
rect 77389 11336 77401 11339
rect 77168 11308 77401 11336
rect 77168 11296 77174 11308
rect 77389 11305 77401 11308
rect 77435 11305 77447 11339
rect 77389 11299 77447 11305
rect 77478 11296 77484 11348
rect 77536 11336 77542 11348
rect 78122 11336 78128 11348
rect 77536 11308 78128 11336
rect 77536 11296 77542 11308
rect 78122 11296 78128 11308
rect 78180 11336 78186 11348
rect 78582 11336 78588 11348
rect 78180 11308 78588 11336
rect 78180 11296 78186 11308
rect 78582 11296 78588 11308
rect 78640 11296 78646 11348
rect 78858 11336 78864 11348
rect 78819 11308 78864 11336
rect 78858 11296 78864 11308
rect 78916 11296 78922 11348
rect 79505 11339 79563 11345
rect 79505 11305 79517 11339
rect 79551 11336 79563 11339
rect 79962 11336 79968 11348
rect 79551 11308 79968 11336
rect 79551 11305 79563 11308
rect 79505 11299 79563 11305
rect 79962 11296 79968 11308
rect 80020 11296 80026 11348
rect 84611 11339 84669 11345
rect 84611 11305 84623 11339
rect 84657 11336 84669 11339
rect 85022 11336 85028 11348
rect 84657 11308 85028 11336
rect 84657 11305 84669 11308
rect 84611 11299 84669 11305
rect 85022 11296 85028 11308
rect 85080 11296 85086 11348
rect 85206 11336 85212 11348
rect 85167 11308 85212 11336
rect 85206 11296 85212 11308
rect 85264 11296 85270 11348
rect 87690 11296 87696 11348
rect 87748 11336 87754 11348
rect 87969 11339 88027 11345
rect 87969 11336 87981 11339
rect 87748 11308 87981 11336
rect 87748 11296 87754 11308
rect 87969 11305 87981 11308
rect 88015 11305 88027 11339
rect 90542 11336 90548 11348
rect 90503 11308 90548 11336
rect 87969 11299 88027 11305
rect 90542 11296 90548 11308
rect 90600 11296 90606 11348
rect 91830 11336 91836 11348
rect 91572 11308 91836 11336
rect 74166 11268 74172 11280
rect 73908 11240 74172 11268
rect 74166 11228 74172 11240
rect 74224 11228 74230 11280
rect 74350 11268 74356 11280
rect 74311 11240 74356 11268
rect 74350 11228 74356 11240
rect 74408 11268 74414 11280
rect 76193 11271 76251 11277
rect 76193 11268 76205 11271
rect 74408 11240 76205 11268
rect 74408 11228 74414 11240
rect 76193 11237 76205 11240
rect 76239 11237 76251 11271
rect 77754 11268 77760 11280
rect 76193 11231 76251 11237
rect 77588 11240 77760 11268
rect 72786 11200 72792 11212
rect 69952 11172 72792 11200
rect 68554 11132 68560 11144
rect 67836 11126 68560 11132
rect 67744 11104 68560 11126
rect 67744 11098 67864 11104
rect 67744 11064 67772 11098
rect 68554 11092 68560 11104
rect 68612 11092 68618 11144
rect 68925 11135 68983 11141
rect 68925 11101 68937 11135
rect 68971 11132 68983 11135
rect 69198 11132 69204 11144
rect 68971 11104 69204 11132
rect 68971 11101 68983 11104
rect 68925 11095 68983 11101
rect 69198 11092 69204 11104
rect 69256 11092 69262 11144
rect 69474 11092 69480 11144
rect 69532 11132 69538 11144
rect 69661 11135 69719 11141
rect 69661 11132 69673 11135
rect 69532 11104 69673 11132
rect 69532 11092 69538 11104
rect 69661 11101 69673 11104
rect 69707 11132 69719 11135
rect 70670 11132 70676 11144
rect 69707 11104 70676 11132
rect 69707 11101 69719 11104
rect 69661 11095 69719 11101
rect 70670 11092 70676 11104
rect 70728 11092 70734 11144
rect 71130 11132 71136 11144
rect 71091 11104 71136 11132
rect 71130 11092 71136 11104
rect 71188 11092 71194 11144
rect 71240 11141 71268 11172
rect 72786 11160 72792 11172
rect 72844 11200 72850 11212
rect 75362 11200 75368 11212
rect 72844 11172 75368 11200
rect 72844 11160 72850 11172
rect 74368 11144 74396 11172
rect 75362 11160 75368 11172
rect 75420 11160 75426 11212
rect 75730 11160 75736 11212
rect 75788 11200 75794 11212
rect 76653 11203 76711 11209
rect 76653 11200 76665 11203
rect 75788 11172 76665 11200
rect 75788 11160 75794 11172
rect 76653 11169 76665 11172
rect 76699 11169 76711 11203
rect 76653 11163 76711 11169
rect 76745 11203 76803 11209
rect 76745 11169 76757 11203
rect 76791 11200 76803 11203
rect 76834 11200 76840 11212
rect 76791 11172 76840 11200
rect 76791 11169 76803 11172
rect 76745 11163 76803 11169
rect 76834 11160 76840 11172
rect 76892 11160 76898 11212
rect 77588 11200 77616 11240
rect 77754 11228 77760 11240
rect 77812 11268 77818 11280
rect 78490 11268 78496 11280
rect 77812 11240 78496 11268
rect 77812 11228 77818 11240
rect 78490 11228 78496 11240
rect 78548 11228 78554 11280
rect 80698 11228 80704 11280
rect 80756 11268 80762 11280
rect 80756 11240 83320 11268
rect 80756 11228 80762 11240
rect 77654 11203 77712 11209
rect 77654 11200 77666 11203
rect 77588 11172 77666 11200
rect 77654 11169 77666 11172
rect 77700 11169 77712 11203
rect 77846 11200 77852 11212
rect 77807 11172 77852 11200
rect 77654 11163 77712 11169
rect 77846 11160 77852 11172
rect 77904 11160 77910 11212
rect 80146 11200 80152 11212
rect 78324 11172 80152 11200
rect 71225 11135 71283 11141
rect 71225 11101 71237 11135
rect 71271 11101 71283 11135
rect 72326 11132 72332 11144
rect 72287 11104 72332 11132
rect 71225 11095 71283 11101
rect 72326 11092 72332 11104
rect 72384 11092 72390 11144
rect 72697 11135 72755 11141
rect 72697 11101 72709 11135
rect 72743 11132 72755 11135
rect 73062 11132 73068 11144
rect 72743 11104 73068 11132
rect 72743 11101 72755 11104
rect 72697 11095 72755 11101
rect 73062 11092 73068 11104
rect 73120 11092 73126 11144
rect 73525 11135 73583 11141
rect 73525 11101 73537 11135
rect 73571 11132 73583 11135
rect 73614 11132 73620 11144
rect 73571 11104 73620 11132
rect 73571 11101 73583 11104
rect 73525 11095 73583 11101
rect 73614 11092 73620 11104
rect 73672 11092 73678 11144
rect 73982 11092 73988 11144
rect 74040 11132 74046 11144
rect 74261 11135 74319 11141
rect 74261 11132 74273 11135
rect 74040 11104 74273 11132
rect 74040 11092 74046 11104
rect 74261 11101 74273 11104
rect 74307 11101 74319 11135
rect 74261 11095 74319 11101
rect 74350 11092 74356 11144
rect 74408 11092 74414 11144
rect 74445 11135 74503 11141
rect 74445 11101 74457 11135
rect 74491 11101 74503 11135
rect 74445 11095 74503 11101
rect 74537 11135 74595 11141
rect 74537 11101 74549 11135
rect 74583 11132 74595 11135
rect 75089 11135 75147 11141
rect 75089 11132 75101 11135
rect 74583 11104 75101 11132
rect 74583 11101 74595 11104
rect 74537 11095 74595 11101
rect 75089 11101 75101 11104
rect 75135 11101 75147 11135
rect 75270 11132 75276 11144
rect 75231 11104 75276 11132
rect 75089 11095 75147 11101
rect 71866 11064 71872 11076
rect 67606 11036 67772 11064
rect 71827 11036 71872 11064
rect 71866 11024 71872 11036
rect 71924 11024 71930 11076
rect 74460 11064 74488 11095
rect 75270 11092 75276 11104
rect 75328 11092 75334 11144
rect 75559 11135 75617 11141
rect 75559 11101 75571 11135
rect 75605 11132 75617 11135
rect 76098 11132 76104 11144
rect 75605 11104 76104 11132
rect 75605 11101 75617 11104
rect 75559 11095 75617 11101
rect 76098 11092 76104 11104
rect 76156 11092 76162 11144
rect 77202 11092 77208 11144
rect 77260 11132 77266 11144
rect 77573 11135 77631 11141
rect 77573 11132 77585 11135
rect 77260 11104 77585 11132
rect 77260 11092 77266 11104
rect 77573 11101 77585 11104
rect 77619 11101 77631 11135
rect 77754 11132 77760 11144
rect 77715 11104 77760 11132
rect 77573 11095 77631 11101
rect 75178 11064 75184 11076
rect 74460 11036 75184 11064
rect 75178 11024 75184 11036
rect 75236 11024 75242 11076
rect 75457 11067 75515 11073
rect 75457 11033 75469 11067
rect 75503 11064 75515 11067
rect 75638 11064 75644 11076
rect 75503 11036 75644 11064
rect 75503 11033 75515 11036
rect 75457 11027 75515 11033
rect 75638 11024 75644 11036
rect 75696 11024 75702 11076
rect 76193 11067 76251 11073
rect 76193 11033 76205 11067
rect 76239 11064 76251 11067
rect 77478 11064 77484 11076
rect 76239 11036 77484 11064
rect 76239 11033 76251 11036
rect 76193 11027 76251 11033
rect 60608 10968 60734 10996
rect 61381 10999 61439 11005
rect 60608 10956 60614 10968
rect 61381 10965 61393 10999
rect 61427 10965 61439 10999
rect 61381 10959 61439 10965
rect 61470 10956 61476 11008
rect 61528 10996 61534 11008
rect 67450 10996 67456 11008
rect 61528 10968 67456 10996
rect 61528 10956 61534 10968
rect 67450 10956 67456 10968
rect 67508 10996 67514 11008
rect 71038 10996 71044 11008
rect 67508 10968 71044 10996
rect 67508 10956 67514 10968
rect 71038 10956 71044 10968
rect 71096 10956 71102 11008
rect 71130 10956 71136 11008
rect 71188 10996 71194 11008
rect 76208 10996 76236 11027
rect 77478 11024 77484 11036
rect 77536 11024 77542 11076
rect 77588 11064 77616 11095
rect 77754 11092 77760 11104
rect 77812 11132 77818 11144
rect 78324 11132 78352 11172
rect 80146 11160 80152 11172
rect 80204 11200 80210 11212
rect 81158 11200 81164 11212
rect 80204 11172 81164 11200
rect 80204 11160 80210 11172
rect 81158 11160 81164 11172
rect 81216 11160 81222 11212
rect 81434 11160 81440 11212
rect 81492 11200 81498 11212
rect 81492 11172 81756 11200
rect 81492 11160 81498 11172
rect 77812 11104 78352 11132
rect 78401 11135 78459 11141
rect 77812 11092 77818 11104
rect 78401 11101 78413 11135
rect 78447 11101 78459 11135
rect 78401 11095 78459 11101
rect 78493 11135 78551 11141
rect 78493 11101 78505 11135
rect 78539 11132 78551 11135
rect 78582 11132 78588 11144
rect 78539 11104 78588 11132
rect 78539 11101 78551 11104
rect 78493 11095 78551 11101
rect 78416 11064 78444 11095
rect 78582 11092 78588 11104
rect 78640 11092 78646 11144
rect 78674 11092 78680 11144
rect 78732 11132 78738 11144
rect 79594 11132 79600 11144
rect 78732 11104 78777 11132
rect 79555 11104 79600 11132
rect 78732 11092 78738 11104
rect 79594 11092 79600 11104
rect 79652 11092 79658 11144
rect 81728 11141 81756 11172
rect 80517 11135 80575 11141
rect 80517 11101 80529 11135
rect 80563 11132 80575 11135
rect 81713 11135 81771 11141
rect 80563 11104 81664 11132
rect 80563 11101 80575 11104
rect 80517 11095 80575 11101
rect 77588 11036 78444 11064
rect 78858 11024 78864 11076
rect 78916 11064 78922 11076
rect 79686 11064 79692 11076
rect 78916 11036 79692 11064
rect 78916 11024 78922 11036
rect 79686 11024 79692 11036
rect 79744 11024 79750 11076
rect 81636 11064 81664 11104
rect 81713 11101 81725 11135
rect 81759 11101 81771 11135
rect 82538 11132 82544 11144
rect 82499 11104 82544 11132
rect 81713 11095 81771 11101
rect 82538 11092 82544 11104
rect 82596 11092 82602 11144
rect 83292 11132 83320 11240
rect 84286 11228 84292 11280
rect 84344 11268 84350 11280
rect 84473 11271 84531 11277
rect 84473 11268 84485 11271
rect 84344 11240 84485 11268
rect 84344 11228 84350 11240
rect 84473 11237 84485 11240
rect 84519 11237 84531 11271
rect 85758 11268 85764 11280
rect 85719 11240 85764 11268
rect 84473 11231 84531 11237
rect 85758 11228 85764 11240
rect 85816 11228 85822 11280
rect 85942 11228 85948 11280
rect 86000 11268 86006 11280
rect 88705 11271 88763 11277
rect 88705 11268 88717 11271
rect 86000 11240 88717 11268
rect 86000 11228 86006 11240
rect 88705 11237 88717 11240
rect 88751 11237 88763 11271
rect 91572 11268 91600 11308
rect 91830 11296 91836 11308
rect 91888 11336 91894 11348
rect 92290 11336 92296 11348
rect 91888 11308 92296 11336
rect 91888 11296 91894 11308
rect 92290 11296 92296 11308
rect 92348 11296 92354 11348
rect 93302 11336 93308 11348
rect 93263 11308 93308 11336
rect 93302 11296 93308 11308
rect 93360 11296 93366 11348
rect 88705 11231 88763 11237
rect 90008 11240 91600 11268
rect 83734 11160 83740 11212
rect 83792 11200 83798 11212
rect 84010 11200 84016 11212
rect 83792 11172 84016 11200
rect 83792 11160 83798 11172
rect 84010 11160 84016 11172
rect 84068 11160 84074 11212
rect 84102 11160 84108 11212
rect 84160 11200 84166 11212
rect 84381 11203 84439 11209
rect 84381 11200 84393 11203
rect 84160 11172 84393 11200
rect 84160 11160 84166 11172
rect 84381 11169 84393 11172
rect 84427 11169 84439 11203
rect 84381 11163 84439 11169
rect 86218 11160 86224 11212
rect 86276 11200 86282 11212
rect 86589 11203 86647 11209
rect 86589 11200 86601 11203
rect 86276 11172 86601 11200
rect 86276 11160 86282 11172
rect 86589 11169 86601 11172
rect 86635 11169 86647 11203
rect 86589 11163 86647 11169
rect 86862 11160 86868 11212
rect 86920 11200 86926 11212
rect 89257 11203 89315 11209
rect 89257 11200 89269 11203
rect 86920 11172 89269 11200
rect 86920 11160 86926 11172
rect 89257 11169 89269 11172
rect 89303 11169 89315 11203
rect 89257 11163 89315 11169
rect 83292 11104 84792 11132
rect 82170 11064 82176 11076
rect 80256 11036 80560 11064
rect 81636 11036 82176 11064
rect 71188 10968 76236 10996
rect 71188 10956 71194 10968
rect 77110 10956 77116 11008
rect 77168 10996 77174 11008
rect 80256 10996 80284 11036
rect 80422 10996 80428 11008
rect 77168 10968 80284 10996
rect 80383 10968 80428 10996
rect 77168 10956 77174 10968
rect 80422 10956 80428 10968
rect 80480 10956 80486 11008
rect 80532 10996 80560 11036
rect 82170 11024 82176 11036
rect 82228 11024 82234 11076
rect 84010 11064 84016 11076
rect 82556 11036 82662 11064
rect 83971 11036 84016 11064
rect 82556 10996 82584 11036
rect 84010 11024 84016 11036
rect 84068 11024 84074 11076
rect 84764 11073 84792 11104
rect 86034 11092 86040 11144
rect 86092 11132 86098 11144
rect 90008 11141 90036 11240
rect 91833 11203 91891 11209
rect 91833 11169 91845 11203
rect 91879 11200 91891 11203
rect 93857 11203 93915 11209
rect 93857 11200 93869 11203
rect 91879 11172 93869 11200
rect 91879 11169 91891 11172
rect 91833 11163 91891 11169
rect 93857 11169 93869 11172
rect 93903 11169 93915 11203
rect 93857 11163 93915 11169
rect 86681 11135 86739 11141
rect 86681 11132 86693 11135
rect 86092 11104 86693 11132
rect 86092 11092 86098 11104
rect 86681 11101 86693 11104
rect 86727 11101 86739 11135
rect 87969 11135 88027 11141
rect 87969 11132 87981 11135
rect 86681 11095 86739 11101
rect 86926 11104 87981 11132
rect 84749 11067 84807 11073
rect 84749 11033 84761 11067
rect 84795 11064 84807 11067
rect 86586 11064 86592 11076
rect 84795 11036 86592 11064
rect 84795 11033 84807 11036
rect 84749 11027 84807 11033
rect 86586 11024 86592 11036
rect 86644 11024 86650 11076
rect 86696 11064 86724 11095
rect 86926 11064 86954 11104
rect 87969 11101 87981 11104
rect 88015 11101 88027 11135
rect 87969 11095 88027 11101
rect 89993 11135 90051 11141
rect 89993 11101 90005 11135
rect 90039 11101 90051 11135
rect 90450 11132 90456 11144
rect 90411 11104 90456 11132
rect 89993 11095 90051 11101
rect 90450 11092 90456 11104
rect 90508 11092 90514 11144
rect 91557 11135 91615 11141
rect 91557 11101 91569 11135
rect 91603 11101 91615 11135
rect 93762 11132 93768 11144
rect 93723 11104 93768 11132
rect 91557 11095 91615 11101
rect 86696 11036 86954 11064
rect 87509 11067 87567 11073
rect 87509 11033 87521 11067
rect 87555 11064 87567 11067
rect 88150 11064 88156 11076
rect 87555 11036 88156 11064
rect 87555 11033 87567 11036
rect 87509 11027 87567 11033
rect 88150 11024 88156 11036
rect 88208 11024 88214 11076
rect 89622 11024 89628 11076
rect 89680 11064 89686 11076
rect 91572 11064 91600 11095
rect 93762 11092 93768 11104
rect 93820 11092 93826 11144
rect 94222 11064 94228 11076
rect 89680 11036 91600 11064
rect 93058 11036 94228 11064
rect 89680 11024 89686 11036
rect 94222 11024 94228 11036
rect 94280 11024 94286 11076
rect 84102 10996 84108 11008
rect 80532 10968 84108 10996
rect 84102 10956 84108 10968
rect 84160 10956 84166 11008
rect 84286 10956 84292 11008
rect 84344 10996 84350 11008
rect 86862 10996 86868 11008
rect 84344 10968 86868 10996
rect 84344 10956 84350 10968
rect 86862 10956 86868 10968
rect 86920 10956 86926 11008
rect 89898 10996 89904 11008
rect 89859 10968 89904 10996
rect 89898 10956 89904 10968
rect 89956 10956 89962 11008
rect 92474 10956 92480 11008
rect 92532 10996 92538 11008
rect 93762 10996 93768 11008
rect 92532 10968 93768 10996
rect 92532 10956 92538 10968
rect 93762 10956 93768 10968
rect 93820 10956 93826 11008
rect 1104 10906 95011 10928
rect 1104 10854 24386 10906
rect 24438 10854 24450 10906
rect 24502 10854 24514 10906
rect 24566 10854 24578 10906
rect 24630 10854 24642 10906
rect 24694 10854 47823 10906
rect 47875 10854 47887 10906
rect 47939 10854 47951 10906
rect 48003 10854 48015 10906
rect 48067 10854 48079 10906
rect 48131 10854 71260 10906
rect 71312 10854 71324 10906
rect 71376 10854 71388 10906
rect 71440 10854 71452 10906
rect 71504 10854 71516 10906
rect 71568 10854 94697 10906
rect 94749 10854 94761 10906
rect 94813 10854 94825 10906
rect 94877 10854 94889 10906
rect 94941 10854 94953 10906
rect 95005 10854 95011 10906
rect 1104 10832 95011 10854
rect 1762 10792 1768 10804
rect 1723 10764 1768 10792
rect 1762 10752 1768 10764
rect 1820 10752 1826 10804
rect 4065 10795 4123 10801
rect 4065 10761 4077 10795
rect 4111 10792 4123 10795
rect 4982 10792 4988 10804
rect 4111 10764 4988 10792
rect 4111 10761 4123 10764
rect 4065 10755 4123 10761
rect 4982 10752 4988 10764
rect 5040 10752 5046 10804
rect 8018 10792 8024 10804
rect 5276 10764 8024 10792
rect 3970 10724 3976 10736
rect 3818 10696 3976 10724
rect 3970 10684 3976 10696
rect 4028 10684 4034 10736
rect 4522 10656 4528 10668
rect 4483 10628 4528 10656
rect 4522 10616 4528 10628
rect 4580 10616 4586 10668
rect 5276 10656 5304 10764
rect 8018 10752 8024 10764
rect 8076 10752 8082 10804
rect 9217 10795 9275 10801
rect 9217 10761 9229 10795
rect 9263 10792 9275 10795
rect 10134 10792 10140 10804
rect 9263 10764 10140 10792
rect 9263 10761 9275 10764
rect 9217 10755 9275 10761
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 11146 10792 11152 10804
rect 11107 10764 11152 10792
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 12250 10792 12256 10804
rect 12211 10764 12256 10792
rect 12250 10752 12256 10764
rect 12308 10752 12314 10804
rect 12820 10764 15148 10792
rect 7098 10684 7104 10736
rect 7156 10724 7162 10736
rect 7745 10727 7803 10733
rect 7745 10724 7757 10727
rect 7156 10696 7757 10724
rect 7156 10684 7162 10696
rect 7745 10693 7757 10696
rect 7791 10693 7803 10727
rect 12820 10724 12848 10764
rect 12986 10724 12992 10736
rect 7745 10687 7803 10693
rect 9048 10696 12848 10724
rect 12947 10696 12992 10724
rect 6730 10656 6736 10668
rect 4632 10628 5304 10656
rect 6643 10628 6736 10656
rect 2314 10588 2320 10600
rect 2275 10560 2320 10588
rect 2314 10548 2320 10560
rect 2372 10548 2378 10600
rect 2593 10591 2651 10597
rect 2593 10557 2605 10591
rect 2639 10588 2651 10591
rect 4632 10588 4660 10628
rect 6730 10616 6736 10628
rect 6788 10656 6794 10668
rect 7466 10656 7472 10668
rect 6788 10628 7328 10656
rect 7427 10628 7472 10656
rect 6788 10616 6794 10628
rect 4798 10588 4804 10600
rect 2639 10560 4660 10588
rect 4759 10560 4804 10588
rect 2639 10557 2651 10560
rect 2593 10551 2651 10557
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 7300 10588 7328 10628
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 8846 10616 8852 10668
rect 8904 10616 8910 10668
rect 9048 10588 9076 10696
rect 12986 10684 12992 10696
rect 13044 10684 13050 10736
rect 14826 10684 14832 10736
rect 14884 10724 14890 10736
rect 15013 10727 15071 10733
rect 15013 10724 15025 10727
rect 14884 10696 15025 10724
rect 14884 10684 14890 10696
rect 15013 10693 15025 10696
rect 15059 10693 15071 10727
rect 15120 10724 15148 10764
rect 15194 10752 15200 10804
rect 15252 10801 15258 10804
rect 15252 10795 15276 10801
rect 15264 10761 15276 10795
rect 15378 10792 15384 10804
rect 15339 10764 15384 10792
rect 15252 10755 15276 10761
rect 15252 10752 15258 10755
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 18230 10752 18236 10804
rect 18288 10792 18294 10804
rect 18693 10795 18751 10801
rect 18693 10792 18705 10795
rect 18288 10764 18705 10792
rect 18288 10752 18294 10764
rect 18693 10761 18705 10764
rect 18739 10761 18751 10795
rect 18693 10755 18751 10761
rect 18782 10752 18788 10804
rect 18840 10792 18846 10804
rect 24302 10792 24308 10804
rect 18840 10764 24308 10792
rect 18840 10752 18846 10764
rect 24302 10752 24308 10764
rect 24360 10752 24366 10804
rect 24486 10752 24492 10804
rect 24544 10792 24550 10804
rect 24544 10764 28028 10792
rect 24544 10752 24550 10764
rect 15470 10724 15476 10736
rect 15120 10696 15476 10724
rect 15013 10687 15071 10693
rect 15470 10684 15476 10696
rect 15528 10684 15534 10736
rect 16758 10684 16764 10736
rect 16816 10724 16822 10736
rect 20990 10724 20996 10736
rect 16816 10696 20996 10724
rect 16816 10684 16822 10696
rect 20990 10684 20996 10696
rect 21048 10684 21054 10736
rect 21266 10724 21272 10736
rect 21227 10696 21272 10724
rect 21266 10684 21272 10696
rect 21324 10684 21330 10736
rect 22738 10684 22744 10736
rect 22796 10684 22802 10736
rect 24946 10724 24952 10736
rect 24504 10696 24952 10724
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10656 10103 10659
rect 11054 10656 11060 10668
rect 10091 10628 11060 10656
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 11054 10616 11060 10628
rect 11112 10616 11118 10668
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10656 12035 10659
rect 12066 10656 12072 10668
rect 12023 10628 12072 10656
rect 12023 10625 12035 10628
rect 11977 10619 12035 10625
rect 12066 10616 12072 10628
rect 12124 10616 12130 10668
rect 14090 10616 14096 10668
rect 14148 10616 14154 10668
rect 15841 10659 15899 10665
rect 15841 10625 15853 10659
rect 15887 10625 15899 10659
rect 15841 10619 15899 10625
rect 7300 10580 7512 10588
rect 7576 10580 9076 10588
rect 7300 10560 9076 10580
rect 10137 10591 10195 10597
rect 7484 10552 7604 10560
rect 10137 10557 10149 10591
rect 10183 10588 10195 10591
rect 12158 10588 12164 10600
rect 10183 10560 12164 10588
rect 10183 10557 10195 10560
rect 10137 10551 10195 10557
rect 12158 10548 12164 10560
rect 12216 10548 12222 10600
rect 12253 10591 12311 10597
rect 12253 10557 12265 10591
rect 12299 10588 12311 10591
rect 12299 10560 12434 10588
rect 12299 10557 12311 10560
rect 12253 10551 12311 10557
rect 5442 10480 5448 10532
rect 5500 10520 5506 10532
rect 5537 10523 5595 10529
rect 5537 10520 5549 10523
rect 5500 10492 5549 10520
rect 5500 10480 5506 10492
rect 5537 10489 5549 10492
rect 5583 10520 5595 10523
rect 7098 10520 7104 10532
rect 5583 10492 7104 10520
rect 5583 10489 5595 10492
rect 5537 10483 5595 10489
rect 7098 10480 7104 10492
rect 7156 10480 7162 10532
rect 10413 10523 10471 10529
rect 10413 10489 10425 10523
rect 10459 10520 10471 10523
rect 10962 10520 10968 10532
rect 10459 10492 10968 10520
rect 10459 10489 10471 10492
rect 10413 10483 10471 10489
rect 10962 10480 10968 10492
rect 11020 10480 11026 10532
rect 11146 10480 11152 10532
rect 11204 10520 11210 10532
rect 11882 10520 11888 10532
rect 11204 10492 11888 10520
rect 11204 10480 11210 10492
rect 11882 10480 11888 10492
rect 11940 10520 11946 10532
rect 12069 10523 12127 10529
rect 12069 10520 12081 10523
rect 11940 10492 12081 10520
rect 11940 10480 11946 10492
rect 12069 10489 12081 10492
rect 12115 10489 12127 10523
rect 12069 10483 12127 10489
rect 6638 10452 6644 10464
rect 6599 10424 6644 10452
rect 6638 10412 6644 10424
rect 6696 10412 6702 10464
rect 7466 10412 7472 10464
rect 7524 10452 7530 10464
rect 8110 10452 8116 10464
rect 7524 10424 8116 10452
rect 7524 10412 7530 10424
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 12406 10452 12434 10560
rect 12526 10548 12532 10600
rect 12584 10588 12590 10600
rect 12713 10591 12771 10597
rect 12713 10588 12725 10591
rect 12584 10560 12725 10588
rect 12584 10548 12590 10560
rect 12713 10557 12725 10560
rect 12759 10557 12771 10591
rect 12713 10551 12771 10557
rect 14108 10520 14136 10616
rect 14461 10591 14519 10597
rect 14461 10557 14473 10591
rect 14507 10588 14519 10591
rect 15856 10588 15884 10619
rect 16482 10616 16488 10668
rect 16540 10656 16546 10668
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 16540 10628 17049 10656
rect 16540 10616 16546 10628
rect 17037 10625 17049 10628
rect 17083 10656 17095 10659
rect 18046 10656 18052 10668
rect 17083 10628 18052 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 18046 10616 18052 10628
rect 18104 10616 18110 10668
rect 18233 10659 18291 10665
rect 18233 10625 18245 10659
rect 18279 10625 18291 10659
rect 18233 10619 18291 10625
rect 14507 10560 15884 10588
rect 14507 10557 14519 10560
rect 14461 10551 14519 10557
rect 15930 10548 15936 10600
rect 15988 10588 15994 10600
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 15988 10560 16037 10588
rect 15988 10548 15994 10560
rect 16025 10557 16037 10560
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 16114 10548 16120 10600
rect 16172 10588 16178 10600
rect 16945 10591 17003 10597
rect 16945 10588 16957 10591
rect 16172 10560 16957 10588
rect 16172 10548 16178 10560
rect 16945 10557 16957 10560
rect 16991 10557 17003 10591
rect 16945 10551 17003 10557
rect 17954 10548 17960 10600
rect 18012 10588 18018 10600
rect 18248 10588 18276 10619
rect 18322 10616 18328 10668
rect 18380 10656 18386 10668
rect 19058 10656 19064 10668
rect 18380 10628 18736 10656
rect 19019 10628 19064 10656
rect 18380 10616 18386 10628
rect 18598 10588 18604 10600
rect 18012 10560 18604 10588
rect 18012 10548 18018 10560
rect 18598 10548 18604 10560
rect 18656 10548 18662 10600
rect 18708 10588 18736 10628
rect 19058 10616 19064 10628
rect 19116 10616 19122 10668
rect 19702 10656 19708 10668
rect 19663 10628 19708 10656
rect 19702 10616 19708 10628
rect 19760 10616 19766 10668
rect 19153 10591 19211 10597
rect 19153 10588 19165 10591
rect 18708 10560 19165 10588
rect 19153 10557 19165 10560
rect 19199 10588 19211 10591
rect 19886 10588 19892 10600
rect 19199 10560 19892 10588
rect 19199 10557 19211 10560
rect 19153 10551 19211 10557
rect 19886 10548 19892 10560
rect 19944 10548 19950 10600
rect 19978 10548 19984 10600
rect 20036 10588 20042 10600
rect 22005 10591 22063 10597
rect 22005 10588 22017 10591
rect 20036 10560 22017 10588
rect 20036 10548 20042 10560
rect 22005 10557 22017 10560
rect 22051 10557 22063 10591
rect 22005 10551 22063 10557
rect 22281 10591 22339 10597
rect 22281 10557 22293 10591
rect 22327 10588 22339 10591
rect 24504 10588 24532 10696
rect 24946 10684 24952 10696
rect 25004 10684 25010 10736
rect 25130 10684 25136 10736
rect 25188 10724 25194 10736
rect 26605 10727 26663 10733
rect 25188 10696 25346 10724
rect 25188 10684 25194 10696
rect 26605 10693 26617 10727
rect 26651 10724 26663 10727
rect 27522 10724 27528 10736
rect 26651 10696 27528 10724
rect 26651 10693 26663 10696
rect 26605 10687 26663 10693
rect 27522 10684 27528 10696
rect 27580 10684 27586 10736
rect 28000 10733 28028 10764
rect 28902 10752 28908 10804
rect 28960 10792 28966 10804
rect 31202 10792 31208 10804
rect 28960 10764 30696 10792
rect 31115 10764 31208 10792
rect 28960 10752 28966 10764
rect 27985 10727 28043 10733
rect 27985 10693 27997 10727
rect 28031 10693 28043 10727
rect 27985 10687 28043 10693
rect 28994 10684 29000 10736
rect 29052 10684 29058 10736
rect 30668 10733 30696 10764
rect 31202 10752 31208 10764
rect 31260 10792 31266 10804
rect 37458 10792 37464 10804
rect 31260 10764 36308 10792
rect 37419 10764 37464 10792
rect 31260 10752 31266 10764
rect 30653 10727 30711 10733
rect 30653 10693 30665 10727
rect 30699 10724 30711 10727
rect 31294 10724 31300 10736
rect 30699 10696 31300 10724
rect 30699 10693 30711 10696
rect 30653 10687 30711 10693
rect 31294 10684 31300 10696
rect 31352 10684 31358 10736
rect 31404 10696 32904 10724
rect 27249 10659 27307 10665
rect 27249 10625 27261 10659
rect 27295 10656 27307 10659
rect 27430 10656 27436 10668
rect 27295 10628 27436 10656
rect 27295 10625 27307 10628
rect 27249 10619 27307 10625
rect 27430 10616 27436 10628
rect 27488 10616 27494 10668
rect 27706 10656 27712 10668
rect 27667 10628 27712 10656
rect 27706 10616 27712 10628
rect 27764 10616 27770 10668
rect 29638 10616 29644 10668
rect 29696 10656 29702 10668
rect 29733 10659 29791 10665
rect 29733 10656 29745 10659
rect 29696 10628 29745 10656
rect 29696 10616 29702 10628
rect 29733 10625 29745 10628
rect 29779 10656 29791 10659
rect 30282 10656 30288 10668
rect 29779 10628 30288 10656
rect 29779 10625 29791 10628
rect 29733 10619 29791 10625
rect 30282 10616 30288 10628
rect 30340 10616 30346 10668
rect 22327 10560 24532 10588
rect 24581 10591 24639 10597
rect 22327 10557 22339 10560
rect 22281 10551 22339 10557
rect 24581 10557 24593 10591
rect 24627 10557 24639 10591
rect 24854 10588 24860 10600
rect 24815 10560 24860 10588
rect 24581 10551 24639 10557
rect 16758 10520 16764 10532
rect 14108 10492 16764 10520
rect 16758 10480 16764 10492
rect 16816 10480 16822 10532
rect 17405 10523 17463 10529
rect 17405 10489 17417 10523
rect 17451 10520 17463 10523
rect 24486 10520 24492 10532
rect 17451 10492 22140 10520
rect 17451 10489 17463 10492
rect 17405 10483 17463 10489
rect 12986 10452 12992 10464
rect 12406 10424 12992 10452
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 13630 10412 13636 10464
rect 13688 10452 13694 10464
rect 15197 10455 15255 10461
rect 15197 10452 15209 10455
rect 13688 10424 15209 10452
rect 13688 10412 13694 10424
rect 15197 10421 15209 10424
rect 15243 10452 15255 10455
rect 18138 10452 18144 10464
rect 15243 10424 18144 10452
rect 15243 10421 15255 10424
rect 15197 10415 15255 10421
rect 18138 10412 18144 10424
rect 18196 10412 18202 10464
rect 18233 10455 18291 10461
rect 18233 10421 18245 10455
rect 18279 10452 18291 10455
rect 19242 10452 19248 10464
rect 18279 10424 19248 10452
rect 18279 10421 18291 10424
rect 18233 10415 18291 10421
rect 19242 10412 19248 10424
rect 19300 10412 19306 10464
rect 22112 10452 22140 10492
rect 23308 10492 24492 10520
rect 23308 10452 23336 10492
rect 24486 10480 24492 10492
rect 24544 10480 24550 10532
rect 23750 10452 23756 10464
rect 22112 10424 23336 10452
rect 23711 10424 23756 10452
rect 23750 10412 23756 10424
rect 23808 10412 23814 10464
rect 24596 10452 24624 10551
rect 24854 10548 24860 10560
rect 24912 10548 24918 10600
rect 24946 10548 24952 10600
rect 25004 10588 25010 10600
rect 31404 10588 31432 10696
rect 31757 10659 31815 10665
rect 31757 10625 31769 10659
rect 31803 10656 31815 10659
rect 31846 10656 31852 10668
rect 31803 10628 31852 10656
rect 31803 10625 31815 10628
rect 31757 10619 31815 10625
rect 31846 10616 31852 10628
rect 31904 10616 31910 10668
rect 31938 10616 31944 10668
rect 31996 10656 32002 10668
rect 32585 10659 32643 10665
rect 32585 10656 32597 10659
rect 31996 10628 32597 10656
rect 31996 10616 32002 10628
rect 32585 10625 32597 10628
rect 32631 10656 32643 10659
rect 32766 10656 32772 10668
rect 32631 10628 32772 10656
rect 32631 10625 32643 10628
rect 32585 10619 32643 10625
rect 32766 10616 32772 10628
rect 32824 10616 32830 10668
rect 25004 10560 31432 10588
rect 25004 10548 25010 10560
rect 31478 10548 31484 10600
rect 31536 10588 31542 10600
rect 32674 10588 32680 10600
rect 31536 10560 32680 10588
rect 31536 10548 31542 10560
rect 32674 10548 32680 10560
rect 32732 10548 32738 10600
rect 32876 10588 32904 10696
rect 33502 10684 33508 10736
rect 33560 10724 33566 10736
rect 33873 10727 33931 10733
rect 33873 10724 33885 10727
rect 33560 10696 33885 10724
rect 33560 10684 33566 10696
rect 33873 10693 33885 10696
rect 33919 10693 33931 10727
rect 33873 10687 33931 10693
rect 35529 10727 35587 10733
rect 35529 10693 35541 10727
rect 35575 10724 35587 10727
rect 35618 10724 35624 10736
rect 35575 10696 35624 10724
rect 35575 10693 35587 10696
rect 35529 10687 35587 10693
rect 35618 10684 35624 10696
rect 35676 10684 35682 10736
rect 33686 10656 33692 10668
rect 33647 10628 33692 10656
rect 33686 10616 33692 10628
rect 33744 10616 33750 10668
rect 36280 10665 36308 10764
rect 37458 10752 37464 10764
rect 37516 10752 37522 10804
rect 37550 10752 37556 10804
rect 37608 10792 37614 10804
rect 42061 10795 42119 10801
rect 37608 10764 42012 10792
rect 37608 10752 37614 10764
rect 40126 10724 40132 10736
rect 36464 10696 40132 10724
rect 36464 10665 36492 10696
rect 40126 10684 40132 10696
rect 40184 10684 40190 10736
rect 41138 10684 41144 10736
rect 41196 10724 41202 10736
rect 41325 10727 41383 10733
rect 41325 10724 41337 10727
rect 41196 10696 41337 10724
rect 41196 10684 41202 10696
rect 41325 10693 41337 10696
rect 41371 10693 41383 10727
rect 41598 10724 41604 10736
rect 41325 10687 41383 10693
rect 41524 10696 41604 10724
rect 36265 10659 36323 10665
rect 36265 10625 36277 10659
rect 36311 10625 36323 10659
rect 36265 10619 36323 10625
rect 36423 10659 36492 10665
rect 36423 10625 36435 10659
rect 36469 10628 36492 10659
rect 36630 10656 36636 10668
rect 36591 10628 36636 10656
rect 36469 10625 36481 10628
rect 36423 10619 36481 10625
rect 36630 10616 36636 10628
rect 36688 10616 36694 10668
rect 36909 10659 36967 10665
rect 36909 10625 36921 10659
rect 36955 10656 36967 10659
rect 37366 10656 37372 10668
rect 36955 10628 37372 10656
rect 36955 10625 36967 10628
rect 36909 10619 36967 10625
rect 37366 10616 37372 10628
rect 37424 10616 37430 10668
rect 38105 10659 38163 10665
rect 38105 10625 38117 10659
rect 38151 10656 38163 10659
rect 38194 10656 38200 10668
rect 38151 10628 38200 10656
rect 38151 10625 38163 10628
rect 38105 10619 38163 10625
rect 38194 10616 38200 10628
rect 38252 10616 38258 10668
rect 38286 10616 38292 10668
rect 38344 10656 38350 10668
rect 38746 10656 38752 10668
rect 38344 10628 38752 10656
rect 38344 10616 38350 10628
rect 38746 10616 38752 10628
rect 38804 10616 38810 10668
rect 38838 10616 38844 10668
rect 38896 10665 38902 10668
rect 38896 10659 38913 10665
rect 38901 10625 38913 10659
rect 40034 10656 40040 10668
rect 38896 10619 38913 10625
rect 39500 10628 40040 10656
rect 38896 10616 38902 10619
rect 34514 10588 34520 10600
rect 32876 10560 34520 10588
rect 34514 10548 34520 10560
rect 34572 10548 34578 10600
rect 35710 10548 35716 10600
rect 35768 10588 35774 10600
rect 39025 10591 39083 10597
rect 35768 10560 38700 10588
rect 35768 10548 35774 10560
rect 29730 10480 29736 10532
rect 29788 10520 29794 10532
rect 31846 10520 31852 10532
rect 29788 10492 31852 10520
rect 29788 10480 29794 10492
rect 31846 10480 31852 10492
rect 31904 10480 31910 10532
rect 32950 10520 32956 10532
rect 32911 10492 32956 10520
rect 32950 10480 32956 10492
rect 33008 10480 33014 10532
rect 33686 10480 33692 10532
rect 33744 10520 33750 10532
rect 36814 10520 36820 10532
rect 33744 10492 36820 10520
rect 33744 10480 33750 10492
rect 36814 10480 36820 10492
rect 36872 10480 36878 10532
rect 37090 10480 37096 10532
rect 37148 10520 37154 10532
rect 38565 10523 38623 10529
rect 38565 10520 38577 10523
rect 37148 10492 38577 10520
rect 37148 10480 37154 10492
rect 38565 10489 38577 10492
rect 38611 10489 38623 10523
rect 38672 10520 38700 10560
rect 39025 10557 39037 10591
rect 39071 10588 39083 10591
rect 39500 10588 39528 10628
rect 40034 10616 40040 10628
rect 40092 10616 40098 10668
rect 41524 10665 41552 10696
rect 41598 10684 41604 10696
rect 41656 10684 41662 10736
rect 41984 10724 42012 10764
rect 42061 10761 42073 10795
rect 42107 10792 42119 10795
rect 42518 10792 42524 10804
rect 42107 10764 42524 10792
rect 42107 10761 42119 10764
rect 42061 10755 42119 10761
rect 42518 10752 42524 10764
rect 42576 10752 42582 10804
rect 44266 10752 44272 10804
rect 44324 10792 44330 10804
rect 48314 10792 48320 10804
rect 44324 10764 45048 10792
rect 48275 10764 48320 10792
rect 44324 10752 44330 10764
rect 44910 10724 44916 10736
rect 41984 10696 44036 10724
rect 44871 10696 44916 10724
rect 41509 10659 41567 10665
rect 41509 10625 41521 10659
rect 41555 10625 41567 10659
rect 42426 10656 42432 10668
rect 41509 10619 41567 10625
rect 41616 10628 42432 10656
rect 39666 10588 39672 10600
rect 39071 10560 39528 10588
rect 39627 10560 39672 10588
rect 39071 10557 39083 10560
rect 39025 10551 39083 10557
rect 39666 10548 39672 10560
rect 39724 10548 39730 10600
rect 39758 10548 39764 10600
rect 39816 10588 39822 10600
rect 41616 10588 41644 10628
rect 42426 10616 42432 10628
rect 42484 10616 42490 10668
rect 42794 10656 42800 10668
rect 42755 10628 42800 10656
rect 42794 10616 42800 10628
rect 42852 10616 42858 10668
rect 44008 10665 44036 10696
rect 44910 10684 44916 10696
rect 44968 10684 44974 10736
rect 45020 10724 45048 10764
rect 48314 10752 48320 10764
rect 48372 10752 48378 10804
rect 50062 10792 50068 10804
rect 48516 10764 50068 10792
rect 48406 10724 48412 10736
rect 45020 10696 48412 10724
rect 48406 10684 48412 10696
rect 48464 10684 48470 10736
rect 48516 10668 48544 10764
rect 50062 10752 50068 10764
rect 50120 10752 50126 10804
rect 50154 10752 50160 10804
rect 50212 10792 50218 10804
rect 62482 10792 62488 10804
rect 50212 10764 62488 10792
rect 50212 10752 50218 10764
rect 62482 10752 62488 10764
rect 62540 10752 62546 10804
rect 62758 10752 62764 10804
rect 62816 10792 62822 10804
rect 69658 10792 69664 10804
rect 62816 10764 64828 10792
rect 62816 10752 62822 10764
rect 50798 10724 50804 10736
rect 48608 10696 50804 10724
rect 43993 10659 44051 10665
rect 43993 10625 44005 10659
rect 44039 10656 44051 10659
rect 44450 10656 44456 10668
rect 44039 10628 44456 10656
rect 44039 10625 44051 10628
rect 43993 10619 44051 10625
rect 44450 10616 44456 10628
rect 44508 10656 44514 10668
rect 44729 10659 44787 10665
rect 44729 10656 44741 10659
rect 44508 10628 44741 10656
rect 44508 10616 44514 10628
rect 44729 10625 44741 10628
rect 44775 10625 44787 10659
rect 48498 10656 48504 10668
rect 48411 10628 48504 10656
rect 44729 10619 44787 10625
rect 48498 10616 48504 10628
rect 48556 10616 48562 10668
rect 48608 10665 48636 10696
rect 50798 10684 50804 10696
rect 50856 10684 50862 10736
rect 54018 10724 54024 10736
rect 51934 10696 54024 10724
rect 54018 10684 54024 10696
rect 54076 10684 54082 10736
rect 54202 10724 54208 10736
rect 54163 10696 54208 10724
rect 54202 10684 54208 10696
rect 54260 10684 54266 10736
rect 54386 10684 54392 10736
rect 54444 10724 54450 10736
rect 55861 10727 55919 10733
rect 55861 10724 55873 10727
rect 54444 10696 55873 10724
rect 54444 10684 54450 10696
rect 55861 10693 55873 10696
rect 55907 10693 55919 10727
rect 56594 10724 56600 10736
rect 55861 10687 55919 10693
rect 55968 10696 56600 10724
rect 48593 10659 48651 10665
rect 48593 10625 48605 10659
rect 48639 10625 48651 10659
rect 48593 10619 48651 10625
rect 49513 10659 49571 10665
rect 49513 10625 49525 10659
rect 49559 10625 49571 10659
rect 49513 10619 49571 10625
rect 49605 10659 49663 10665
rect 49605 10625 49617 10659
rect 49651 10656 49663 10659
rect 49881 10659 49939 10665
rect 49651 10628 49832 10656
rect 49651 10625 49663 10628
rect 49605 10619 49663 10625
rect 39816 10560 41644 10588
rect 39816 10548 39822 10560
rect 41874 10548 41880 10600
rect 41932 10588 41938 10600
rect 42702 10588 42708 10600
rect 41932 10560 42708 10588
rect 41932 10548 41938 10560
rect 42702 10548 42708 10560
rect 42760 10548 42766 10600
rect 42886 10588 42892 10600
rect 42847 10560 42892 10588
rect 42886 10548 42892 10560
rect 42944 10548 42950 10600
rect 43165 10591 43223 10597
rect 43165 10557 43177 10591
rect 43211 10588 43223 10591
rect 43254 10588 43260 10600
rect 43211 10560 43260 10588
rect 43211 10557 43223 10560
rect 43165 10551 43223 10557
rect 43254 10548 43260 10560
rect 43312 10548 43318 10600
rect 43898 10588 43904 10600
rect 43859 10560 43904 10588
rect 43898 10548 43904 10560
rect 43956 10548 43962 10600
rect 45186 10588 45192 10600
rect 45147 10560 45192 10588
rect 45186 10548 45192 10560
rect 45244 10548 45250 10600
rect 47213 10591 47271 10597
rect 47213 10557 47225 10591
rect 47259 10588 47271 10591
rect 48869 10591 48927 10597
rect 48869 10588 48881 10591
rect 47259 10560 48881 10588
rect 47259 10557 47271 10560
rect 47213 10551 47271 10557
rect 48869 10557 48881 10560
rect 48915 10588 48927 10591
rect 49528 10588 49556 10619
rect 49694 10588 49700 10600
rect 48915 10560 49464 10588
rect 49528 10560 49700 10588
rect 48915 10557 48927 10560
rect 48869 10551 48927 10557
rect 43625 10523 43683 10529
rect 43625 10520 43637 10523
rect 38672 10492 43637 10520
rect 38565 10483 38623 10489
rect 43625 10489 43637 10492
rect 43671 10489 43683 10523
rect 43625 10483 43683 10489
rect 48774 10480 48780 10532
rect 48832 10520 48838 10532
rect 49436 10520 49464 10560
rect 49694 10548 49700 10560
rect 49752 10548 49758 10600
rect 49804 10588 49832 10628
rect 49881 10625 49893 10659
rect 49927 10656 49939 10659
rect 50338 10656 50344 10668
rect 49927 10628 50344 10656
rect 49927 10625 49939 10628
rect 49881 10619 49939 10625
rect 50338 10616 50344 10628
rect 50396 10616 50402 10668
rect 53193 10659 53251 10665
rect 53193 10625 53205 10659
rect 53239 10625 53251 10659
rect 53193 10619 53251 10625
rect 50430 10588 50436 10600
rect 49804 10560 50436 10588
rect 49804 10520 49832 10560
rect 50430 10548 50436 10560
rect 50488 10548 50494 10600
rect 50706 10588 50712 10600
rect 50667 10560 50712 10588
rect 50706 10548 50712 10560
rect 50764 10548 50770 10600
rect 53098 10548 53104 10600
rect 53156 10588 53162 10600
rect 53208 10588 53236 10619
rect 53282 10616 53288 10668
rect 53340 10656 53346 10668
rect 53466 10656 53472 10668
rect 53340 10628 53385 10656
rect 53427 10628 53472 10656
rect 53340 10616 53346 10628
rect 53466 10616 53472 10628
rect 53524 10616 53530 10668
rect 53558 10616 53564 10668
rect 53616 10656 53622 10668
rect 53653 10659 53711 10665
rect 53653 10656 53665 10659
rect 53616 10628 53665 10656
rect 53616 10616 53622 10628
rect 53653 10625 53665 10628
rect 53699 10625 53711 10659
rect 53653 10619 53711 10625
rect 53742 10616 53748 10668
rect 53800 10656 53806 10668
rect 54113 10659 54171 10665
rect 54113 10656 54125 10659
rect 53800 10628 54125 10656
rect 53800 10616 53806 10628
rect 54113 10625 54125 10628
rect 54159 10625 54171 10659
rect 54113 10619 54171 10625
rect 54297 10659 54355 10665
rect 54297 10625 54309 10659
rect 54343 10625 54355 10659
rect 54297 10619 54355 10625
rect 53156 10560 53512 10588
rect 53156 10548 53162 10560
rect 53009 10523 53067 10529
rect 53009 10520 53021 10523
rect 48832 10492 48877 10520
rect 49436 10492 49832 10520
rect 52012 10492 53021 10520
rect 48832 10480 48838 10492
rect 25866 10452 25872 10464
rect 24596 10424 25872 10452
rect 25866 10412 25872 10424
rect 25924 10412 25930 10464
rect 26694 10412 26700 10464
rect 26752 10452 26758 10464
rect 27522 10452 27528 10464
rect 26752 10424 27528 10452
rect 26752 10412 26758 10424
rect 27522 10412 27528 10424
rect 27580 10412 27586 10464
rect 28074 10412 28080 10464
rect 28132 10452 28138 10464
rect 31202 10452 31208 10464
rect 28132 10424 31208 10452
rect 28132 10412 28138 10424
rect 31202 10412 31208 10424
rect 31260 10412 31266 10464
rect 33042 10412 33048 10464
rect 33100 10452 33106 10464
rect 35710 10452 35716 10464
rect 33100 10424 35716 10452
rect 33100 10412 33106 10424
rect 35710 10412 35716 10424
rect 35768 10412 35774 10464
rect 36633 10455 36691 10461
rect 36633 10421 36645 10455
rect 36679 10452 36691 10455
rect 37274 10452 37280 10464
rect 36679 10424 37280 10452
rect 36679 10421 36691 10424
rect 36633 10415 36691 10421
rect 37274 10412 37280 10424
rect 37332 10412 37338 10464
rect 37366 10412 37372 10464
rect 37424 10452 37430 10464
rect 41874 10452 41880 10464
rect 37424 10424 41880 10452
rect 37424 10412 37430 10424
rect 41874 10412 41880 10424
rect 41932 10412 41938 10464
rect 41966 10412 41972 10464
rect 42024 10452 42030 10464
rect 45186 10452 45192 10464
rect 42024 10424 45192 10452
rect 42024 10412 42030 10424
rect 45186 10412 45192 10424
rect 45244 10412 45250 10464
rect 48314 10412 48320 10464
rect 48372 10452 48378 10464
rect 49329 10455 49387 10461
rect 49329 10452 49341 10455
rect 48372 10424 49341 10452
rect 48372 10412 48378 10424
rect 49329 10421 49341 10424
rect 49375 10421 49387 10455
rect 49329 10415 49387 10421
rect 49789 10455 49847 10461
rect 49789 10421 49801 10455
rect 49835 10452 49847 10455
rect 49878 10452 49884 10464
rect 49835 10424 49884 10452
rect 49835 10421 49847 10424
rect 49789 10415 49847 10421
rect 49878 10412 49884 10424
rect 49936 10412 49942 10464
rect 50062 10412 50068 10464
rect 50120 10452 50126 10464
rect 52012 10452 52040 10492
rect 53009 10489 53021 10492
rect 53055 10489 53067 10523
rect 53374 10520 53380 10532
rect 53335 10492 53380 10520
rect 53009 10483 53067 10489
rect 53374 10480 53380 10492
rect 53432 10480 53438 10532
rect 53484 10520 53512 10560
rect 54202 10520 54208 10532
rect 53484 10492 54208 10520
rect 54202 10480 54208 10492
rect 54260 10480 54266 10532
rect 54312 10520 54340 10619
rect 54478 10616 54484 10668
rect 54536 10656 54542 10668
rect 54938 10656 54944 10668
rect 54536 10628 54944 10656
rect 54536 10616 54542 10628
rect 54938 10616 54944 10628
rect 54996 10616 55002 10668
rect 55766 10656 55772 10668
rect 55727 10628 55772 10656
rect 55766 10616 55772 10628
rect 55824 10616 55830 10668
rect 55968 10665 55996 10696
rect 56594 10684 56600 10696
rect 56652 10724 56658 10736
rect 57790 10724 57796 10736
rect 56652 10696 57796 10724
rect 56652 10684 56658 10696
rect 57790 10684 57796 10696
rect 57848 10684 57854 10736
rect 58802 10684 58808 10736
rect 58860 10684 58866 10736
rect 59630 10684 59636 10736
rect 59688 10724 59694 10736
rect 61654 10724 61660 10736
rect 59688 10696 61660 10724
rect 59688 10684 59694 10696
rect 61654 10684 61660 10696
rect 61712 10724 61718 10736
rect 61712 10696 62436 10724
rect 61712 10684 61718 10696
rect 55953 10659 56011 10665
rect 55953 10625 55965 10659
rect 55999 10625 56011 10659
rect 56502 10656 56508 10668
rect 56463 10628 56508 10656
rect 55953 10619 56011 10625
rect 56502 10616 56508 10628
rect 56560 10616 56566 10668
rect 57330 10656 57336 10668
rect 57291 10628 57336 10656
rect 57330 10616 57336 10628
rect 57388 10616 57394 10668
rect 60737 10659 60795 10665
rect 60737 10625 60749 10659
rect 60783 10656 60795 10659
rect 62301 10659 62359 10665
rect 60783 10628 62252 10656
rect 60783 10625 60795 10628
rect 60737 10619 60795 10625
rect 54570 10548 54576 10600
rect 54628 10588 54634 10600
rect 54849 10591 54907 10597
rect 54849 10588 54861 10591
rect 54628 10560 54861 10588
rect 54628 10548 54634 10560
rect 54849 10557 54861 10560
rect 54895 10557 54907 10591
rect 54849 10551 54907 10557
rect 55490 10548 55496 10600
rect 55548 10588 55554 10600
rect 57422 10588 57428 10600
rect 55548 10560 57100 10588
rect 57383 10560 57428 10588
rect 55548 10548 55554 10560
rect 54312 10492 56272 10520
rect 52178 10452 52184 10464
rect 50120 10424 52040 10452
rect 52139 10424 52184 10452
rect 50120 10412 50126 10424
rect 52178 10412 52184 10424
rect 52236 10412 52242 10464
rect 52270 10412 52276 10464
rect 52328 10452 52334 10464
rect 54312 10452 54340 10492
rect 55306 10452 55312 10464
rect 52328 10424 54340 10452
rect 55267 10424 55312 10452
rect 52328 10412 52334 10424
rect 55306 10412 55312 10424
rect 55364 10412 55370 10464
rect 56244 10452 56272 10492
rect 56318 10480 56324 10532
rect 56376 10520 56382 10532
rect 56965 10523 57023 10529
rect 56965 10520 56977 10523
rect 56376 10492 56977 10520
rect 56376 10480 56382 10492
rect 56965 10489 56977 10492
rect 57011 10489 57023 10523
rect 57072 10520 57100 10560
rect 57422 10548 57428 10560
rect 57480 10548 57486 10600
rect 58069 10591 58127 10597
rect 58069 10557 58081 10591
rect 58115 10557 58127 10591
rect 58069 10551 58127 10557
rect 58345 10591 58403 10597
rect 58345 10557 58357 10591
rect 58391 10588 58403 10591
rect 60645 10591 60703 10597
rect 60645 10588 60657 10591
rect 58391 10560 60657 10588
rect 58391 10557 58403 10560
rect 58345 10551 58403 10557
rect 60645 10557 60657 10560
rect 60691 10557 60703 10591
rect 61562 10588 61568 10600
rect 61523 10560 61568 10588
rect 60645 10551 60703 10557
rect 58084 10520 58112 10551
rect 61562 10548 61568 10560
rect 61620 10548 61626 10600
rect 62114 10588 62120 10600
rect 62075 10560 62120 10588
rect 62114 10548 62120 10560
rect 62172 10548 62178 10600
rect 57072 10492 58112 10520
rect 59817 10523 59875 10529
rect 56965 10483 57023 10489
rect 59817 10489 59829 10523
rect 59863 10520 59875 10523
rect 61930 10520 61936 10532
rect 59863 10492 61936 10520
rect 59863 10489 59875 10492
rect 59817 10483 59875 10489
rect 61930 10480 61936 10492
rect 61988 10480 61994 10532
rect 62224 10520 62252 10628
rect 62301 10625 62313 10659
rect 62347 10625 62359 10659
rect 62408 10656 62436 10696
rect 62666 10684 62672 10736
rect 62724 10724 62730 10736
rect 62724 10696 63986 10724
rect 62724 10684 62730 10696
rect 63218 10656 63224 10668
rect 62408 10628 63224 10656
rect 62301 10619 62359 10625
rect 62316 10588 62344 10619
rect 63218 10616 63224 10628
rect 63276 10616 63282 10668
rect 64800 10656 64828 10764
rect 67192 10764 69664 10792
rect 65426 10724 65432 10736
rect 65387 10696 65432 10724
rect 65426 10684 65432 10696
rect 65484 10684 65490 10736
rect 67192 10733 67220 10764
rect 69658 10752 69664 10764
rect 69716 10792 69722 10804
rect 69716 10764 70624 10792
rect 69716 10752 69722 10764
rect 67177 10727 67235 10733
rect 67177 10693 67189 10727
rect 67223 10693 67235 10727
rect 68738 10724 68744 10736
rect 67177 10687 67235 10693
rect 67284 10696 68744 10724
rect 67284 10656 67312 10696
rect 68738 10684 68744 10696
rect 68796 10684 68802 10736
rect 70302 10724 70308 10736
rect 69874 10696 70308 10724
rect 70302 10684 70308 10696
rect 70360 10684 70366 10736
rect 70596 10733 70624 10764
rect 71038 10752 71044 10804
rect 71096 10792 71102 10804
rect 79502 10792 79508 10804
rect 71096 10764 79508 10792
rect 71096 10752 71102 10764
rect 79502 10752 79508 10764
rect 79560 10752 79566 10804
rect 80422 10792 80428 10804
rect 79612 10764 80428 10792
rect 70581 10727 70639 10733
rect 70581 10693 70593 10727
rect 70627 10693 70639 10727
rect 70581 10687 70639 10693
rect 70670 10684 70676 10736
rect 70728 10724 70734 10736
rect 72234 10724 72240 10736
rect 70728 10696 72240 10724
rect 70728 10684 70734 10696
rect 72234 10684 72240 10696
rect 72292 10684 72298 10736
rect 72329 10727 72387 10733
rect 72329 10693 72341 10727
rect 72375 10724 72387 10727
rect 73522 10724 73528 10736
rect 72375 10696 73528 10724
rect 72375 10693 72387 10696
rect 72329 10687 72387 10693
rect 73522 10684 73528 10696
rect 73580 10684 73586 10736
rect 76006 10684 76012 10736
rect 76064 10684 76070 10736
rect 79612 10733 79640 10764
rect 80422 10752 80428 10764
rect 80480 10752 80486 10804
rect 82262 10752 82268 10804
rect 82320 10792 82326 10804
rect 88429 10795 88487 10801
rect 88429 10792 88441 10795
rect 82320 10764 88441 10792
rect 82320 10752 82326 10764
rect 88429 10761 88441 10764
rect 88475 10761 88487 10795
rect 88429 10755 88487 10761
rect 91649 10795 91707 10801
rect 91649 10761 91661 10795
rect 91695 10792 91707 10795
rect 92106 10792 92112 10804
rect 91695 10764 92112 10792
rect 91695 10761 91707 10764
rect 91649 10755 91707 10761
rect 92106 10752 92112 10764
rect 92164 10752 92170 10804
rect 94222 10792 94228 10804
rect 94183 10764 94228 10792
rect 94222 10752 94228 10764
rect 94280 10752 94286 10804
rect 79597 10727 79655 10733
rect 79597 10693 79609 10727
rect 79643 10693 79655 10727
rect 81342 10724 81348 10736
rect 80822 10696 81348 10724
rect 79597 10687 79655 10693
rect 81342 10684 81348 10696
rect 81400 10684 81406 10736
rect 86129 10727 86187 10733
rect 82004 10696 86080 10724
rect 64800 10628 67312 10656
rect 67726 10616 67732 10668
rect 67784 10656 67790 10668
rect 67821 10659 67879 10665
rect 67821 10656 67833 10659
rect 67784 10628 67833 10656
rect 67784 10616 67790 10628
rect 67821 10625 67833 10628
rect 67867 10656 67879 10659
rect 68278 10656 68284 10668
rect 67867 10628 68284 10656
rect 67867 10625 67879 10628
rect 67821 10619 67879 10625
rect 68278 10616 68284 10628
rect 68336 10616 68342 10668
rect 71774 10656 71780 10668
rect 69860 10628 71780 10656
rect 62390 10588 62396 10600
rect 62316 10560 62396 10588
rect 62390 10548 62396 10560
rect 62448 10588 62454 10600
rect 64969 10591 65027 10597
rect 62448 10560 64552 10588
rect 62448 10548 62454 10560
rect 63126 10520 63132 10532
rect 62224 10492 63132 10520
rect 63126 10480 63132 10492
rect 63184 10480 63190 10532
rect 64524 10520 64552 10560
rect 64969 10557 64981 10591
rect 65015 10588 65027 10591
rect 67358 10588 67364 10600
rect 65015 10560 67364 10588
rect 65015 10557 65027 10560
rect 64969 10551 65027 10557
rect 67358 10548 67364 10560
rect 67416 10548 67422 10600
rect 68370 10588 68376 10600
rect 68331 10560 68376 10588
rect 68370 10548 68376 10560
rect 68428 10548 68434 10600
rect 68646 10588 68652 10600
rect 68607 10560 68652 10588
rect 68646 10548 68652 10560
rect 68704 10548 68710 10600
rect 68738 10548 68744 10600
rect 68796 10588 68802 10600
rect 69860 10588 69888 10628
rect 71774 10616 71780 10628
rect 71832 10656 71838 10668
rect 72973 10659 73031 10665
rect 72973 10656 72985 10659
rect 71832 10628 72985 10656
rect 71832 10616 71838 10628
rect 72973 10625 72985 10628
rect 73019 10625 73031 10659
rect 72973 10619 73031 10625
rect 73709 10659 73767 10665
rect 73709 10625 73721 10659
rect 73755 10656 73767 10659
rect 74074 10656 74080 10668
rect 73755 10628 74080 10656
rect 73755 10625 73767 10628
rect 73709 10619 73767 10625
rect 74074 10616 74080 10628
rect 74132 10616 74138 10668
rect 76742 10616 76748 10668
rect 76800 10656 76806 10668
rect 77110 10656 77116 10668
rect 76800 10628 77116 10656
rect 76800 10616 76806 10628
rect 77110 10616 77116 10628
rect 77168 10656 77174 10668
rect 77573 10659 77631 10665
rect 77573 10656 77585 10659
rect 77168 10628 77585 10656
rect 77168 10616 77174 10628
rect 77573 10625 77585 10628
rect 77619 10625 77631 10659
rect 77573 10619 77631 10625
rect 78490 10616 78496 10668
rect 78548 10656 78554 10668
rect 78677 10659 78735 10665
rect 78677 10656 78689 10659
rect 78548 10628 78689 10656
rect 78548 10616 78554 10628
rect 78677 10625 78689 10628
rect 78723 10625 78735 10659
rect 78677 10619 78735 10625
rect 78769 10659 78827 10665
rect 78769 10625 78781 10659
rect 78815 10656 78827 10659
rect 78858 10656 78864 10668
rect 78815 10628 78864 10656
rect 78815 10625 78827 10628
rect 78769 10619 78827 10625
rect 78858 10616 78864 10628
rect 78916 10616 78922 10668
rect 82004 10665 82032 10696
rect 81989 10659 82047 10665
rect 81989 10656 82001 10659
rect 81084 10628 82001 10656
rect 68796 10560 69888 10588
rect 68796 10548 68802 10560
rect 70394 10548 70400 10600
rect 70452 10588 70458 10600
rect 74442 10588 74448 10600
rect 70452 10560 74448 10588
rect 70452 10548 70458 10560
rect 74442 10548 74448 10560
rect 74500 10548 74506 10600
rect 75181 10591 75239 10597
rect 75181 10557 75193 10591
rect 75227 10557 75239 10591
rect 75181 10551 75239 10557
rect 75457 10591 75515 10597
rect 75457 10557 75469 10591
rect 75503 10588 75515 10591
rect 79321 10591 79379 10597
rect 75503 10560 78904 10588
rect 75503 10557 75515 10560
rect 75457 10551 75515 10557
rect 66070 10520 66076 10532
rect 64524 10492 66076 10520
rect 66070 10480 66076 10492
rect 66128 10480 66134 10532
rect 68388 10520 68416 10548
rect 66180 10492 68416 10520
rect 59078 10452 59084 10464
rect 56244 10424 59084 10452
rect 59078 10412 59084 10424
rect 59136 10412 59142 10464
rect 63310 10412 63316 10464
rect 63368 10452 63374 10464
rect 63478 10455 63536 10461
rect 63478 10452 63490 10455
rect 63368 10424 63490 10452
rect 63368 10412 63374 10424
rect 63478 10421 63490 10424
rect 63524 10421 63536 10455
rect 63478 10415 63536 10421
rect 63862 10412 63868 10464
rect 63920 10452 63926 10464
rect 66180 10452 66208 10492
rect 69658 10480 69664 10532
rect 69716 10520 69722 10532
rect 73522 10520 73528 10532
rect 69716 10492 73528 10520
rect 69716 10480 69722 10492
rect 73522 10480 73528 10492
rect 73580 10480 73586 10532
rect 63920 10424 66208 10452
rect 63920 10412 63926 10424
rect 67634 10412 67640 10464
rect 67692 10452 67698 10464
rect 67729 10455 67787 10461
rect 67729 10452 67741 10455
rect 67692 10424 67741 10452
rect 67692 10412 67698 10424
rect 67729 10421 67741 10424
rect 67775 10421 67787 10455
rect 67729 10415 67787 10421
rect 67818 10412 67824 10464
rect 67876 10452 67882 10464
rect 70121 10455 70179 10461
rect 70121 10452 70133 10455
rect 67876 10424 70133 10452
rect 67876 10412 67882 10424
rect 70121 10421 70133 10424
rect 70167 10421 70179 10455
rect 70121 10415 70179 10421
rect 70486 10412 70492 10464
rect 70544 10452 70550 10464
rect 72881 10455 72939 10461
rect 72881 10452 72893 10455
rect 70544 10424 72893 10452
rect 70544 10412 70550 10424
rect 72881 10421 72893 10424
rect 72927 10421 72939 10455
rect 72881 10415 72939 10421
rect 72970 10412 72976 10464
rect 73028 10452 73034 10464
rect 73617 10455 73675 10461
rect 73617 10452 73629 10455
rect 73028 10424 73629 10452
rect 73028 10412 73034 10424
rect 73617 10421 73629 10424
rect 73663 10421 73675 10455
rect 74166 10452 74172 10464
rect 74127 10424 74172 10452
rect 73617 10415 73675 10421
rect 74166 10412 74172 10424
rect 74224 10412 74230 10464
rect 75196 10452 75224 10551
rect 77938 10520 77944 10532
rect 76484 10492 77944 10520
rect 76484 10452 76512 10492
rect 77938 10480 77944 10492
rect 77996 10520 78002 10532
rect 78766 10520 78772 10532
rect 77996 10492 78772 10520
rect 77996 10480 78002 10492
rect 78766 10480 78772 10492
rect 78824 10480 78830 10532
rect 76926 10452 76932 10464
rect 75196 10424 76512 10452
rect 76887 10424 76932 10452
rect 76926 10412 76932 10424
rect 76984 10412 76990 10464
rect 77570 10412 77576 10464
rect 77628 10452 77634 10464
rect 77665 10455 77723 10461
rect 77665 10452 77677 10455
rect 77628 10424 77677 10452
rect 77628 10412 77634 10424
rect 77665 10421 77677 10424
rect 77711 10421 77723 10455
rect 78876 10452 78904 10560
rect 79321 10557 79333 10591
rect 79367 10588 79379 10591
rect 79594 10588 79600 10600
rect 79367 10560 79600 10588
rect 79367 10557 79379 10560
rect 79321 10551 79379 10557
rect 79594 10548 79600 10560
rect 79652 10548 79658 10600
rect 81084 10597 81112 10628
rect 81989 10625 82001 10628
rect 82035 10625 82047 10659
rect 82262 10656 82268 10668
rect 82223 10628 82268 10656
rect 81989 10619 82047 10625
rect 82262 10616 82268 10628
rect 82320 10616 82326 10668
rect 83277 10659 83335 10665
rect 83277 10625 83289 10659
rect 83323 10656 83335 10659
rect 83366 10656 83372 10668
rect 83323 10628 83372 10656
rect 83323 10625 83335 10628
rect 83277 10619 83335 10625
rect 83366 10616 83372 10628
rect 83424 10616 83430 10668
rect 83550 10616 83556 10668
rect 83608 10656 83614 10668
rect 83829 10659 83887 10665
rect 83829 10656 83841 10659
rect 83608 10628 83841 10656
rect 83608 10616 83614 10628
rect 83829 10625 83841 10628
rect 83875 10625 83887 10659
rect 83829 10619 83887 10625
rect 83921 10659 83979 10665
rect 83921 10625 83933 10659
rect 83967 10656 83979 10659
rect 83967 10628 84148 10656
rect 83967 10625 83979 10628
rect 83921 10619 83979 10625
rect 81069 10591 81127 10597
rect 81069 10557 81081 10591
rect 81115 10557 81127 10591
rect 81069 10551 81127 10557
rect 82633 10591 82691 10597
rect 82633 10557 82645 10591
rect 82679 10588 82691 10591
rect 84010 10588 84016 10600
rect 82679 10560 84016 10588
rect 82679 10557 82691 10560
rect 82633 10551 82691 10557
rect 84010 10548 84016 10560
rect 84068 10548 84074 10600
rect 84120 10588 84148 10628
rect 84194 10616 84200 10668
rect 84252 10656 84258 10668
rect 84654 10656 84660 10668
rect 84252 10628 84297 10656
rect 84615 10628 84660 10656
rect 84252 10616 84258 10628
rect 84654 10616 84660 10628
rect 84712 10616 84718 10668
rect 86052 10665 86080 10696
rect 86129 10693 86141 10727
rect 86175 10724 86187 10727
rect 86957 10727 87015 10733
rect 86957 10724 86969 10727
rect 86175 10696 86969 10724
rect 86175 10693 86187 10696
rect 86129 10687 86187 10693
rect 86957 10693 86969 10696
rect 87003 10693 87015 10727
rect 89073 10727 89131 10733
rect 89073 10724 89085 10727
rect 88182 10696 89085 10724
rect 86957 10687 87015 10693
rect 89073 10693 89085 10696
rect 89119 10693 89131 10727
rect 89073 10687 89131 10693
rect 89898 10684 89904 10736
rect 89956 10724 89962 10736
rect 90177 10727 90235 10733
rect 90177 10724 90189 10727
rect 89956 10696 90189 10724
rect 89956 10684 89962 10696
rect 90177 10693 90189 10696
rect 90223 10693 90235 10727
rect 90177 10687 90235 10693
rect 90634 10684 90640 10736
rect 90692 10684 90698 10736
rect 86037 10659 86095 10665
rect 86037 10625 86049 10659
rect 86083 10625 86095 10659
rect 86037 10619 86095 10625
rect 88978 10616 88984 10668
rect 89036 10656 89042 10668
rect 89162 10656 89168 10668
rect 89036 10628 89168 10656
rect 89036 10616 89042 10628
rect 89162 10616 89168 10628
rect 89220 10616 89226 10668
rect 92569 10659 92627 10665
rect 92569 10625 92581 10659
rect 92615 10656 92627 10659
rect 93302 10656 93308 10668
rect 92615 10628 93308 10656
rect 92615 10625 92627 10628
rect 92569 10619 92627 10625
rect 93302 10616 93308 10628
rect 93360 10616 93366 10668
rect 94130 10656 94136 10668
rect 94091 10628 94136 10656
rect 94130 10616 94136 10628
rect 94188 10616 94194 10668
rect 84286 10588 84292 10600
rect 84120 10560 84292 10588
rect 84286 10548 84292 10560
rect 84344 10588 84350 10600
rect 84562 10588 84568 10600
rect 84344 10560 84568 10588
rect 84344 10548 84350 10560
rect 84562 10548 84568 10560
rect 84620 10548 84626 10600
rect 86494 10548 86500 10600
rect 86552 10588 86558 10600
rect 86681 10591 86739 10597
rect 86681 10588 86693 10591
rect 86552 10560 86693 10588
rect 86552 10548 86558 10560
rect 86681 10557 86693 10560
rect 86727 10588 86739 10591
rect 89901 10591 89959 10597
rect 89901 10588 89913 10591
rect 86727 10560 89913 10588
rect 86727 10557 86739 10560
rect 86681 10551 86739 10557
rect 89901 10557 89913 10560
rect 89947 10588 89959 10591
rect 90726 10588 90732 10600
rect 89947 10560 90732 10588
rect 89947 10557 89959 10560
rect 89901 10551 89959 10557
rect 90726 10548 90732 10560
rect 90784 10548 90790 10600
rect 92474 10588 92480 10600
rect 92435 10560 92480 10588
rect 92474 10548 92480 10560
rect 92532 10548 92538 10600
rect 93210 10588 93216 10600
rect 93171 10560 93216 10588
rect 93210 10548 93216 10560
rect 93268 10548 93274 10600
rect 83185 10523 83243 10529
rect 83185 10520 83197 10523
rect 80992 10492 83197 10520
rect 80992 10452 81020 10492
rect 83185 10489 83197 10492
rect 83231 10489 83243 10523
rect 84838 10520 84844 10532
rect 83185 10483 83243 10489
rect 83292 10492 84844 10520
rect 78876 10424 81020 10452
rect 77665 10415 77723 10421
rect 82354 10412 82360 10464
rect 82412 10452 82418 10464
rect 83292 10452 83320 10492
rect 84838 10480 84844 10492
rect 84896 10480 84902 10532
rect 84746 10452 84752 10464
rect 82412 10424 83320 10452
rect 84707 10424 84752 10452
rect 82412 10412 82418 10424
rect 84746 10412 84752 10424
rect 84804 10412 84810 10464
rect 85298 10452 85304 10464
rect 85259 10424 85304 10452
rect 85298 10412 85304 10424
rect 85356 10412 85362 10464
rect 1104 10362 94852 10384
rect 1104 10310 12668 10362
rect 12720 10310 12732 10362
rect 12784 10310 12796 10362
rect 12848 10310 12860 10362
rect 12912 10310 12924 10362
rect 12976 10310 36105 10362
rect 36157 10310 36169 10362
rect 36221 10310 36233 10362
rect 36285 10310 36297 10362
rect 36349 10310 36361 10362
rect 36413 10310 59542 10362
rect 59594 10310 59606 10362
rect 59658 10310 59670 10362
rect 59722 10310 59734 10362
rect 59786 10310 59798 10362
rect 59850 10310 82979 10362
rect 83031 10310 83043 10362
rect 83095 10310 83107 10362
rect 83159 10310 83171 10362
rect 83223 10310 83235 10362
rect 83287 10310 94852 10362
rect 1104 10288 94852 10310
rect 1765 10251 1823 10257
rect 1765 10217 1777 10251
rect 1811 10248 1823 10251
rect 4522 10248 4528 10260
rect 1811 10220 4528 10248
rect 1811 10217 1823 10220
rect 1765 10211 1823 10217
rect 4522 10208 4528 10220
rect 4580 10208 4586 10260
rect 5074 10248 5080 10260
rect 4632 10220 5080 10248
rect 3418 10180 3424 10192
rect 3379 10152 3424 10180
rect 3418 10140 3424 10152
rect 3476 10140 3482 10192
rect 4062 10180 4068 10192
rect 4023 10152 4068 10180
rect 4062 10140 4068 10152
rect 4120 10140 4126 10192
rect 4522 10112 4528 10124
rect 4172 10084 4528 10112
rect 1578 10044 1584 10056
rect 1539 10016 1584 10044
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 2222 10044 2228 10056
rect 2183 10016 2228 10044
rect 2222 10004 2228 10016
rect 2280 10004 2286 10056
rect 2498 10044 2504 10056
rect 2459 10016 2504 10044
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10044 3295 10047
rect 3878 10044 3884 10056
rect 3283 10016 3884 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 4172 10053 4200 10084
rect 4522 10072 4528 10084
rect 4580 10112 4586 10124
rect 4632 10112 4660 10220
rect 5074 10208 5080 10220
rect 5132 10208 5138 10260
rect 11790 10248 11796 10260
rect 10796 10220 11796 10248
rect 4580 10084 4660 10112
rect 4893 10115 4951 10121
rect 4580 10072 4586 10084
rect 4893 10081 4905 10115
rect 4939 10112 4951 10115
rect 6638 10112 6644 10124
rect 4939 10084 6644 10112
rect 4939 10081 4951 10084
rect 4893 10075 4951 10081
rect 6638 10072 6644 10084
rect 6696 10072 6702 10124
rect 10796 10121 10824 10220
rect 11790 10208 11796 10220
rect 11848 10208 11854 10260
rect 18690 10248 18696 10260
rect 15948 10220 18696 10248
rect 10781 10115 10839 10121
rect 10781 10081 10793 10115
rect 10827 10081 10839 10115
rect 10781 10075 10839 10081
rect 12526 10072 12532 10124
rect 12584 10112 12590 10124
rect 13538 10112 13544 10124
rect 12584 10084 13544 10112
rect 12584 10072 12590 10084
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 15102 10112 15108 10124
rect 15063 10084 15108 10112
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10013 4031 10047
rect 3973 10007 4031 10013
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10013 4215 10047
rect 4614 10044 4620 10056
rect 4575 10016 4620 10044
rect 4157 10007 4215 10013
rect 3988 9920 4016 10007
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 5994 10004 6000 10056
rect 6052 10044 6058 10056
rect 7285 10047 7343 10053
rect 6052 10016 6868 10044
rect 6052 10004 6058 10016
rect 6641 9979 6699 9985
rect 6641 9945 6653 9979
rect 6687 9976 6699 9979
rect 6730 9976 6736 9988
rect 6687 9948 6736 9976
rect 6687 9945 6699 9948
rect 6641 9939 6699 9945
rect 6730 9936 6736 9948
rect 6788 9936 6794 9988
rect 6840 9976 6868 10016
rect 7285 10013 7297 10047
rect 7331 10044 7343 10047
rect 7650 10044 7656 10056
rect 7331 10016 7656 10044
rect 7331 10013 7343 10016
rect 7285 10007 7343 10013
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 8018 10044 8024 10056
rect 7979 10016 8024 10044
rect 8018 10004 8024 10016
rect 8076 10004 8082 10056
rect 8110 10004 8116 10056
rect 8168 10044 8174 10056
rect 8294 10044 8300 10056
rect 8168 10016 8300 10044
rect 8168 10004 8174 10016
rect 8294 10004 8300 10016
rect 8352 10004 8358 10056
rect 10873 10047 10931 10053
rect 10873 10013 10885 10047
rect 10919 10044 10931 10047
rect 11054 10044 11060 10056
rect 10919 10016 11060 10044
rect 10919 10013 10931 10016
rect 10873 10007 10931 10013
rect 11054 10004 11060 10016
rect 11112 10044 11118 10056
rect 11974 10044 11980 10056
rect 11112 10016 11980 10044
rect 11112 10004 11118 10016
rect 11974 10004 11980 10016
rect 12032 10004 12038 10056
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 15013 10047 15071 10053
rect 15013 10044 15025 10047
rect 13872 10016 15025 10044
rect 13872 10004 13878 10016
rect 15013 10013 15025 10016
rect 15059 10044 15071 10047
rect 15948 10044 15976 10220
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 18785 10251 18843 10257
rect 18785 10217 18797 10251
rect 18831 10248 18843 10251
rect 20714 10248 20720 10260
rect 18831 10220 20720 10248
rect 18831 10217 18843 10220
rect 18785 10211 18843 10217
rect 20714 10208 20720 10220
rect 20772 10208 20778 10260
rect 22554 10248 22560 10260
rect 22515 10220 22560 10248
rect 22554 10208 22560 10220
rect 22612 10208 22618 10260
rect 23750 10208 23756 10260
rect 23808 10248 23814 10260
rect 30374 10248 30380 10260
rect 23808 10220 30380 10248
rect 23808 10208 23814 10220
rect 30374 10208 30380 10220
rect 30432 10208 30438 10260
rect 32539 10251 32597 10257
rect 32539 10217 32551 10251
rect 32585 10248 32597 10251
rect 33686 10248 33692 10260
rect 32585 10220 33692 10248
rect 32585 10217 32597 10220
rect 32539 10211 32597 10217
rect 33686 10208 33692 10220
rect 33744 10208 33750 10260
rect 34330 10208 34336 10260
rect 34388 10248 34394 10260
rect 35158 10248 35164 10260
rect 34388 10220 35164 10248
rect 34388 10208 34394 10220
rect 35158 10208 35164 10220
rect 35216 10208 35222 10260
rect 36538 10248 36544 10260
rect 36499 10220 36544 10248
rect 36538 10208 36544 10220
rect 36596 10208 36602 10260
rect 41874 10248 41880 10260
rect 38304 10220 41880 10248
rect 18046 10140 18052 10192
rect 18104 10180 18110 10192
rect 19058 10180 19064 10192
rect 18104 10152 19064 10180
rect 18104 10140 18110 10152
rect 19058 10140 19064 10152
rect 19116 10180 19122 10192
rect 19429 10183 19487 10189
rect 19429 10180 19441 10183
rect 19116 10152 19441 10180
rect 19116 10140 19122 10152
rect 19429 10149 19441 10152
rect 19475 10149 19487 10183
rect 19429 10143 19487 10149
rect 26786 10140 26792 10192
rect 26844 10180 26850 10192
rect 29086 10180 29092 10192
rect 26844 10152 27660 10180
rect 29047 10152 29092 10180
rect 26844 10140 26850 10152
rect 17954 10072 17960 10124
rect 18012 10112 18018 10124
rect 18233 10115 18291 10121
rect 18233 10112 18245 10115
rect 18012 10084 18245 10112
rect 18012 10072 18018 10084
rect 18233 10081 18245 10084
rect 18279 10112 18291 10115
rect 19150 10112 19156 10124
rect 18279 10084 19156 10112
rect 18279 10081 18291 10084
rect 18233 10075 18291 10081
rect 19150 10072 19156 10084
rect 19208 10072 19214 10124
rect 19978 10112 19984 10124
rect 19939 10084 19984 10112
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 20257 10115 20315 10121
rect 20257 10081 20269 10115
rect 20303 10112 20315 10115
rect 22002 10112 22008 10124
rect 20303 10084 21496 10112
rect 21963 10084 22008 10112
rect 20303 10081 20315 10084
rect 20257 10075 20315 10081
rect 15059 10016 15976 10044
rect 17405 10047 17463 10053
rect 15059 10013 15071 10016
rect 15013 10007 15071 10013
rect 17405 10013 17417 10047
rect 17451 10044 17463 10047
rect 19702 10044 19708 10056
rect 17451 10016 19708 10044
rect 17451 10013 17463 10016
rect 17405 10007 17463 10013
rect 19702 10004 19708 10016
rect 19760 10004 19766 10056
rect 21468 10044 21496 10084
rect 22002 10072 22008 10084
rect 22060 10072 22066 10124
rect 25409 10115 25467 10121
rect 25409 10081 25421 10115
rect 25455 10112 25467 10115
rect 25774 10112 25780 10124
rect 25455 10084 25780 10112
rect 25455 10081 25467 10084
rect 25409 10075 25467 10081
rect 25774 10072 25780 10084
rect 25832 10072 25838 10124
rect 27632 10112 27660 10152
rect 29086 10140 29092 10152
rect 29144 10140 29150 10192
rect 33134 10180 33140 10192
rect 31726 10152 33140 10180
rect 29638 10112 29644 10124
rect 27632 10084 29644 10112
rect 29638 10072 29644 10084
rect 29696 10072 29702 10124
rect 30561 10115 30619 10121
rect 30561 10081 30573 10115
rect 30607 10112 30619 10115
rect 31726 10112 31754 10152
rect 33134 10140 33140 10152
rect 33192 10140 33198 10192
rect 35066 10140 35072 10192
rect 35124 10180 35130 10192
rect 36446 10180 36452 10192
rect 35124 10152 36452 10180
rect 35124 10140 35130 10152
rect 36446 10140 36452 10152
rect 36504 10140 36510 10192
rect 38197 10183 38255 10189
rect 38197 10180 38209 10183
rect 36556 10152 38209 10180
rect 30607 10084 31754 10112
rect 30607 10081 30619 10084
rect 30561 10075 30619 10081
rect 32490 10072 32496 10124
rect 32548 10112 32554 10124
rect 34333 10115 34391 10121
rect 34333 10112 34345 10115
rect 32548 10084 34345 10112
rect 32548 10072 32554 10084
rect 34333 10081 34345 10084
rect 34379 10081 34391 10115
rect 34333 10075 34391 10081
rect 35710 10072 35716 10124
rect 35768 10112 35774 10124
rect 36556 10112 36584 10152
rect 38197 10149 38209 10152
rect 38243 10149 38255 10183
rect 38197 10143 38255 10149
rect 35768 10084 36584 10112
rect 36909 10115 36967 10121
rect 35768 10072 35774 10084
rect 36909 10081 36921 10115
rect 36955 10112 36967 10115
rect 38304 10112 38332 10220
rect 41874 10208 41880 10220
rect 41932 10208 41938 10260
rect 41969 10251 42027 10257
rect 41969 10217 41981 10251
rect 42015 10248 42027 10251
rect 42058 10248 42064 10260
rect 42015 10220 42064 10248
rect 42015 10217 42027 10220
rect 41969 10211 42027 10217
rect 42058 10208 42064 10220
rect 42116 10208 42122 10260
rect 42797 10251 42855 10257
rect 42797 10217 42809 10251
rect 42843 10248 42855 10251
rect 43898 10248 43904 10260
rect 42843 10220 43904 10248
rect 42843 10217 42855 10220
rect 42797 10211 42855 10217
rect 43898 10208 43904 10220
rect 43956 10208 43962 10260
rect 44450 10248 44456 10260
rect 44411 10220 44456 10248
rect 44450 10208 44456 10220
rect 44508 10208 44514 10260
rect 47026 10248 47032 10260
rect 46987 10220 47032 10248
rect 47026 10208 47032 10220
rect 47084 10208 47090 10260
rect 47578 10208 47584 10260
rect 47636 10248 47642 10260
rect 48041 10251 48099 10257
rect 48041 10248 48053 10251
rect 47636 10220 48053 10248
rect 47636 10208 47642 10220
rect 48041 10217 48053 10220
rect 48087 10217 48099 10251
rect 48041 10211 48099 10217
rect 48593 10251 48651 10257
rect 48593 10217 48605 10251
rect 48639 10248 48651 10251
rect 49694 10248 49700 10260
rect 48639 10220 49700 10248
rect 48639 10217 48651 10220
rect 48593 10211 48651 10217
rect 49694 10208 49700 10220
rect 49752 10208 49758 10260
rect 49789 10251 49847 10257
rect 49789 10217 49801 10251
rect 49835 10248 49847 10251
rect 50706 10248 50712 10260
rect 49835 10220 50712 10248
rect 49835 10217 49847 10220
rect 49789 10211 49847 10217
rect 50706 10208 50712 10220
rect 50764 10208 50770 10260
rect 50798 10208 50804 10260
rect 50856 10248 50862 10260
rect 53282 10248 53288 10260
rect 50856 10220 53288 10248
rect 50856 10208 50862 10220
rect 53282 10208 53288 10220
rect 53340 10208 53346 10260
rect 53466 10248 53472 10260
rect 53427 10220 53472 10248
rect 53466 10208 53472 10220
rect 53524 10208 53530 10260
rect 53650 10208 53656 10260
rect 53708 10248 53714 10260
rect 53745 10251 53803 10257
rect 53745 10248 53757 10251
rect 53708 10220 53757 10248
rect 53708 10208 53714 10220
rect 53745 10217 53757 10220
rect 53791 10217 53803 10251
rect 53745 10211 53803 10217
rect 54018 10208 54024 10260
rect 54076 10248 54082 10260
rect 54389 10251 54447 10257
rect 54389 10248 54401 10251
rect 54076 10220 54401 10248
rect 54076 10208 54082 10220
rect 54389 10217 54401 10220
rect 54435 10217 54447 10251
rect 54389 10211 54447 10217
rect 54570 10208 54576 10260
rect 54628 10248 54634 10260
rect 54628 10220 57284 10248
rect 54628 10208 54634 10220
rect 40129 10183 40187 10189
rect 40129 10180 40141 10183
rect 38488 10152 40141 10180
rect 38488 10121 38516 10152
rect 40129 10149 40141 10152
rect 40175 10149 40187 10183
rect 40129 10143 40187 10149
rect 40218 10140 40224 10192
rect 40276 10180 40282 10192
rect 41782 10180 41788 10192
rect 40276 10152 41788 10180
rect 40276 10140 40282 10152
rect 41782 10140 41788 10152
rect 41840 10140 41846 10192
rect 42426 10140 42432 10192
rect 42484 10180 42490 10192
rect 42484 10152 42932 10180
rect 42484 10140 42490 10152
rect 42904 10121 42932 10152
rect 44910 10140 44916 10192
rect 44968 10180 44974 10192
rect 44968 10152 47348 10180
rect 44968 10140 44974 10152
rect 36955 10084 38332 10112
rect 38473 10115 38531 10121
rect 36955 10081 36967 10084
rect 36909 10075 36967 10081
rect 38473 10081 38485 10115
rect 38519 10081 38531 10115
rect 41233 10115 41291 10121
rect 38473 10075 38531 10081
rect 40037 10085 40095 10091
rect 22554 10044 22560 10056
rect 21468 10016 22560 10044
rect 22554 10004 22560 10016
rect 22612 10004 22618 10056
rect 22646 10004 22652 10056
rect 22704 10044 22710 10056
rect 27430 10044 27436 10056
rect 22704 10016 24992 10044
rect 27343 10016 27436 10044
rect 22704 10004 22710 10016
rect 8846 9976 8852 9988
rect 6840 9948 8852 9976
rect 8846 9936 8852 9948
rect 8904 9976 8910 9988
rect 13265 9979 13323 9985
rect 8904 9948 12098 9976
rect 8904 9936 8910 9948
rect 13265 9945 13277 9979
rect 13311 9945 13323 9979
rect 13265 9939 13323 9945
rect 3970 9868 3976 9920
rect 4028 9868 4034 9920
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7101 9911 7159 9917
rect 7101 9908 7113 9911
rect 6972 9880 7113 9908
rect 6972 9868 6978 9880
rect 7101 9877 7113 9880
rect 7147 9908 7159 9911
rect 7834 9908 7840 9920
rect 7147 9880 7840 9908
rect 7147 9877 7159 9880
rect 7101 9871 7159 9877
rect 7834 9868 7840 9880
rect 7892 9908 7898 9920
rect 8938 9908 8944 9920
rect 7892 9880 8944 9908
rect 7892 9868 7898 9880
rect 8938 9868 8944 9880
rect 8996 9868 9002 9920
rect 9217 9911 9275 9917
rect 9217 9877 9229 9911
rect 9263 9908 9275 9911
rect 9398 9908 9404 9920
rect 9263 9880 9404 9908
rect 9263 9877 9275 9880
rect 9217 9871 9275 9877
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 9766 9908 9772 9920
rect 9727 9880 9772 9908
rect 9766 9868 9772 9880
rect 9824 9868 9830 9920
rect 10502 9908 10508 9920
rect 10463 9880 10508 9908
rect 10502 9868 10508 9880
rect 10560 9868 10566 9920
rect 10962 9868 10968 9920
rect 11020 9908 11026 9920
rect 13280 9908 13308 9939
rect 13906 9936 13912 9988
rect 13964 9976 13970 9988
rect 15657 9979 15715 9985
rect 15657 9976 15669 9979
rect 13964 9948 15669 9976
rect 13964 9936 13970 9948
rect 15657 9945 15669 9948
rect 15703 9945 15715 9979
rect 15657 9939 15715 9945
rect 18046 9936 18052 9988
rect 18104 9976 18110 9988
rect 18417 9979 18475 9985
rect 18417 9976 18429 9979
rect 18104 9948 18429 9976
rect 18104 9936 18110 9948
rect 18417 9945 18429 9948
rect 18463 9945 18475 9979
rect 22462 9976 22468 9988
rect 21482 9948 22468 9976
rect 18417 9939 18475 9945
rect 22462 9936 22468 9948
rect 22520 9976 22526 9988
rect 22830 9976 22836 9988
rect 22520 9948 22836 9976
rect 22520 9936 22526 9948
rect 22830 9936 22836 9948
rect 22888 9936 22894 9988
rect 23937 9979 23995 9985
rect 23937 9945 23949 9979
rect 23983 9976 23995 9979
rect 24670 9976 24676 9988
rect 23983 9948 24676 9976
rect 23983 9945 23995 9948
rect 23937 9939 23995 9945
rect 24670 9936 24676 9948
rect 24728 9936 24734 9988
rect 24857 9979 24915 9985
rect 24857 9945 24869 9979
rect 24903 9945 24915 9979
rect 24964 9976 24992 10016
rect 27430 10004 27436 10016
rect 27488 10044 27494 10056
rect 29822 10044 29828 10056
rect 27488 10016 29828 10044
rect 27488 10004 27494 10016
rect 29822 10004 29828 10016
rect 29880 10004 29886 10056
rect 29914 10004 29920 10056
rect 29972 10044 29978 10056
rect 30193 10047 30251 10053
rect 30193 10044 30205 10047
rect 29972 10016 30205 10044
rect 29972 10004 29978 10016
rect 30193 10013 30205 10016
rect 30239 10013 30251 10047
rect 30193 10007 30251 10013
rect 31987 10047 32045 10053
rect 31987 10013 31999 10047
rect 32033 10044 32045 10047
rect 33134 10044 33140 10056
rect 32033 10016 33140 10044
rect 32033 10013 32045 10016
rect 31987 10007 32045 10013
rect 33134 10004 33140 10016
rect 33192 10004 33198 10056
rect 33965 10047 34023 10053
rect 33965 10013 33977 10047
rect 34011 10044 34023 10047
rect 36538 10044 36544 10056
rect 34011 10016 36544 10044
rect 34011 10013 34023 10016
rect 33965 10007 34023 10013
rect 36538 10004 36544 10016
rect 36596 10004 36602 10056
rect 36722 10004 36728 10056
rect 36780 10053 36786 10056
rect 36780 10047 36797 10053
rect 36785 10013 36797 10047
rect 38562 10044 38568 10056
rect 38523 10016 38568 10044
rect 36780 10007 36797 10013
rect 36780 10004 36786 10007
rect 38562 10004 38568 10016
rect 38620 10004 38626 10056
rect 39942 10044 39948 10056
rect 39316 10016 39948 10044
rect 25685 9979 25743 9985
rect 25685 9976 25697 9979
rect 24964 9948 25697 9976
rect 24857 9939 24915 9945
rect 25685 9945 25697 9948
rect 25731 9945 25743 9979
rect 25685 9939 25743 9945
rect 26068 9948 26174 9976
rect 11020 9880 13308 9908
rect 11020 9868 11026 9880
rect 13538 9868 13544 9920
rect 13596 9908 13602 9920
rect 14645 9911 14703 9917
rect 14645 9908 14657 9911
rect 13596 9880 14657 9908
rect 13596 9868 13602 9880
rect 14645 9877 14657 9880
rect 14691 9877 14703 9911
rect 14645 9871 14703 9877
rect 15378 9868 15384 9920
rect 15436 9908 15442 9920
rect 16390 9908 16396 9920
rect 15436 9880 16396 9908
rect 15436 9868 15442 9880
rect 16390 9868 16396 9880
rect 16448 9868 16454 9920
rect 18322 9868 18328 9920
rect 18380 9908 18386 9920
rect 18509 9911 18567 9917
rect 18509 9908 18521 9911
rect 18380 9880 18521 9908
rect 18380 9868 18386 9880
rect 18509 9877 18521 9880
rect 18555 9877 18567 9911
rect 18509 9871 18567 9877
rect 18598 9868 18604 9920
rect 18656 9908 18662 9920
rect 18656 9880 18701 9908
rect 18656 9868 18662 9880
rect 19058 9868 19064 9920
rect 19116 9908 19122 9920
rect 23109 9911 23167 9917
rect 23109 9908 23121 9911
rect 19116 9880 23121 9908
rect 19116 9868 19122 9880
rect 23109 9877 23121 9880
rect 23155 9908 23167 9911
rect 23382 9908 23388 9920
rect 23155 9880 23388 9908
rect 23155 9877 23167 9880
rect 23109 9871 23167 9877
rect 23382 9868 23388 9880
rect 23440 9868 23446 9920
rect 23845 9911 23903 9917
rect 23845 9877 23857 9911
rect 23891 9908 23903 9911
rect 24578 9908 24584 9920
rect 23891 9880 24584 9908
rect 23891 9877 23903 9880
rect 23845 9871 23903 9877
rect 24578 9868 24584 9880
rect 24636 9868 24642 9920
rect 24872 9908 24900 9939
rect 26068 9920 26096 9948
rect 27982 9936 27988 9988
rect 28040 9976 28046 9988
rect 32766 9976 32772 9988
rect 28040 9948 28085 9976
rect 31602 9948 32772 9976
rect 28040 9936 28046 9948
rect 32766 9936 32772 9948
rect 32824 9936 32830 9988
rect 33410 9936 33416 9988
rect 33468 9936 33474 9988
rect 34256 9948 35112 9976
rect 25314 9908 25320 9920
rect 24872 9880 25320 9908
rect 25314 9868 25320 9880
rect 25372 9868 25378 9920
rect 26050 9868 26056 9920
rect 26108 9908 26114 9920
rect 28077 9911 28135 9917
rect 28077 9908 28089 9911
rect 26108 9880 28089 9908
rect 26108 9868 26114 9880
rect 28077 9877 28089 9880
rect 28123 9908 28135 9911
rect 28994 9908 29000 9920
rect 28123 9880 29000 9908
rect 28123 9877 28135 9880
rect 28077 9871 28135 9877
rect 28994 9868 29000 9880
rect 29052 9868 29058 9920
rect 33134 9868 33140 9920
rect 33192 9908 33198 9920
rect 34256 9908 34284 9948
rect 33192 9880 34284 9908
rect 33192 9868 33198 9880
rect 34606 9868 34612 9920
rect 34664 9908 34670 9920
rect 34977 9911 35035 9917
rect 34977 9908 34989 9911
rect 34664 9880 34989 9908
rect 34664 9868 34670 9880
rect 34977 9877 34989 9880
rect 35023 9877 35035 9911
rect 35084 9908 35112 9948
rect 35158 9936 35164 9988
rect 35216 9976 35222 9988
rect 35253 9979 35311 9985
rect 35253 9976 35265 9979
rect 35216 9948 35265 9976
rect 35216 9936 35222 9948
rect 35253 9945 35265 9948
rect 35299 9945 35311 9979
rect 39316 9976 39344 10016
rect 39942 10004 39948 10016
rect 40000 10004 40006 10056
rect 40037 10051 40049 10085
rect 40083 10051 40095 10085
rect 41233 10081 41245 10115
rect 41279 10112 41291 10115
rect 42705 10115 42763 10121
rect 42705 10112 42717 10115
rect 41279 10084 42104 10112
rect 41279 10081 41291 10084
rect 41233 10075 41291 10081
rect 40037 10045 40095 10051
rect 40221 10047 40279 10053
rect 39758 9976 39764 9988
rect 35253 9939 35311 9945
rect 35360 9948 39344 9976
rect 39408 9948 39764 9976
rect 35360 9908 35388 9948
rect 35986 9908 35992 9920
rect 35084 9880 35388 9908
rect 35947 9880 35992 9908
rect 34977 9871 35035 9877
rect 35986 9868 35992 9880
rect 36044 9908 36050 9920
rect 37645 9911 37703 9917
rect 37645 9908 37657 9911
rect 36044 9880 37657 9908
rect 36044 9868 36050 9880
rect 37645 9877 37657 9880
rect 37691 9908 37703 9911
rect 39408 9908 39436 9948
rect 39758 9936 39764 9948
rect 39816 9976 39822 9988
rect 40052 9976 40080 10045
rect 40221 10013 40233 10047
rect 40267 10013 40279 10047
rect 40221 10007 40279 10013
rect 39816 9948 40080 9976
rect 39816 9936 39822 9948
rect 40236 9920 40264 10007
rect 40310 10004 40316 10056
rect 40368 10044 40374 10056
rect 41138 10044 41144 10056
rect 40368 10016 40413 10044
rect 41099 10016 41144 10044
rect 40368 10004 40374 10016
rect 41138 10004 41144 10016
rect 41196 10004 41202 10056
rect 41319 10047 41377 10053
rect 41319 10044 41331 10047
rect 41248 10016 41331 10044
rect 41248 9988 41276 10016
rect 41319 10013 41331 10016
rect 41365 10013 41377 10047
rect 41966 10044 41972 10056
rect 41319 10007 41377 10013
rect 41432 10016 41972 10044
rect 40586 9936 40592 9988
rect 40644 9976 40650 9988
rect 41230 9976 41236 9988
rect 40644 9948 41236 9976
rect 40644 9936 40650 9948
rect 41230 9936 41236 9948
rect 41288 9936 41294 9988
rect 37691 9880 39436 9908
rect 39485 9911 39543 9917
rect 37691 9877 37703 9880
rect 37645 9871 37703 9877
rect 39485 9877 39497 9911
rect 39531 9908 39543 9911
rect 39850 9908 39856 9920
rect 39531 9880 39856 9908
rect 39531 9877 39543 9880
rect 39485 9871 39543 9877
rect 39850 9868 39856 9880
rect 39908 9868 39914 9920
rect 40218 9868 40224 9920
rect 40276 9868 40282 9920
rect 40310 9868 40316 9920
rect 40368 9908 40374 9920
rect 41432 9908 41460 10016
rect 41966 10004 41972 10016
rect 42024 10004 42030 10056
rect 42076 10038 42104 10084
rect 42352 10084 42717 10112
rect 42352 10038 42380 10084
rect 42705 10081 42717 10084
rect 42751 10081 42763 10115
rect 42705 10075 42763 10081
rect 42889 10115 42947 10121
rect 42889 10081 42901 10115
rect 42935 10112 42947 10115
rect 43346 10112 43352 10124
rect 42935 10084 43352 10112
rect 42935 10081 42947 10084
rect 42889 10075 42947 10081
rect 43346 10072 43352 10084
rect 43404 10072 43410 10124
rect 44542 10112 44548 10124
rect 43548 10084 44548 10112
rect 43548 10056 43576 10084
rect 44542 10072 44548 10084
rect 44600 10072 44606 10124
rect 44726 10072 44732 10124
rect 44784 10112 44790 10124
rect 45833 10115 45891 10121
rect 44784 10084 45692 10112
rect 44784 10072 44790 10084
rect 42610 10044 42616 10056
rect 42076 10010 42380 10038
rect 42571 10016 42616 10044
rect 42610 10004 42616 10016
rect 42668 10004 42674 10056
rect 43530 10004 43536 10056
rect 43588 10044 43594 10056
rect 43806 10044 43812 10056
rect 43588 10016 43681 10044
rect 43767 10016 43812 10044
rect 43588 10004 43594 10016
rect 43806 10004 43812 10016
rect 43864 10004 43870 10056
rect 44358 10004 44364 10056
rect 44416 10044 44422 10056
rect 44453 10047 44511 10053
rect 44453 10044 44465 10047
rect 44416 10016 44465 10044
rect 44416 10004 44422 10016
rect 44453 10013 44465 10016
rect 44499 10013 44511 10047
rect 44453 10007 44511 10013
rect 44637 10047 44695 10053
rect 44637 10013 44649 10047
rect 44683 10044 44695 10047
rect 44818 10044 44824 10056
rect 44683 10016 44824 10044
rect 44683 10013 44695 10016
rect 44637 10007 44695 10013
rect 41782 9976 41788 9988
rect 41743 9948 41788 9976
rect 41782 9936 41788 9948
rect 41840 9936 41846 9988
rect 44468 9976 44496 10007
rect 44818 10004 44824 10016
rect 44876 10044 44882 10056
rect 45664 10053 45692 10084
rect 45833 10081 45845 10115
rect 45879 10112 45891 10115
rect 47213 10115 47271 10121
rect 47213 10112 47225 10115
rect 45879 10084 47225 10112
rect 45879 10081 45891 10084
rect 45833 10075 45891 10081
rect 47213 10081 47225 10084
rect 47259 10081 47271 10115
rect 47213 10075 47271 10081
rect 45373 10047 45431 10053
rect 45373 10044 45385 10047
rect 44876 10016 45385 10044
rect 44876 10004 44882 10016
rect 45373 10013 45385 10016
rect 45419 10013 45431 10047
rect 45373 10007 45431 10013
rect 45649 10047 45707 10053
rect 45649 10013 45661 10047
rect 45695 10044 45707 10047
rect 46106 10044 46112 10056
rect 45695 10016 46112 10044
rect 45695 10013 45707 10016
rect 45649 10007 45707 10013
rect 46106 10004 46112 10016
rect 46164 10004 46170 10056
rect 46290 10044 46296 10056
rect 46251 10016 46296 10044
rect 46290 10004 46296 10016
rect 46348 10004 46354 10056
rect 47320 10053 47348 10152
rect 48774 10140 48780 10192
rect 48832 10180 48838 10192
rect 49878 10180 49884 10192
rect 48832 10152 49884 10180
rect 48832 10140 48838 10152
rect 49878 10140 49884 10152
rect 49936 10180 49942 10192
rect 54754 10180 54760 10192
rect 49936 10152 54760 10180
rect 49936 10140 49942 10152
rect 54754 10140 54760 10152
rect 54812 10140 54818 10192
rect 54846 10140 54852 10192
rect 54904 10180 54910 10192
rect 56594 10180 56600 10192
rect 54904 10152 56600 10180
rect 54904 10140 54910 10152
rect 56594 10140 56600 10152
rect 56652 10140 56658 10192
rect 57256 10180 57284 10220
rect 57330 10208 57336 10260
rect 57388 10248 57394 10260
rect 59173 10251 59231 10257
rect 59173 10248 59185 10251
rect 57388 10220 59185 10248
rect 57388 10208 57394 10220
rect 59173 10217 59185 10220
rect 59219 10248 59231 10251
rect 60734 10248 60740 10260
rect 59219 10220 60740 10248
rect 59219 10217 59231 10220
rect 59173 10211 59231 10217
rect 60734 10208 60740 10220
rect 60792 10208 60798 10260
rect 62666 10248 62672 10260
rect 62627 10220 62672 10248
rect 62666 10208 62672 10220
rect 62724 10208 62730 10260
rect 63310 10248 63316 10260
rect 63271 10220 63316 10248
rect 63310 10208 63316 10220
rect 63368 10208 63374 10260
rect 67450 10248 67456 10260
rect 67411 10220 67456 10248
rect 67450 10208 67456 10220
rect 67508 10208 67514 10260
rect 68097 10251 68155 10257
rect 68097 10217 68109 10251
rect 68143 10248 68155 10251
rect 68646 10248 68652 10260
rect 68143 10220 68652 10248
rect 68143 10217 68155 10220
rect 68097 10211 68155 10217
rect 68646 10208 68652 10220
rect 68704 10208 68710 10260
rect 71682 10248 71688 10260
rect 68756 10220 71688 10248
rect 60366 10180 60372 10192
rect 57256 10152 60372 10180
rect 60366 10140 60372 10152
rect 60424 10140 60430 10192
rect 60458 10140 60464 10192
rect 60516 10180 60522 10192
rect 65426 10180 65432 10192
rect 60516 10152 65432 10180
rect 60516 10140 60522 10152
rect 65426 10140 65432 10152
rect 65484 10140 65490 10192
rect 67818 10180 67824 10192
rect 66088 10152 67824 10180
rect 48961 10115 49019 10121
rect 48961 10081 48973 10115
rect 49007 10112 49019 10115
rect 49602 10112 49608 10124
rect 49007 10084 49608 10112
rect 49007 10081 49019 10084
rect 48961 10075 49019 10081
rect 49602 10072 49608 10084
rect 49660 10112 49666 10124
rect 52270 10112 52276 10124
rect 49660 10084 52276 10112
rect 49660 10072 49666 10084
rect 52270 10072 52276 10084
rect 52328 10072 52334 10124
rect 53282 10072 53288 10124
rect 53340 10112 53346 10124
rect 53561 10115 53619 10121
rect 53561 10112 53573 10115
rect 53340 10084 53573 10112
rect 53340 10072 53346 10084
rect 53561 10081 53573 10084
rect 53607 10081 53619 10115
rect 53561 10075 53619 10081
rect 53650 10072 53656 10124
rect 53708 10112 53714 10124
rect 55769 10115 55827 10121
rect 55769 10112 55781 10115
rect 53708 10084 55781 10112
rect 53708 10072 53714 10084
rect 55769 10081 55781 10084
rect 55815 10081 55827 10115
rect 56962 10112 56968 10124
rect 56923 10084 56968 10112
rect 55769 10075 55827 10081
rect 56962 10072 56968 10084
rect 57020 10072 57026 10124
rect 59354 10112 59360 10124
rect 59315 10084 59360 10112
rect 59354 10072 59360 10084
rect 59412 10072 59418 10124
rect 62390 10112 62396 10124
rect 59464 10084 62396 10112
rect 46477 10047 46535 10053
rect 46477 10013 46489 10047
rect 46523 10013 46535 10047
rect 46477 10007 46535 10013
rect 47305 10047 47363 10053
rect 47305 10013 47317 10047
rect 47351 10013 47363 10047
rect 48774 10044 48780 10056
rect 48735 10016 48780 10044
rect 47305 10007 47363 10013
rect 44910 9976 44916 9988
rect 44468 9948 44916 9976
rect 44910 9936 44916 9948
rect 44968 9936 44974 9988
rect 45465 9979 45523 9985
rect 45465 9945 45477 9979
rect 45511 9976 45523 9979
rect 46385 9979 46443 9985
rect 46385 9976 46397 9979
rect 45511 9948 46397 9976
rect 45511 9945 45523 9948
rect 45465 9939 45523 9945
rect 46385 9945 46397 9948
rect 46431 9945 46443 9979
rect 46492 9976 46520 10007
rect 48774 10004 48780 10016
rect 48832 10004 48838 10056
rect 49053 10047 49111 10053
rect 49053 10013 49065 10047
rect 49099 10044 49111 10047
rect 49234 10044 49240 10056
rect 49099 10016 49240 10044
rect 49099 10013 49111 10016
rect 49053 10007 49111 10013
rect 49234 10004 49240 10016
rect 49292 10044 49298 10056
rect 49510 10044 49516 10056
rect 49292 10016 49516 10044
rect 49292 10004 49298 10016
rect 49510 10004 49516 10016
rect 49568 10004 49574 10056
rect 49786 10044 49792 10056
rect 49747 10016 49792 10044
rect 49786 10004 49792 10016
rect 49844 10004 49850 10056
rect 50246 10004 50252 10056
rect 50304 10044 50310 10056
rect 50341 10047 50399 10053
rect 50341 10044 50353 10047
rect 50304 10016 50353 10044
rect 50304 10004 50310 10016
rect 50341 10013 50353 10016
rect 50387 10013 50399 10047
rect 50341 10007 50399 10013
rect 52733 10047 52791 10053
rect 52733 10013 52745 10047
rect 52779 10044 52791 10047
rect 53374 10044 53380 10056
rect 52779 10016 53380 10044
rect 52779 10013 52791 10016
rect 52733 10007 52791 10013
rect 53374 10004 53380 10016
rect 53432 10004 53438 10056
rect 53469 10047 53527 10053
rect 53469 10013 53481 10047
rect 53515 10044 53527 10047
rect 53742 10044 53748 10056
rect 53515 10016 53748 10044
rect 53515 10013 53527 10016
rect 53469 10007 53527 10013
rect 46566 9976 46572 9988
rect 46492 9948 46572 9976
rect 46385 9939 46443 9945
rect 46566 9936 46572 9948
rect 46624 9936 46630 9988
rect 49418 9936 49424 9988
rect 49476 9976 49482 9988
rect 50798 9976 50804 9988
rect 49476 9948 50804 9976
rect 49476 9936 49482 9948
rect 50798 9936 50804 9948
rect 50856 9936 50862 9988
rect 50893 9979 50951 9985
rect 50893 9945 50905 9979
rect 50939 9976 50951 9979
rect 51258 9976 51264 9988
rect 50939 9948 51264 9976
rect 50939 9945 50951 9948
rect 50893 9939 50951 9945
rect 51258 9936 51264 9948
rect 51316 9936 51322 9988
rect 52546 9976 52552 9988
rect 52507 9948 52552 9976
rect 52546 9936 52552 9948
rect 52604 9936 52610 9988
rect 53006 9936 53012 9988
rect 53064 9976 53070 9988
rect 53484 9976 53512 10007
rect 53742 10004 53748 10016
rect 53800 10004 53806 10056
rect 53837 10047 53895 10053
rect 53837 10013 53849 10047
rect 53883 10013 53895 10047
rect 53837 10007 53895 10013
rect 54481 10047 54539 10053
rect 54481 10013 54493 10047
rect 54527 10044 54539 10047
rect 55674 10044 55680 10056
rect 54527 10016 55680 10044
rect 54527 10013 54539 10016
rect 54481 10007 54539 10013
rect 53064 9948 53512 9976
rect 53064 9936 53070 9948
rect 40368 9880 41460 9908
rect 40368 9868 40374 9880
rect 41966 9868 41972 9920
rect 42024 9917 42030 9920
rect 42024 9911 42043 9917
rect 42031 9877 42043 9911
rect 42024 9871 42043 9877
rect 42153 9911 42211 9917
rect 42153 9877 42165 9911
rect 42199 9908 42211 9911
rect 42610 9908 42616 9920
rect 42199 9880 42616 9908
rect 42199 9877 42211 9880
rect 42153 9871 42211 9877
rect 42024 9868 42030 9871
rect 42610 9868 42616 9880
rect 42668 9868 42674 9920
rect 42702 9868 42708 9920
rect 42760 9908 42766 9920
rect 43349 9911 43407 9917
rect 43349 9908 43361 9911
rect 42760 9880 43361 9908
rect 42760 9868 42766 9880
rect 43349 9877 43361 9880
rect 43395 9877 43407 9911
rect 43349 9871 43407 9877
rect 43717 9911 43775 9917
rect 43717 9877 43729 9911
rect 43763 9908 43775 9911
rect 43898 9908 43904 9920
rect 43763 9880 43904 9908
rect 43763 9877 43775 9880
rect 43717 9871 43775 9877
rect 43898 9868 43904 9880
rect 43956 9908 43962 9920
rect 44269 9911 44327 9917
rect 44269 9908 44281 9911
rect 43956 9880 44281 9908
rect 43956 9868 43962 9880
rect 44269 9877 44281 9880
rect 44315 9877 44327 9911
rect 44269 9871 44327 9877
rect 49326 9868 49332 9920
rect 49384 9908 49390 9920
rect 53852 9908 53880 10007
rect 55674 10004 55680 10016
rect 55732 10004 55738 10056
rect 55858 10044 55864 10056
rect 55819 10016 55864 10044
rect 55858 10004 55864 10016
rect 55916 10004 55922 10056
rect 56778 10044 56784 10056
rect 56739 10016 56784 10044
rect 56778 10004 56784 10016
rect 56836 10004 56842 10056
rect 59464 10053 59492 10084
rect 62390 10072 62396 10084
rect 62448 10072 62454 10124
rect 62482 10072 62488 10124
rect 62540 10112 62546 10124
rect 63402 10112 63408 10124
rect 62540 10084 63408 10112
rect 62540 10072 62546 10084
rect 63402 10072 63408 10084
rect 63460 10072 63466 10124
rect 66088 10112 66116 10152
rect 67818 10140 67824 10152
rect 67876 10140 67882 10192
rect 68756 10112 68784 10220
rect 71682 10208 71688 10220
rect 71740 10208 71746 10260
rect 72234 10208 72240 10260
rect 72292 10248 72298 10260
rect 74166 10248 74172 10260
rect 72292 10220 74172 10248
rect 72292 10208 72298 10220
rect 74166 10208 74172 10220
rect 74224 10208 74230 10260
rect 75457 10251 75515 10257
rect 75457 10217 75469 10251
rect 75503 10248 75515 10251
rect 75914 10248 75920 10260
rect 75503 10220 75920 10248
rect 75503 10217 75515 10220
rect 75457 10211 75515 10217
rect 75914 10208 75920 10220
rect 75972 10208 75978 10260
rect 77110 10248 77116 10260
rect 76208 10220 77116 10248
rect 69658 10112 69664 10124
rect 63512 10084 66116 10112
rect 66180 10084 68784 10112
rect 68848 10084 69664 10112
rect 59449 10047 59507 10053
rect 59449 10013 59461 10047
rect 59495 10013 59507 10047
rect 59449 10007 59507 10013
rect 60737 10047 60795 10053
rect 60737 10013 60749 10047
rect 60783 10013 60795 10047
rect 61102 10044 61108 10056
rect 61063 10016 61108 10044
rect 60737 10007 60795 10013
rect 58618 9976 58624 9988
rect 58579 9948 58624 9976
rect 58618 9936 58624 9948
rect 58676 9936 58682 9988
rect 58894 9936 58900 9988
rect 58952 9976 58958 9988
rect 60752 9976 60780 10007
rect 61102 10004 61108 10016
rect 61160 10004 61166 10056
rect 62577 10047 62635 10053
rect 62577 10044 62589 10047
rect 61672 10016 62589 10044
rect 58952 9948 60780 9976
rect 58952 9936 58958 9948
rect 54478 9908 54484 9920
rect 49384 9880 54484 9908
rect 49384 9868 49390 9880
rect 54478 9868 54484 9880
rect 54536 9908 54542 9920
rect 54846 9908 54852 9920
rect 54536 9880 54852 9908
rect 54536 9868 54542 9880
rect 54846 9868 54852 9880
rect 54904 9868 54910 9920
rect 55490 9908 55496 9920
rect 55451 9880 55496 9908
rect 55490 9868 55496 9880
rect 55548 9868 55554 9920
rect 57790 9868 57796 9920
rect 57848 9908 57854 9920
rect 60366 9908 60372 9920
rect 57848 9880 60372 9908
rect 57848 9868 57854 9880
rect 60366 9868 60372 9880
rect 60424 9868 60430 9920
rect 60458 9868 60464 9920
rect 60516 9908 60522 9920
rect 61672 9908 61700 10016
rect 62577 10013 62589 10016
rect 62623 10044 62635 10047
rect 62758 10044 62764 10056
rect 62623 10016 62764 10044
rect 62623 10013 62635 10016
rect 62577 10007 62635 10013
rect 62758 10004 62764 10016
rect 62816 10004 62822 10056
rect 63512 10053 63540 10084
rect 63497 10047 63555 10053
rect 63497 10013 63509 10047
rect 63543 10013 63555 10047
rect 63497 10007 63555 10013
rect 63678 10004 63684 10056
rect 63736 10044 63742 10056
rect 66180 10053 66208 10084
rect 64417 10047 64475 10053
rect 64417 10044 64429 10047
rect 63736 10016 64429 10044
rect 63736 10004 63742 10016
rect 64417 10013 64429 10016
rect 64463 10013 64475 10047
rect 64417 10007 64475 10013
rect 66165 10047 66223 10053
rect 66165 10013 66177 10047
rect 66211 10013 66223 10047
rect 66165 10007 66223 10013
rect 66533 10047 66591 10053
rect 66533 10013 66545 10047
rect 66579 10044 66591 10047
rect 66579 10016 66852 10044
rect 66579 10013 66591 10016
rect 66533 10007 66591 10013
rect 61749 9979 61807 9985
rect 61749 9945 61761 9979
rect 61795 9976 61807 9979
rect 64690 9976 64696 9988
rect 61795 9948 63632 9976
rect 64651 9948 64696 9976
rect 61795 9945 61807 9948
rect 61749 9939 61807 9945
rect 60516 9880 61700 9908
rect 60516 9868 60522 9880
rect 61930 9868 61936 9920
rect 61988 9908 61994 9920
rect 63494 9908 63500 9920
rect 61988 9880 63500 9908
rect 61988 9868 61994 9880
rect 63494 9868 63500 9880
rect 63552 9868 63558 9920
rect 63604 9908 63632 9948
rect 64690 9936 64696 9948
rect 64748 9936 64754 9988
rect 66622 9976 66628 9988
rect 65168 9948 66628 9976
rect 65168 9908 65196 9948
rect 66622 9936 66628 9948
rect 66680 9936 66686 9988
rect 63604 9880 65196 9908
rect 65245 9911 65303 9917
rect 65245 9877 65257 9911
rect 65291 9908 65303 9911
rect 65426 9908 65432 9920
rect 65291 9880 65432 9908
rect 65291 9877 65303 9880
rect 65245 9871 65303 9877
rect 65426 9868 65432 9880
rect 65484 9868 65490 9920
rect 66824 9908 66852 10016
rect 67358 10004 67364 10056
rect 67416 10044 67422 10056
rect 67913 10047 67971 10053
rect 67913 10044 67925 10047
rect 67416 10016 67925 10044
rect 67416 10004 67422 10016
rect 67913 10013 67925 10016
rect 67959 10013 67971 10047
rect 67913 10007 67971 10013
rect 68370 10004 68376 10056
rect 68428 10044 68434 10056
rect 68848 10044 68876 10084
rect 69658 10072 69664 10084
rect 69716 10072 69722 10124
rect 70118 10072 70124 10124
rect 70176 10112 70182 10124
rect 71225 10115 71283 10121
rect 71225 10112 71237 10115
rect 70176 10084 71237 10112
rect 70176 10072 70182 10084
rect 71225 10081 71237 10084
rect 71271 10081 71283 10115
rect 71225 10075 71283 10081
rect 71682 10072 71688 10124
rect 71740 10112 71746 10124
rect 72697 10115 72755 10121
rect 72697 10112 72709 10115
rect 71740 10084 72709 10112
rect 71740 10072 71746 10084
rect 72697 10081 72709 10084
rect 72743 10081 72755 10115
rect 76208 10112 76236 10220
rect 77110 10208 77116 10220
rect 77168 10208 77174 10260
rect 81342 10248 81348 10260
rect 81303 10220 81348 10248
rect 81342 10208 81348 10220
rect 81400 10208 81406 10260
rect 81989 10251 82047 10257
rect 81989 10217 82001 10251
rect 82035 10248 82047 10251
rect 85298 10248 85304 10260
rect 82035 10220 85304 10248
rect 82035 10217 82047 10220
rect 81989 10211 82047 10217
rect 78674 10140 78680 10192
rect 78732 10180 78738 10192
rect 82004 10180 82032 10211
rect 85298 10208 85304 10220
rect 85356 10208 85362 10260
rect 85390 10208 85396 10260
rect 85448 10248 85454 10260
rect 88613 10251 88671 10257
rect 88613 10248 88625 10251
rect 85448 10220 88625 10248
rect 85448 10208 85454 10220
rect 88613 10217 88625 10220
rect 88659 10217 88671 10251
rect 88613 10211 88671 10217
rect 89901 10251 89959 10257
rect 89901 10217 89913 10251
rect 89947 10248 89959 10251
rect 90634 10248 90640 10260
rect 89947 10220 90640 10248
rect 89947 10217 89959 10220
rect 89901 10211 89959 10217
rect 90634 10208 90640 10220
rect 90692 10208 90698 10260
rect 78732 10152 82032 10180
rect 78732 10140 78738 10152
rect 87874 10140 87880 10192
rect 87932 10180 87938 10192
rect 90453 10183 90511 10189
rect 90453 10180 90465 10183
rect 87932 10152 90465 10180
rect 87932 10140 87938 10152
rect 90453 10149 90465 10152
rect 90499 10149 90511 10183
rect 90453 10143 90511 10149
rect 72697 10075 72755 10081
rect 73172 10084 76236 10112
rect 76377 10115 76435 10121
rect 73172 10056 73200 10084
rect 76377 10081 76389 10115
rect 76423 10112 76435 10115
rect 79045 10115 79103 10121
rect 79045 10112 79057 10115
rect 76423 10084 79057 10112
rect 76423 10081 76435 10084
rect 76377 10075 76435 10081
rect 79045 10081 79057 10084
rect 79091 10081 79103 10115
rect 79778 10112 79784 10124
rect 79739 10084 79784 10112
rect 79045 10075 79103 10081
rect 79778 10072 79784 10084
rect 79836 10072 79842 10124
rect 80790 10072 80796 10124
rect 80848 10112 80854 10124
rect 81710 10112 81716 10124
rect 80848 10084 81716 10112
rect 80848 10072 80854 10084
rect 81710 10072 81716 10084
rect 81768 10072 81774 10124
rect 82449 10115 82507 10121
rect 82449 10081 82461 10115
rect 82495 10112 82507 10115
rect 83366 10112 83372 10124
rect 82495 10084 83372 10112
rect 82495 10081 82507 10084
rect 82449 10075 82507 10081
rect 83366 10072 83372 10084
rect 83424 10072 83430 10124
rect 83921 10115 83979 10121
rect 83921 10081 83933 10115
rect 83967 10112 83979 10115
rect 84746 10112 84752 10124
rect 83967 10084 84752 10112
rect 83967 10081 83979 10084
rect 83921 10075 83979 10081
rect 84746 10072 84752 10084
rect 84804 10072 84810 10124
rect 85482 10072 85488 10124
rect 85540 10112 85546 10124
rect 89165 10115 89223 10121
rect 89165 10112 89177 10115
rect 85540 10084 89177 10112
rect 85540 10072 85546 10084
rect 89165 10081 89177 10084
rect 89211 10081 89223 10115
rect 91557 10115 91615 10121
rect 91557 10112 91569 10115
rect 89165 10075 89223 10081
rect 89272 10084 91569 10112
rect 68428 10016 68876 10044
rect 70397 10047 70455 10053
rect 68428 10004 68434 10016
rect 70397 10013 70409 10047
rect 70443 10044 70455 10047
rect 70670 10044 70676 10056
rect 70443 10016 70676 10044
rect 70443 10013 70455 10016
rect 70397 10007 70455 10013
rect 70670 10004 70676 10016
rect 70728 10004 70734 10056
rect 70946 10044 70952 10056
rect 70907 10016 70952 10044
rect 70946 10004 70952 10016
rect 71004 10004 71010 10056
rect 72970 10044 72976 10056
rect 72358 10016 72976 10044
rect 72970 10004 72976 10016
rect 73028 10004 73034 10056
rect 73154 10044 73160 10056
rect 73115 10016 73160 10044
rect 73154 10004 73160 10016
rect 73212 10004 73218 10056
rect 75365 10047 75423 10053
rect 75365 10013 75377 10047
rect 75411 10044 75423 10047
rect 75914 10044 75920 10056
rect 75411 10016 75920 10044
rect 75411 10013 75423 10016
rect 75365 10007 75423 10013
rect 75914 10004 75920 10016
rect 75972 10004 75978 10056
rect 76098 10044 76104 10056
rect 76059 10016 76104 10044
rect 76098 10004 76104 10016
rect 76156 10004 76162 10056
rect 77662 10004 77668 10056
rect 77720 10044 77726 10056
rect 78309 10047 78367 10053
rect 78309 10044 78321 10047
rect 77720 10016 78321 10044
rect 77720 10004 77726 10016
rect 78309 10013 78321 10016
rect 78355 10013 78367 10047
rect 79134 10044 79140 10056
rect 79095 10016 79140 10044
rect 78309 10007 78367 10013
rect 79134 10004 79140 10016
rect 79192 10004 79198 10056
rect 79962 10053 79968 10056
rect 79951 10047 79968 10053
rect 79951 10013 79963 10047
rect 79951 10007 79968 10013
rect 79962 10004 79968 10007
rect 80020 10004 80026 10056
rect 81437 10047 81495 10053
rect 81437 10013 81449 10047
rect 81483 10044 81495 10047
rect 82354 10044 82360 10056
rect 81483 10016 82360 10044
rect 81483 10013 81495 10016
rect 81437 10007 81495 10013
rect 66901 9979 66959 9985
rect 66901 9945 66913 9979
rect 66947 9976 66959 9979
rect 68462 9976 68468 9988
rect 66947 9948 68468 9976
rect 66947 9945 66959 9948
rect 66901 9939 66959 9945
rect 68462 9936 68468 9948
rect 68520 9936 68526 9988
rect 70121 9979 70179 9985
rect 69690 9948 69796 9976
rect 68649 9911 68707 9917
rect 68649 9908 68661 9911
rect 66824 9880 68661 9908
rect 68649 9877 68661 9880
rect 68695 9908 68707 9911
rect 68830 9908 68836 9920
rect 68695 9880 68836 9908
rect 68695 9877 68707 9880
rect 68649 9871 68707 9877
rect 68830 9868 68836 9880
rect 68888 9868 68894 9920
rect 69768 9908 69796 9948
rect 70121 9945 70133 9979
rect 70167 9976 70179 9979
rect 70854 9976 70860 9988
rect 70167 9948 70860 9976
rect 70167 9945 70179 9948
rect 70121 9939 70179 9945
rect 70854 9936 70860 9948
rect 70912 9936 70918 9988
rect 73430 9976 73436 9988
rect 73391 9948 73436 9976
rect 73430 9936 73436 9948
rect 73488 9936 73494 9988
rect 75270 9976 75276 9988
rect 74658 9948 75276 9976
rect 75270 9936 75276 9948
rect 75328 9936 75334 9988
rect 71590 9908 71596 9920
rect 69768 9880 71596 9908
rect 71590 9868 71596 9880
rect 71648 9868 71654 9920
rect 74810 9868 74816 9920
rect 74868 9908 74874 9920
rect 74905 9911 74963 9917
rect 74905 9908 74917 9911
rect 74868 9880 74917 9908
rect 74868 9868 74874 9880
rect 74905 9877 74917 9880
rect 74951 9877 74963 9911
rect 76116 9908 76144 10004
rect 77386 9936 77392 9988
rect 77444 9936 77450 9988
rect 77754 9936 77760 9988
rect 77812 9976 77818 9988
rect 81452 9976 81480 10007
rect 82354 10004 82360 10016
rect 82412 10004 82418 10056
rect 84194 10004 84200 10056
rect 84252 10044 84258 10056
rect 84838 10044 84844 10056
rect 84252 10016 84297 10044
rect 84799 10016 84844 10044
rect 84252 10004 84258 10016
rect 84838 10004 84844 10016
rect 84896 10004 84902 10056
rect 85758 10044 85764 10056
rect 85719 10016 85764 10044
rect 85758 10004 85764 10016
rect 85816 10004 85822 10056
rect 86402 10044 86408 10056
rect 86363 10016 86408 10044
rect 86402 10004 86408 10016
rect 86460 10004 86466 10056
rect 87782 10004 87788 10056
rect 87840 10004 87846 10056
rect 88518 10004 88524 10056
rect 88576 10044 88582 10056
rect 89272 10044 89300 10084
rect 91557 10081 91569 10084
rect 91603 10081 91615 10115
rect 91557 10075 91615 10081
rect 93305 10115 93363 10121
rect 93305 10081 93317 10115
rect 93351 10112 93363 10115
rect 93854 10112 93860 10124
rect 93351 10084 93860 10112
rect 93351 10081 93363 10084
rect 93305 10075 93363 10081
rect 93854 10072 93860 10084
rect 93912 10072 93918 10124
rect 89806 10044 89812 10056
rect 88576 10016 89300 10044
rect 89767 10016 89812 10044
rect 88576 10004 88582 10016
rect 89806 10004 89812 10016
rect 89864 10044 89870 10056
rect 90450 10044 90456 10056
rect 89864 10016 90456 10044
rect 89864 10004 89870 10016
rect 90450 10004 90456 10016
rect 90508 10004 90514 10056
rect 93949 10047 94007 10053
rect 93949 10013 93961 10047
rect 93995 10044 94007 10047
rect 94130 10044 94136 10056
rect 93995 10016 94136 10044
rect 93995 10013 94007 10016
rect 93949 10007 94007 10013
rect 94130 10004 94136 10016
rect 94188 10004 94194 10056
rect 83826 9976 83832 9988
rect 77812 9948 81480 9976
rect 83490 9948 83832 9976
rect 77812 9936 77818 9948
rect 83826 9936 83832 9948
rect 83884 9936 83890 9988
rect 85853 9979 85911 9985
rect 85853 9945 85865 9979
rect 85899 9976 85911 9979
rect 86681 9979 86739 9985
rect 86681 9976 86693 9979
rect 85899 9948 86693 9976
rect 85899 9945 85911 9948
rect 85853 9939 85911 9945
rect 86681 9945 86693 9948
rect 86727 9945 86739 9979
rect 86681 9939 86739 9945
rect 90637 9979 90695 9985
rect 90637 9945 90649 9979
rect 90683 9976 90695 9979
rect 90726 9976 90732 9988
rect 90683 9948 90732 9976
rect 90683 9945 90695 9948
rect 90637 9939 90695 9945
rect 90726 9936 90732 9948
rect 90784 9936 90790 9988
rect 91094 9936 91100 9988
rect 91152 9976 91158 9988
rect 91833 9979 91891 9985
rect 91833 9976 91845 9979
rect 91152 9948 91845 9976
rect 91152 9936 91158 9948
rect 91833 9945 91845 9948
rect 91879 9945 91891 9979
rect 94222 9976 94228 9988
rect 93058 9948 94228 9976
rect 91833 9939 91891 9945
rect 94222 9936 94228 9948
rect 94280 9936 94286 9988
rect 77662 9908 77668 9920
rect 76116 9880 77668 9908
rect 74905 9871 74963 9877
rect 77662 9868 77668 9880
rect 77720 9868 77726 9920
rect 77849 9911 77907 9917
rect 77849 9877 77861 9911
rect 77895 9908 77907 9911
rect 78122 9908 78128 9920
rect 77895 9880 78128 9908
rect 77895 9877 77907 9880
rect 77849 9871 77907 9877
rect 78122 9868 78128 9880
rect 78180 9868 78186 9920
rect 78401 9911 78459 9917
rect 78401 9877 78413 9911
rect 78447 9908 78459 9911
rect 79042 9908 79048 9920
rect 78447 9880 79048 9908
rect 78447 9877 78459 9880
rect 78401 9871 78459 9877
rect 79042 9868 79048 9880
rect 79100 9908 79106 9920
rect 79410 9908 79416 9920
rect 79100 9880 79416 9908
rect 79100 9868 79106 9880
rect 79410 9868 79416 9880
rect 79468 9868 79474 9920
rect 80238 9908 80244 9920
rect 80199 9880 80244 9908
rect 80238 9868 80244 9880
rect 80296 9868 80302 9920
rect 84746 9908 84752 9920
rect 84707 9880 84752 9908
rect 84746 9868 84752 9880
rect 84804 9868 84810 9920
rect 87690 9868 87696 9920
rect 87748 9908 87754 9920
rect 88153 9911 88211 9917
rect 88153 9908 88165 9911
rect 87748 9880 88165 9908
rect 87748 9868 87754 9880
rect 88153 9877 88165 9880
rect 88199 9877 88211 9911
rect 88153 9871 88211 9877
rect 93762 9868 93768 9920
rect 93820 9908 93826 9920
rect 93857 9911 93915 9917
rect 93857 9908 93869 9911
rect 93820 9880 93869 9908
rect 93820 9868 93826 9880
rect 93857 9877 93869 9880
rect 93903 9877 93915 9911
rect 93857 9871 93915 9877
rect 1104 9818 95011 9840
rect 1104 9766 24386 9818
rect 24438 9766 24450 9818
rect 24502 9766 24514 9818
rect 24566 9766 24578 9818
rect 24630 9766 24642 9818
rect 24694 9766 47823 9818
rect 47875 9766 47887 9818
rect 47939 9766 47951 9818
rect 48003 9766 48015 9818
rect 48067 9766 48079 9818
rect 48131 9766 71260 9818
rect 71312 9766 71324 9818
rect 71376 9766 71388 9818
rect 71440 9766 71452 9818
rect 71504 9766 71516 9818
rect 71568 9766 94697 9818
rect 94749 9766 94761 9818
rect 94813 9766 94825 9818
rect 94877 9766 94889 9818
rect 94941 9766 94953 9818
rect 95005 9766 95011 9818
rect 1104 9744 95011 9766
rect 4798 9664 4804 9716
rect 4856 9704 4862 9716
rect 14918 9704 14924 9716
rect 4856 9676 14924 9704
rect 4856 9664 4862 9676
rect 14918 9664 14924 9676
rect 14976 9664 14982 9716
rect 17862 9704 17868 9716
rect 17823 9676 17868 9704
rect 17862 9664 17868 9676
rect 17920 9664 17926 9716
rect 18414 9664 18420 9716
rect 18472 9704 18478 9716
rect 20714 9704 20720 9716
rect 18472 9676 19380 9704
rect 18472 9664 18478 9676
rect 2314 9596 2320 9648
rect 2372 9636 2378 9648
rect 4614 9636 4620 9648
rect 2372 9608 4620 9636
rect 2372 9596 2378 9608
rect 2130 9568 2136 9580
rect 2091 9540 2136 9568
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 2608 9577 2636 9608
rect 4614 9596 4620 9608
rect 4672 9636 4678 9648
rect 7466 9636 7472 9648
rect 4672 9608 7472 9636
rect 4672 9596 4678 9608
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9537 2651 9571
rect 2593 9531 2651 9537
rect 2869 9571 2927 9577
rect 2869 9537 2881 9571
rect 2915 9568 2927 9571
rect 3605 9571 3663 9577
rect 2915 9540 3556 9568
rect 2915 9537 2927 9540
rect 2869 9531 2927 9537
rect 3528 9500 3556 9540
rect 3605 9537 3617 9571
rect 3651 9568 3663 9571
rect 3878 9568 3884 9580
rect 3651 9540 3884 9568
rect 3651 9537 3663 9540
rect 3605 9531 3663 9537
rect 3878 9528 3884 9540
rect 3936 9528 3942 9580
rect 4338 9568 4344 9580
rect 4251 9540 4344 9568
rect 4338 9528 4344 9540
rect 4396 9568 4402 9580
rect 5077 9571 5135 9577
rect 5077 9568 5089 9571
rect 4396 9540 5089 9568
rect 4396 9528 4402 9540
rect 5077 9537 5089 9540
rect 5123 9568 5135 9571
rect 5442 9568 5448 9580
rect 5123 9540 5448 9568
rect 5123 9537 5135 9540
rect 5077 9531 5135 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5810 9568 5816 9580
rect 5771 9540 5816 9568
rect 5810 9528 5816 9540
rect 5868 9528 5874 9580
rect 6748 9578 6776 9608
rect 7466 9596 7472 9608
rect 7524 9596 7530 9648
rect 8018 9636 8024 9648
rect 7576 9608 8024 9636
rect 7098 9578 7104 9580
rect 6656 9577 6776 9578
rect 6932 9577 7104 9578
rect 6641 9571 6776 9577
rect 6641 9537 6653 9571
rect 6687 9550 6776 9571
rect 6917 9571 7104 9577
rect 6687 9537 6699 9550
rect 6641 9531 6699 9537
rect 6917 9537 6929 9571
rect 6963 9550 7104 9571
rect 6963 9537 6975 9550
rect 6917 9531 6975 9537
rect 7098 9528 7104 9550
rect 7156 9578 7162 9580
rect 7156 9568 7420 9578
rect 7576 9568 7604 9608
rect 8018 9596 8024 9608
rect 8076 9596 8082 9648
rect 9493 9639 9551 9645
rect 9493 9636 9505 9639
rect 8128 9608 9505 9636
rect 7156 9550 7604 9568
rect 7156 9528 7162 9550
rect 7392 9540 7604 9550
rect 7650 9528 7656 9580
rect 7708 9568 7714 9580
rect 8128 9568 8156 9608
rect 9493 9605 9505 9608
rect 9539 9605 9551 9639
rect 9493 9599 9551 9605
rect 11149 9639 11207 9645
rect 11149 9605 11161 9639
rect 11195 9636 11207 9639
rect 11238 9636 11244 9648
rect 11195 9608 11244 9636
rect 11195 9605 11207 9608
rect 11149 9599 11207 9605
rect 11238 9596 11244 9608
rect 11296 9596 11302 9648
rect 12621 9639 12679 9645
rect 11348 9608 12434 9636
rect 7708 9540 7801 9568
rect 7944 9540 8156 9568
rect 8573 9571 8631 9577
rect 7708 9528 7714 9540
rect 4356 9500 4384 9528
rect 3528 9472 4384 9500
rect 4614 9460 4620 9512
rect 4672 9500 4678 9512
rect 4801 9503 4859 9509
rect 4801 9500 4813 9503
rect 4672 9472 4813 9500
rect 4672 9460 4678 9472
rect 4801 9469 4813 9472
rect 4847 9469 4859 9503
rect 7668 9500 7696 9528
rect 7944 9500 7972 9540
rect 8573 9537 8585 9571
rect 8619 9568 8631 9571
rect 9214 9568 9220 9580
rect 8619 9540 9220 9568
rect 8619 9537 8631 9540
rect 8573 9531 8631 9537
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9568 9367 9571
rect 10042 9568 10048 9580
rect 9355 9540 10048 9568
rect 9355 9537 9367 9540
rect 9309 9531 9367 9537
rect 8294 9500 8300 9512
rect 7668 9472 7788 9500
rect 4801 9463 4859 9469
rect 3789 9435 3847 9441
rect 3789 9401 3801 9435
rect 3835 9401 3847 9435
rect 3789 9395 3847 9401
rect 1949 9367 2007 9373
rect 1949 9333 1961 9367
rect 1995 9364 2007 9367
rect 3234 9364 3240 9376
rect 1995 9336 3240 9364
rect 1995 9333 2007 9336
rect 1949 9327 2007 9333
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 3804 9364 3832 9395
rect 5997 9367 6055 9373
rect 5997 9364 6009 9367
rect 3476 9336 6009 9364
rect 3476 9324 3482 9336
rect 5997 9333 6009 9336
rect 6043 9364 6055 9367
rect 6914 9364 6920 9376
rect 6043 9336 6920 9364
rect 6043 9333 6055 9336
rect 5997 9327 6055 9333
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 7006 9324 7012 9376
rect 7064 9364 7070 9376
rect 7760 9364 7788 9472
rect 7852 9472 7972 9500
rect 8255 9472 8300 9500
rect 7852 9444 7880 9472
rect 8294 9460 8300 9472
rect 8352 9460 8358 9512
rect 7834 9392 7840 9444
rect 7892 9432 7898 9444
rect 7892 9404 7937 9432
rect 7892 9392 7898 9404
rect 9324 9364 9352 9531
rect 10042 9528 10048 9540
rect 10100 9528 10106 9580
rect 11348 9568 11376 9608
rect 11698 9568 11704 9580
rect 10152 9540 11376 9568
rect 11659 9540 11704 9568
rect 9398 9460 9404 9512
rect 9456 9500 9462 9512
rect 9953 9503 10011 9509
rect 9953 9500 9965 9503
rect 9456 9472 9965 9500
rect 9456 9460 9462 9472
rect 9953 9469 9965 9472
rect 9999 9500 10011 9503
rect 10152 9500 10180 9540
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 12406 9568 12434 9608
rect 12621 9605 12633 9639
rect 12667 9636 12679 9639
rect 12986 9636 12992 9648
rect 12667 9608 12992 9636
rect 12667 9605 12679 9608
rect 12621 9599 12679 9605
rect 12986 9596 12992 9608
rect 13044 9596 13050 9648
rect 13541 9639 13599 9645
rect 13541 9605 13553 9639
rect 13587 9636 13599 9639
rect 13630 9636 13636 9648
rect 13587 9608 13636 9636
rect 13587 9605 13599 9608
rect 13541 9599 13599 9605
rect 13630 9596 13636 9608
rect 13688 9596 13694 9648
rect 15841 9639 15899 9645
rect 15841 9605 15853 9639
rect 15887 9636 15899 9639
rect 16114 9636 16120 9648
rect 15887 9608 16120 9636
rect 15887 9605 15899 9608
rect 15841 9599 15899 9605
rect 16114 9596 16120 9608
rect 16172 9596 16178 9648
rect 17034 9596 17040 9648
rect 17092 9636 17098 9648
rect 19242 9636 19248 9648
rect 17092 9608 19248 9636
rect 17092 9596 17098 9608
rect 12897 9571 12955 9577
rect 12406 9540 12848 9568
rect 9999 9472 10180 9500
rect 9999 9469 10011 9472
rect 9953 9463 10011 9469
rect 10502 9460 10508 9512
rect 10560 9500 10566 9512
rect 12066 9500 12072 9512
rect 10560 9472 12072 9500
rect 10560 9460 10566 9472
rect 12066 9460 12072 9472
rect 12124 9500 12130 9512
rect 12621 9503 12679 9509
rect 12621 9500 12633 9503
rect 12124 9472 12633 9500
rect 12124 9460 12130 9472
rect 12621 9469 12633 9472
rect 12667 9469 12679 9503
rect 12820 9500 12848 9540
rect 12897 9537 12909 9571
rect 12943 9568 12955 9571
rect 13446 9568 13452 9580
rect 12943 9540 13452 9568
rect 12943 9537 12955 9540
rect 12897 9531 12955 9537
rect 13446 9528 13452 9540
rect 13504 9528 13510 9580
rect 14182 9568 14188 9580
rect 14143 9540 14188 9568
rect 14182 9528 14188 9540
rect 14240 9528 14246 9580
rect 16022 9568 16028 9580
rect 15983 9540 16028 9568
rect 16022 9528 16028 9540
rect 16080 9528 16086 9580
rect 16206 9568 16212 9580
rect 16167 9540 16212 9568
rect 16206 9528 16212 9540
rect 16264 9528 16270 9580
rect 16298 9528 16304 9580
rect 16356 9568 16362 9580
rect 17497 9571 17555 9577
rect 17497 9568 17509 9571
rect 16356 9540 16401 9568
rect 16500 9540 17509 9568
rect 16356 9528 16362 9540
rect 14277 9503 14335 9509
rect 12820 9472 13584 9500
rect 12621 9463 12679 9469
rect 10597 9435 10655 9441
rect 10597 9401 10609 9435
rect 10643 9432 10655 9435
rect 11974 9432 11980 9444
rect 10643 9404 11980 9432
rect 10643 9401 10655 9404
rect 10597 9395 10655 9401
rect 11974 9392 11980 9404
rect 12032 9432 12038 9444
rect 12805 9435 12863 9441
rect 12805 9432 12817 9435
rect 12032 9404 12817 9432
rect 12032 9392 12038 9404
rect 12805 9401 12817 9404
rect 12851 9401 12863 9435
rect 12805 9395 12863 9401
rect 11882 9364 11888 9376
rect 7064 9336 9352 9364
rect 11843 9336 11888 9364
rect 7064 9324 7070 9336
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 13556 9364 13584 9472
rect 14277 9469 14289 9503
rect 14323 9500 14335 9503
rect 14642 9500 14648 9512
rect 14323 9472 14648 9500
rect 14323 9469 14335 9472
rect 14277 9463 14335 9469
rect 14642 9460 14648 9472
rect 14700 9460 14706 9512
rect 16114 9460 16120 9512
rect 16172 9500 16178 9512
rect 16500 9500 16528 9540
rect 17497 9537 17509 9540
rect 17543 9568 17555 9571
rect 17954 9568 17960 9580
rect 17543 9540 17960 9568
rect 17543 9537 17555 9540
rect 17497 9531 17555 9537
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 18891 9577 18919 9608
rect 19242 9596 19248 9608
rect 19300 9596 19306 9648
rect 18877 9571 18935 9577
rect 18877 9537 18889 9571
rect 18923 9537 18935 9571
rect 18877 9531 18935 9537
rect 19153 9571 19211 9577
rect 19153 9537 19165 9571
rect 19199 9568 19211 9571
rect 19352 9568 19380 9676
rect 19812 9676 20720 9704
rect 19812 9645 19840 9676
rect 20714 9664 20720 9676
rect 20772 9664 20778 9716
rect 21085 9707 21143 9713
rect 21085 9673 21097 9707
rect 21131 9704 21143 9707
rect 22646 9704 22652 9716
rect 21131 9676 22652 9704
rect 21131 9673 21143 9676
rect 21085 9667 21143 9673
rect 22646 9664 22652 9676
rect 22704 9664 22710 9716
rect 25866 9704 25872 9716
rect 24688 9676 25872 9704
rect 19797 9639 19855 9645
rect 19797 9605 19809 9639
rect 19843 9605 19855 9639
rect 20990 9636 20996 9648
rect 19797 9599 19855 9605
rect 19996 9608 20996 9636
rect 19996 9577 20024 9608
rect 20990 9596 20996 9608
rect 21048 9596 21054 9648
rect 21174 9596 21180 9648
rect 21232 9636 21238 9648
rect 23201 9639 23259 9645
rect 21232 9608 22692 9636
rect 21232 9596 21238 9608
rect 19199 9540 19380 9568
rect 19981 9571 20039 9577
rect 19199 9537 19211 9540
rect 19153 9531 19211 9537
rect 19981 9537 19993 9571
rect 20027 9537 20039 9571
rect 19981 9531 20039 9537
rect 20070 9528 20076 9580
rect 20128 9568 20134 9580
rect 20717 9571 20775 9577
rect 20717 9568 20729 9571
rect 20128 9540 20173 9568
rect 20272 9540 20729 9568
rect 20128 9528 20134 9540
rect 16172 9472 16528 9500
rect 16172 9460 16178 9472
rect 16942 9460 16948 9512
rect 17000 9500 17006 9512
rect 17405 9503 17463 9509
rect 17405 9500 17417 9503
rect 17000 9472 17417 9500
rect 17000 9460 17006 9472
rect 17405 9469 17417 9472
rect 17451 9469 17463 9503
rect 17972 9500 18000 9528
rect 18969 9503 19027 9509
rect 18969 9500 18981 9503
rect 17972 9472 18981 9500
rect 17405 9463 17463 9469
rect 18969 9469 18981 9472
rect 19015 9469 19027 9503
rect 18969 9463 19027 9469
rect 19058 9460 19064 9512
rect 19116 9500 19122 9512
rect 19334 9500 19340 9512
rect 19116 9472 19161 9500
rect 19295 9472 19340 9500
rect 19116 9460 19122 9472
rect 19334 9460 19340 9472
rect 19392 9460 19398 9512
rect 20272 9500 20300 9540
rect 20717 9537 20729 9540
rect 20763 9568 20775 9571
rect 20763 9540 22094 9568
rect 20763 9537 20775 9540
rect 20717 9531 20775 9537
rect 22066 9512 22094 9540
rect 20806 9500 20812 9512
rect 19996 9472 20300 9500
rect 20767 9472 20812 9500
rect 14550 9432 14556 9444
rect 14511 9404 14556 9432
rect 14550 9392 14556 9404
rect 14608 9392 14614 9444
rect 15381 9435 15439 9441
rect 15381 9401 15393 9435
rect 15427 9432 15439 9435
rect 18322 9432 18328 9444
rect 15427 9404 18328 9432
rect 15427 9401 15439 9404
rect 15381 9395 15439 9401
rect 18322 9392 18328 9404
rect 18380 9432 18386 9444
rect 19996 9432 20024 9472
rect 20806 9460 20812 9472
rect 20864 9460 20870 9512
rect 20990 9460 20996 9512
rect 21048 9500 21054 9512
rect 21818 9500 21824 9512
rect 21048 9472 21824 9500
rect 21048 9460 21054 9472
rect 21818 9460 21824 9472
rect 21876 9460 21882 9512
rect 22066 9472 22100 9512
rect 22094 9460 22100 9472
rect 22152 9500 22158 9512
rect 22664 9500 22692 9608
rect 23201 9605 23213 9639
rect 23247 9636 23259 9639
rect 23382 9636 23388 9648
rect 23247 9608 23388 9636
rect 23247 9605 23259 9608
rect 23201 9599 23259 9605
rect 23382 9596 23388 9608
rect 23440 9596 23446 9648
rect 24688 9636 24716 9676
rect 25866 9664 25872 9676
rect 25924 9704 25930 9716
rect 25924 9676 26188 9704
rect 25924 9664 25930 9676
rect 24596 9608 24716 9636
rect 24596 9577 24624 9608
rect 24854 9596 24860 9648
rect 24912 9636 24918 9648
rect 26160 9636 26188 9676
rect 26234 9664 26240 9716
rect 26292 9704 26298 9716
rect 33134 9704 33140 9716
rect 26292 9676 33140 9704
rect 26292 9664 26298 9676
rect 33134 9664 33140 9676
rect 33192 9664 33198 9716
rect 35710 9704 35716 9716
rect 33244 9676 35716 9704
rect 27706 9636 27712 9648
rect 24912 9608 25346 9636
rect 26160 9608 27712 9636
rect 24912 9596 24918 9608
rect 24581 9571 24639 9577
rect 24581 9537 24593 9571
rect 24627 9537 24639 9571
rect 24581 9531 24639 9537
rect 26605 9571 26663 9577
rect 26605 9537 26617 9571
rect 26651 9568 26663 9571
rect 27062 9568 27068 9580
rect 26651 9540 27068 9568
rect 26651 9537 26663 9540
rect 26605 9531 26663 9537
rect 27062 9528 27068 9540
rect 27120 9528 27126 9580
rect 27172 9577 27200 9608
rect 27706 9596 27712 9608
rect 27764 9596 27770 9648
rect 30190 9636 30196 9648
rect 30151 9608 30196 9636
rect 30190 9596 30196 9608
rect 30248 9596 30254 9648
rect 33244 9645 33272 9676
rect 35710 9664 35716 9676
rect 35768 9664 35774 9716
rect 36188 9676 36400 9704
rect 33236 9639 33294 9645
rect 33236 9605 33248 9639
rect 33282 9605 33294 9639
rect 33236 9599 33294 9605
rect 33502 9596 33508 9648
rect 33560 9636 33566 9648
rect 33686 9636 33692 9648
rect 33560 9608 33692 9636
rect 33560 9596 33566 9608
rect 33686 9596 33692 9608
rect 33744 9596 33750 9648
rect 35342 9636 35348 9648
rect 35303 9608 35348 9636
rect 35342 9596 35348 9608
rect 35400 9596 35406 9648
rect 35529 9639 35587 9645
rect 35529 9605 35541 9639
rect 35575 9636 35587 9639
rect 36188 9636 36216 9676
rect 35575 9608 35664 9636
rect 35575 9605 35587 9608
rect 35529 9599 35587 9605
rect 27157 9571 27215 9577
rect 27157 9537 27169 9571
rect 27203 9537 27215 9571
rect 27157 9531 27215 9537
rect 24857 9503 24915 9509
rect 24857 9500 24869 9503
rect 22152 9472 22197 9500
rect 22664 9472 24869 9500
rect 22152 9460 22158 9472
rect 24857 9469 24869 9472
rect 24903 9469 24915 9503
rect 24857 9463 24915 9469
rect 25314 9460 25320 9512
rect 25372 9500 25378 9512
rect 26050 9500 26056 9512
rect 25372 9472 26056 9500
rect 25372 9460 25378 9472
rect 26050 9460 26056 9472
rect 26108 9460 26114 9512
rect 27433 9503 27491 9509
rect 27433 9500 27445 9503
rect 26252 9472 27445 9500
rect 18380 9404 20024 9432
rect 20073 9435 20131 9441
rect 18380 9392 18386 9404
rect 20073 9401 20085 9435
rect 20119 9432 20131 9435
rect 22922 9432 22928 9444
rect 20119 9404 22928 9432
rect 20119 9401 20131 9404
rect 20073 9395 20131 9401
rect 22922 9392 22928 9404
rect 22980 9392 22986 9444
rect 21910 9364 21916 9376
rect 13556 9336 21916 9364
rect 21910 9324 21916 9336
rect 21968 9324 21974 9376
rect 22646 9364 22652 9376
rect 22607 9336 22652 9364
rect 22646 9324 22652 9336
rect 22704 9324 22710 9376
rect 23382 9324 23388 9376
rect 23440 9364 23446 9376
rect 26252 9364 26280 9472
rect 27433 9469 27445 9472
rect 27479 9469 27491 9503
rect 27433 9463 27491 9469
rect 27522 9460 27528 9512
rect 27580 9500 27586 9512
rect 28552 9500 28580 9554
rect 29914 9500 29920 9512
rect 27580 9472 28580 9500
rect 29875 9472 29920 9500
rect 27580 9460 27586 9472
rect 26602 9392 26608 9444
rect 26660 9392 26666 9444
rect 28552 9432 28580 9472
rect 29914 9460 29920 9472
rect 29972 9460 29978 9512
rect 30650 9500 30656 9512
rect 30024 9472 30656 9500
rect 30024 9432 30052 9472
rect 30650 9460 30656 9472
rect 30708 9500 30714 9512
rect 31312 9500 31340 9554
rect 32490 9528 32496 9580
rect 32548 9568 32554 9580
rect 32953 9571 33011 9577
rect 32953 9568 32965 9571
rect 32548 9540 32965 9568
rect 32548 9528 32554 9540
rect 32953 9537 32965 9540
rect 32999 9537 33011 9571
rect 32953 9531 33011 9537
rect 32401 9503 32459 9509
rect 32401 9500 32413 9503
rect 30708 9472 31340 9500
rect 31404 9472 32413 9500
rect 30708 9460 30714 9472
rect 28552 9404 30052 9432
rect 23440 9336 26280 9364
rect 26620 9364 26648 9392
rect 28905 9367 28963 9373
rect 28905 9364 28917 9367
rect 26620 9336 28917 9364
rect 23440 9324 23446 9336
rect 28905 9333 28917 9336
rect 28951 9333 28963 9367
rect 28905 9327 28963 9333
rect 28994 9324 29000 9376
rect 29052 9364 29058 9376
rect 31404 9364 31432 9472
rect 32401 9469 32413 9472
rect 32447 9500 32459 9503
rect 34514 9500 34520 9512
rect 32447 9472 34520 9500
rect 32447 9469 32459 9472
rect 32401 9463 32459 9469
rect 34514 9460 34520 9472
rect 34572 9460 34578 9512
rect 35360 9500 35388 9596
rect 35636 9578 35664 9608
rect 36096 9608 36216 9636
rect 36372 9636 36400 9676
rect 36446 9664 36452 9716
rect 36504 9704 36510 9716
rect 38378 9704 38384 9716
rect 36504 9676 38384 9704
rect 36504 9664 36510 9676
rect 38378 9664 38384 9676
rect 38436 9704 38442 9716
rect 39301 9707 39359 9713
rect 38436 9676 39160 9704
rect 38436 9664 38442 9676
rect 36372 9608 36492 9636
rect 36096 9578 36124 9608
rect 35636 9550 36124 9578
rect 36173 9571 36231 9577
rect 36173 9537 36185 9571
rect 36219 9537 36231 9571
rect 36173 9531 36231 9537
rect 36365 9571 36423 9577
rect 36365 9537 36377 9571
rect 36411 9568 36423 9571
rect 36464 9568 36492 9608
rect 36998 9596 37004 9648
rect 37056 9636 37062 9648
rect 39022 9636 39028 9648
rect 37056 9608 39028 9636
rect 37056 9596 37062 9608
rect 39022 9596 39028 9608
rect 39080 9596 39086 9648
rect 39132 9636 39160 9676
rect 39301 9673 39313 9707
rect 39347 9704 39359 9707
rect 39347 9676 40172 9704
rect 39347 9673 39359 9676
rect 39301 9667 39359 9673
rect 39853 9639 39911 9645
rect 39853 9636 39865 9639
rect 39132 9608 39865 9636
rect 39853 9605 39865 9608
rect 39899 9605 39911 9639
rect 40144 9636 40172 9676
rect 40218 9664 40224 9716
rect 40276 9704 40282 9716
rect 40313 9707 40371 9713
rect 40313 9704 40325 9707
rect 40276 9676 40325 9704
rect 40276 9664 40282 9676
rect 40313 9673 40325 9676
rect 40359 9673 40371 9707
rect 40313 9667 40371 9673
rect 41782 9664 41788 9716
rect 41840 9704 41846 9716
rect 44266 9704 44272 9716
rect 41840 9676 44272 9704
rect 41840 9664 41846 9676
rect 44266 9664 44272 9676
rect 44324 9704 44330 9716
rect 46290 9704 46296 9716
rect 44324 9676 46296 9704
rect 44324 9664 44330 9676
rect 46290 9664 46296 9676
rect 46348 9664 46354 9716
rect 48774 9704 48780 9716
rect 48148 9676 48780 9704
rect 40586 9636 40592 9648
rect 40144 9608 40592 9636
rect 39853 9599 39911 9605
rect 40586 9596 40592 9608
rect 40644 9596 40650 9648
rect 41874 9596 41880 9648
rect 41932 9636 41938 9648
rect 43625 9639 43683 9645
rect 43625 9636 43637 9639
rect 41932 9608 43637 9636
rect 41932 9596 41938 9608
rect 43625 9605 43637 9608
rect 43671 9605 43683 9639
rect 44634 9636 44640 9648
rect 43625 9599 43683 9605
rect 44192 9608 44640 9636
rect 36538 9568 36544 9580
rect 36411 9540 36544 9568
rect 36411 9537 36423 9540
rect 36365 9531 36423 9537
rect 36188 9500 36216 9531
rect 36538 9528 36544 9540
rect 36596 9528 36602 9580
rect 36814 9568 36820 9580
rect 36775 9540 36820 9568
rect 36814 9528 36820 9540
rect 36872 9528 36878 9580
rect 37458 9568 37464 9580
rect 36924 9540 37464 9568
rect 35360 9472 36216 9500
rect 36446 9460 36452 9512
rect 36504 9500 36510 9512
rect 36924 9500 36952 9540
rect 37458 9528 37464 9540
rect 37516 9528 37522 9580
rect 37734 9568 37740 9580
rect 37695 9540 37740 9568
rect 37734 9528 37740 9540
rect 37792 9528 37798 9580
rect 38746 9528 38752 9580
rect 38804 9568 38810 9580
rect 38841 9571 38899 9577
rect 38841 9568 38853 9571
rect 38804 9540 38853 9568
rect 38804 9528 38810 9540
rect 38841 9537 38853 9540
rect 38887 9537 38899 9571
rect 38841 9531 38899 9537
rect 39117 9571 39175 9577
rect 39117 9537 39129 9571
rect 39163 9568 39175 9571
rect 41141 9571 41199 9577
rect 39163 9540 39344 9568
rect 39163 9537 39175 9540
rect 39117 9531 39175 9537
rect 36504 9472 36952 9500
rect 36504 9460 36510 9472
rect 37366 9460 37372 9512
rect 37424 9500 37430 9512
rect 38562 9500 38568 9512
rect 37424 9472 38568 9500
rect 37424 9460 37430 9472
rect 38562 9460 38568 9472
rect 38620 9500 38626 9512
rect 38930 9500 38936 9512
rect 38620 9472 38936 9500
rect 38620 9460 38626 9472
rect 38930 9460 38936 9472
rect 38988 9460 38994 9512
rect 39316 9500 39344 9540
rect 41141 9537 41153 9571
rect 41187 9568 41199 9571
rect 41506 9568 41512 9580
rect 41187 9540 41512 9568
rect 41187 9537 41199 9540
rect 41141 9531 41199 9537
rect 41506 9528 41512 9540
rect 41564 9528 41570 9580
rect 41969 9571 42027 9577
rect 41969 9537 41981 9571
rect 42015 9568 42027 9571
rect 42150 9568 42156 9580
rect 42015 9540 42156 9568
rect 42015 9537 42027 9540
rect 41969 9531 42027 9537
rect 42150 9528 42156 9540
rect 42208 9528 42214 9580
rect 42794 9528 42800 9580
rect 42852 9568 42858 9580
rect 43165 9571 43223 9577
rect 43165 9568 43177 9571
rect 42852 9540 43177 9568
rect 42852 9528 42858 9540
rect 43165 9537 43177 9540
rect 43211 9568 43223 9571
rect 43530 9568 43536 9580
rect 43211 9540 43536 9568
rect 43211 9537 43223 9540
rect 43165 9531 43223 9537
rect 43530 9528 43536 9540
rect 43588 9528 43594 9580
rect 43806 9568 43812 9580
rect 43767 9540 43812 9568
rect 43806 9528 43812 9540
rect 43864 9528 43870 9580
rect 43898 9528 43904 9580
rect 43956 9568 43962 9580
rect 44192 9577 44220 9608
rect 44634 9596 44640 9608
rect 44692 9636 44698 9648
rect 47118 9636 47124 9648
rect 44692 9608 46336 9636
rect 47079 9608 47124 9636
rect 44692 9596 44698 9608
rect 44085 9571 44143 9577
rect 43956 9540 44001 9568
rect 43956 9528 43962 9540
rect 44085 9537 44097 9571
rect 44131 9537 44143 9571
rect 44085 9531 44143 9537
rect 44177 9571 44235 9577
rect 44177 9537 44189 9571
rect 44223 9537 44235 9571
rect 44177 9531 44235 9537
rect 39390 9500 39396 9512
rect 39316 9472 39396 9500
rect 39390 9460 39396 9472
rect 39448 9460 39454 9512
rect 41046 9500 41052 9512
rect 39960 9472 41052 9500
rect 31478 9392 31484 9444
rect 31536 9432 31542 9444
rect 34698 9432 34704 9444
rect 31536 9404 33088 9432
rect 34659 9404 34704 9432
rect 31536 9392 31542 9404
rect 33060 9376 33088 9404
rect 34698 9392 34704 9404
rect 34756 9392 34762 9444
rect 35526 9392 35532 9444
rect 35584 9392 35590 9444
rect 35618 9392 35624 9444
rect 35676 9432 35682 9444
rect 36078 9432 36084 9444
rect 35676 9404 36084 9432
rect 35676 9392 35682 9404
rect 36078 9392 36084 9404
rect 36136 9392 36142 9444
rect 36538 9392 36544 9444
rect 36596 9432 36602 9444
rect 37918 9432 37924 9444
rect 36596 9404 37924 9432
rect 36596 9392 36602 9404
rect 37918 9392 37924 9404
rect 37976 9432 37982 9444
rect 39960 9432 39988 9472
rect 41046 9460 41052 9472
rect 41104 9460 41110 9512
rect 41230 9500 41236 9512
rect 41191 9472 41236 9500
rect 41230 9460 41236 9472
rect 41288 9460 41294 9512
rect 42058 9460 42064 9512
rect 42116 9500 42122 9512
rect 44100 9500 44128 9531
rect 44358 9528 44364 9580
rect 44416 9568 44422 9580
rect 45373 9571 45431 9577
rect 45373 9568 45385 9571
rect 44416 9540 45385 9568
rect 44416 9528 44422 9540
rect 45373 9537 45385 9540
rect 45419 9537 45431 9571
rect 45373 9531 45431 9537
rect 46308 9512 46336 9608
rect 47118 9596 47124 9608
rect 47176 9636 47182 9648
rect 48148 9636 48176 9676
rect 48774 9664 48780 9676
rect 48832 9664 48838 9716
rect 49145 9707 49203 9713
rect 49145 9673 49157 9707
rect 49191 9674 49203 9707
rect 49191 9673 49280 9674
rect 49145 9667 49280 9673
rect 48314 9636 48320 9648
rect 47176 9608 48176 9636
rect 48275 9608 48320 9636
rect 47176 9596 47182 9608
rect 48314 9596 48320 9608
rect 48372 9596 48378 9648
rect 48498 9636 48504 9648
rect 48459 9608 48504 9636
rect 48498 9596 48504 9608
rect 48556 9596 48562 9648
rect 49160 9646 49280 9667
rect 50338 9664 50344 9716
rect 50396 9704 50402 9716
rect 50396 9676 53236 9704
rect 50396 9664 50402 9676
rect 49252 9636 49280 9646
rect 49602 9636 49608 9648
rect 49252 9608 49608 9636
rect 49602 9596 49608 9608
rect 49660 9596 49666 9648
rect 49970 9636 49976 9648
rect 49931 9608 49976 9636
rect 49970 9596 49976 9608
rect 50028 9596 50034 9648
rect 51350 9596 51356 9648
rect 51408 9636 51414 9648
rect 52917 9639 52975 9645
rect 52917 9636 52929 9639
rect 51408 9608 52929 9636
rect 51408 9596 51414 9608
rect 52917 9605 52929 9608
rect 52963 9605 52975 9639
rect 53098 9636 53104 9648
rect 53059 9608 53104 9636
rect 52917 9599 52975 9605
rect 53098 9596 53104 9608
rect 53156 9596 53162 9648
rect 53208 9636 53236 9676
rect 62390 9664 62396 9716
rect 62448 9664 62454 9716
rect 62500 9676 63540 9704
rect 53834 9636 53840 9648
rect 53208 9608 53840 9636
rect 53834 9596 53840 9608
rect 53892 9596 53898 9648
rect 61102 9636 61108 9648
rect 57348 9608 61108 9636
rect 49237 9571 49295 9577
rect 49237 9537 49249 9571
rect 49283 9537 49295 9571
rect 49237 9531 49295 9537
rect 42116 9472 44128 9500
rect 45465 9503 45523 9509
rect 42116 9460 42122 9472
rect 45465 9469 45477 9503
rect 45511 9500 45523 9503
rect 46198 9500 46204 9512
rect 45511 9472 46204 9500
rect 45511 9469 45523 9472
rect 45465 9463 45523 9469
rect 46198 9460 46204 9472
rect 46256 9460 46262 9512
rect 46290 9460 46296 9512
rect 46348 9460 46354 9512
rect 46566 9500 46572 9512
rect 46527 9472 46572 9500
rect 46566 9460 46572 9472
rect 46624 9500 46630 9512
rect 48222 9500 48228 9512
rect 46624 9472 48228 9500
rect 46624 9460 46630 9472
rect 48222 9460 48228 9472
rect 48280 9500 48286 9512
rect 48280 9460 48314 9500
rect 48682 9460 48688 9512
rect 48740 9500 48746 9512
rect 48961 9503 49019 9509
rect 48961 9500 48973 9503
rect 48740 9472 48973 9500
rect 48740 9460 48746 9472
rect 48961 9469 48973 9472
rect 49007 9469 49019 9503
rect 49252 9500 49280 9531
rect 49326 9528 49332 9580
rect 49384 9568 49390 9580
rect 49384 9540 49429 9568
rect 49384 9528 49390 9540
rect 51442 9528 51448 9580
rect 51500 9568 51506 9580
rect 52178 9568 52184 9580
rect 51500 9540 52184 9568
rect 51500 9528 51506 9540
rect 52178 9528 52184 9540
rect 52236 9528 52242 9580
rect 52270 9528 52276 9580
rect 52328 9568 52334 9580
rect 52365 9571 52423 9577
rect 52365 9568 52377 9571
rect 52328 9540 52377 9568
rect 52328 9528 52334 9540
rect 52365 9537 52377 9540
rect 52411 9537 52423 9571
rect 52365 9531 52423 9537
rect 52454 9528 52460 9580
rect 52512 9568 52518 9580
rect 53282 9568 53288 9580
rect 52512 9540 53288 9568
rect 52512 9528 52518 9540
rect 53282 9528 53288 9540
rect 53340 9528 53346 9580
rect 57348 9577 57376 9608
rect 61102 9596 61108 9608
rect 61160 9596 61166 9648
rect 62408 9636 62436 9664
rect 61948 9608 62436 9636
rect 57333 9571 57391 9577
rect 57333 9537 57345 9571
rect 57379 9537 57391 9571
rect 58066 9568 58072 9580
rect 58027 9540 58072 9568
rect 57333 9531 57391 9537
rect 58066 9528 58072 9540
rect 58124 9528 58130 9580
rect 58161 9571 58219 9577
rect 58161 9537 58173 9571
rect 58207 9568 58219 9571
rect 58802 9568 58808 9580
rect 58207 9540 58808 9568
rect 58207 9537 58219 9540
rect 58161 9531 58219 9537
rect 58802 9528 58808 9540
rect 58860 9528 58866 9580
rect 58897 9571 58955 9577
rect 58897 9537 58909 9571
rect 58943 9568 58955 9571
rect 58986 9568 58992 9580
rect 58943 9540 58992 9568
rect 58943 9537 58955 9540
rect 58897 9531 58955 9537
rect 58986 9528 58992 9540
rect 59044 9528 59050 9580
rect 61948 9577 61976 9608
rect 61933 9571 61991 9577
rect 61933 9537 61945 9571
rect 61979 9537 61991 9571
rect 62390 9568 62396 9580
rect 62351 9540 62396 9568
rect 61933 9531 61991 9537
rect 62390 9528 62396 9540
rect 62448 9568 62454 9580
rect 62500 9568 62528 9676
rect 63512 9665 63540 9676
rect 63310 9636 63316 9648
rect 63271 9608 63316 9636
rect 63310 9596 63316 9608
rect 63368 9596 63374 9648
rect 63512 9637 63724 9665
rect 65426 9664 65432 9716
rect 65484 9704 65490 9716
rect 70394 9704 70400 9716
rect 65484 9676 70400 9704
rect 65484 9664 65490 9676
rect 70394 9664 70400 9676
rect 70452 9664 70458 9716
rect 73154 9704 73160 9716
rect 71976 9676 73160 9704
rect 63696 9636 63724 9637
rect 64322 9636 64328 9648
rect 63696 9608 64328 9636
rect 62448 9540 62528 9568
rect 62577 9571 62635 9577
rect 62448 9528 62454 9540
rect 62577 9537 62589 9571
rect 62623 9568 62635 9571
rect 63034 9568 63040 9580
rect 62623 9540 63040 9568
rect 62623 9537 62635 9540
rect 62577 9531 62635 9537
rect 63034 9528 63040 9540
rect 63092 9528 63098 9580
rect 63218 9568 63224 9580
rect 63179 9540 63224 9568
rect 63218 9528 63224 9540
rect 63276 9528 63282 9580
rect 63435 9571 63493 9577
rect 63435 9537 63447 9571
rect 63481 9568 63493 9571
rect 63696 9568 63724 9608
rect 64322 9596 64328 9608
rect 64380 9596 64386 9648
rect 64690 9596 64696 9648
rect 64748 9636 64754 9648
rect 64785 9639 64843 9645
rect 64785 9636 64797 9639
rect 64748 9608 64797 9636
rect 64748 9596 64754 9608
rect 64785 9605 64797 9608
rect 64831 9605 64843 9639
rect 67634 9636 67640 9648
rect 66010 9608 67640 9636
rect 64785 9599 64843 9605
rect 67634 9596 67640 9608
rect 67692 9596 67698 9648
rect 67729 9639 67787 9645
rect 67729 9605 67741 9639
rect 67775 9636 67787 9639
rect 67910 9636 67916 9648
rect 67775 9608 67916 9636
rect 67775 9605 67787 9608
rect 67729 9599 67787 9605
rect 67910 9596 67916 9608
rect 67968 9596 67974 9648
rect 70486 9636 70492 9648
rect 70334 9608 70492 9636
rect 70486 9596 70492 9608
rect 70544 9596 70550 9648
rect 71976 9636 72004 9676
rect 73154 9664 73160 9676
rect 73212 9664 73218 9716
rect 73614 9664 73620 9716
rect 73672 9704 73678 9716
rect 75914 9704 75920 9716
rect 73672 9676 75920 9704
rect 73672 9664 73678 9676
rect 75914 9664 75920 9676
rect 75972 9704 75978 9716
rect 76834 9704 76840 9716
rect 75972 9676 76840 9704
rect 75972 9664 75978 9676
rect 76834 9664 76840 9676
rect 76892 9664 76898 9716
rect 76926 9664 76932 9716
rect 76984 9704 76990 9716
rect 84470 9704 84476 9716
rect 76984 9676 84476 9704
rect 76984 9664 76990 9676
rect 84470 9664 84476 9676
rect 84528 9704 84534 9716
rect 84654 9704 84660 9716
rect 84528 9676 84660 9704
rect 84528 9664 84534 9676
rect 84654 9664 84660 9676
rect 84712 9664 84718 9716
rect 84838 9664 84844 9716
rect 84896 9704 84902 9716
rect 84896 9676 87920 9704
rect 84896 9664 84902 9676
rect 71884 9608 72004 9636
rect 72973 9639 73031 9645
rect 71884 9590 71912 9608
rect 72973 9605 72985 9639
rect 73019 9636 73031 9639
rect 73430 9636 73436 9648
rect 73019 9608 73436 9636
rect 73019 9605 73031 9608
rect 72973 9599 73031 9605
rect 73430 9596 73436 9608
rect 73488 9596 73494 9648
rect 74166 9596 74172 9648
rect 74224 9636 74230 9648
rect 74224 9608 75224 9636
rect 74224 9596 74230 9608
rect 63481 9540 63724 9568
rect 63481 9537 63493 9540
rect 63435 9531 63493 9537
rect 66438 9528 66444 9580
rect 66496 9568 66502 9580
rect 67545 9571 67603 9577
rect 67545 9568 67557 9571
rect 66496 9540 67557 9568
rect 66496 9528 66502 9540
rect 67545 9537 67557 9540
rect 67591 9537 67603 9571
rect 67818 9568 67824 9580
rect 67779 9540 67824 9568
rect 67545 9531 67603 9537
rect 67818 9528 67824 9540
rect 67876 9528 67882 9580
rect 70394 9528 70400 9580
rect 70452 9568 70458 9580
rect 71581 9577 71639 9583
rect 71700 9577 71912 9590
rect 71581 9574 71593 9577
rect 71424 9568 71593 9574
rect 70452 9546 71593 9568
rect 70452 9540 71452 9546
rect 71581 9543 71593 9546
rect 71627 9543 71639 9577
rect 70452 9528 70458 9540
rect 71581 9537 71639 9543
rect 71685 9571 71912 9577
rect 71685 9537 71697 9571
rect 71731 9562 71912 9571
rect 72694 9568 72700 9580
rect 71731 9537 71743 9562
rect 72655 9540 72700 9568
rect 71685 9531 71743 9537
rect 72694 9528 72700 9540
rect 72752 9528 72758 9580
rect 73614 9528 73620 9580
rect 73672 9568 73678 9580
rect 73893 9571 73951 9577
rect 73893 9568 73905 9571
rect 73672 9540 73905 9568
rect 73672 9528 73678 9540
rect 73893 9537 73905 9540
rect 73939 9537 73951 9571
rect 74810 9568 74816 9580
rect 74771 9540 74816 9568
rect 73893 9531 73951 9537
rect 74810 9528 74816 9540
rect 74868 9528 74874 9580
rect 49252 9472 49372 9500
rect 48961 9463 49019 9469
rect 37976 9404 39988 9432
rect 37976 9392 37982 9404
rect 40034 9392 40040 9444
rect 40092 9432 40098 9444
rect 40129 9435 40187 9441
rect 40129 9432 40141 9435
rect 40092 9404 40141 9432
rect 40092 9392 40098 9404
rect 40129 9401 40141 9404
rect 40175 9401 40187 9435
rect 40129 9395 40187 9401
rect 40218 9392 40224 9444
rect 40276 9432 40282 9444
rect 40773 9435 40831 9441
rect 40773 9432 40785 9435
rect 40276 9404 40785 9432
rect 40276 9392 40282 9404
rect 40773 9401 40785 9404
rect 40819 9401 40831 9435
rect 45002 9432 45008 9444
rect 44963 9404 45008 9432
rect 40773 9395 40831 9401
rect 45002 9392 45008 9404
rect 45060 9392 45066 9444
rect 47486 9392 47492 9444
rect 47544 9432 47550 9444
rect 48133 9435 48191 9441
rect 48133 9432 48145 9435
rect 47544 9404 48145 9432
rect 47544 9392 47550 9404
rect 48133 9401 48145 9404
rect 48179 9401 48191 9435
rect 48286 9432 48314 9460
rect 49344 9432 49372 9472
rect 49694 9460 49700 9512
rect 49752 9500 49758 9512
rect 49789 9503 49847 9509
rect 49789 9500 49801 9503
rect 49752 9472 49801 9500
rect 49752 9460 49758 9472
rect 49789 9469 49801 9472
rect 49835 9469 49847 9503
rect 49789 9463 49847 9469
rect 51350 9460 51356 9512
rect 51408 9500 51414 9512
rect 51629 9503 51687 9509
rect 51629 9500 51641 9503
rect 51408 9472 51641 9500
rect 51408 9460 51414 9472
rect 51629 9469 51641 9472
rect 51675 9500 51687 9503
rect 55766 9500 55772 9512
rect 51675 9472 55772 9500
rect 51675 9469 51687 9472
rect 51629 9463 51687 9469
rect 55766 9460 55772 9472
rect 55824 9460 55830 9512
rect 56042 9500 56048 9512
rect 56003 9472 56048 9500
rect 56042 9460 56048 9472
rect 56100 9460 56106 9512
rect 56229 9503 56287 9509
rect 56229 9469 56241 9503
rect 56275 9500 56287 9503
rect 56502 9500 56508 9512
rect 56275 9472 56508 9500
rect 56275 9469 56287 9472
rect 56229 9463 56287 9469
rect 56502 9460 56508 9472
rect 56560 9460 56566 9512
rect 58618 9460 58624 9512
rect 58676 9500 58682 9512
rect 60642 9500 60648 9512
rect 58676 9472 60648 9500
rect 58676 9460 58682 9472
rect 60642 9460 60648 9472
rect 60700 9460 60706 9512
rect 61105 9503 61163 9509
rect 61105 9469 61117 9503
rect 61151 9469 61163 9503
rect 61286 9500 61292 9512
rect 61247 9472 61292 9500
rect 61105 9463 61163 9469
rect 48286 9404 49372 9432
rect 48133 9395 48191 9401
rect 31662 9364 31668 9376
rect 29052 9336 31432 9364
rect 31623 9336 31668 9364
rect 29052 9324 29058 9336
rect 31662 9324 31668 9336
rect 31720 9324 31726 9376
rect 33042 9324 33048 9376
rect 33100 9324 33106 9376
rect 33318 9324 33324 9376
rect 33376 9364 33382 9376
rect 35158 9364 35164 9376
rect 33376 9336 35164 9364
rect 33376 9324 33382 9336
rect 35158 9324 35164 9336
rect 35216 9324 35222 9376
rect 35544 9364 35572 9392
rect 35713 9367 35771 9373
rect 35713 9364 35725 9367
rect 35544 9336 35725 9364
rect 35713 9333 35725 9336
rect 35759 9333 35771 9367
rect 36262 9364 36268 9376
rect 36223 9336 36268 9364
rect 35713 9327 35771 9333
rect 36262 9324 36268 9336
rect 36320 9324 36326 9376
rect 38194 9324 38200 9376
rect 38252 9364 38258 9376
rect 38289 9367 38347 9373
rect 38289 9364 38301 9367
rect 38252 9336 38301 9364
rect 38252 9324 38258 9336
rect 38289 9333 38301 9336
rect 38335 9333 38347 9367
rect 38289 9327 38347 9333
rect 38378 9324 38384 9376
rect 38436 9364 38442 9376
rect 38841 9367 38899 9373
rect 38841 9364 38853 9367
rect 38436 9336 38853 9364
rect 38436 9324 38442 9336
rect 38841 9333 38853 9336
rect 38887 9333 38899 9367
rect 38841 9327 38899 9333
rect 38930 9324 38936 9376
rect 38988 9364 38994 9376
rect 41782 9364 41788 9376
rect 38988 9336 41788 9364
rect 38988 9324 38994 9336
rect 41782 9324 41788 9336
rect 41840 9324 41846 9376
rect 45554 9324 45560 9376
rect 45612 9364 45618 9376
rect 46017 9367 46075 9373
rect 46017 9364 46029 9367
rect 45612 9336 46029 9364
rect 45612 9324 45618 9336
rect 46017 9333 46029 9336
rect 46063 9364 46075 9367
rect 48866 9364 48872 9376
rect 46063 9336 48872 9364
rect 46063 9333 46075 9336
rect 46017 9327 46075 9333
rect 48866 9324 48872 9336
rect 48924 9324 48930 9376
rect 49050 9364 49056 9376
rect 49011 9336 49056 9364
rect 49050 9324 49056 9336
rect 49108 9324 49114 9376
rect 49344 9364 49372 9404
rect 49418 9392 49424 9444
rect 49476 9432 49482 9444
rect 61010 9432 61016 9444
rect 49476 9404 61016 9432
rect 49476 9392 49482 9404
rect 61010 9392 61016 9404
rect 61068 9392 61074 9444
rect 61120 9432 61148 9463
rect 61286 9460 61292 9472
rect 61344 9460 61350 9512
rect 62114 9460 62120 9512
rect 62172 9500 62178 9512
rect 63589 9503 63647 9509
rect 63589 9500 63601 9503
rect 62172 9472 63601 9500
rect 62172 9460 62178 9472
rect 63589 9469 63601 9472
rect 63635 9500 63647 9503
rect 64138 9500 64144 9512
rect 63635 9472 64144 9500
rect 63635 9469 63647 9472
rect 63589 9463 63647 9469
rect 64138 9460 64144 9472
rect 64196 9460 64202 9512
rect 64414 9460 64420 9512
rect 64472 9500 64478 9512
rect 64509 9503 64567 9509
rect 64509 9500 64521 9503
rect 64472 9472 64521 9500
rect 64472 9460 64478 9472
rect 64509 9469 64521 9472
rect 64555 9469 64567 9503
rect 67836 9500 67864 9528
rect 68830 9500 68836 9512
rect 64509 9463 64567 9469
rect 64616 9472 67864 9500
rect 68791 9472 68836 9500
rect 63126 9432 63132 9444
rect 61120 9404 63132 9432
rect 63126 9392 63132 9404
rect 63184 9392 63190 9444
rect 63497 9435 63555 9441
rect 63497 9401 63509 9435
rect 63543 9432 63555 9435
rect 64616 9432 64644 9472
rect 68830 9460 68836 9472
rect 68888 9460 68894 9512
rect 69109 9503 69167 9509
rect 69109 9469 69121 9503
rect 69155 9500 69167 9503
rect 70581 9503 70639 9509
rect 69155 9472 70532 9500
rect 69155 9469 69167 9472
rect 69109 9463 69167 9469
rect 63543 9404 64644 9432
rect 63543 9401 63555 9404
rect 63497 9395 63555 9401
rect 65794 9392 65800 9444
rect 65852 9432 65858 9444
rect 70504 9432 70532 9472
rect 70581 9469 70593 9503
rect 70627 9500 70639 9503
rect 71406 9500 71412 9512
rect 70627 9472 71412 9500
rect 70627 9469 70639 9472
rect 70581 9463 70639 9469
rect 71406 9460 71412 9472
rect 71464 9460 71470 9512
rect 74721 9503 74779 9509
rect 74721 9500 74733 9503
rect 71700 9472 74733 9500
rect 71700 9432 71728 9472
rect 74721 9469 74733 9472
rect 74767 9469 74779 9503
rect 75196 9500 75224 9608
rect 75270 9596 75276 9648
rect 75328 9636 75334 9648
rect 75365 9639 75423 9645
rect 75365 9636 75377 9639
rect 75328 9608 75377 9636
rect 75328 9596 75334 9608
rect 75365 9605 75377 9608
rect 75411 9605 75423 9639
rect 76006 9636 76012 9648
rect 75967 9608 76012 9636
rect 75365 9599 75423 9605
rect 76006 9596 76012 9608
rect 76064 9596 76070 9648
rect 78950 9636 78956 9648
rect 76116 9608 78956 9636
rect 75454 9528 75460 9580
rect 75512 9568 75518 9580
rect 75917 9571 75975 9577
rect 75917 9568 75929 9571
rect 75512 9540 75557 9568
rect 75749 9540 75929 9568
rect 75512 9528 75518 9540
rect 75749 9500 75777 9540
rect 75917 9537 75929 9540
rect 75963 9568 75975 9571
rect 76116 9568 76144 9608
rect 78950 9596 78956 9608
rect 79008 9596 79014 9648
rect 79226 9596 79232 9648
rect 79284 9636 79290 9648
rect 82449 9639 82507 9645
rect 79284 9608 80054 9636
rect 79284 9596 79290 9608
rect 75963 9540 76144 9568
rect 76653 9571 76711 9577
rect 75963 9537 75975 9540
rect 75917 9531 75975 9537
rect 76653 9537 76665 9571
rect 76699 9537 76711 9571
rect 78122 9568 78128 9580
rect 78035 9540 78128 9568
rect 76653 9531 76711 9537
rect 76668 9500 76696 9531
rect 78122 9528 78128 9540
rect 78180 9528 78186 9580
rect 79134 9528 79140 9580
rect 79192 9568 79198 9580
rect 79505 9571 79563 9577
rect 79505 9568 79517 9571
rect 79192 9540 79517 9568
rect 79192 9528 79198 9540
rect 79505 9537 79517 9540
rect 79551 9537 79563 9571
rect 79505 9531 79563 9537
rect 76926 9500 76932 9512
rect 75196 9472 75777 9500
rect 75932 9472 76696 9500
rect 76887 9472 76932 9500
rect 74721 9463 74779 9469
rect 75932 9444 75960 9472
rect 65852 9404 67634 9432
rect 70504 9404 71728 9432
rect 71792 9404 74212 9432
rect 65852 9392 65858 9404
rect 55858 9364 55864 9376
rect 49344 9336 55864 9364
rect 55858 9324 55864 9336
rect 55916 9324 55922 9376
rect 57146 9364 57152 9376
rect 57107 9336 57152 9364
rect 57146 9324 57152 9336
rect 57204 9324 57210 9376
rect 58802 9364 58808 9376
rect 58763 9336 58808 9364
rect 58802 9324 58808 9336
rect 58860 9324 58866 9376
rect 58986 9324 58992 9376
rect 59044 9364 59050 9376
rect 61746 9364 61752 9376
rect 59044 9336 61752 9364
rect 59044 9324 59050 9336
rect 61746 9324 61752 9336
rect 61804 9324 61810 9376
rect 61841 9367 61899 9373
rect 61841 9333 61853 9367
rect 61887 9364 61899 9367
rect 61930 9364 61936 9376
rect 61887 9336 61936 9364
rect 61887 9333 61899 9336
rect 61841 9327 61899 9333
rect 61930 9324 61936 9336
rect 61988 9324 61994 9376
rect 62574 9364 62580 9376
rect 62535 9336 62580 9364
rect 62574 9324 62580 9336
rect 62632 9324 62638 9376
rect 63770 9324 63776 9376
rect 63828 9364 63834 9376
rect 66257 9367 66315 9373
rect 66257 9364 66269 9367
rect 63828 9336 66269 9364
rect 63828 9324 63834 9336
rect 66257 9333 66269 9336
rect 66303 9333 66315 9367
rect 66714 9364 66720 9376
rect 66675 9336 66720 9364
rect 66257 9327 66315 9333
rect 66714 9324 66720 9336
rect 66772 9324 66778 9376
rect 67358 9364 67364 9376
rect 67319 9336 67364 9364
rect 67358 9324 67364 9336
rect 67416 9324 67422 9376
rect 67606 9364 67634 9404
rect 70394 9364 70400 9376
rect 67606 9336 70400 9364
rect 70394 9324 70400 9336
rect 70452 9324 70458 9376
rect 71038 9364 71044 9376
rect 70999 9336 71044 9364
rect 71038 9324 71044 9336
rect 71096 9324 71102 9376
rect 71130 9324 71136 9376
rect 71188 9364 71194 9376
rect 71792 9373 71820 9404
rect 71777 9367 71835 9373
rect 71777 9364 71789 9367
rect 71188 9336 71789 9364
rect 71188 9324 71194 9336
rect 71777 9333 71789 9336
rect 71823 9333 71835 9367
rect 71777 9327 71835 9333
rect 71961 9367 72019 9373
rect 71961 9333 71973 9367
rect 72007 9364 72019 9367
rect 72142 9364 72148 9376
rect 72007 9336 72148 9364
rect 72007 9333 72019 9336
rect 71961 9327 72019 9333
rect 72142 9324 72148 9336
rect 72200 9324 72206 9376
rect 74074 9364 74080 9376
rect 74035 9336 74080 9364
rect 74074 9324 74080 9336
rect 74132 9324 74138 9376
rect 74184 9364 74212 9404
rect 75914 9392 75920 9444
rect 75972 9392 75978 9444
rect 76668 9432 76696 9472
rect 76926 9460 76932 9472
rect 76984 9500 76990 9512
rect 77754 9500 77760 9512
rect 76984 9472 77760 9500
rect 76984 9460 76990 9472
rect 77754 9460 77760 9472
rect 77812 9460 77818 9512
rect 77849 9503 77907 9509
rect 77849 9469 77861 9503
rect 77895 9500 77907 9503
rect 77938 9500 77944 9512
rect 77895 9472 77944 9500
rect 77895 9469 77907 9472
rect 77849 9463 77907 9469
rect 77938 9460 77944 9472
rect 77996 9460 78002 9512
rect 78140 9500 78168 9528
rect 79413 9503 79471 9509
rect 79413 9500 79425 9503
rect 78140 9472 79425 9500
rect 79413 9469 79425 9472
rect 79459 9469 79471 9503
rect 79413 9463 79471 9469
rect 79226 9432 79232 9444
rect 76668 9404 79232 9432
rect 79226 9392 79232 9404
rect 79284 9392 79290 9444
rect 78122 9364 78128 9376
rect 74184 9336 78128 9364
rect 78122 9324 78128 9336
rect 78180 9364 78186 9376
rect 78769 9367 78827 9373
rect 78769 9364 78781 9367
rect 78180 9336 78781 9364
rect 78180 9324 78186 9336
rect 78769 9333 78781 9336
rect 78815 9364 78827 9367
rect 78858 9364 78864 9376
rect 78815 9336 78864 9364
rect 78815 9333 78827 9336
rect 78769 9327 78827 9333
rect 78858 9324 78864 9336
rect 78916 9364 78922 9376
rect 79594 9364 79600 9376
rect 78916 9336 79600 9364
rect 78916 9324 78922 9336
rect 79594 9324 79600 9336
rect 79652 9324 79658 9376
rect 80026 9364 80054 9608
rect 82449 9605 82461 9639
rect 82495 9636 82507 9639
rect 85574 9636 85580 9648
rect 82495 9608 85580 9636
rect 82495 9605 82507 9608
rect 82449 9599 82507 9605
rect 85574 9596 85580 9608
rect 85632 9596 85638 9648
rect 85942 9596 85948 9648
rect 86000 9596 86006 9648
rect 87782 9636 87788 9648
rect 87743 9608 87788 9636
rect 87782 9596 87788 9608
rect 87840 9596 87846 9648
rect 82814 9528 82820 9580
rect 82872 9568 82878 9580
rect 83093 9571 83151 9577
rect 83093 9568 83105 9571
rect 82872 9540 83105 9568
rect 82872 9528 82878 9540
rect 83093 9537 83105 9540
rect 83139 9537 83151 9571
rect 83093 9531 83151 9537
rect 83366 9528 83372 9580
rect 83424 9568 83430 9580
rect 84197 9571 84255 9577
rect 84197 9568 84209 9571
rect 83424 9540 84209 9568
rect 83424 9528 83430 9540
rect 84197 9537 84209 9540
rect 84243 9537 84255 9571
rect 84470 9568 84476 9580
rect 84431 9540 84476 9568
rect 84197 9531 84255 9537
rect 84470 9528 84476 9540
rect 84528 9528 84534 9580
rect 87892 9577 87920 9676
rect 91186 9636 91192 9648
rect 90192 9608 91192 9636
rect 87877 9571 87935 9577
rect 87877 9537 87889 9571
rect 87923 9568 87935 9571
rect 88242 9568 88248 9580
rect 87923 9540 88248 9568
rect 87923 9537 87935 9540
rect 87877 9531 87935 9537
rect 88242 9528 88248 9540
rect 88300 9528 88306 9580
rect 90192 9577 90220 9608
rect 91186 9596 91192 9608
rect 91244 9596 91250 9648
rect 93762 9636 93768 9648
rect 92138 9608 93768 9636
rect 93762 9596 93768 9608
rect 93820 9596 93826 9648
rect 94222 9636 94228 9648
rect 94183 9608 94228 9636
rect 94222 9596 94228 9608
rect 94280 9596 94286 9648
rect 88981 9571 89039 9577
rect 88981 9537 88993 9571
rect 89027 9537 89039 9571
rect 88981 9531 89039 9537
rect 90177 9571 90235 9577
rect 90177 9537 90189 9571
rect 90223 9537 90235 9571
rect 90177 9531 90235 9537
rect 80333 9503 80391 9509
rect 80333 9469 80345 9503
rect 80379 9500 80391 9503
rect 80698 9500 80704 9512
rect 80379 9472 80704 9500
rect 80379 9469 80391 9472
rect 80333 9463 80391 9469
rect 80698 9460 80704 9472
rect 80756 9460 80762 9512
rect 80793 9503 80851 9509
rect 80793 9469 80805 9503
rect 80839 9469 80851 9503
rect 80793 9463 80851 9469
rect 82633 9503 82691 9509
rect 82633 9469 82645 9503
rect 82679 9500 82691 9503
rect 82722 9500 82728 9512
rect 82679 9472 82728 9500
rect 82679 9469 82691 9472
rect 82633 9463 82691 9469
rect 80606 9392 80612 9444
rect 80664 9432 80670 9444
rect 80808 9432 80836 9463
rect 82722 9460 82728 9472
rect 82780 9460 82786 9512
rect 83826 9500 83832 9512
rect 83787 9472 83832 9500
rect 83826 9460 83832 9472
rect 83884 9460 83890 9512
rect 86957 9503 87015 9509
rect 86957 9469 86969 9503
rect 87003 9500 87015 9503
rect 87003 9472 87184 9500
rect 87003 9469 87015 9472
rect 86957 9463 87015 9469
rect 81434 9432 81440 9444
rect 80664 9404 81440 9432
rect 80664 9392 80670 9404
rect 81434 9392 81440 9404
rect 81492 9392 81498 9444
rect 83185 9435 83243 9441
rect 83185 9401 83197 9435
rect 83231 9432 83243 9435
rect 85390 9432 85396 9444
rect 83231 9404 85396 9432
rect 83231 9401 83243 9404
rect 83185 9395 83243 9401
rect 85390 9392 85396 9404
rect 85448 9392 85454 9444
rect 87156 9432 87184 9472
rect 87230 9460 87236 9512
rect 87288 9500 87294 9512
rect 87288 9472 87333 9500
rect 87288 9460 87294 9472
rect 87690 9460 87696 9512
rect 87748 9500 87754 9512
rect 88996 9500 89024 9531
rect 92842 9528 92848 9580
rect 92900 9568 92906 9580
rect 93213 9571 93271 9577
rect 93213 9568 93225 9571
rect 92900 9540 93225 9568
rect 92900 9528 92906 9540
rect 93213 9537 93225 9540
rect 93259 9537 93271 9571
rect 93213 9531 93271 9537
rect 94038 9528 94044 9580
rect 94096 9568 94102 9580
rect 94133 9571 94191 9577
rect 94133 9568 94145 9571
rect 94096 9540 94145 9568
rect 94096 9528 94102 9540
rect 94133 9537 94145 9540
rect 94179 9537 94191 9571
rect 94133 9531 94191 9537
rect 87748 9472 89024 9500
rect 87748 9460 87754 9472
rect 89714 9460 89720 9512
rect 89772 9500 89778 9512
rect 90634 9500 90640 9512
rect 89772 9472 90640 9500
rect 89772 9460 89778 9472
rect 90634 9460 90640 9472
rect 90692 9460 90698 9512
rect 90913 9503 90971 9509
rect 90913 9469 90925 9503
rect 90959 9500 90971 9503
rect 93946 9500 93952 9512
rect 90959 9472 93952 9500
rect 90959 9469 90971 9472
rect 90913 9463 90971 9469
rect 93946 9460 93952 9472
rect 94004 9460 94010 9512
rect 89073 9435 89131 9441
rect 89073 9432 89085 9435
rect 87156 9404 89085 9432
rect 89073 9401 89085 9404
rect 89119 9401 89131 9435
rect 89073 9395 89131 9401
rect 84102 9364 84108 9376
rect 80026 9336 84108 9364
rect 84102 9324 84108 9336
rect 84160 9324 84166 9376
rect 85485 9367 85543 9373
rect 85485 9333 85497 9367
rect 85531 9364 85543 9367
rect 85758 9364 85764 9376
rect 85531 9336 85764 9364
rect 85531 9333 85543 9336
rect 85485 9327 85543 9333
rect 85758 9324 85764 9336
rect 85816 9364 85822 9376
rect 86494 9364 86500 9376
rect 85816 9336 86500 9364
rect 85816 9324 85822 9336
rect 86494 9324 86500 9336
rect 86552 9324 86558 9376
rect 86586 9324 86592 9376
rect 86644 9364 86650 9376
rect 88058 9364 88064 9376
rect 86644 9336 88064 9364
rect 86644 9324 86650 9336
rect 88058 9324 88064 9336
rect 88116 9324 88122 9376
rect 88242 9324 88248 9376
rect 88300 9364 88306 9376
rect 88337 9367 88395 9373
rect 88337 9364 88349 9367
rect 88300 9336 88349 9364
rect 88300 9324 88306 9336
rect 88337 9333 88349 9336
rect 88383 9333 88395 9367
rect 88337 9327 88395 9333
rect 90177 9367 90235 9373
rect 90177 9333 90189 9367
rect 90223 9364 90235 9367
rect 91094 9364 91100 9376
rect 90223 9336 91100 9364
rect 90223 9333 90235 9336
rect 90177 9327 90235 9333
rect 91094 9324 91100 9336
rect 91152 9324 91158 9376
rect 91278 9324 91284 9376
rect 91336 9364 91342 9376
rect 92382 9364 92388 9376
rect 91336 9336 92388 9364
rect 91336 9324 91342 9336
rect 92382 9324 92388 9336
rect 92440 9324 92446 9376
rect 92474 9324 92480 9376
rect 92532 9364 92538 9376
rect 92937 9367 92995 9373
rect 92937 9364 92949 9367
rect 92532 9336 92949 9364
rect 92532 9324 92538 9336
rect 92937 9333 92949 9336
rect 92983 9333 92995 9367
rect 92937 9327 92995 9333
rect 1104 9274 94852 9296
rect 1104 9222 12668 9274
rect 12720 9222 12732 9274
rect 12784 9222 12796 9274
rect 12848 9222 12860 9274
rect 12912 9222 12924 9274
rect 12976 9222 36105 9274
rect 36157 9222 36169 9274
rect 36221 9222 36233 9274
rect 36285 9222 36297 9274
rect 36349 9222 36361 9274
rect 36413 9222 59542 9274
rect 59594 9222 59606 9274
rect 59658 9222 59670 9274
rect 59722 9222 59734 9274
rect 59786 9222 59798 9274
rect 59850 9222 82979 9274
rect 83031 9222 83043 9274
rect 83095 9222 83107 9274
rect 83159 9222 83171 9274
rect 83223 9222 83235 9274
rect 83287 9222 94852 9274
rect 1104 9200 94852 9222
rect 1765 9163 1823 9169
rect 1765 9129 1777 9163
rect 1811 9160 1823 9163
rect 2498 9160 2504 9172
rect 1811 9132 2504 9160
rect 1811 9129 1823 9132
rect 1765 9123 1823 9129
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 3418 9160 3424 9172
rect 3379 9132 3424 9160
rect 3418 9120 3424 9132
rect 3476 9120 3482 9172
rect 5810 9120 5816 9172
rect 5868 9160 5874 9172
rect 7006 9160 7012 9172
rect 5868 9132 7012 9160
rect 5868 9120 5874 9132
rect 7006 9120 7012 9132
rect 7064 9120 7070 9172
rect 14642 9160 14648 9172
rect 7576 9132 14136 9160
rect 14603 9132 14648 9160
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 5828 9092 5856 9120
rect 4120 9064 5856 9092
rect 4120 9052 4126 9064
rect 2222 9024 2228 9036
rect 2183 8996 2228 9024
rect 2222 8984 2228 8996
rect 2280 8984 2286 9036
rect 4246 9024 4252 9036
rect 4207 8996 4252 9024
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 5077 9027 5135 9033
rect 5077 8993 5089 9027
rect 5123 9024 5135 9027
rect 7576 9024 7604 9132
rect 8018 9052 8024 9104
rect 8076 9092 8082 9104
rect 8389 9095 8447 9101
rect 8389 9092 8401 9095
rect 8076 9064 8401 9092
rect 8076 9052 8082 9064
rect 8389 9061 8401 9064
rect 8435 9092 8447 9095
rect 9214 9092 9220 9104
rect 8435 9064 9220 9092
rect 8435 9061 8447 9064
rect 8389 9055 8447 9061
rect 9214 9052 9220 9064
rect 9272 9052 9278 9104
rect 13446 9092 13452 9104
rect 12176 9064 13452 9092
rect 5123 8996 7604 9024
rect 7745 9027 7803 9033
rect 5123 8993 5135 8996
rect 5077 8987 5135 8993
rect 7745 8993 7757 9027
rect 7791 9024 7803 9027
rect 9122 9024 9128 9036
rect 7791 8996 9128 9024
rect 7791 8993 7803 8996
rect 7745 8987 7803 8993
rect 9122 8984 9128 8996
rect 9180 8984 9186 9036
rect 9398 9024 9404 9036
rect 9359 8996 9404 9024
rect 9398 8984 9404 8996
rect 9456 9024 9462 9036
rect 9766 9024 9772 9036
rect 9456 8996 9772 9024
rect 9456 8984 9462 8996
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 11238 8984 11244 9036
rect 11296 9024 11302 9036
rect 12176 9024 12204 9064
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 14108 9092 14136 9132
rect 14642 9120 14648 9132
rect 14700 9120 14706 9172
rect 15657 9163 15715 9169
rect 15657 9129 15669 9163
rect 15703 9160 15715 9163
rect 16022 9160 16028 9172
rect 15703 9132 16028 9160
rect 15703 9129 15715 9132
rect 15657 9123 15715 9129
rect 16022 9120 16028 9132
rect 16080 9120 16086 9172
rect 16206 9160 16212 9172
rect 16167 9132 16212 9160
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 16942 9160 16948 9172
rect 16903 9132 16948 9160
rect 16942 9120 16948 9132
rect 17000 9120 17006 9172
rect 17218 9120 17224 9172
rect 17276 9160 17282 9172
rect 17681 9163 17739 9169
rect 17681 9160 17693 9163
rect 17276 9132 17693 9160
rect 17276 9120 17282 9132
rect 17681 9129 17693 9132
rect 17727 9160 17739 9163
rect 17770 9160 17776 9172
rect 17727 9132 17776 9160
rect 17727 9129 17739 9132
rect 17681 9123 17739 9129
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 18141 9163 18199 9169
rect 18141 9160 18153 9163
rect 17880 9132 18153 9160
rect 14826 9092 14832 9104
rect 14108 9064 14832 9092
rect 14826 9052 14832 9064
rect 14884 9052 14890 9104
rect 14918 9052 14924 9104
rect 14976 9092 14982 9104
rect 14976 9064 16528 9092
rect 14976 9052 14982 9064
rect 16500 9036 16528 9064
rect 16758 9052 16764 9104
rect 16816 9092 16822 9104
rect 17880 9092 17908 9132
rect 18141 9129 18153 9132
rect 18187 9160 18199 9163
rect 18414 9160 18420 9172
rect 18187 9132 18420 9160
rect 18187 9129 18199 9132
rect 18141 9123 18199 9129
rect 18414 9120 18420 9132
rect 18472 9120 18478 9172
rect 18506 9120 18512 9172
rect 18564 9160 18570 9172
rect 19702 9160 19708 9172
rect 18564 9132 19708 9160
rect 18564 9120 18570 9132
rect 19702 9120 19708 9132
rect 19760 9120 19766 9172
rect 19886 9160 19892 9172
rect 19847 9132 19892 9160
rect 19886 9120 19892 9132
rect 19944 9120 19950 9172
rect 20901 9163 20959 9169
rect 20901 9129 20913 9163
rect 20947 9160 20959 9163
rect 21174 9160 21180 9172
rect 20947 9132 21180 9160
rect 20947 9129 20959 9132
rect 20901 9123 20959 9129
rect 21174 9120 21180 9132
rect 21232 9120 21238 9172
rect 21818 9160 21824 9172
rect 21779 9132 21824 9160
rect 21818 9120 21824 9132
rect 21876 9120 21882 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 27430 9160 27436 9172
rect 22152 9132 27436 9160
rect 22152 9120 22158 9132
rect 27430 9120 27436 9132
rect 27488 9120 27494 9172
rect 27522 9120 27528 9172
rect 27580 9160 27586 9172
rect 28994 9160 29000 9172
rect 27580 9132 29000 9160
rect 27580 9120 27586 9132
rect 28994 9120 29000 9132
rect 29052 9120 29058 9172
rect 29362 9120 29368 9172
rect 29420 9160 29426 9172
rect 29825 9163 29883 9169
rect 29825 9160 29837 9163
rect 29420 9132 29837 9160
rect 29420 9120 29426 9132
rect 29825 9129 29837 9132
rect 29871 9129 29883 9163
rect 29825 9123 29883 9129
rect 31662 9120 31668 9172
rect 31720 9160 31726 9172
rect 41230 9160 41236 9172
rect 31720 9132 41236 9160
rect 31720 9120 31726 9132
rect 41230 9120 41236 9132
rect 41288 9120 41294 9172
rect 41322 9120 41328 9172
rect 41380 9160 41386 9172
rect 42886 9160 42892 9172
rect 41380 9132 42892 9160
rect 41380 9120 41386 9132
rect 42886 9120 42892 9132
rect 42944 9120 42950 9172
rect 43806 9120 43812 9172
rect 43864 9160 43870 9172
rect 44361 9163 44419 9169
rect 44361 9160 44373 9163
rect 43864 9132 44373 9160
rect 43864 9120 43870 9132
rect 44361 9129 44373 9132
rect 44407 9129 44419 9163
rect 44361 9123 44419 9129
rect 45094 9120 45100 9172
rect 45152 9160 45158 9172
rect 45189 9163 45247 9169
rect 45189 9160 45201 9163
rect 45152 9132 45201 9160
rect 45152 9120 45158 9132
rect 45189 9129 45201 9132
rect 45235 9129 45247 9163
rect 46198 9160 46204 9172
rect 46159 9132 46204 9160
rect 45189 9123 45247 9129
rect 46198 9120 46204 9132
rect 46256 9120 46262 9172
rect 46290 9120 46296 9172
rect 46348 9160 46354 9172
rect 49418 9160 49424 9172
rect 46348 9132 49424 9160
rect 46348 9120 46354 9132
rect 49418 9120 49424 9132
rect 49476 9120 49482 9172
rect 49789 9163 49847 9169
rect 49789 9129 49801 9163
rect 49835 9160 49847 9163
rect 50614 9160 50620 9172
rect 49835 9132 50620 9160
rect 49835 9129 49847 9132
rect 49789 9123 49847 9129
rect 50614 9120 50620 9132
rect 50672 9120 50678 9172
rect 55214 9160 55220 9172
rect 51460 9132 55220 9160
rect 16816 9064 17908 9092
rect 16816 9052 16822 9064
rect 18046 9052 18052 9104
rect 18104 9092 18110 9104
rect 21453 9095 21511 9101
rect 18104 9064 19104 9092
rect 18104 9052 18110 9064
rect 11296 8996 12204 9024
rect 12253 9027 12311 9033
rect 11296 8984 11302 8996
rect 12253 8993 12265 9027
rect 12299 9024 12311 9027
rect 12526 9024 12532 9036
rect 12299 8996 12532 9024
rect 12299 8993 12311 8996
rect 12253 8987 12311 8993
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 13538 9024 13544 9036
rect 12636 8996 13544 9024
rect 2498 8956 2504 8968
rect 2459 8928 2504 8956
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 3234 8956 3240 8968
rect 3147 8928 3240 8956
rect 3234 8916 3240 8928
rect 3292 8956 3298 8968
rect 4062 8956 4068 8968
rect 3292 8928 4068 8956
rect 3292 8916 3298 8928
rect 4062 8916 4068 8928
rect 4120 8916 4126 8968
rect 4430 8956 4436 8968
rect 4391 8928 4436 8956
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 4706 8916 4712 8968
rect 4764 8956 4770 8968
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 4764 8928 6009 8956
rect 4764 8916 4770 8928
rect 5997 8925 6009 8928
rect 6043 8925 6055 8959
rect 8294 8956 8300 8968
rect 7406 8928 8300 8956
rect 5997 8919 6055 8925
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 9493 8959 9551 8965
rect 9493 8925 9505 8959
rect 9539 8956 9551 8959
rect 10502 8956 10508 8968
rect 9539 8928 10508 8956
rect 9539 8925 9551 8928
rect 9493 8919 9551 8925
rect 10502 8916 10508 8928
rect 10560 8916 10566 8968
rect 10870 8916 10876 8968
rect 10928 8916 10934 8968
rect 6270 8888 6276 8900
rect 6231 8860 6276 8888
rect 6270 8848 6276 8860
rect 6328 8848 6334 8900
rect 11977 8891 12035 8897
rect 7576 8860 9168 8888
rect 2130 8780 2136 8832
rect 2188 8820 2194 8832
rect 5534 8820 5540 8832
rect 2188 8792 5540 8820
rect 2188 8780 2194 8792
rect 5534 8780 5540 8792
rect 5592 8780 5598 8832
rect 7098 8780 7104 8832
rect 7156 8820 7162 8832
rect 7576 8820 7604 8860
rect 7156 8792 7604 8820
rect 7156 8780 7162 8792
rect 7650 8780 7656 8832
rect 7708 8820 7714 8832
rect 8570 8820 8576 8832
rect 7708 8792 8576 8820
rect 7708 8780 7714 8792
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 9140 8829 9168 8860
rect 11977 8857 11989 8891
rect 12023 8888 12035 8891
rect 12636 8888 12664 8996
rect 13538 8984 13544 8996
rect 13596 8984 13602 9036
rect 13725 9027 13783 9033
rect 13725 8993 13737 9027
rect 13771 9024 13783 9027
rect 15102 9024 15108 9036
rect 13771 8996 15108 9024
rect 13771 8993 13783 8996
rect 13725 8987 13783 8993
rect 15102 8984 15108 8996
rect 15160 8984 15166 9036
rect 16500 8996 16534 9036
rect 16528 8984 16534 8996
rect 16586 9024 16592 9036
rect 16586 8996 16633 9024
rect 16586 8984 16592 8996
rect 16666 8984 16672 9036
rect 16724 9024 16730 9036
rect 16942 9024 16948 9036
rect 16724 8996 16948 9024
rect 16724 8984 16730 8996
rect 16942 8984 16948 8996
rect 17000 9024 17006 9036
rect 17037 9027 17095 9033
rect 17037 9024 17049 9027
rect 17000 8996 17049 9024
rect 17000 8984 17006 8996
rect 17037 8993 17049 8996
rect 17083 8993 17095 9027
rect 17586 9024 17592 9036
rect 17499 8996 17592 9024
rect 17037 8987 17095 8993
rect 12713 8959 12771 8965
rect 12713 8925 12725 8959
rect 12759 8925 12771 8959
rect 12713 8919 12771 8925
rect 12989 8959 13047 8965
rect 12989 8925 13001 8959
rect 13035 8956 13047 8959
rect 13814 8956 13820 8968
rect 13035 8928 13820 8956
rect 13035 8925 13047 8928
rect 12989 8919 13047 8925
rect 12023 8860 12664 8888
rect 12023 8857 12035 8860
rect 11977 8851 12035 8857
rect 9125 8823 9183 8829
rect 9125 8789 9137 8823
rect 9171 8789 9183 8823
rect 9125 8783 9183 8789
rect 10505 8823 10563 8829
rect 10505 8789 10517 8823
rect 10551 8820 10563 8823
rect 12728 8820 12756 8919
rect 13556 8900 13584 8928
rect 13814 8916 13820 8928
rect 13872 8916 13878 8968
rect 14553 8959 14611 8965
rect 14553 8925 14565 8959
rect 14599 8925 14611 8959
rect 14553 8919 14611 8925
rect 14737 8959 14795 8965
rect 14737 8925 14749 8959
rect 14783 8925 14795 8959
rect 16114 8956 16120 8968
rect 16075 8928 16120 8956
rect 14737 8919 14795 8925
rect 13538 8848 13544 8900
rect 13596 8848 13602 8900
rect 10551 8792 12756 8820
rect 14568 8820 14596 8919
rect 14752 8888 14780 8919
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 16301 8959 16359 8965
rect 16301 8925 16313 8959
rect 16347 8956 16359 8959
rect 16758 8956 16764 8968
rect 16347 8928 16764 8956
rect 16347 8925 16359 8928
rect 16301 8919 16359 8925
rect 16758 8916 16764 8928
rect 16816 8916 16822 8968
rect 16850 8916 16856 8968
rect 16908 8956 16914 8968
rect 16908 8928 16953 8956
rect 16908 8916 16914 8928
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 17512 8965 17540 8996
rect 17586 8984 17592 8996
rect 17644 9024 17650 9036
rect 17644 8996 18552 9024
rect 17644 8984 17650 8996
rect 17497 8959 17555 8965
rect 17497 8956 17509 8959
rect 17368 8928 17509 8956
rect 17368 8916 17374 8928
rect 17497 8925 17509 8928
rect 17543 8925 17555 8959
rect 17497 8919 17555 8925
rect 17681 8959 17739 8965
rect 17681 8925 17693 8959
rect 17727 8956 17739 8959
rect 18046 8956 18052 8968
rect 17727 8928 18052 8956
rect 17727 8925 17739 8928
rect 17681 8919 17739 8925
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 16666 8888 16672 8900
rect 14752 8860 16672 8888
rect 16666 8848 16672 8860
rect 16724 8848 16730 8900
rect 18322 8888 18328 8900
rect 17512 8860 17954 8888
rect 18283 8860 18328 8888
rect 15286 8820 15292 8832
rect 14568 8792 15292 8820
rect 10551 8789 10563 8792
rect 10505 8783 10563 8789
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 15838 8780 15844 8832
rect 15896 8820 15902 8832
rect 17512 8820 17540 8860
rect 15896 8792 17540 8820
rect 17926 8820 17954 8860
rect 18322 8848 18328 8860
rect 18380 8848 18386 8900
rect 18414 8820 18420 8832
rect 17926 8792 18420 8820
rect 15896 8780 15902 8792
rect 18414 8780 18420 8792
rect 18472 8780 18478 8832
rect 18524 8829 18552 8996
rect 19076 8956 19104 9064
rect 19628 9064 20668 9092
rect 19150 8984 19156 9036
rect 19208 9024 19214 9036
rect 19521 9027 19579 9033
rect 19521 9024 19533 9027
rect 19208 8996 19533 9024
rect 19208 8984 19214 8996
rect 19521 8993 19533 8996
rect 19567 8993 19579 9027
rect 19521 8987 19579 8993
rect 19628 8968 19656 9064
rect 20530 9024 20536 9036
rect 20491 8996 20536 9024
rect 20530 8984 20536 8996
rect 20588 8984 20594 9036
rect 20640 9024 20668 9064
rect 21453 9061 21465 9095
rect 21499 9061 21511 9095
rect 21453 9055 21511 9061
rect 24765 9095 24823 9101
rect 24765 9061 24777 9095
rect 24811 9092 24823 9095
rect 25314 9092 25320 9104
rect 24811 9064 25320 9092
rect 24811 9061 24823 9064
rect 24765 9055 24823 9061
rect 21468 9024 21496 9055
rect 25314 9052 25320 9064
rect 25372 9052 25378 9104
rect 27062 9052 27068 9104
rect 27120 9092 27126 9104
rect 27120 9064 28994 9092
rect 27120 9052 27126 9064
rect 22094 9024 22100 9036
rect 20640 8996 21496 9024
rect 21652 8996 22100 9024
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 19076 8928 19441 8956
rect 19429 8925 19441 8928
rect 19475 8956 19487 8959
rect 19610 8956 19616 8968
rect 19475 8928 19616 8956
rect 19475 8925 19487 8928
rect 19429 8919 19487 8925
rect 19610 8916 19616 8928
rect 19668 8916 19674 8968
rect 19702 8916 19708 8968
rect 19760 8956 19766 8968
rect 20622 8956 20628 8968
rect 19760 8928 20628 8956
rect 19760 8916 19766 8928
rect 20622 8916 20628 8928
rect 20680 8916 20686 8968
rect 20714 8916 20720 8968
rect 20772 8956 20778 8968
rect 21652 8965 21680 8996
rect 22094 8984 22100 8996
rect 22152 8984 22158 9036
rect 22186 8984 22192 9036
rect 22244 9024 22250 9036
rect 25038 9024 25044 9036
rect 22244 8996 25044 9024
rect 22244 8984 22250 8996
rect 25038 8984 25044 8996
rect 25096 8984 25102 9036
rect 25774 9024 25780 9036
rect 25735 8996 25780 9024
rect 25774 8984 25780 8996
rect 25832 8984 25838 9036
rect 26053 9027 26111 9033
rect 26053 8993 26065 9027
rect 26099 9024 26111 9027
rect 28534 9024 28540 9036
rect 26099 8996 28304 9024
rect 28495 8996 28540 9024
rect 26099 8993 26111 8996
rect 26053 8987 26111 8993
rect 21637 8959 21695 8965
rect 21637 8956 21649 8959
rect 20772 8928 21649 8956
rect 20772 8916 20778 8928
rect 21637 8925 21649 8928
rect 21683 8925 21695 8959
rect 21637 8919 21695 8925
rect 21729 8959 21787 8965
rect 21729 8925 21741 8959
rect 21775 8956 21787 8959
rect 22370 8956 22376 8968
rect 21775 8928 22376 8956
rect 21775 8925 21787 8928
rect 21729 8919 21787 8925
rect 18690 8848 18696 8900
rect 18748 8888 18754 8900
rect 19518 8888 19524 8900
rect 18748 8860 19524 8888
rect 18748 8848 18754 8860
rect 19518 8848 19524 8860
rect 19576 8848 19582 8900
rect 19794 8848 19800 8900
rect 19852 8888 19858 8900
rect 21744 8888 21772 8919
rect 22370 8916 22376 8928
rect 22428 8916 22434 8968
rect 22554 8956 22560 8968
rect 22515 8928 22560 8956
rect 22554 8916 22560 8928
rect 22612 8916 22618 8968
rect 21910 8888 21916 8900
rect 19852 8860 21772 8888
rect 21871 8860 21916 8888
rect 19852 8848 19858 8860
rect 21910 8848 21916 8860
rect 21968 8848 21974 8900
rect 26510 8848 26516 8900
rect 26568 8848 26574 8900
rect 27801 8891 27859 8897
rect 27801 8857 27813 8891
rect 27847 8857 27859 8891
rect 28276 8888 28304 8996
rect 28534 8984 28540 8996
rect 28592 8984 28598 9036
rect 28442 8956 28448 8968
rect 28403 8928 28448 8956
rect 28442 8916 28448 8928
rect 28500 8916 28506 8968
rect 28966 8956 28994 9064
rect 29730 9052 29736 9104
rect 29788 9092 29794 9104
rect 31021 9095 31079 9101
rect 31021 9092 31033 9095
rect 29788 9064 31033 9092
rect 29788 9052 29794 9064
rect 31021 9061 31033 9064
rect 31067 9092 31079 9095
rect 31478 9092 31484 9104
rect 31067 9064 31484 9092
rect 31067 9061 31079 9064
rect 31021 9055 31079 9061
rect 31478 9052 31484 9064
rect 31536 9052 31542 9104
rect 33226 9052 33232 9104
rect 33284 9092 33290 9104
rect 36633 9095 36691 9101
rect 33284 9064 35020 9092
rect 33284 9052 33290 9064
rect 29914 8984 29920 9036
rect 29972 9024 29978 9036
rect 31573 9027 31631 9033
rect 31573 9024 31585 9027
rect 29972 8996 31585 9024
rect 29972 8984 29978 8996
rect 31573 8993 31585 8996
rect 31619 9024 31631 9027
rect 32490 9024 32496 9036
rect 31619 8996 32496 9024
rect 31619 8993 31631 8996
rect 31573 8987 31631 8993
rect 32490 8984 32496 8996
rect 32548 9024 32554 9036
rect 34885 9027 34943 9033
rect 34885 9024 34897 9027
rect 32548 8996 34897 9024
rect 32548 8984 32554 8996
rect 34885 8993 34897 8996
rect 34931 8993 34943 9027
rect 34992 9024 35020 9064
rect 36633 9061 36645 9095
rect 36679 9092 36691 9095
rect 38838 9092 38844 9104
rect 36679 9064 38844 9092
rect 36679 9061 36691 9064
rect 36633 9055 36691 9061
rect 38838 9052 38844 9064
rect 38896 9052 38902 9104
rect 41506 9092 41512 9104
rect 38948 9064 41512 9092
rect 37645 9027 37703 9033
rect 34992 8996 37504 9024
rect 34885 8987 34943 8993
rect 28966 8928 31616 8956
rect 31478 8888 31484 8900
rect 28276 8860 31484 8888
rect 27801 8851 27859 8857
rect 18509 8823 18567 8829
rect 18509 8789 18521 8823
rect 18555 8820 18567 8823
rect 19702 8820 19708 8832
rect 18555 8792 19708 8820
rect 18555 8789 18567 8792
rect 18509 8783 18567 8789
rect 19702 8780 19708 8792
rect 19760 8780 19766 8832
rect 20254 8780 20260 8832
rect 20312 8820 20318 8832
rect 22373 8823 22431 8829
rect 22373 8820 22385 8823
rect 20312 8792 22385 8820
rect 20312 8780 20318 8792
rect 22373 8789 22385 8792
rect 22419 8789 22431 8823
rect 22373 8783 22431 8789
rect 22646 8780 22652 8832
rect 22704 8820 22710 8832
rect 23109 8823 23167 8829
rect 23109 8820 23121 8823
rect 22704 8792 23121 8820
rect 22704 8780 22710 8792
rect 23109 8789 23121 8792
rect 23155 8820 23167 8823
rect 27062 8820 27068 8832
rect 23155 8792 27068 8820
rect 23155 8789 23167 8792
rect 23109 8783 23167 8789
rect 27062 8780 27068 8792
rect 27120 8780 27126 8832
rect 27816 8820 27844 8851
rect 31478 8848 31484 8860
rect 31536 8848 31542 8900
rect 31588 8888 31616 8928
rect 32858 8916 32864 8968
rect 32916 8956 32922 8968
rect 33502 8956 33508 8968
rect 32916 8928 33508 8956
rect 32916 8916 32922 8928
rect 33502 8916 33508 8928
rect 33560 8916 33566 8968
rect 33686 8916 33692 8968
rect 33744 8956 33750 8968
rect 33962 8956 33968 8968
rect 33744 8928 33968 8956
rect 33744 8916 33750 8928
rect 33962 8916 33968 8928
rect 34020 8956 34026 8968
rect 34057 8959 34115 8965
rect 34057 8956 34069 8959
rect 34020 8928 34069 8956
rect 34020 8916 34026 8928
rect 34057 8925 34069 8928
rect 34103 8925 34115 8959
rect 34330 8956 34336 8968
rect 34291 8928 34336 8956
rect 34057 8919 34115 8925
rect 34330 8916 34336 8928
rect 34388 8916 34394 8968
rect 31754 8888 31760 8900
rect 31588 8860 31760 8888
rect 31754 8848 31760 8860
rect 31812 8848 31818 8900
rect 31849 8891 31907 8897
rect 31849 8857 31861 8891
rect 31895 8857 31907 8891
rect 34514 8888 34520 8900
rect 31849 8851 31907 8857
rect 33152 8860 34520 8888
rect 28718 8820 28724 8832
rect 27816 8792 28724 8820
rect 28718 8780 28724 8792
rect 28776 8780 28782 8832
rect 28813 8823 28871 8829
rect 28813 8789 28825 8823
rect 28859 8820 28871 8823
rect 29638 8820 29644 8832
rect 28859 8792 29644 8820
rect 28859 8789 28871 8792
rect 28813 8783 28871 8789
rect 29638 8780 29644 8792
rect 29696 8780 29702 8832
rect 30006 8780 30012 8832
rect 30064 8820 30070 8832
rect 30469 8823 30527 8829
rect 30469 8820 30481 8823
rect 30064 8792 30481 8820
rect 30064 8780 30070 8792
rect 30469 8789 30481 8792
rect 30515 8820 30527 8823
rect 31662 8820 31668 8832
rect 30515 8792 31668 8820
rect 30515 8789 30527 8792
rect 30469 8783 30527 8789
rect 31662 8780 31668 8792
rect 31720 8780 31726 8832
rect 31864 8820 31892 8851
rect 33152 8820 33180 8860
rect 34514 8848 34520 8860
rect 34572 8848 34578 8900
rect 35158 8888 35164 8900
rect 35119 8860 35164 8888
rect 35158 8848 35164 8860
rect 35216 8848 35222 8900
rect 35618 8848 35624 8900
rect 35676 8848 35682 8900
rect 36814 8848 36820 8900
rect 36872 8888 36878 8900
rect 37476 8888 37504 8996
rect 37645 8993 37657 9027
rect 37691 9024 37703 9027
rect 38289 9027 38347 9033
rect 38289 9024 38301 9027
rect 37691 8996 38301 9024
rect 37691 8993 37703 8996
rect 37645 8987 37703 8993
rect 38289 8993 38301 8996
rect 38335 8993 38347 9027
rect 38289 8987 38347 8993
rect 37550 8916 37556 8968
rect 37608 8956 37614 8968
rect 37608 8928 37653 8956
rect 37608 8916 37614 8928
rect 38102 8916 38108 8968
rect 38160 8956 38166 8968
rect 38197 8959 38255 8965
rect 38197 8956 38209 8959
rect 38160 8928 38209 8956
rect 38160 8916 38166 8928
rect 38197 8925 38209 8928
rect 38243 8925 38255 8959
rect 38378 8956 38384 8968
rect 38339 8928 38384 8956
rect 38197 8919 38255 8925
rect 38378 8916 38384 8928
rect 38436 8916 38442 8968
rect 38948 8888 38976 9064
rect 41506 9052 41512 9064
rect 41564 9052 41570 9104
rect 41598 9052 41604 9104
rect 41656 9092 41662 9104
rect 43530 9092 43536 9104
rect 41656 9064 43536 9092
rect 41656 9052 41662 9064
rect 43530 9052 43536 9064
rect 43588 9052 43594 9104
rect 51460 9092 51488 9132
rect 55214 9120 55220 9132
rect 55272 9120 55278 9172
rect 56134 9120 56140 9172
rect 56192 9160 56198 9172
rect 57882 9160 57888 9172
rect 56192 9132 57888 9160
rect 56192 9120 56198 9132
rect 57882 9120 57888 9132
rect 57940 9120 57946 9172
rect 58158 9120 58164 9172
rect 58216 9160 58222 9172
rect 58986 9160 58992 9172
rect 58216 9132 58992 9160
rect 58216 9120 58222 9132
rect 58986 9120 58992 9132
rect 59044 9120 59050 9172
rect 59909 9163 59967 9169
rect 59909 9129 59921 9163
rect 59955 9160 59967 9163
rect 62390 9160 62396 9172
rect 59955 9132 62396 9160
rect 59955 9129 59967 9132
rect 59909 9123 59967 9129
rect 62390 9120 62396 9132
rect 62448 9120 62454 9172
rect 67266 9120 67272 9172
rect 67324 9160 67330 9172
rect 70210 9160 70216 9172
rect 67324 9132 70216 9160
rect 67324 9120 67330 9132
rect 70210 9120 70216 9132
rect 70268 9120 70274 9172
rect 70302 9120 70308 9172
rect 70360 9160 70366 9172
rect 71038 9160 71044 9172
rect 70360 9132 71044 9160
rect 70360 9120 70366 9132
rect 71038 9120 71044 9132
rect 71096 9120 71102 9172
rect 71590 9120 71596 9172
rect 71648 9160 71654 9172
rect 71685 9163 71743 9169
rect 71685 9160 71697 9163
rect 71648 9132 71697 9160
rect 71648 9120 71654 9132
rect 71685 9129 71697 9132
rect 71731 9129 71743 9163
rect 74810 9160 74816 9172
rect 71685 9123 71743 9129
rect 73172 9132 74816 9160
rect 52454 9092 52460 9104
rect 43640 9064 51488 9092
rect 51552 9064 52460 9092
rect 39298 9024 39304 9036
rect 39259 8996 39304 9024
rect 39298 8984 39304 8996
rect 39356 8984 39362 9036
rect 39758 8984 39764 9036
rect 39816 9024 39822 9036
rect 43349 9027 43407 9033
rect 39816 8996 40816 9024
rect 39816 8984 39822 8996
rect 39022 8916 39028 8968
rect 39080 8956 39086 8968
rect 39209 8959 39267 8965
rect 39209 8956 39221 8959
rect 39080 8928 39221 8956
rect 39080 8916 39086 8928
rect 39209 8925 39221 8928
rect 39255 8925 39267 8959
rect 40494 8956 40500 8968
rect 40455 8928 40500 8956
rect 39209 8919 39267 8925
rect 36872 8860 37412 8888
rect 37476 8860 38976 8888
rect 39224 8888 39252 8919
rect 40494 8916 40500 8928
rect 40552 8916 40558 8968
rect 40678 8956 40684 8968
rect 40639 8928 40684 8956
rect 40678 8916 40684 8928
rect 40736 8916 40742 8968
rect 40788 8956 40816 8996
rect 43349 8993 43361 9027
rect 43395 9024 43407 9027
rect 43438 9024 43444 9036
rect 43395 8996 43444 9024
rect 43395 8993 43407 8996
rect 43349 8987 43407 8993
rect 43438 8984 43444 8996
rect 43496 8984 43502 9036
rect 43640 9033 43668 9064
rect 43625 9027 43683 9033
rect 43625 8993 43637 9027
rect 43671 8993 43683 9027
rect 44266 9024 44272 9036
rect 44227 8996 44272 9024
rect 43625 8987 43683 8993
rect 44266 8984 44272 8996
rect 44324 8984 44330 9036
rect 49050 9024 49056 9036
rect 45388 8996 46520 9024
rect 40788 8928 42380 8956
rect 41598 8888 41604 8900
rect 39224 8860 41604 8888
rect 36872 8848 36878 8860
rect 33318 8820 33324 8832
rect 31864 8792 33180 8820
rect 33279 8792 33324 8820
rect 33318 8780 33324 8792
rect 33376 8780 33382 8832
rect 33870 8820 33876 8832
rect 33831 8792 33876 8820
rect 33870 8780 33876 8792
rect 33928 8780 33934 8832
rect 34146 8780 34152 8832
rect 34204 8820 34210 8832
rect 34241 8823 34299 8829
rect 34241 8820 34253 8823
rect 34204 8792 34253 8820
rect 34204 8780 34210 8792
rect 34241 8789 34253 8792
rect 34287 8789 34299 8823
rect 34241 8783 34299 8789
rect 34882 8780 34888 8832
rect 34940 8820 34946 8832
rect 36722 8820 36728 8832
rect 34940 8792 36728 8820
rect 34940 8780 34946 8792
rect 36722 8780 36728 8792
rect 36780 8780 36786 8832
rect 37182 8820 37188 8832
rect 37143 8792 37188 8820
rect 37182 8780 37188 8792
rect 37240 8780 37246 8832
rect 37384 8820 37412 8860
rect 41598 8848 41604 8860
rect 41656 8848 41662 8900
rect 38654 8820 38660 8832
rect 37384 8792 38660 8820
rect 38654 8780 38660 8792
rect 38712 8780 38718 8832
rect 38838 8820 38844 8832
rect 38799 8792 38844 8820
rect 38838 8780 38844 8792
rect 38896 8780 38902 8832
rect 40681 8823 40739 8829
rect 40681 8789 40693 8823
rect 40727 8820 40739 8823
rect 40954 8820 40960 8832
rect 40727 8792 40960 8820
rect 40727 8789 40739 8792
rect 40681 8783 40739 8789
rect 40954 8780 40960 8792
rect 41012 8780 41018 8832
rect 41414 8780 41420 8832
rect 41472 8820 41478 8832
rect 42352 8820 42380 8928
rect 43806 8916 43812 8968
rect 43864 8956 43870 8968
rect 43864 8928 43909 8956
rect 43864 8916 43870 8928
rect 44450 8916 44456 8968
rect 44508 8956 44514 8968
rect 44545 8959 44603 8965
rect 44545 8956 44557 8959
rect 44508 8928 44557 8956
rect 44508 8916 44514 8928
rect 44545 8925 44557 8928
rect 44591 8925 44603 8959
rect 44545 8919 44603 8925
rect 44637 8959 44695 8965
rect 44637 8925 44649 8959
rect 44683 8956 44695 8959
rect 44726 8956 44732 8968
rect 44683 8928 44732 8956
rect 44683 8925 44695 8928
rect 44637 8919 44695 8925
rect 44726 8916 44732 8928
rect 44784 8956 44790 8968
rect 45186 8956 45192 8968
rect 44784 8928 45192 8956
rect 44784 8916 44790 8928
rect 45186 8916 45192 8928
rect 45244 8916 45250 8968
rect 45388 8965 45416 8996
rect 45373 8959 45431 8965
rect 45373 8925 45385 8959
rect 45419 8925 45431 8959
rect 45373 8919 45431 8925
rect 45462 8916 45468 8968
rect 45520 8956 45526 8968
rect 45646 8956 45652 8968
rect 45520 8928 45565 8956
rect 45607 8928 45652 8956
rect 45520 8916 45526 8928
rect 45646 8916 45652 8928
rect 45704 8916 45710 8968
rect 45741 8959 45799 8965
rect 45741 8925 45753 8959
rect 45787 8956 45799 8959
rect 46198 8956 46204 8968
rect 45787 8928 46204 8956
rect 45787 8925 45799 8928
rect 45741 8919 45799 8925
rect 46198 8916 46204 8928
rect 46256 8916 46262 8968
rect 46382 8956 46388 8968
rect 46343 8928 46388 8956
rect 46382 8916 46388 8928
rect 46440 8916 46446 8968
rect 46492 8956 46520 8996
rect 46860 8996 49056 9024
rect 46661 8959 46719 8965
rect 46661 8956 46673 8959
rect 46492 8928 46673 8956
rect 46661 8925 46673 8928
rect 46707 8956 46719 8959
rect 46860 8956 46888 8996
rect 49050 8984 49056 8996
rect 49108 8984 49114 9036
rect 50706 8984 50712 9036
rect 50764 9024 50770 9036
rect 51552 9024 51580 9064
rect 52454 9052 52460 9064
rect 52512 9052 52518 9104
rect 58526 9092 58532 9104
rect 53944 9064 58532 9092
rect 53944 9033 53972 9064
rect 58526 9052 58532 9064
rect 58584 9092 58590 9104
rect 59630 9092 59636 9104
rect 58584 9064 59636 9092
rect 58584 9052 58590 9064
rect 59630 9052 59636 9064
rect 59688 9052 59694 9104
rect 60090 9052 60096 9104
rect 60148 9092 60154 9104
rect 61286 9092 61292 9104
rect 60148 9064 61292 9092
rect 60148 9052 60154 9064
rect 61286 9052 61292 9064
rect 61344 9052 61350 9104
rect 61746 9052 61752 9104
rect 61804 9092 61810 9104
rect 64693 9095 64751 9101
rect 64693 9092 64705 9095
rect 61804 9064 64705 9092
rect 61804 9052 61810 9064
rect 64693 9061 64705 9064
rect 64739 9092 64751 9095
rect 66714 9092 66720 9104
rect 64739 9064 66720 9092
rect 64739 9061 64751 9064
rect 64693 9055 64751 9061
rect 66714 9052 66720 9064
rect 66772 9092 66778 9104
rect 66772 9064 73108 9092
rect 66772 9052 66778 9064
rect 50764 8996 51580 9024
rect 51629 9027 51687 9033
rect 50764 8984 50770 8996
rect 51629 8993 51641 9027
rect 51675 9024 51687 9027
rect 53745 9027 53803 9033
rect 53745 9024 53757 9027
rect 51675 8996 53757 9024
rect 51675 8993 51687 8996
rect 51629 8987 51687 8993
rect 53745 8993 53757 8996
rect 53791 8993 53803 9027
rect 53745 8987 53803 8993
rect 53929 9027 53987 9033
rect 53929 8993 53941 9027
rect 53975 8993 53987 9027
rect 53929 8987 53987 8993
rect 55766 8984 55772 9036
rect 55824 9024 55830 9036
rect 57333 9027 57391 9033
rect 57333 9024 57345 9027
rect 55824 8996 57345 9024
rect 55824 8984 55830 8996
rect 57333 8993 57345 8996
rect 57379 9024 57391 9027
rect 58618 9024 58624 9036
rect 57379 8996 58624 9024
rect 57379 8993 57391 8996
rect 57333 8987 57391 8993
rect 58618 8984 58624 8996
rect 58676 8984 58682 9036
rect 59906 9024 59912 9036
rect 58728 8996 59912 9024
rect 47394 8956 47400 8968
rect 46707 8928 46888 8956
rect 47355 8928 47400 8956
rect 46707 8925 46719 8928
rect 46661 8919 46719 8925
rect 47394 8916 47400 8928
rect 47452 8916 47458 8968
rect 49786 8916 49792 8968
rect 49844 8956 49850 8968
rect 50614 8956 50620 8968
rect 49844 8928 50620 8956
rect 49844 8916 49850 8928
rect 50614 8916 50620 8928
rect 50672 8956 50678 8968
rect 50801 8959 50859 8965
rect 50801 8956 50813 8959
rect 50672 8928 50813 8956
rect 50672 8916 50678 8928
rect 50801 8925 50813 8928
rect 50847 8925 50859 8959
rect 50801 8919 50859 8925
rect 51261 8959 51319 8965
rect 51261 8925 51273 8959
rect 51307 8956 51319 8959
rect 51442 8956 51448 8968
rect 51307 8928 51448 8956
rect 51307 8925 51319 8928
rect 51261 8919 51319 8925
rect 51442 8916 51448 8928
rect 51500 8916 51506 8968
rect 52089 8959 52147 8965
rect 52089 8925 52101 8959
rect 52135 8956 52147 8959
rect 52270 8956 52276 8968
rect 52135 8928 52276 8956
rect 52135 8925 52147 8928
rect 52089 8919 52147 8925
rect 52270 8916 52276 8928
rect 52328 8916 52334 8968
rect 54573 8959 54631 8965
rect 54573 8925 54585 8959
rect 54619 8956 54631 8959
rect 54938 8956 54944 8968
rect 54619 8928 54944 8956
rect 54619 8925 54631 8928
rect 54573 8919 54631 8925
rect 54938 8916 54944 8928
rect 54996 8916 55002 8968
rect 57793 8959 57851 8965
rect 57793 8925 57805 8959
rect 57839 8925 57851 8959
rect 57793 8919 57851 8925
rect 47578 8888 47584 8900
rect 47539 8860 47584 8888
rect 47578 8848 47584 8860
rect 47636 8848 47642 8900
rect 49237 8891 49295 8897
rect 49237 8857 49249 8891
rect 49283 8888 49295 8891
rect 51350 8888 51356 8900
rect 49283 8860 51356 8888
rect 49283 8857 49295 8860
rect 49237 8851 49295 8857
rect 44358 8820 44364 8832
rect 41472 8792 41517 8820
rect 42352 8792 44364 8820
rect 41472 8780 41478 8792
rect 44358 8780 44364 8792
rect 44416 8780 44422 8832
rect 44453 8823 44511 8829
rect 44453 8789 44465 8823
rect 44499 8820 44511 8823
rect 44910 8820 44916 8832
rect 44499 8792 44916 8820
rect 44499 8789 44511 8792
rect 44453 8783 44511 8789
rect 44910 8780 44916 8792
rect 44968 8780 44974 8832
rect 45462 8780 45468 8832
rect 45520 8820 45526 8832
rect 46566 8820 46572 8832
rect 45520 8792 46572 8820
rect 45520 8780 45526 8792
rect 46566 8780 46572 8792
rect 46624 8780 46630 8832
rect 46750 8780 46756 8832
rect 46808 8820 46814 8832
rect 49252 8820 49280 8851
rect 51350 8848 51356 8860
rect 51408 8848 51414 8900
rect 51552 8860 57560 8888
rect 46808 8792 49280 8820
rect 46808 8780 46814 8792
rect 49418 8780 49424 8832
rect 49476 8820 49482 8832
rect 51552 8820 51580 8860
rect 49476 8792 51580 8820
rect 49476 8780 49482 8792
rect 51626 8780 51632 8832
rect 51684 8820 51690 8832
rect 54481 8823 54539 8829
rect 54481 8820 54493 8823
rect 51684 8792 54493 8820
rect 51684 8780 51690 8792
rect 54481 8789 54493 8792
rect 54527 8789 54539 8823
rect 57532 8820 57560 8860
rect 57606 8848 57612 8900
rect 57664 8888 57670 8900
rect 57664 8860 57709 8888
rect 57664 8848 57670 8860
rect 57808 8820 57836 8919
rect 57882 8916 57888 8968
rect 57940 8956 57946 8968
rect 58345 8959 58403 8965
rect 58345 8956 58357 8959
rect 57940 8928 58357 8956
rect 57940 8916 57946 8928
rect 58345 8925 58357 8928
rect 58391 8956 58403 8959
rect 58728 8956 58756 8996
rect 59906 8984 59912 8996
rect 59964 8984 59970 9036
rect 60642 9024 60648 9036
rect 60603 8996 60648 9024
rect 60642 8984 60648 8996
rect 60700 8984 60706 9036
rect 62114 9024 62120 9036
rect 61120 8996 62120 9024
rect 58894 8956 58900 8968
rect 58391 8928 58756 8956
rect 58855 8928 58900 8956
rect 58391 8925 58403 8928
rect 58345 8919 58403 8925
rect 58894 8916 58900 8928
rect 58952 8916 58958 8968
rect 58989 8959 59047 8965
rect 58989 8925 59001 8959
rect 59035 8956 59047 8959
rect 60016 8956 60136 8958
rect 60918 8956 60924 8968
rect 59035 8930 60924 8956
rect 59035 8928 60044 8930
rect 60108 8928 60924 8930
rect 59035 8925 59047 8928
rect 58989 8919 59047 8925
rect 60918 8916 60924 8928
rect 60976 8916 60982 8968
rect 59630 8848 59636 8900
rect 59688 8888 59694 8900
rect 60093 8891 60151 8897
rect 60093 8888 60105 8891
rect 59688 8860 60105 8888
rect 59688 8848 59694 8860
rect 60093 8857 60105 8860
rect 60139 8888 60151 8891
rect 61120 8888 61148 8996
rect 62114 8984 62120 8996
rect 62172 8984 62178 9036
rect 62298 9024 62304 9036
rect 62259 8996 62304 9024
rect 62298 8984 62304 8996
rect 62356 8984 62362 9036
rect 63494 9024 63500 9036
rect 63455 8996 63500 9024
rect 63494 8984 63500 8996
rect 63552 8984 63558 9036
rect 66162 9024 66168 9036
rect 66123 8996 66168 9024
rect 66162 8984 66168 8996
rect 66220 8984 66226 9036
rect 66254 8984 66260 9036
rect 66312 9024 66318 9036
rect 66441 9027 66499 9033
rect 66441 9024 66453 9027
rect 66312 8996 66453 9024
rect 66312 8984 66318 8996
rect 66441 8993 66453 8996
rect 66487 9024 66499 9027
rect 68186 9024 68192 9036
rect 66487 8996 68192 9024
rect 66487 8993 66499 8996
rect 66441 8987 66499 8993
rect 68186 8984 68192 8996
rect 68244 8984 68250 9036
rect 68462 9024 68468 9036
rect 68423 8996 68468 9024
rect 68462 8984 68468 8996
rect 68520 8984 68526 9036
rect 70854 8984 70860 9036
rect 70912 9024 70918 9036
rect 71041 9027 71099 9033
rect 71041 9024 71053 9027
rect 70912 8996 71053 9024
rect 70912 8984 70918 8996
rect 71041 8993 71053 8996
rect 71087 8993 71099 9027
rect 71041 8987 71099 8993
rect 71406 8984 71412 9036
rect 71464 9024 71470 9036
rect 72694 9024 72700 9036
rect 71464 8996 72700 9024
rect 71464 8984 71470 8996
rect 72694 8984 72700 8996
rect 72752 9024 72758 9036
rect 72752 8996 72924 9024
rect 72752 8984 72758 8996
rect 62485 8959 62543 8965
rect 62485 8925 62497 8959
rect 62531 8925 62543 8959
rect 62485 8919 62543 8925
rect 63589 8959 63647 8965
rect 63589 8925 63601 8959
rect 63635 8956 63647 8959
rect 63770 8956 63776 8968
rect 63635 8928 63776 8956
rect 63635 8925 63647 8928
rect 63589 8919 63647 8925
rect 60139 8860 61148 8888
rect 60139 8857 60151 8860
rect 60093 8851 60151 8857
rect 61286 8848 61292 8900
rect 61344 8888 61350 8900
rect 62500 8888 62528 8919
rect 63770 8916 63776 8928
rect 63828 8916 63834 8968
rect 64230 8956 64236 8968
rect 64191 8928 64236 8956
rect 64230 8916 64236 8928
rect 64288 8916 64294 8968
rect 64322 8916 64328 8968
rect 64380 8956 64386 8968
rect 65981 8959 66039 8965
rect 65981 8956 65993 8959
rect 64380 8928 65993 8956
rect 64380 8916 64386 8928
rect 65981 8925 65993 8928
rect 66027 8925 66039 8959
rect 68281 8959 68339 8965
rect 68281 8956 68293 8959
rect 65981 8919 66039 8925
rect 67560 8950 67680 8956
rect 67744 8950 68293 8956
rect 67560 8928 68293 8950
rect 61344 8860 62528 8888
rect 65996 8888 66024 8919
rect 66530 8888 66536 8900
rect 65996 8860 66536 8888
rect 61344 8848 61350 8860
rect 66530 8848 66536 8860
rect 66588 8848 66594 8900
rect 66990 8848 66996 8900
rect 67048 8888 67054 8900
rect 67560 8888 67588 8928
rect 67652 8922 67772 8928
rect 68281 8925 68293 8928
rect 68327 8925 68339 8959
rect 68281 8919 68339 8925
rect 69934 8916 69940 8968
rect 69992 8956 69998 8968
rect 71133 8959 71191 8965
rect 69992 8928 70900 8956
rect 69992 8916 69998 8928
rect 67048 8860 67588 8888
rect 67048 8848 67054 8860
rect 68186 8848 68192 8900
rect 68244 8888 68250 8900
rect 70121 8891 70179 8897
rect 70121 8888 70133 8891
rect 68244 8860 70133 8888
rect 68244 8848 68250 8860
rect 70121 8857 70133 8860
rect 70167 8888 70179 8891
rect 70762 8888 70768 8900
rect 70167 8860 70768 8888
rect 70167 8857 70179 8860
rect 70121 8851 70179 8857
rect 70762 8848 70768 8860
rect 70820 8848 70826 8900
rect 70872 8888 70900 8928
rect 71133 8925 71145 8959
rect 71179 8956 71191 8959
rect 71682 8956 71688 8968
rect 71179 8928 71688 8956
rect 71179 8925 71191 8928
rect 71133 8919 71191 8925
rect 71682 8916 71688 8928
rect 71740 8916 71746 8968
rect 71774 8916 71780 8968
rect 71832 8956 71838 8968
rect 72896 8965 72924 8996
rect 72881 8959 72939 8965
rect 71832 8928 72740 8956
rect 71832 8916 71838 8928
rect 72237 8891 72295 8897
rect 72237 8888 72249 8891
rect 70872 8860 72249 8888
rect 72237 8857 72249 8860
rect 72283 8857 72295 8891
rect 72712 8888 72740 8928
rect 72881 8925 72893 8959
rect 72927 8925 72939 8959
rect 73080 8956 73108 9064
rect 73172 9033 73200 9132
rect 74810 9120 74816 9132
rect 74868 9120 74874 9172
rect 77021 9163 77079 9169
rect 77021 9129 77033 9163
rect 77067 9160 77079 9163
rect 77386 9160 77392 9172
rect 77067 9132 77392 9160
rect 77067 9129 77079 9132
rect 77021 9123 77079 9129
rect 77386 9120 77392 9132
rect 77444 9120 77450 9172
rect 77496 9132 78904 9160
rect 76650 9092 76656 9104
rect 75104 9064 76656 9092
rect 73157 9027 73215 9033
rect 73157 8993 73169 9027
rect 73203 8993 73215 9027
rect 74074 9024 74080 9036
rect 74035 8996 74080 9024
rect 73157 8987 73215 8993
rect 74074 8984 74080 8996
rect 74132 8984 74138 9036
rect 74534 8984 74540 9036
rect 74592 9024 74598 9036
rect 75104 9024 75132 9064
rect 76650 9052 76656 9064
rect 76708 9052 76714 9104
rect 74592 8996 75132 9024
rect 74592 8984 74598 8996
rect 75270 8984 75276 9036
rect 75328 9024 75334 9036
rect 76190 9024 76196 9036
rect 75328 8996 76196 9024
rect 75328 8984 75334 8996
rect 76190 8984 76196 8996
rect 76248 9024 76254 9036
rect 76248 8996 76696 9024
rect 76248 8984 76254 8996
rect 73798 8956 73804 8968
rect 73080 8928 73660 8956
rect 73759 8928 73804 8956
rect 72881 8919 72939 8925
rect 73062 8888 73068 8900
rect 72712 8860 73068 8888
rect 72237 8851 72295 8857
rect 73062 8848 73068 8860
rect 73120 8848 73126 8900
rect 73632 8888 73660 8928
rect 73798 8916 73804 8928
rect 73856 8916 73862 8968
rect 75178 8916 75184 8968
rect 75236 8916 75242 8968
rect 76377 8959 76435 8965
rect 76377 8925 76389 8959
rect 76423 8956 76435 8959
rect 76558 8956 76564 8968
rect 76423 8928 76564 8956
rect 76423 8925 76435 8928
rect 76377 8919 76435 8925
rect 76558 8916 76564 8928
rect 76616 8916 76622 8968
rect 76668 8956 76696 8996
rect 76926 8956 76932 8968
rect 76668 8928 76932 8956
rect 76926 8916 76932 8928
rect 76984 8916 76990 8968
rect 74350 8888 74356 8900
rect 73632 8860 74356 8888
rect 74350 8848 74356 8860
rect 74408 8848 74414 8900
rect 77496 8888 77524 9132
rect 78876 9092 78904 9132
rect 79134 9120 79140 9172
rect 79192 9160 79198 9172
rect 79321 9163 79379 9169
rect 79321 9160 79333 9163
rect 79192 9132 79333 9160
rect 79192 9120 79198 9132
rect 79321 9129 79333 9132
rect 79367 9129 79379 9163
rect 79321 9123 79379 9129
rect 79410 9120 79416 9172
rect 79468 9160 79474 9172
rect 79468 9132 83688 9160
rect 79468 9120 79474 9132
rect 80606 9092 80612 9104
rect 78876 9064 80612 9092
rect 80606 9052 80612 9064
rect 80664 9052 80670 9104
rect 83660 9092 83688 9132
rect 85666 9120 85672 9172
rect 85724 9160 85730 9172
rect 86586 9160 86592 9172
rect 85724 9132 86592 9160
rect 85724 9120 85730 9132
rect 86586 9120 86592 9132
rect 86644 9120 86650 9172
rect 88058 9120 88064 9172
rect 88116 9160 88122 9172
rect 88426 9160 88432 9172
rect 88116 9132 88432 9160
rect 88116 9120 88122 9132
rect 88426 9120 88432 9132
rect 88484 9120 88490 9172
rect 93946 9160 93952 9172
rect 93907 9132 93952 9160
rect 93946 9120 93952 9132
rect 94004 9120 94010 9172
rect 87230 9092 87236 9104
rect 83660 9064 87236 9092
rect 87230 9052 87236 9064
rect 87288 9052 87294 9104
rect 94130 9092 94136 9104
rect 87340 9064 89714 9092
rect 77846 9024 77852 9036
rect 77807 8996 77852 9024
rect 77846 8984 77852 8996
rect 77904 8984 77910 9036
rect 77938 8984 77944 9036
rect 77996 9024 78002 9036
rect 84013 9027 84071 9033
rect 77996 8996 83964 9024
rect 77996 8984 78002 8996
rect 83936 8990 83964 8996
rect 84013 8993 84025 9027
rect 84059 8993 84071 9027
rect 84013 8990 84071 8993
rect 83936 8987 84071 8990
rect 77573 8959 77631 8965
rect 77573 8925 77585 8959
rect 77619 8925 77631 8959
rect 77573 8919 77631 8925
rect 75380 8860 77524 8888
rect 77588 8888 77616 8919
rect 79134 8916 79140 8968
rect 79192 8956 79198 8968
rect 79965 8959 80023 8965
rect 79965 8956 79977 8959
rect 79192 8928 79977 8956
rect 79192 8916 79198 8928
rect 79965 8925 79977 8928
rect 80011 8925 80023 8959
rect 79965 8919 80023 8925
rect 80514 8916 80520 8968
rect 80572 8958 80578 8968
rect 80572 8930 80615 8958
rect 81250 8956 81256 8968
rect 80572 8916 80578 8930
rect 81211 8928 81256 8956
rect 81250 8916 81256 8928
rect 81308 8916 81314 8968
rect 83936 8962 84044 8987
rect 86034 8984 86040 9036
rect 86092 9024 86098 9036
rect 87340 9024 87368 9064
rect 88150 9024 88156 9036
rect 86092 8996 87368 9024
rect 88111 8996 88156 9024
rect 86092 8984 86098 8996
rect 88150 8984 88156 8996
rect 88208 8984 88214 9036
rect 88426 9024 88432 9036
rect 88387 8996 88432 9024
rect 88426 8984 88432 8996
rect 88484 8984 88490 9036
rect 89686 9024 89714 9064
rect 90836 9064 94136 9092
rect 89806 9024 89812 9036
rect 89686 8996 89812 9024
rect 89806 8984 89812 8996
rect 89864 9024 89870 9036
rect 90836 9033 90864 9064
rect 94130 9052 94136 9064
rect 94188 9052 94194 9104
rect 90821 9027 90879 9033
rect 90821 9024 90833 9027
rect 89864 8996 90833 9024
rect 89864 8984 89870 8996
rect 90821 8993 90833 8996
rect 90867 8993 90879 9027
rect 93210 9024 93216 9036
rect 93171 8996 93216 9024
rect 90821 8987 90879 8993
rect 93210 8984 93216 8996
rect 93268 8984 93274 9036
rect 86494 8956 86500 8968
rect 86455 8928 86500 8956
rect 86494 8916 86500 8928
rect 86552 8916 86558 8968
rect 86865 8959 86923 8965
rect 86865 8925 86877 8959
rect 86911 8956 86923 8959
rect 87690 8956 87696 8968
rect 86911 8928 87696 8956
rect 86911 8925 86923 8928
rect 86865 8919 86923 8925
rect 87690 8916 87696 8928
rect 87748 8916 87754 8968
rect 87874 8916 87880 8968
rect 87932 8956 87938 8968
rect 87969 8959 88027 8965
rect 87969 8956 87981 8959
rect 87932 8928 87981 8956
rect 87932 8916 87938 8928
rect 87969 8925 87981 8928
rect 88015 8925 88027 8959
rect 87969 8919 88027 8925
rect 89438 8916 89444 8968
rect 89496 8956 89502 8968
rect 91005 8959 91063 8965
rect 91005 8956 91017 8959
rect 89496 8928 91017 8956
rect 89496 8916 89502 8928
rect 91005 8925 91017 8928
rect 91051 8956 91063 8959
rect 91278 8956 91284 8968
rect 91051 8928 91284 8956
rect 91051 8925 91063 8928
rect 91005 8919 91063 8925
rect 91278 8916 91284 8928
rect 91336 8916 91342 8968
rect 93397 8959 93455 8965
rect 93397 8925 93409 8959
rect 93443 8925 93455 8959
rect 93854 8956 93860 8968
rect 93815 8928 93860 8956
rect 93397 8919 93455 8925
rect 78122 8888 78128 8900
rect 77588 8860 78128 8888
rect 58434 8820 58440 8832
rect 57532 8792 58440 8820
rect 54481 8783 54539 8789
rect 58434 8780 58440 8792
rect 58492 8780 58498 8832
rect 59354 8780 59360 8832
rect 59412 8820 59418 8832
rect 59725 8823 59783 8829
rect 59725 8820 59737 8823
rect 59412 8792 59737 8820
rect 59412 8780 59418 8792
rect 59725 8789 59737 8792
rect 59771 8789 59783 8823
rect 59725 8783 59783 8789
rect 59893 8823 59951 8829
rect 59893 8789 59905 8823
rect 59939 8820 59951 8823
rect 60550 8820 60556 8832
rect 59939 8792 60556 8820
rect 59939 8789 59951 8792
rect 59893 8783 59951 8789
rect 60550 8780 60556 8792
rect 60608 8820 60614 8832
rect 63218 8820 63224 8832
rect 60608 8792 63224 8820
rect 60608 8780 60614 8792
rect 63218 8780 63224 8792
rect 63276 8780 63282 8832
rect 66622 8780 66628 8832
rect 66680 8820 66686 8832
rect 67542 8820 67548 8832
rect 66680 8792 67548 8820
rect 66680 8780 66686 8792
rect 67542 8780 67548 8792
rect 67600 8780 67606 8832
rect 67634 8780 67640 8832
rect 67692 8820 67698 8832
rect 69934 8820 69940 8832
rect 67692 8792 69940 8820
rect 67692 8780 67698 8792
rect 69934 8780 69940 8792
rect 69992 8780 69998 8832
rect 72510 8780 72516 8832
rect 72568 8820 72574 8832
rect 75380 8820 75408 8860
rect 78122 8848 78128 8860
rect 78180 8848 78186 8900
rect 79873 8891 79931 8897
rect 79873 8888 79885 8891
rect 79074 8860 79885 8888
rect 79873 8857 79885 8860
rect 79919 8857 79931 8891
rect 81526 8888 81532 8900
rect 81487 8860 81532 8888
rect 79873 8851 79931 8857
rect 81526 8848 81532 8860
rect 81584 8848 81590 8900
rect 81636 8860 82018 8888
rect 75546 8820 75552 8832
rect 72568 8792 75408 8820
rect 75507 8792 75552 8820
rect 72568 8780 72574 8792
rect 75546 8780 75552 8792
rect 75604 8780 75610 8832
rect 75730 8780 75736 8832
rect 75788 8820 75794 8832
rect 76193 8823 76251 8829
rect 76193 8820 76205 8823
rect 75788 8792 76205 8820
rect 75788 8780 75794 8792
rect 76193 8789 76205 8792
rect 76239 8789 76251 8823
rect 76193 8783 76251 8789
rect 80609 8823 80667 8829
rect 80609 8789 80621 8823
rect 80655 8820 80667 8823
rect 81636 8820 81664 8860
rect 84010 8848 84016 8900
rect 84068 8888 84074 8900
rect 84197 8891 84255 8897
rect 84197 8888 84209 8891
rect 84068 8860 84209 8888
rect 84068 8848 84074 8860
rect 84197 8857 84209 8860
rect 84243 8857 84255 8891
rect 84197 8851 84255 8857
rect 85666 8848 85672 8900
rect 85724 8888 85730 8900
rect 85853 8891 85911 8897
rect 85853 8888 85865 8891
rect 85724 8860 85865 8888
rect 85724 8848 85730 8860
rect 85853 8857 85865 8860
rect 85899 8857 85911 8891
rect 90174 8888 90180 8900
rect 85853 8851 85911 8857
rect 85960 8860 90180 8888
rect 80655 8792 81664 8820
rect 80655 8789 80667 8792
rect 80609 8783 80667 8789
rect 82814 8780 82820 8832
rect 82872 8820 82878 8832
rect 83001 8823 83059 8829
rect 83001 8820 83013 8823
rect 82872 8792 83013 8820
rect 82872 8780 82878 8792
rect 83001 8789 83013 8792
rect 83047 8789 83059 8823
rect 83001 8783 83059 8789
rect 83458 8780 83464 8832
rect 83516 8820 83522 8832
rect 85960 8820 85988 8860
rect 90174 8848 90180 8860
rect 90232 8848 90238 8900
rect 91557 8891 91615 8897
rect 91557 8857 91569 8891
rect 91603 8857 91615 8891
rect 91557 8851 91615 8857
rect 83516 8792 85988 8820
rect 87509 8823 87567 8829
rect 83516 8780 83522 8792
rect 87509 8789 87521 8823
rect 87555 8820 87567 8823
rect 89162 8820 89168 8832
rect 87555 8792 89168 8820
rect 87555 8789 87567 8792
rect 87509 8783 87567 8789
rect 89162 8780 89168 8792
rect 89220 8780 89226 8832
rect 91002 8780 91008 8832
rect 91060 8820 91066 8832
rect 91572 8820 91600 8851
rect 93118 8848 93124 8900
rect 93176 8888 93182 8900
rect 93412 8888 93440 8919
rect 93854 8916 93860 8928
rect 93912 8916 93918 8968
rect 93176 8860 93440 8888
rect 93176 8848 93182 8860
rect 91060 8792 91600 8820
rect 91060 8780 91066 8792
rect 1104 8730 95011 8752
rect 1104 8678 24386 8730
rect 24438 8678 24450 8730
rect 24502 8678 24514 8730
rect 24566 8678 24578 8730
rect 24630 8678 24642 8730
rect 24694 8678 47823 8730
rect 47875 8678 47887 8730
rect 47939 8678 47951 8730
rect 48003 8678 48015 8730
rect 48067 8678 48079 8730
rect 48131 8678 71260 8730
rect 71312 8678 71324 8730
rect 71376 8678 71388 8730
rect 71440 8678 71452 8730
rect 71504 8678 71516 8730
rect 71568 8678 94697 8730
rect 94749 8678 94761 8730
rect 94813 8678 94825 8730
rect 94877 8678 94889 8730
rect 94941 8678 94953 8730
rect 95005 8678 95011 8730
rect 1104 8656 95011 8678
rect 2130 8616 2136 8628
rect 2091 8588 2136 8616
rect 2130 8576 2136 8588
rect 2188 8576 2194 8628
rect 4706 8616 4712 8628
rect 4667 8588 4712 8616
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 6270 8576 6276 8628
rect 6328 8616 6334 8628
rect 8481 8619 8539 8625
rect 8481 8616 8493 8619
rect 6328 8588 8493 8616
rect 6328 8576 6334 8588
rect 8481 8585 8493 8588
rect 8527 8585 8539 8619
rect 8481 8579 8539 8585
rect 8570 8576 8576 8628
rect 8628 8616 8634 8628
rect 8628 8588 11836 8616
rect 8628 8576 8634 8588
rect 4430 8548 4436 8560
rect 4343 8520 4436 8548
rect 4356 8489 4384 8520
rect 4430 8508 4436 8520
rect 4488 8548 4494 8560
rect 5074 8548 5080 8560
rect 4488 8520 5080 8548
rect 4488 8508 4494 8520
rect 5074 8508 5080 8520
rect 5132 8548 5138 8560
rect 5132 8520 5488 8548
rect 5132 8508 5138 8520
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8480 3019 8483
rect 4341 8483 4399 8489
rect 3007 8452 4292 8480
rect 3007 8449 3019 8452
rect 2961 8443 3019 8449
rect 4264 8424 4292 8452
rect 4341 8449 4353 8483
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 3053 8415 3111 8421
rect 3053 8381 3065 8415
rect 3099 8381 3111 8415
rect 3053 8375 3111 8381
rect 3697 8415 3755 8421
rect 3697 8381 3709 8415
rect 3743 8412 3755 8415
rect 3970 8412 3976 8424
rect 3743 8384 3976 8412
rect 3743 8381 3755 8384
rect 3697 8375 3755 8381
rect 2222 8304 2228 8356
rect 2280 8344 2286 8356
rect 2593 8347 2651 8353
rect 2593 8344 2605 8347
rect 2280 8316 2605 8344
rect 2280 8304 2286 8316
rect 2593 8313 2605 8316
rect 2639 8313 2651 8347
rect 2593 8307 2651 8313
rect 2866 8304 2872 8356
rect 2924 8344 2930 8356
rect 3068 8344 3096 8375
rect 3970 8372 3976 8384
rect 4028 8372 4034 8424
rect 4246 8412 4252 8424
rect 4207 8384 4252 8412
rect 4246 8372 4252 8384
rect 4304 8372 4310 8424
rect 4522 8344 4528 8356
rect 2924 8316 4528 8344
rect 2924 8304 2930 8316
rect 4522 8304 4528 8316
rect 4580 8304 4586 8356
rect 5368 8344 5396 8443
rect 5460 8412 5488 8520
rect 5718 8508 5724 8560
rect 5776 8548 5782 8560
rect 5776 8520 7972 8548
rect 5776 8508 5782 8520
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8480 6699 8483
rect 6730 8480 6736 8492
rect 6687 8452 6736 8480
rect 6687 8449 6699 8452
rect 6641 8443 6699 8449
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8480 6975 8483
rect 7006 8480 7012 8492
rect 6963 8452 7012 8480
rect 6963 8449 6975 8452
rect 6917 8443 6975 8449
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 7466 8480 7472 8492
rect 7116 8452 7472 8480
rect 5905 8415 5963 8421
rect 5905 8412 5917 8415
rect 5460 8384 5917 8412
rect 5905 8381 5917 8384
rect 5951 8412 5963 8415
rect 7116 8412 7144 8452
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 7558 8440 7564 8492
rect 7616 8480 7622 8492
rect 7616 8452 7661 8480
rect 7616 8440 7622 8452
rect 5951 8384 7144 8412
rect 7837 8415 7895 8421
rect 5951 8381 5963 8384
rect 5905 8375 5963 8381
rect 7837 8381 7849 8415
rect 7883 8412 7895 8415
rect 7944 8412 7972 8520
rect 8588 8520 9536 8548
rect 8202 8440 8208 8492
rect 8260 8480 8266 8492
rect 8588 8489 8616 8520
rect 8573 8483 8631 8489
rect 8573 8480 8585 8483
rect 8260 8452 8585 8480
rect 8260 8440 8266 8452
rect 8573 8449 8585 8452
rect 8619 8449 8631 8483
rect 9122 8480 9128 8492
rect 9083 8452 9128 8480
rect 8573 8443 8631 8449
rect 9122 8440 9128 8452
rect 9180 8440 9186 8492
rect 9508 8489 9536 8520
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8449 9551 8483
rect 9493 8443 9551 8449
rect 10870 8412 10876 8424
rect 7883 8384 7972 8412
rect 10831 8384 10876 8412
rect 7883 8381 7895 8384
rect 7837 8375 7895 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 11701 8415 11759 8421
rect 11701 8381 11713 8415
rect 11747 8381 11759 8415
rect 11808 8412 11836 8588
rect 11882 8576 11888 8628
rect 11940 8616 11946 8628
rect 15010 8616 15016 8628
rect 11940 8588 13492 8616
rect 11940 8576 11946 8588
rect 13464 8557 13492 8588
rect 13924 8588 15016 8616
rect 13449 8551 13507 8557
rect 13449 8517 13461 8551
rect 13495 8517 13507 8551
rect 13449 8511 13507 8517
rect 12342 8440 12348 8492
rect 12400 8440 12406 8492
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 13780 8452 13825 8480
rect 13780 8440 13786 8452
rect 13924 8412 13952 8588
rect 15010 8576 15016 8588
rect 15068 8576 15074 8628
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 16850 8616 16856 8628
rect 16347 8588 16856 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 16850 8576 16856 8588
rect 16908 8576 16914 8628
rect 17034 8616 17040 8628
rect 16995 8588 17040 8616
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 20530 8576 20536 8628
rect 20588 8616 20594 8628
rect 20625 8619 20683 8625
rect 20625 8616 20637 8619
rect 20588 8588 20637 8616
rect 20588 8576 20594 8588
rect 20625 8585 20637 8588
rect 20671 8585 20683 8619
rect 20625 8579 20683 8585
rect 22557 8619 22615 8625
rect 22557 8585 22569 8619
rect 22603 8616 22615 8619
rect 27617 8619 27675 8625
rect 22603 8588 26280 8616
rect 22603 8585 22615 8588
rect 22557 8579 22615 8585
rect 14182 8508 14188 8560
rect 14240 8548 14246 8560
rect 15838 8548 15844 8560
rect 14240 8520 15844 8548
rect 14240 8508 14246 8520
rect 15838 8508 15844 8520
rect 15896 8508 15902 8560
rect 16022 8508 16028 8560
rect 16080 8548 16086 8560
rect 17126 8548 17132 8560
rect 16080 8520 17132 8548
rect 16080 8508 16086 8520
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 20254 8548 20260 8560
rect 20215 8520 20260 8548
rect 20254 8508 20260 8520
rect 20312 8508 20318 8560
rect 21450 8548 21456 8560
rect 21284 8520 21456 8548
rect 14737 8483 14795 8489
rect 14737 8449 14749 8483
rect 14783 8449 14795 8483
rect 17494 8480 17500 8492
rect 14737 8443 14795 8449
rect 14844 8452 17500 8480
rect 11808 8384 13952 8412
rect 11701 8375 11759 8381
rect 11330 8344 11336 8356
rect 5368 8316 7328 8344
rect 5258 8276 5264 8288
rect 5219 8248 5264 8276
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 7300 8276 7328 8316
rect 7760 8316 11336 8344
rect 7760 8276 7788 8316
rect 11330 8304 11336 8316
rect 11388 8344 11394 8356
rect 11716 8344 11744 8375
rect 11388 8316 11744 8344
rect 14752 8344 14780 8443
rect 14844 8421 14872 8452
rect 17494 8440 17500 8452
rect 17552 8440 17558 8492
rect 17586 8440 17592 8492
rect 17644 8440 17650 8492
rect 17678 8440 17684 8492
rect 17736 8480 17742 8492
rect 17865 8483 17923 8489
rect 17736 8452 17781 8480
rect 17736 8440 17742 8452
rect 17865 8449 17877 8483
rect 17911 8480 17923 8483
rect 18690 8480 18696 8492
rect 17911 8452 18696 8480
rect 17911 8449 17923 8452
rect 17865 8443 17923 8449
rect 18690 8440 18696 8452
rect 18748 8440 18754 8492
rect 19153 8483 19211 8489
rect 19153 8449 19165 8483
rect 19199 8449 19211 8483
rect 19153 8443 19211 8449
rect 14829 8415 14887 8421
rect 14829 8381 14841 8415
rect 14875 8381 14887 8415
rect 17402 8412 17408 8424
rect 14829 8375 14887 8381
rect 14936 8384 17408 8412
rect 14936 8344 14964 8384
rect 17402 8372 17408 8384
rect 17460 8372 17466 8424
rect 17604 8412 17632 8440
rect 17773 8415 17831 8421
rect 17773 8412 17785 8415
rect 17604 8384 17785 8412
rect 17773 8381 17785 8384
rect 17819 8381 17831 8415
rect 17773 8375 17831 8381
rect 17954 8372 17960 8424
rect 18012 8412 18018 8424
rect 18012 8384 18057 8412
rect 18012 8372 18018 8384
rect 18322 8372 18328 8424
rect 18380 8412 18386 8424
rect 19061 8415 19119 8421
rect 19061 8412 19073 8415
rect 18380 8384 19073 8412
rect 18380 8372 18386 8384
rect 19061 8381 19073 8384
rect 19107 8381 19119 8415
rect 19168 8412 19196 8443
rect 19610 8440 19616 8492
rect 19668 8480 19674 8492
rect 20165 8483 20223 8489
rect 20165 8480 20177 8483
rect 19668 8452 20177 8480
rect 19668 8440 19674 8452
rect 20165 8449 20177 8452
rect 20211 8449 20223 8483
rect 20438 8480 20444 8492
rect 20399 8452 20444 8480
rect 20165 8443 20223 8449
rect 20438 8440 20444 8452
rect 20496 8480 20502 8492
rect 21284 8480 21312 8520
rect 21450 8508 21456 8520
rect 21508 8508 21514 8560
rect 22370 8548 22376 8560
rect 22204 8520 22376 8548
rect 20496 8452 21312 8480
rect 21361 8483 21419 8489
rect 20496 8440 20502 8452
rect 21361 8449 21373 8483
rect 21407 8480 21419 8483
rect 22094 8480 22100 8492
rect 21407 8452 22100 8480
rect 21407 8449 21419 8452
rect 21361 8443 21419 8449
rect 22094 8440 22100 8452
rect 22152 8440 22158 8492
rect 22204 8489 22232 8520
rect 22370 8508 22376 8520
rect 22428 8548 22434 8560
rect 22428 8520 23428 8548
rect 22428 8508 22434 8520
rect 22189 8483 22247 8489
rect 22189 8449 22201 8483
rect 22235 8449 22247 8483
rect 22189 8443 22247 8449
rect 22554 8440 22560 8492
rect 22612 8480 22618 8492
rect 23017 8483 23075 8489
rect 23017 8480 23029 8483
rect 22612 8452 23029 8480
rect 22612 8440 22618 8452
rect 23017 8449 23029 8452
rect 23063 8449 23075 8483
rect 23017 8443 23075 8449
rect 21818 8412 21824 8424
rect 19168 8384 21824 8412
rect 19061 8375 19119 8381
rect 21818 8372 21824 8384
rect 21876 8372 21882 8424
rect 22281 8415 22339 8421
rect 22281 8381 22293 8415
rect 22327 8381 22339 8415
rect 22281 8375 22339 8381
rect 15102 8344 15108 8356
rect 14752 8316 14964 8344
rect 15063 8316 15108 8344
rect 11388 8304 11394 8316
rect 15102 8304 15108 8316
rect 15160 8304 15166 8356
rect 16209 8347 16267 8353
rect 16209 8313 16221 8347
rect 16255 8344 16267 8347
rect 17218 8344 17224 8356
rect 16255 8316 17224 8344
rect 16255 8313 16267 8316
rect 16209 8307 16267 8313
rect 17218 8304 17224 8316
rect 17276 8304 17282 8356
rect 17497 8347 17555 8353
rect 17497 8313 17509 8347
rect 17543 8344 17555 8347
rect 17586 8344 17592 8356
rect 17543 8316 17592 8344
rect 17543 8313 17555 8316
rect 17497 8307 17555 8313
rect 17586 8304 17592 8316
rect 17644 8304 17650 8356
rect 19521 8347 19579 8353
rect 19521 8313 19533 8347
rect 19567 8344 19579 8347
rect 22296 8344 22324 8375
rect 22922 8372 22928 8424
rect 22980 8412 22986 8424
rect 23109 8415 23167 8421
rect 23109 8412 23121 8415
rect 22980 8384 23121 8412
rect 22980 8372 22986 8384
rect 23109 8381 23121 8384
rect 23155 8381 23167 8415
rect 23290 8412 23296 8424
rect 23251 8384 23296 8412
rect 23109 8375 23167 8381
rect 23290 8372 23296 8384
rect 23348 8372 23354 8424
rect 23400 8412 23428 8520
rect 24854 8508 24860 8560
rect 24912 8548 24918 8560
rect 26252 8557 26280 8588
rect 27617 8585 27629 8619
rect 27663 8616 27675 8619
rect 27706 8616 27712 8628
rect 27663 8588 27712 8616
rect 27663 8585 27675 8588
rect 27617 8579 27675 8585
rect 26237 8551 26295 8557
rect 24912 8520 25070 8548
rect 24912 8508 24918 8520
rect 26237 8517 26249 8551
rect 26283 8517 26295 8551
rect 26237 8511 26295 8517
rect 23750 8480 23756 8492
rect 23711 8452 23756 8480
rect 23750 8440 23756 8452
rect 23808 8480 23814 8492
rect 26513 8483 26571 8489
rect 23808 8452 24900 8480
rect 23808 8440 23814 8452
rect 24765 8415 24823 8421
rect 24765 8412 24777 8415
rect 23400 8384 24777 8412
rect 24765 8381 24777 8384
rect 24811 8381 24823 8415
rect 24872 8412 24900 8452
rect 26513 8449 26525 8483
rect 26559 8480 26571 8483
rect 27632 8480 27660 8579
rect 27706 8576 27712 8588
rect 27764 8576 27770 8628
rect 28534 8576 28540 8628
rect 28592 8616 28598 8628
rect 33870 8616 33876 8628
rect 28592 8588 33876 8616
rect 28592 8576 28598 8588
rect 33870 8576 33876 8588
rect 33928 8576 33934 8628
rect 34256 8588 35204 8616
rect 28905 8551 28963 8557
rect 28905 8517 28917 8551
rect 28951 8548 28963 8551
rect 29822 8548 29828 8560
rect 28951 8520 29828 8548
rect 28951 8517 28963 8520
rect 28905 8511 28963 8517
rect 29822 8508 29828 8520
rect 29880 8508 29886 8560
rect 30650 8508 30656 8560
rect 30708 8508 30714 8560
rect 31478 8508 31484 8560
rect 31536 8548 31542 8560
rect 34256 8548 34284 8588
rect 31536 8520 34284 8548
rect 31536 8508 31542 8520
rect 34514 8508 34520 8560
rect 34572 8508 34578 8560
rect 35176 8548 35204 8588
rect 35710 8576 35716 8628
rect 35768 8616 35774 8628
rect 36262 8616 36268 8628
rect 35768 8588 36268 8616
rect 35768 8576 35774 8588
rect 36262 8576 36268 8588
rect 36320 8576 36326 8628
rect 36446 8616 36452 8628
rect 36407 8588 36452 8616
rect 36446 8576 36452 8588
rect 36504 8576 36510 8628
rect 37090 8576 37096 8628
rect 37148 8616 37154 8628
rect 37829 8619 37887 8625
rect 37829 8616 37841 8619
rect 37148 8588 37841 8616
rect 37148 8576 37154 8588
rect 37829 8585 37841 8588
rect 37875 8585 37887 8619
rect 37829 8579 37887 8585
rect 38378 8576 38384 8628
rect 38436 8616 38442 8628
rect 40313 8619 40371 8625
rect 40313 8616 40325 8619
rect 38436 8588 40325 8616
rect 38436 8576 38442 8588
rect 40313 8585 40325 8588
rect 40359 8585 40371 8619
rect 40313 8579 40371 8585
rect 42426 8576 42432 8628
rect 42484 8616 42490 8628
rect 42981 8619 43039 8625
rect 42981 8616 42993 8619
rect 42484 8588 42993 8616
rect 42484 8576 42490 8588
rect 42981 8585 42993 8588
rect 43027 8585 43039 8619
rect 44174 8616 44180 8628
rect 42981 8579 43039 8585
rect 43088 8588 44180 8616
rect 37182 8548 37188 8560
rect 35176 8520 37188 8548
rect 37182 8508 37188 8520
rect 37240 8508 37246 8560
rect 37550 8508 37556 8560
rect 37608 8548 37614 8560
rect 41322 8548 41328 8560
rect 37608 8520 41328 8548
rect 37608 8508 37614 8520
rect 41322 8508 41328 8520
rect 41380 8508 41386 8560
rect 29914 8480 29920 8492
rect 26559 8452 27660 8480
rect 29875 8452 29920 8480
rect 26559 8449 26571 8452
rect 26513 8443 26571 8449
rect 29914 8440 29920 8452
rect 29972 8440 29978 8492
rect 32490 8440 32496 8492
rect 32548 8480 32554 8492
rect 33318 8480 33324 8492
rect 32548 8452 33324 8480
rect 32548 8440 32554 8452
rect 33318 8440 33324 8452
rect 33376 8480 33382 8492
rect 33597 8483 33655 8489
rect 33597 8480 33609 8483
rect 33376 8452 33609 8480
rect 33376 8440 33382 8452
rect 33597 8449 33609 8452
rect 33643 8449 33655 8483
rect 36265 8483 36323 8489
rect 36265 8480 36277 8483
rect 33597 8443 33655 8449
rect 35544 8452 36277 8480
rect 29730 8412 29736 8424
rect 24872 8384 29736 8412
rect 24765 8375 24823 8381
rect 29730 8372 29736 8384
rect 29788 8372 29794 8424
rect 30193 8415 30251 8421
rect 30193 8381 30205 8415
rect 30239 8412 30251 8415
rect 33870 8412 33876 8424
rect 30239 8384 33732 8412
rect 33831 8384 33876 8412
rect 30239 8381 30251 8384
rect 30193 8375 30251 8381
rect 23201 8347 23259 8353
rect 23201 8344 23213 8347
rect 19567 8316 22232 8344
rect 22296 8316 23213 8344
rect 19567 8313 19579 8316
rect 19521 8307 19579 8313
rect 7300 8248 7788 8276
rect 16298 8236 16304 8288
rect 16356 8276 16362 8288
rect 19886 8276 19892 8288
rect 16356 8248 19892 8276
rect 16356 8236 16362 8248
rect 19886 8236 19892 8248
rect 19944 8236 19950 8288
rect 22204 8276 22232 8316
rect 23201 8313 23213 8316
rect 23247 8313 23259 8347
rect 29454 8344 29460 8356
rect 23201 8307 23259 8313
rect 23308 8316 24900 8344
rect 29415 8316 29460 8344
rect 23308 8276 23336 8316
rect 22204 8248 23336 8276
rect 24872 8276 24900 8316
rect 29454 8304 29460 8316
rect 29512 8344 29518 8356
rect 29914 8344 29920 8356
rect 29512 8316 29920 8344
rect 29512 8304 29518 8316
rect 29914 8304 29920 8316
rect 29972 8304 29978 8356
rect 31846 8304 31852 8356
rect 31904 8344 31910 8356
rect 32398 8344 32404 8356
rect 31904 8316 32404 8344
rect 31904 8304 31910 8316
rect 32398 8304 32404 8316
rect 32456 8344 32462 8356
rect 32585 8347 32643 8353
rect 32585 8344 32597 8347
rect 32456 8316 32597 8344
rect 32456 8304 32462 8316
rect 32585 8313 32597 8316
rect 32631 8344 32643 8347
rect 33410 8344 33416 8356
rect 32631 8316 33416 8344
rect 32631 8313 32643 8316
rect 32585 8307 32643 8313
rect 33410 8304 33416 8316
rect 33468 8304 33474 8356
rect 26142 8276 26148 8288
rect 24872 8248 26148 8276
rect 26142 8236 26148 8248
rect 26200 8236 26206 8288
rect 31662 8276 31668 8288
rect 31623 8248 31668 8276
rect 31662 8236 31668 8248
rect 31720 8236 31726 8288
rect 32766 8236 32772 8288
rect 32824 8276 32830 8288
rect 33045 8279 33103 8285
rect 33045 8276 33057 8279
rect 32824 8248 33057 8276
rect 32824 8236 32830 8248
rect 33045 8245 33057 8248
rect 33091 8245 33103 8279
rect 33704 8276 33732 8384
rect 33870 8372 33876 8384
rect 33928 8372 33934 8424
rect 33962 8372 33968 8424
rect 34020 8412 34026 8424
rect 35544 8412 35572 8452
rect 36265 8449 36277 8452
rect 36311 8480 36323 8483
rect 36354 8480 36360 8492
rect 36311 8452 36360 8480
rect 36311 8449 36323 8452
rect 36265 8443 36323 8449
rect 36354 8440 36360 8452
rect 36412 8440 36418 8492
rect 36541 8483 36599 8489
rect 36541 8449 36553 8483
rect 36587 8480 36599 8483
rect 37461 8483 37519 8489
rect 37461 8480 37473 8483
rect 36587 8452 37473 8480
rect 36587 8449 36599 8452
rect 36541 8443 36599 8449
rect 37461 8449 37473 8452
rect 37507 8449 37519 8483
rect 37461 8443 37519 8449
rect 34020 8384 35572 8412
rect 35621 8415 35679 8421
rect 34020 8372 34026 8384
rect 35621 8381 35633 8415
rect 35667 8381 35679 8415
rect 35621 8375 35679 8381
rect 35636 8344 35664 8375
rect 35802 8372 35808 8424
rect 35860 8412 35866 8424
rect 36556 8412 36584 8443
rect 37642 8440 37648 8492
rect 37700 8480 37706 8492
rect 37700 8452 37745 8480
rect 37700 8440 37706 8452
rect 38654 8440 38660 8492
rect 38712 8480 38718 8492
rect 39301 8483 39359 8489
rect 39301 8480 39313 8483
rect 38712 8452 39313 8480
rect 38712 8440 38718 8452
rect 39301 8449 39313 8452
rect 39347 8480 39359 8483
rect 40310 8480 40316 8492
rect 39347 8452 40316 8480
rect 39347 8449 39359 8452
rect 39301 8443 39359 8449
rect 40310 8440 40316 8452
rect 40368 8440 40374 8492
rect 40494 8480 40500 8492
rect 40455 8452 40500 8480
rect 40494 8440 40500 8452
rect 40552 8440 40558 8492
rect 40770 8480 40776 8492
rect 40731 8452 40776 8480
rect 40770 8440 40776 8452
rect 40828 8440 40834 8492
rect 41046 8440 41052 8492
rect 41104 8480 41110 8492
rect 41693 8483 41751 8489
rect 41693 8480 41705 8483
rect 41104 8452 41705 8480
rect 41104 8440 41110 8452
rect 41693 8449 41705 8452
rect 41739 8449 41751 8483
rect 41693 8443 41751 8449
rect 42797 8483 42855 8489
rect 42797 8449 42809 8483
rect 42843 8449 42855 8483
rect 42797 8443 42855 8449
rect 40402 8412 40408 8424
rect 35860 8384 36584 8412
rect 37752 8384 40408 8412
rect 35860 8372 35866 8384
rect 37752 8344 37780 8384
rect 40402 8372 40408 8384
rect 40460 8372 40466 8424
rect 40589 8415 40647 8421
rect 40589 8381 40601 8415
rect 40635 8381 40647 8415
rect 40589 8375 40647 8381
rect 35636 8316 37780 8344
rect 37826 8304 37832 8356
rect 37884 8344 37890 8356
rect 39758 8344 39764 8356
rect 37884 8316 39764 8344
rect 37884 8304 37890 8316
rect 39758 8304 39764 8316
rect 39816 8304 39822 8356
rect 40604 8344 40632 8375
rect 40678 8372 40684 8424
rect 40736 8412 40742 8424
rect 41598 8412 41604 8424
rect 40736 8384 40781 8412
rect 41559 8384 41604 8412
rect 40736 8372 40742 8384
rect 41598 8372 41604 8384
rect 41656 8372 41662 8424
rect 42058 8412 42064 8424
rect 42019 8384 42064 8412
rect 42058 8372 42064 8384
rect 42116 8372 42122 8424
rect 42613 8415 42671 8421
rect 42613 8381 42625 8415
rect 42659 8412 42671 8415
rect 42702 8412 42708 8424
rect 42659 8384 42708 8412
rect 42659 8381 42671 8384
rect 42613 8375 42671 8381
rect 42702 8372 42708 8384
rect 42760 8372 42766 8424
rect 42812 8412 42840 8443
rect 42886 8440 42892 8492
rect 42944 8480 42950 8492
rect 43088 8480 43116 8588
rect 44174 8576 44180 8588
rect 44232 8576 44238 8628
rect 45186 8616 45192 8628
rect 45147 8588 45192 8616
rect 45186 8576 45192 8588
rect 45244 8576 45250 8628
rect 45370 8576 45376 8628
rect 45428 8616 45434 8628
rect 47394 8616 47400 8628
rect 45428 8588 47400 8616
rect 45428 8576 45434 8588
rect 47394 8576 47400 8588
rect 47452 8576 47458 8628
rect 47857 8619 47915 8625
rect 47857 8616 47869 8619
rect 47504 8588 47869 8616
rect 46566 8508 46572 8560
rect 46624 8548 46630 8560
rect 47504 8548 47532 8588
rect 47857 8585 47869 8588
rect 47903 8585 47915 8619
rect 49510 8616 49516 8628
rect 49471 8588 49516 8616
rect 47857 8579 47915 8585
rect 49510 8576 49516 8588
rect 49568 8576 49574 8628
rect 50614 8616 50620 8628
rect 50575 8588 50620 8616
rect 50614 8576 50620 8588
rect 50672 8576 50678 8628
rect 53469 8619 53527 8625
rect 50816 8588 52224 8616
rect 48501 8551 48559 8557
rect 48501 8548 48513 8551
rect 46624 8520 47532 8548
rect 47780 8520 48513 8548
rect 46624 8508 46630 8520
rect 42944 8452 43116 8480
rect 42944 8440 42950 8452
rect 43162 8440 43168 8492
rect 43220 8480 43226 8492
rect 43901 8483 43959 8489
rect 43901 8480 43913 8483
rect 43220 8452 43913 8480
rect 43220 8440 43226 8452
rect 43901 8449 43913 8452
rect 43947 8449 43959 8483
rect 43901 8443 43959 8449
rect 44910 8440 44916 8492
rect 44968 8480 44974 8492
rect 46201 8483 46259 8489
rect 46201 8480 46213 8483
rect 44968 8452 46213 8480
rect 44968 8440 44974 8452
rect 46201 8449 46213 8452
rect 46247 8449 46259 8483
rect 46201 8443 46259 8449
rect 46842 8440 46848 8492
rect 46900 8480 46906 8492
rect 47780 8489 47808 8520
rect 48501 8517 48513 8520
rect 48547 8517 48559 8551
rect 48501 8511 48559 8517
rect 47765 8483 47823 8489
rect 47765 8480 47777 8483
rect 46900 8452 47777 8480
rect 46900 8440 46906 8452
rect 47765 8449 47777 8452
rect 47811 8449 47823 8483
rect 47765 8443 47823 8449
rect 47949 8483 48007 8489
rect 47949 8449 47961 8483
rect 47995 8480 48007 8483
rect 48777 8483 48835 8489
rect 48777 8480 48789 8483
rect 47995 8452 48789 8480
rect 47995 8449 48007 8452
rect 47949 8443 48007 8449
rect 48777 8449 48789 8452
rect 48823 8480 48835 8483
rect 49418 8480 49424 8492
rect 48823 8452 49424 8480
rect 48823 8449 48835 8452
rect 48777 8443 48835 8449
rect 43438 8412 43444 8424
rect 42812 8384 43444 8412
rect 42812 8344 42840 8384
rect 43438 8372 43444 8384
rect 43496 8372 43502 8424
rect 43530 8372 43536 8424
rect 43588 8412 43594 8424
rect 43993 8415 44051 8421
rect 43993 8412 44005 8415
rect 43588 8384 44005 8412
rect 43588 8372 43594 8384
rect 43993 8381 44005 8384
rect 44039 8412 44051 8415
rect 44082 8412 44088 8424
rect 44039 8384 44088 8412
rect 44039 8381 44051 8384
rect 43993 8375 44051 8381
rect 44082 8372 44088 8384
rect 44140 8372 44146 8424
rect 44269 8415 44327 8421
rect 44269 8381 44281 8415
rect 44315 8412 44327 8415
rect 45646 8412 45652 8424
rect 44315 8384 45652 8412
rect 44315 8381 44327 8384
rect 44269 8375 44327 8381
rect 45646 8372 45652 8384
rect 45704 8372 45710 8424
rect 46753 8415 46811 8421
rect 46753 8381 46765 8415
rect 46799 8412 46811 8415
rect 47026 8412 47032 8424
rect 46799 8384 47032 8412
rect 46799 8381 46811 8384
rect 46753 8375 46811 8381
rect 47026 8372 47032 8384
rect 47084 8372 47090 8424
rect 47213 8415 47271 8421
rect 47213 8381 47225 8415
rect 47259 8381 47271 8415
rect 47213 8375 47271 8381
rect 40604 8316 42840 8344
rect 43165 8347 43223 8353
rect 43165 8313 43177 8347
rect 43211 8344 43223 8347
rect 43211 8316 46520 8344
rect 43211 8313 43223 8316
rect 43165 8307 43223 8313
rect 35802 8276 35808 8288
rect 33704 8248 35808 8276
rect 33045 8239 33103 8245
rect 35802 8236 35808 8248
rect 35860 8236 35866 8288
rect 35894 8236 35900 8288
rect 35952 8276 35958 8288
rect 36081 8279 36139 8285
rect 36081 8276 36093 8279
rect 35952 8248 36093 8276
rect 35952 8236 35958 8248
rect 36081 8245 36093 8248
rect 36127 8245 36139 8279
rect 36081 8239 36139 8245
rect 36262 8236 36268 8288
rect 36320 8276 36326 8288
rect 37550 8276 37556 8288
rect 36320 8248 37556 8276
rect 36320 8236 36326 8248
rect 37550 8236 37556 8248
rect 37608 8236 37614 8288
rect 38746 8276 38752 8288
rect 38707 8248 38752 8276
rect 38746 8236 38752 8248
rect 38804 8236 38810 8288
rect 40678 8236 40684 8288
rect 40736 8276 40742 8288
rect 42886 8276 42892 8288
rect 40736 8248 42892 8276
rect 40736 8236 40742 8248
rect 42886 8236 42892 8248
rect 42944 8236 42950 8288
rect 45738 8276 45744 8288
rect 45699 8248 45744 8276
rect 45738 8236 45744 8248
rect 45796 8236 45802 8288
rect 46492 8276 46520 8316
rect 46566 8304 46572 8356
rect 46624 8344 46630 8356
rect 46937 8347 46995 8353
rect 46937 8344 46949 8347
rect 46624 8316 46949 8344
rect 46624 8304 46630 8316
rect 46937 8313 46949 8316
rect 46983 8313 46995 8347
rect 46937 8307 46995 8313
rect 46750 8276 46756 8288
rect 46492 8248 46756 8276
rect 46750 8236 46756 8248
rect 46808 8236 46814 8288
rect 47228 8276 47256 8375
rect 47302 8372 47308 8424
rect 47360 8412 47366 8424
rect 47964 8412 47992 8443
rect 49418 8440 49424 8452
rect 49476 8440 49482 8492
rect 49602 8440 49608 8492
rect 49660 8480 49666 8492
rect 49881 8483 49939 8489
rect 49881 8480 49893 8483
rect 49660 8452 49893 8480
rect 49660 8440 49666 8452
rect 49881 8449 49893 8452
rect 49927 8480 49939 8483
rect 50816 8480 50844 8588
rect 52196 8560 52224 8588
rect 53469 8585 53481 8619
rect 53515 8616 53527 8619
rect 53650 8616 53656 8628
rect 53515 8588 53656 8616
rect 53515 8585 53527 8588
rect 53469 8579 53527 8585
rect 53650 8576 53656 8588
rect 53708 8576 53714 8628
rect 53742 8576 53748 8628
rect 53800 8616 53806 8628
rect 54573 8619 54631 8625
rect 54573 8616 54585 8619
rect 53800 8588 54585 8616
rect 53800 8576 53806 8588
rect 54573 8585 54585 8588
rect 54619 8616 54631 8619
rect 57238 8616 57244 8628
rect 54619 8588 57244 8616
rect 54619 8585 54631 8588
rect 54573 8579 54631 8585
rect 57238 8576 57244 8588
rect 57296 8616 57302 8628
rect 57425 8619 57483 8625
rect 57425 8616 57437 8619
rect 57296 8588 57437 8616
rect 57296 8576 57302 8588
rect 57425 8585 57437 8588
rect 57471 8585 57483 8619
rect 57425 8579 57483 8585
rect 59262 8576 59268 8628
rect 59320 8616 59326 8628
rect 62574 8616 62580 8628
rect 59320 8588 62580 8616
rect 59320 8576 59326 8588
rect 62574 8576 62580 8588
rect 62632 8576 62638 8628
rect 64049 8619 64107 8625
rect 64049 8585 64061 8619
rect 64095 8616 64107 8619
rect 73798 8616 73804 8628
rect 64095 8588 73804 8616
rect 64095 8585 64107 8588
rect 64049 8579 64107 8585
rect 73798 8576 73804 8588
rect 73856 8576 73862 8628
rect 75178 8616 75184 8628
rect 75139 8588 75184 8616
rect 75178 8576 75184 8588
rect 75236 8576 75242 8628
rect 78125 8619 78183 8625
rect 78125 8616 78137 8619
rect 75840 8588 78137 8616
rect 51626 8508 51632 8560
rect 51684 8508 51690 8560
rect 52086 8548 52092 8560
rect 52047 8520 52092 8548
rect 52086 8508 52092 8520
rect 52144 8508 52150 8560
rect 52178 8508 52184 8560
rect 52236 8548 52242 8560
rect 58618 8548 58624 8560
rect 52236 8520 53328 8548
rect 56718 8520 58624 8548
rect 52236 8508 52242 8520
rect 53190 8480 53196 8492
rect 49927 8452 50844 8480
rect 53151 8452 53196 8480
rect 49927 8449 49939 8452
rect 49881 8443 49939 8449
rect 53190 8440 53196 8452
rect 53248 8440 53254 8492
rect 53300 8480 53328 8520
rect 58618 8508 58624 8520
rect 58676 8508 58682 8560
rect 60090 8548 60096 8560
rect 58912 8520 60096 8548
rect 53926 8480 53932 8492
rect 53300 8452 53604 8480
rect 53887 8452 53932 8480
rect 48682 8412 48688 8424
rect 47360 8384 47992 8412
rect 48643 8384 48688 8412
rect 47360 8372 47366 8384
rect 48682 8372 48688 8384
rect 48740 8372 48746 8424
rect 49970 8412 49976 8424
rect 49931 8384 49976 8412
rect 49970 8372 49976 8384
rect 50028 8372 50034 8424
rect 52362 8412 52368 8424
rect 52323 8384 52368 8412
rect 52362 8372 52368 8384
rect 52420 8372 52426 8424
rect 52638 8372 52644 8424
rect 52696 8412 52702 8424
rect 53466 8412 53472 8424
rect 52696 8384 53472 8412
rect 52696 8372 52702 8384
rect 53466 8372 53472 8384
rect 53524 8372 53530 8424
rect 53576 8412 53604 8452
rect 53926 8440 53932 8452
rect 53984 8440 53990 8492
rect 54113 8483 54171 8489
rect 54113 8449 54125 8483
rect 54159 8449 54171 8483
rect 54113 8443 54171 8449
rect 58069 8483 58127 8489
rect 58069 8449 58081 8483
rect 58115 8480 58127 8483
rect 58158 8480 58164 8492
rect 58115 8452 58164 8480
rect 58115 8449 58127 8452
rect 58069 8443 58127 8449
rect 54128 8412 54156 8443
rect 58158 8440 58164 8452
rect 58216 8440 58222 8492
rect 55214 8412 55220 8424
rect 53576 8384 54156 8412
rect 55175 8384 55220 8412
rect 48314 8304 48320 8356
rect 48372 8344 48378 8356
rect 53285 8347 53343 8353
rect 48372 8316 49004 8344
rect 48372 8304 48378 8316
rect 48777 8279 48835 8285
rect 48777 8276 48789 8279
rect 47228 8248 48789 8276
rect 48777 8245 48789 8248
rect 48823 8276 48835 8279
rect 48866 8276 48872 8288
rect 48823 8248 48872 8276
rect 48823 8245 48835 8248
rect 48777 8239 48835 8245
rect 48866 8236 48872 8248
rect 48924 8236 48930 8288
rect 48976 8285 49004 8316
rect 53285 8313 53297 8347
rect 53331 8344 53343 8347
rect 53331 8316 53420 8344
rect 53331 8313 53343 8316
rect 53285 8307 53343 8313
rect 48961 8279 49019 8285
rect 48961 8245 48973 8279
rect 49007 8276 49019 8279
rect 51442 8276 51448 8288
rect 49007 8248 51448 8276
rect 49007 8245 49019 8248
rect 48961 8239 49019 8245
rect 51442 8236 51448 8248
rect 51500 8236 51506 8288
rect 53392 8276 53420 8316
rect 53929 8279 53987 8285
rect 53929 8276 53941 8279
rect 53392 8248 53941 8276
rect 53929 8245 53941 8248
rect 53975 8245 53987 8279
rect 54128 8276 54156 8384
rect 55214 8372 55220 8384
rect 55272 8372 55278 8424
rect 55490 8412 55496 8424
rect 55451 8384 55496 8412
rect 55490 8372 55496 8384
rect 55548 8372 55554 8424
rect 55858 8372 55864 8424
rect 55916 8412 55922 8424
rect 58250 8412 58256 8424
rect 55916 8384 58256 8412
rect 55916 8372 55922 8384
rect 58250 8372 58256 8384
rect 58308 8412 58314 8424
rect 58912 8412 58940 8520
rect 60090 8508 60096 8520
rect 60148 8508 60154 8560
rect 66806 8508 66812 8560
rect 66864 8508 66870 8560
rect 67542 8508 67548 8560
rect 67600 8548 67606 8560
rect 69017 8551 69075 8557
rect 69017 8548 69029 8551
rect 67600 8520 69029 8548
rect 67600 8508 67606 8520
rect 69017 8517 69029 8520
rect 69063 8517 69075 8551
rect 69017 8511 69075 8517
rect 69750 8508 69756 8560
rect 69808 8548 69814 8560
rect 75546 8548 75552 8560
rect 69808 8520 75552 8548
rect 69808 8508 69814 8520
rect 59354 8480 59360 8492
rect 59315 8452 59360 8480
rect 59354 8440 59360 8452
rect 59412 8440 59418 8492
rect 62206 8480 62212 8492
rect 59078 8412 59084 8424
rect 58308 8384 58940 8412
rect 59039 8384 59084 8412
rect 58308 8372 58314 8384
rect 59078 8372 59084 8384
rect 59136 8372 59142 8424
rect 59262 8412 59268 8424
rect 59223 8384 59268 8412
rect 59262 8372 59268 8384
rect 59320 8372 59326 8424
rect 59814 8412 59820 8424
rect 59775 8384 59820 8412
rect 59814 8372 59820 8384
rect 59872 8372 59878 8424
rect 60090 8412 60096 8424
rect 60051 8384 60096 8412
rect 60090 8372 60096 8384
rect 60148 8372 60154 8424
rect 58161 8347 58219 8353
rect 58161 8313 58173 8347
rect 58207 8344 58219 8347
rect 59354 8344 59360 8356
rect 58207 8316 59360 8344
rect 58207 8313 58219 8316
rect 58161 8307 58219 8313
rect 59354 8304 59360 8316
rect 59412 8304 59418 8356
rect 61212 8344 61240 8466
rect 62167 8452 62212 8480
rect 62206 8440 62212 8452
rect 62264 8440 62270 8492
rect 63678 8440 63684 8492
rect 63736 8480 63742 8492
rect 64506 8480 64512 8492
rect 63736 8452 63781 8480
rect 64467 8452 64512 8480
rect 63736 8440 63742 8452
rect 64506 8440 64512 8452
rect 64564 8440 64570 8492
rect 73614 8480 73620 8492
rect 73575 8452 73620 8480
rect 73614 8440 73620 8452
rect 73672 8440 73678 8492
rect 73816 8489 73844 8520
rect 75546 8508 75552 8520
rect 75604 8508 75610 8560
rect 73801 8483 73859 8489
rect 73801 8449 73813 8483
rect 73847 8449 73859 8483
rect 73801 8443 73859 8449
rect 74350 8440 74356 8492
rect 74408 8480 74414 8492
rect 75270 8480 75276 8492
rect 74408 8452 75276 8480
rect 74408 8440 74414 8452
rect 75270 8440 75276 8452
rect 75328 8440 75334 8492
rect 75730 8480 75736 8492
rect 75380 8452 75736 8480
rect 63770 8412 63776 8424
rect 63731 8384 63776 8412
rect 63770 8372 63776 8384
rect 63828 8372 63834 8424
rect 64782 8412 64788 8424
rect 64743 8384 64788 8412
rect 64782 8372 64788 8384
rect 64840 8372 64846 8424
rect 67542 8412 67548 8424
rect 67503 8384 67548 8412
rect 67542 8372 67548 8384
rect 67600 8372 67606 8424
rect 67821 8415 67879 8421
rect 67821 8381 67833 8415
rect 67867 8412 67879 8415
rect 68186 8412 68192 8424
rect 67867 8384 68192 8412
rect 67867 8381 67879 8384
rect 67821 8375 67879 8381
rect 68186 8372 68192 8384
rect 68244 8372 68250 8424
rect 68554 8372 68560 8424
rect 68612 8412 68618 8424
rect 68833 8415 68891 8421
rect 68833 8412 68845 8415
rect 68612 8384 68845 8412
rect 68612 8372 68618 8384
rect 68833 8381 68845 8384
rect 68879 8381 68891 8415
rect 68833 8375 68891 8381
rect 70673 8415 70731 8421
rect 70673 8381 70685 8415
rect 70719 8381 70731 8415
rect 70673 8375 70731 8381
rect 62485 8347 62543 8353
rect 62485 8344 62497 8347
rect 61212 8316 62497 8344
rect 62485 8313 62497 8316
rect 62531 8344 62543 8347
rect 63402 8344 63408 8356
rect 62531 8316 63408 8344
rect 62531 8313 62543 8316
rect 62485 8307 62543 8313
rect 63402 8304 63408 8316
rect 63460 8304 63466 8356
rect 70688 8344 70716 8375
rect 70762 8372 70768 8424
rect 70820 8412 70826 8424
rect 72510 8412 72516 8424
rect 70820 8384 72516 8412
rect 70820 8372 70826 8384
rect 72510 8372 72516 8384
rect 72568 8372 72574 8424
rect 72786 8412 72792 8424
rect 72747 8384 72792 8412
rect 72786 8372 72792 8384
rect 72844 8372 72850 8424
rect 72970 8412 72976 8424
rect 72931 8384 72976 8412
rect 72970 8372 72976 8384
rect 73028 8372 73034 8424
rect 73062 8372 73068 8424
rect 73120 8412 73126 8424
rect 74629 8415 74687 8421
rect 73120 8384 73568 8412
rect 73120 8372 73126 8384
rect 73154 8344 73160 8356
rect 70688 8316 73160 8344
rect 73154 8304 73160 8316
rect 73212 8304 73218 8356
rect 73540 8344 73568 8384
rect 74629 8381 74641 8415
rect 74675 8412 74687 8415
rect 74718 8412 74724 8424
rect 74675 8384 74724 8412
rect 74675 8381 74687 8384
rect 74629 8375 74687 8381
rect 74718 8372 74724 8384
rect 74776 8372 74782 8424
rect 74810 8372 74816 8424
rect 74868 8412 74874 8424
rect 75380 8412 75408 8452
rect 75730 8440 75736 8452
rect 75788 8440 75794 8492
rect 75840 8412 75868 8588
rect 78125 8585 78137 8588
rect 78171 8616 78183 8619
rect 80514 8616 80520 8628
rect 78171 8588 80520 8616
rect 78171 8585 78183 8588
rect 78125 8579 78183 8585
rect 80514 8576 80520 8588
rect 80572 8576 80578 8628
rect 81526 8576 81532 8628
rect 81584 8616 81590 8628
rect 82173 8619 82231 8625
rect 82173 8616 82185 8619
rect 81584 8588 82185 8616
rect 81584 8576 81590 8588
rect 82173 8585 82185 8588
rect 82219 8585 82231 8619
rect 82173 8579 82231 8585
rect 82630 8576 82636 8628
rect 82688 8616 82694 8628
rect 86865 8619 86923 8625
rect 86865 8616 86877 8619
rect 82688 8588 86877 8616
rect 82688 8576 82694 8588
rect 86865 8585 86877 8588
rect 86911 8585 86923 8619
rect 88978 8616 88984 8628
rect 86865 8579 86923 8585
rect 87892 8588 88984 8616
rect 76466 8508 76472 8560
rect 76524 8508 76530 8560
rect 77527 8551 77585 8557
rect 77527 8548 77539 8551
rect 77266 8520 77539 8548
rect 76098 8412 76104 8424
rect 74868 8384 75408 8412
rect 75748 8384 75868 8412
rect 76059 8384 76104 8412
rect 74868 8372 74874 8384
rect 75748 8344 75776 8384
rect 76098 8372 76104 8384
rect 76156 8372 76162 8424
rect 76374 8372 76380 8424
rect 76432 8412 76438 8424
rect 77266 8412 77294 8520
rect 77527 8517 77539 8520
rect 77573 8548 77585 8551
rect 77938 8548 77944 8560
rect 77573 8520 77944 8548
rect 77573 8517 77585 8520
rect 77527 8511 77585 8517
rect 77938 8508 77944 8520
rect 77996 8508 78002 8560
rect 78858 8548 78864 8560
rect 78819 8520 78864 8548
rect 78858 8508 78864 8520
rect 78916 8508 78922 8560
rect 83550 8548 83556 8560
rect 82924 8520 83556 8548
rect 80238 8440 80244 8492
rect 80296 8480 80302 8492
rect 81253 8483 81311 8489
rect 81253 8480 81265 8483
rect 80296 8452 81265 8480
rect 80296 8440 80302 8452
rect 81253 8449 81265 8452
rect 81299 8480 81311 8483
rect 82265 8483 82323 8489
rect 81299 8452 82124 8480
rect 81299 8449 81311 8452
rect 81253 8443 81311 8449
rect 78674 8412 78680 8424
rect 76432 8384 77294 8412
rect 78635 8384 78680 8412
rect 76432 8372 76438 8384
rect 78674 8372 78680 8384
rect 78732 8372 78738 8424
rect 78858 8372 78864 8424
rect 78916 8412 78922 8424
rect 79137 8415 79195 8421
rect 79137 8412 79149 8415
rect 78916 8384 79149 8412
rect 78916 8372 78922 8384
rect 79137 8381 79149 8384
rect 79183 8412 79195 8415
rect 81710 8412 81716 8424
rect 79183 8384 81716 8412
rect 79183 8381 79195 8384
rect 79137 8375 79195 8381
rect 81710 8372 81716 8384
rect 81768 8372 81774 8424
rect 73540 8316 75776 8344
rect 77956 8316 78168 8344
rect 56502 8276 56508 8288
rect 54128 8248 56508 8276
rect 53929 8239 53987 8245
rect 56502 8236 56508 8248
rect 56560 8236 56566 8288
rect 56965 8279 57023 8285
rect 56965 8245 56977 8279
rect 57011 8276 57023 8279
rect 57238 8276 57244 8288
rect 57011 8248 57244 8276
rect 57011 8245 57023 8248
rect 56965 8239 57023 8245
rect 57238 8236 57244 8248
rect 57296 8236 57302 8288
rect 59170 8276 59176 8288
rect 59131 8248 59176 8276
rect 59170 8236 59176 8248
rect 59228 8236 59234 8288
rect 60182 8236 60188 8288
rect 60240 8276 60246 8288
rect 61565 8279 61623 8285
rect 61565 8276 61577 8279
rect 60240 8248 61577 8276
rect 60240 8236 60246 8248
rect 61565 8245 61577 8248
rect 61611 8276 61623 8279
rect 63310 8276 63316 8288
rect 61611 8248 63316 8276
rect 61611 8245 61623 8248
rect 61565 8239 61623 8245
rect 63310 8236 63316 8248
rect 63368 8236 63374 8288
rect 64138 8236 64144 8288
rect 64196 8276 64202 8288
rect 65429 8279 65487 8285
rect 65429 8276 65441 8279
rect 64196 8248 65441 8276
rect 64196 8236 64202 8248
rect 65429 8245 65441 8248
rect 65475 8245 65487 8279
rect 66070 8276 66076 8288
rect 65983 8248 66076 8276
rect 65429 8239 65487 8245
rect 66070 8236 66076 8248
rect 66128 8276 66134 8288
rect 66990 8276 66996 8288
rect 66128 8248 66996 8276
rect 66128 8236 66134 8248
rect 66990 8236 66996 8248
rect 67048 8276 67054 8288
rect 67450 8276 67456 8288
rect 67048 8248 67456 8276
rect 67048 8236 67054 8248
rect 67450 8236 67456 8248
rect 67508 8236 67514 8288
rect 69106 8236 69112 8288
rect 69164 8276 69170 8288
rect 73614 8276 73620 8288
rect 69164 8248 73620 8276
rect 69164 8236 69170 8248
rect 73614 8236 73620 8248
rect 73672 8236 73678 8288
rect 74350 8236 74356 8288
rect 74408 8276 74414 8288
rect 77956 8276 77984 8316
rect 74408 8248 77984 8276
rect 78140 8276 78168 8316
rect 80992 8316 81204 8344
rect 80992 8276 81020 8316
rect 78140 8248 81020 8276
rect 81176 8276 81204 8316
rect 81250 8304 81256 8356
rect 81308 8344 81314 8356
rect 82096 8344 82124 8452
rect 82265 8449 82277 8483
rect 82311 8480 82323 8483
rect 82630 8480 82636 8492
rect 82311 8452 82636 8480
rect 82311 8449 82323 8452
rect 82265 8443 82323 8449
rect 82630 8440 82636 8452
rect 82688 8440 82694 8492
rect 82924 8489 82952 8520
rect 83550 8508 83556 8520
rect 83608 8508 83614 8560
rect 84286 8508 84292 8560
rect 84344 8548 84350 8560
rect 87892 8557 87920 8588
rect 88978 8576 88984 8588
rect 89036 8576 89042 8628
rect 87877 8551 87935 8557
rect 87877 8548 87889 8551
rect 84344 8520 85882 8548
rect 87432 8520 87889 8548
rect 84344 8508 84350 8520
rect 82909 8483 82967 8489
rect 82909 8449 82921 8483
rect 82955 8449 82967 8483
rect 83366 8480 83372 8492
rect 82909 8443 82967 8449
rect 83016 8452 83372 8480
rect 83016 8421 83044 8452
rect 83366 8440 83372 8452
rect 83424 8440 83430 8492
rect 83642 8440 83648 8492
rect 83700 8480 83706 8492
rect 84105 8483 84163 8489
rect 84105 8480 84117 8483
rect 83700 8452 84117 8480
rect 83700 8440 83706 8452
rect 84105 8449 84117 8452
rect 84151 8480 84163 8483
rect 84194 8480 84200 8492
rect 84151 8452 84200 8480
rect 84151 8449 84163 8452
rect 84105 8443 84163 8449
rect 84194 8440 84200 8452
rect 84252 8440 84258 8492
rect 83001 8415 83059 8421
rect 83001 8381 83013 8415
rect 83047 8381 83059 8415
rect 85117 8415 85175 8421
rect 85117 8412 85129 8415
rect 83001 8375 83059 8381
rect 83108 8384 85129 8412
rect 83108 8344 83136 8384
rect 85117 8381 85129 8384
rect 85163 8381 85175 8415
rect 85390 8412 85396 8424
rect 85351 8384 85396 8412
rect 85117 8375 85175 8381
rect 85390 8372 85396 8384
rect 85448 8372 85454 8424
rect 85482 8372 85488 8424
rect 85540 8412 85546 8424
rect 87432 8412 87460 8520
rect 87877 8517 87889 8520
rect 87923 8517 87935 8551
rect 87877 8511 87935 8517
rect 88334 8508 88340 8560
rect 88392 8548 88398 8560
rect 93394 8548 93400 8560
rect 88392 8520 90772 8548
rect 93355 8520 93400 8548
rect 88392 8508 88398 8520
rect 87509 8483 87567 8489
rect 87509 8449 87521 8483
rect 87555 8480 87567 8483
rect 89254 8480 89260 8492
rect 87555 8452 88196 8480
rect 89215 8452 89260 8480
rect 87555 8449 87567 8452
rect 87509 8443 87567 8449
rect 85540 8384 87460 8412
rect 85540 8372 85546 8384
rect 81308 8316 81353 8344
rect 82096 8316 83136 8344
rect 83277 8347 83335 8353
rect 81308 8304 81314 8316
rect 83277 8313 83289 8347
rect 83323 8344 83335 8347
rect 84654 8344 84660 8356
rect 83323 8316 84660 8344
rect 83323 8313 83335 8316
rect 83277 8307 83335 8313
rect 84654 8304 84660 8316
rect 84712 8304 84718 8356
rect 82722 8276 82728 8288
rect 81176 8248 82728 8276
rect 74408 8236 74414 8248
rect 82722 8236 82728 8248
rect 82780 8236 82786 8288
rect 84197 8279 84255 8285
rect 84197 8245 84209 8279
rect 84243 8276 84255 8279
rect 84286 8276 84292 8288
rect 84243 8248 84292 8276
rect 84243 8245 84255 8248
rect 84197 8239 84255 8245
rect 84286 8236 84292 8248
rect 84344 8236 84350 8288
rect 86678 8236 86684 8288
rect 86736 8276 86742 8288
rect 87524 8276 87552 8443
rect 88168 8412 88196 8452
rect 89254 8440 89260 8452
rect 89312 8440 89318 8492
rect 89714 8440 89720 8492
rect 89772 8480 89778 8492
rect 89901 8483 89959 8489
rect 89901 8480 89913 8483
rect 89772 8452 89913 8480
rect 89772 8440 89778 8452
rect 89901 8449 89913 8452
rect 89947 8480 89959 8483
rect 89947 8452 90680 8480
rect 89947 8449 89959 8452
rect 89901 8443 89959 8449
rect 89438 8412 89444 8424
rect 88168 8384 89444 8412
rect 89438 8372 89444 8384
rect 89496 8372 89502 8424
rect 90174 8372 90180 8424
rect 90232 8412 90238 8424
rect 90232 8384 90277 8412
rect 90232 8372 90238 8384
rect 90652 8344 90680 8452
rect 90744 8421 90772 8520
rect 93394 8508 93400 8520
rect 93452 8508 93458 8560
rect 90821 8483 90879 8489
rect 90821 8449 90833 8483
rect 90867 8480 90879 8483
rect 90867 8452 92244 8480
rect 90867 8449 90879 8452
rect 90821 8443 90879 8449
rect 90729 8415 90787 8421
rect 90729 8381 90741 8415
rect 90775 8381 90787 8415
rect 90729 8375 90787 8381
rect 91002 8372 91008 8424
rect 91060 8412 91066 8424
rect 91741 8415 91799 8421
rect 91741 8412 91753 8415
rect 91060 8384 91753 8412
rect 91060 8372 91066 8384
rect 91741 8381 91753 8384
rect 91787 8381 91799 8415
rect 92216 8412 92244 8452
rect 93578 8412 93584 8424
rect 92216 8384 93584 8412
rect 91741 8375 91799 8381
rect 93578 8372 93584 8384
rect 93636 8372 93642 8424
rect 91020 8344 91048 8372
rect 91186 8344 91192 8356
rect 90652 8316 91048 8344
rect 91147 8316 91192 8344
rect 91186 8304 91192 8316
rect 91244 8304 91250 8356
rect 94130 8344 94136 8356
rect 94091 8316 94136 8344
rect 94130 8304 94136 8316
rect 94188 8304 94194 8356
rect 86736 8248 87552 8276
rect 88981 8279 89039 8285
rect 86736 8236 86742 8248
rect 88981 8245 88993 8279
rect 89027 8276 89039 8279
rect 89806 8276 89812 8288
rect 89027 8248 89812 8276
rect 89027 8245 89039 8248
rect 88981 8239 89039 8245
rect 89806 8236 89812 8248
rect 89864 8236 89870 8288
rect 1104 8186 94852 8208
rect 1104 8134 12668 8186
rect 12720 8134 12732 8186
rect 12784 8134 12796 8186
rect 12848 8134 12860 8186
rect 12912 8134 12924 8186
rect 12976 8134 36105 8186
rect 36157 8134 36169 8186
rect 36221 8134 36233 8186
rect 36285 8134 36297 8186
rect 36349 8134 36361 8186
rect 36413 8134 59542 8186
rect 59594 8134 59606 8186
rect 59658 8134 59670 8186
rect 59722 8134 59734 8186
rect 59786 8134 59798 8186
rect 59850 8134 82979 8186
rect 83031 8134 83043 8186
rect 83095 8134 83107 8186
rect 83159 8134 83171 8186
rect 83223 8134 83235 8186
rect 83287 8134 94852 8186
rect 1104 8112 94852 8134
rect 2866 8072 2872 8084
rect 2827 8044 2872 8072
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 3421 8075 3479 8081
rect 3421 8041 3433 8075
rect 3467 8072 3479 8075
rect 4338 8072 4344 8084
rect 3467 8044 4344 8072
rect 3467 8041 3479 8044
rect 3421 8035 3479 8041
rect 4338 8032 4344 8044
rect 4396 8032 4402 8084
rect 6822 8072 6828 8084
rect 5000 8044 6828 8072
rect 5000 7945 5028 8044
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 11698 8072 11704 8084
rect 7024 8044 11704 8072
rect 4985 7939 5043 7945
rect 4985 7905 4997 7939
rect 5031 7905 5043 7939
rect 5258 7936 5264 7948
rect 5219 7908 5264 7936
rect 4985 7899 5043 7905
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 7024 7945 7052 8044
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 12526 8032 12532 8084
rect 12584 8072 12590 8084
rect 15565 8075 15623 8081
rect 15565 8072 15577 8075
rect 12584 8044 15577 8072
rect 12584 8032 12590 8044
rect 15565 8041 15577 8044
rect 15611 8041 15623 8075
rect 15565 8035 15623 8041
rect 17310 8032 17316 8084
rect 17368 8072 17374 8084
rect 17405 8075 17463 8081
rect 17405 8072 17417 8075
rect 17368 8044 17417 8072
rect 17368 8032 17374 8044
rect 17405 8041 17417 8044
rect 17451 8041 17463 8075
rect 17405 8035 17463 8041
rect 17494 8032 17500 8084
rect 17552 8072 17558 8084
rect 18601 8075 18659 8081
rect 18601 8072 18613 8075
rect 17552 8044 18613 8072
rect 17552 8032 17558 8044
rect 18601 8041 18613 8044
rect 18647 8041 18659 8075
rect 18601 8035 18659 8041
rect 18874 8032 18880 8084
rect 18932 8072 18938 8084
rect 20625 8075 20683 8081
rect 20625 8072 20637 8075
rect 18932 8044 20637 8072
rect 18932 8032 18938 8044
rect 20625 8041 20637 8044
rect 20671 8041 20683 8075
rect 21634 8072 21640 8084
rect 21595 8044 21640 8072
rect 20625 8035 20683 8041
rect 21634 8032 21640 8044
rect 21692 8032 21698 8084
rect 21818 8072 21824 8084
rect 21779 8044 21824 8072
rect 21818 8032 21824 8044
rect 21876 8032 21882 8084
rect 21910 8032 21916 8084
rect 21968 8072 21974 8084
rect 28537 8075 28595 8081
rect 28537 8072 28549 8075
rect 21968 8044 28549 8072
rect 21968 8032 21974 8044
rect 28537 8041 28549 8044
rect 28583 8041 28595 8075
rect 28537 8035 28595 8041
rect 28626 8032 28632 8084
rect 28684 8072 28690 8084
rect 33134 8072 33140 8084
rect 28684 8044 33140 8072
rect 28684 8032 28690 8044
rect 33134 8032 33140 8044
rect 33192 8032 33198 8084
rect 33318 8072 33324 8084
rect 33279 8044 33324 8072
rect 33318 8032 33324 8044
rect 33376 8032 33382 8084
rect 35710 8072 35716 8084
rect 34256 8044 35716 8072
rect 7650 8004 7656 8016
rect 7611 7976 7656 8004
rect 7650 7964 7656 7976
rect 7708 7964 7714 8016
rect 13538 7964 13544 8016
rect 13596 8004 13602 8016
rect 13633 8007 13691 8013
rect 13633 8004 13645 8007
rect 13596 7976 13645 8004
rect 13596 7964 13602 7976
rect 13633 7973 13645 7976
rect 13679 7973 13691 8007
rect 13633 7967 13691 7973
rect 15102 7964 15108 8016
rect 15160 8004 15166 8016
rect 27801 8007 27859 8013
rect 15160 7976 22048 8004
rect 15160 7964 15166 7976
rect 7009 7939 7067 7945
rect 7009 7905 7021 7939
rect 7055 7905 7067 7939
rect 7009 7899 7067 7905
rect 17954 7896 17960 7948
rect 18012 7936 18018 7948
rect 18509 7939 18567 7945
rect 18509 7936 18521 7939
rect 18012 7908 18521 7936
rect 18012 7896 18018 7908
rect 18509 7905 18521 7908
rect 18555 7905 18567 7939
rect 18509 7899 18567 7905
rect 20073 7939 20131 7945
rect 20073 7905 20085 7939
rect 20119 7936 20131 7939
rect 20714 7936 20720 7948
rect 20119 7908 20720 7936
rect 20119 7905 20131 7908
rect 20073 7899 20131 7905
rect 20714 7896 20720 7908
rect 20772 7896 20778 7948
rect 20898 7936 20904 7948
rect 20859 7908 20904 7936
rect 20898 7896 20904 7908
rect 20956 7896 20962 7948
rect 21910 7944 21916 7948
rect 21744 7916 21916 7944
rect 3694 7828 3700 7880
rect 3752 7868 3758 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3752 7840 3985 7868
rect 3752 7828 3758 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7868 8447 7871
rect 9122 7868 9128 7880
rect 8435 7840 9128 7868
rect 8435 7837 8447 7840
rect 8389 7831 8447 7837
rect 9122 7828 9128 7840
rect 9180 7828 9186 7880
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7868 9459 7871
rect 9674 7868 9680 7880
rect 9447 7840 9680 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7868 10103 7871
rect 10134 7868 10140 7880
rect 10091 7840 10140 7868
rect 10091 7837 10103 7840
rect 10045 7831 10103 7837
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7837 10379 7871
rect 11330 7868 11336 7880
rect 11291 7840 11336 7868
rect 10321 7831 10379 7837
rect 5718 7760 5724 7812
rect 5776 7760 5782 7812
rect 8297 7803 8355 7809
rect 8297 7800 8309 7803
rect 7116 7772 8309 7800
rect 4157 7735 4215 7741
rect 4157 7701 4169 7735
rect 4203 7732 4215 7735
rect 4246 7732 4252 7744
rect 4203 7704 4252 7732
rect 4203 7701 4215 7704
rect 4157 7695 4215 7701
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 4430 7692 4436 7744
rect 4488 7732 4494 7744
rect 7116 7732 7144 7772
rect 8297 7769 8309 7772
rect 8343 7769 8355 7803
rect 10336 7800 10364 7831
rect 11330 7828 11336 7840
rect 11388 7828 11394 7880
rect 11698 7868 11704 7880
rect 11659 7840 11704 7868
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7868 18107 7871
rect 18138 7868 18144 7880
rect 18095 7840 18144 7868
rect 18095 7837 18107 7840
rect 18049 7831 18107 7837
rect 18138 7828 18144 7840
rect 18196 7828 18202 7880
rect 18690 7868 18696 7880
rect 18651 7840 18696 7868
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 18785 7871 18843 7877
rect 18785 7837 18797 7871
rect 18831 7868 18843 7871
rect 18831 7840 19932 7868
rect 18831 7837 18843 7840
rect 18785 7831 18843 7837
rect 12342 7800 12348 7812
rect 10336 7772 12348 7800
rect 8297 7763 8355 7769
rect 12342 7760 12348 7772
rect 12400 7760 12406 7812
rect 13170 7800 13176 7812
rect 13131 7772 13176 7800
rect 13170 7760 13176 7772
rect 13228 7760 13234 7812
rect 13722 7760 13728 7812
rect 13780 7800 13786 7812
rect 14277 7803 14335 7809
rect 14277 7800 14289 7803
rect 13780 7772 14289 7800
rect 13780 7760 13786 7772
rect 14277 7769 14289 7772
rect 14323 7769 14335 7803
rect 18708 7800 18736 7828
rect 19904 7809 19932 7840
rect 20254 7828 20260 7880
rect 20312 7868 20318 7880
rect 20993 7871 21051 7877
rect 20993 7868 21005 7871
rect 20312 7840 21005 7868
rect 20312 7828 20318 7840
rect 20993 7837 21005 7840
rect 21039 7868 21051 7871
rect 21266 7868 21272 7880
rect 21039 7840 21272 7868
rect 21039 7837 21051 7840
rect 20993 7831 21051 7837
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 19797 7803 19855 7809
rect 19797 7800 19809 7803
rect 18708 7772 19809 7800
rect 14277 7763 14335 7769
rect 19797 7769 19809 7772
rect 19843 7769 19855 7803
rect 19797 7763 19855 7769
rect 19889 7803 19947 7809
rect 19889 7769 19901 7803
rect 19935 7800 19947 7803
rect 21744 7800 21772 7916
rect 21910 7896 21916 7916
rect 21968 7896 21974 7948
rect 22020 7936 22048 7976
rect 27801 7973 27813 8007
rect 27847 8004 27859 8007
rect 27982 8004 27988 8016
rect 27847 7976 27988 8004
rect 27847 7973 27859 7976
rect 27801 7967 27859 7973
rect 27982 7964 27988 7976
rect 28040 7964 28046 8016
rect 28994 7964 29000 8016
rect 29052 8004 29058 8016
rect 34256 8013 34284 8044
rect 35710 8032 35716 8044
rect 35768 8032 35774 8084
rect 35802 8032 35808 8084
rect 35860 8072 35866 8084
rect 40405 8075 40463 8081
rect 40405 8072 40417 8075
rect 35860 8044 40417 8072
rect 35860 8032 35866 8044
rect 40405 8041 40417 8044
rect 40451 8041 40463 8075
rect 42981 8075 43039 8081
rect 42981 8072 42993 8075
rect 40405 8035 40463 8041
rect 41248 8044 42993 8072
rect 34241 8007 34299 8013
rect 34241 8004 34253 8007
rect 29052 7976 34253 8004
rect 29052 7964 29058 7976
rect 34241 7973 34253 7976
rect 34287 7973 34299 8007
rect 37277 8007 37335 8013
rect 37277 8004 37289 8007
rect 34241 7967 34299 7973
rect 36372 7976 37289 8004
rect 22020 7908 22140 7936
rect 22112 7868 22140 7908
rect 24854 7896 24860 7948
rect 24912 7936 24918 7948
rect 26234 7936 26240 7948
rect 24912 7908 26240 7936
rect 24912 7896 24918 7908
rect 22112 7840 25544 7868
rect 25792 7854 25820 7908
rect 26234 7896 26240 7908
rect 26292 7936 26298 7948
rect 26510 7936 26516 7948
rect 26292 7908 26516 7936
rect 26292 7896 26298 7908
rect 26510 7896 26516 7908
rect 26568 7896 26574 7948
rect 27154 7936 27160 7948
rect 27115 7908 27160 7936
rect 27154 7896 27160 7908
rect 27212 7896 27218 7948
rect 27246 7896 27252 7948
rect 27304 7936 27310 7948
rect 33042 7936 33048 7948
rect 27304 7908 33048 7936
rect 27304 7896 27310 7908
rect 33042 7896 33048 7908
rect 33100 7896 33106 7948
rect 33134 7896 33140 7948
rect 33192 7936 33198 7948
rect 36372 7936 36400 7976
rect 37277 7973 37289 7976
rect 37323 8004 37335 8007
rect 40034 8004 40040 8016
rect 37323 7976 40040 8004
rect 37323 7973 37335 7976
rect 37277 7967 37335 7973
rect 40034 7964 40040 7976
rect 40092 7964 40098 8016
rect 40678 8004 40684 8016
rect 40144 7976 40684 8004
rect 40144 7948 40172 7976
rect 40678 7964 40684 7976
rect 40736 7964 40742 8016
rect 33192 7908 36400 7936
rect 36633 7939 36691 7945
rect 33192 7896 33198 7908
rect 36633 7905 36645 7939
rect 36679 7936 36691 7939
rect 40126 7936 40132 7948
rect 36679 7908 40132 7936
rect 36679 7905 36691 7908
rect 36633 7899 36691 7905
rect 40126 7896 40132 7908
rect 40184 7896 40190 7948
rect 40770 7936 40776 7948
rect 40731 7908 40776 7936
rect 40770 7896 40776 7908
rect 40828 7896 40834 7948
rect 21800 7803 21858 7809
rect 21800 7800 21812 7803
rect 19935 7772 21812 7800
rect 19935 7769 19947 7772
rect 19889 7763 19947 7769
rect 21800 7769 21812 7772
rect 21846 7769 21858 7803
rect 21800 7763 21858 7769
rect 22005 7803 22063 7809
rect 22005 7769 22017 7803
rect 22051 7800 22063 7803
rect 22186 7800 22192 7812
rect 22051 7772 22192 7800
rect 22051 7769 22063 7772
rect 22005 7763 22063 7769
rect 22186 7760 22192 7772
rect 22244 7800 22250 7812
rect 22244 7772 25452 7800
rect 22244 7760 22250 7772
rect 4488 7704 7144 7732
rect 4488 7692 4494 7704
rect 8570 7692 8576 7744
rect 8628 7732 8634 7744
rect 9125 7735 9183 7741
rect 9125 7732 9137 7735
rect 8628 7704 9137 7732
rect 8628 7692 8634 7704
rect 9125 7701 9137 7704
rect 9171 7701 9183 7735
rect 16942 7732 16948 7744
rect 16903 7704 16948 7732
rect 9125 7695 9183 7701
rect 16942 7692 16948 7704
rect 17000 7692 17006 7744
rect 18598 7692 18604 7744
rect 18656 7732 18662 7744
rect 19429 7735 19487 7741
rect 19429 7732 19441 7735
rect 18656 7704 19441 7732
rect 18656 7692 18662 7704
rect 19429 7701 19441 7704
rect 19475 7701 19487 7735
rect 22922 7732 22928 7744
rect 22883 7704 22928 7732
rect 19429 7695 19487 7701
rect 22922 7692 22928 7704
rect 22980 7732 22986 7744
rect 23290 7732 23296 7744
rect 22980 7704 23296 7732
rect 22980 7692 22986 7704
rect 23290 7692 23296 7704
rect 23348 7692 23354 7744
rect 25424 7741 25452 7772
rect 25409 7735 25467 7741
rect 25409 7701 25421 7735
rect 25455 7701 25467 7735
rect 25516 7732 25544 7840
rect 28442 7828 28448 7880
rect 28500 7868 28506 7880
rect 28721 7871 28779 7877
rect 28721 7868 28733 7871
rect 28500 7840 28733 7868
rect 28500 7828 28506 7840
rect 28721 7837 28733 7840
rect 28767 7837 28779 7871
rect 29089 7871 29147 7877
rect 29089 7868 29101 7871
rect 28721 7831 28779 7837
rect 28966 7840 29101 7868
rect 26881 7803 26939 7809
rect 26881 7769 26893 7803
rect 26927 7769 26939 7803
rect 26881 7763 26939 7769
rect 26896 7732 26924 7763
rect 27706 7760 27712 7812
rect 27764 7800 27770 7812
rect 28966 7800 28994 7840
rect 29089 7837 29101 7840
rect 29135 7868 29147 7871
rect 30466 7868 30472 7880
rect 29135 7840 30472 7868
rect 29135 7837 29147 7840
rect 29089 7831 29147 7837
rect 30466 7828 30472 7840
rect 30524 7828 30530 7880
rect 31573 7871 31631 7877
rect 31573 7837 31585 7871
rect 31619 7868 31631 7871
rect 33594 7868 33600 7880
rect 31619 7840 33600 7868
rect 31619 7837 31631 7840
rect 31573 7831 31631 7837
rect 33594 7828 33600 7840
rect 33652 7828 33658 7880
rect 34882 7868 34888 7880
rect 34843 7840 34888 7868
rect 34882 7828 34888 7840
rect 34940 7828 34946 7880
rect 37734 7828 37740 7880
rect 37792 7868 37798 7880
rect 39393 7871 39451 7877
rect 39393 7868 39405 7871
rect 37792 7840 39405 7868
rect 37792 7828 37798 7840
rect 39393 7837 39405 7840
rect 39439 7837 39451 7871
rect 39393 7831 39451 7837
rect 40034 7828 40040 7880
rect 40092 7868 40098 7880
rect 40681 7871 40739 7877
rect 40681 7868 40693 7871
rect 40092 7840 40693 7868
rect 40092 7828 40098 7840
rect 40681 7837 40693 7840
rect 40727 7868 40739 7871
rect 41248 7868 41276 8044
rect 42981 8041 42993 8044
rect 43027 8072 43039 8075
rect 43070 8072 43076 8084
rect 43027 8044 43076 8072
rect 43027 8041 43039 8044
rect 42981 8035 43039 8041
rect 43070 8032 43076 8044
rect 43128 8072 43134 8084
rect 45646 8072 45652 8084
rect 43128 8044 45652 8072
rect 43128 8032 43134 8044
rect 45646 8032 45652 8044
rect 45704 8032 45710 8084
rect 47210 8032 47216 8084
rect 47268 8072 47274 8084
rect 47949 8075 48007 8081
rect 47949 8072 47961 8075
rect 47268 8044 47961 8072
rect 47268 8032 47274 8044
rect 47949 8041 47961 8044
rect 47995 8041 48007 8075
rect 48222 8072 48228 8084
rect 48183 8044 48228 8072
rect 47949 8035 48007 8041
rect 48222 8032 48228 8044
rect 48280 8032 48286 8084
rect 49234 8072 49240 8084
rect 49195 8044 49240 8072
rect 49234 8032 49240 8044
rect 49292 8032 49298 8084
rect 49694 8072 49700 8084
rect 49655 8044 49700 8072
rect 49694 8032 49700 8044
rect 49752 8032 49758 8084
rect 49970 8032 49976 8084
rect 50028 8072 50034 8084
rect 50985 8075 51043 8081
rect 50985 8072 50997 8075
rect 50028 8044 50997 8072
rect 50028 8032 50034 8044
rect 50985 8041 50997 8044
rect 51031 8041 51043 8075
rect 52178 8072 52184 8084
rect 52139 8044 52184 8072
rect 50985 8035 51043 8041
rect 52178 8032 52184 8044
rect 52236 8032 52242 8084
rect 52365 8075 52423 8081
rect 52365 8041 52377 8075
rect 52411 8072 52423 8075
rect 53190 8072 53196 8084
rect 52411 8044 53196 8072
rect 52411 8041 52423 8044
rect 52365 8035 52423 8041
rect 53190 8032 53196 8044
rect 53248 8032 53254 8084
rect 54849 8075 54907 8081
rect 54849 8041 54861 8075
rect 54895 8072 54907 8075
rect 55490 8072 55496 8084
rect 54895 8044 55496 8072
rect 54895 8041 54907 8044
rect 54849 8035 54907 8041
rect 55490 8032 55496 8044
rect 55548 8032 55554 8084
rect 58069 8075 58127 8081
rect 58069 8041 58081 8075
rect 58115 8072 58127 8075
rect 58894 8072 58900 8084
rect 58115 8044 58900 8072
rect 58115 8041 58127 8044
rect 58069 8035 58127 8041
rect 58894 8032 58900 8044
rect 58952 8032 58958 8084
rect 61010 8072 61016 8084
rect 59832 8044 61016 8072
rect 42610 7964 42616 8016
rect 42668 8004 42674 8016
rect 45281 8007 45339 8013
rect 45281 8004 45293 8007
rect 42668 7976 45293 8004
rect 42668 7964 42674 7976
rect 45281 7973 45293 7976
rect 45327 7973 45339 8007
rect 46937 8007 46995 8013
rect 46937 8004 46949 8007
rect 45281 7967 45339 7973
rect 45756 7976 46949 8004
rect 41340 7908 42840 7936
rect 41340 7877 41368 7908
rect 40727 7840 41276 7868
rect 41325 7871 41383 7877
rect 40727 7837 40739 7840
rect 40681 7831 40739 7837
rect 41325 7837 41337 7871
rect 41371 7837 41383 7871
rect 41598 7868 41604 7880
rect 41511 7840 41604 7868
rect 41325 7831 41383 7837
rect 41598 7828 41604 7840
rect 41656 7868 41662 7880
rect 42518 7868 42524 7880
rect 41656 7840 42524 7868
rect 41656 7828 41662 7840
rect 42518 7828 42524 7840
rect 42576 7828 42582 7880
rect 29822 7800 29828 7812
rect 27764 7772 28994 7800
rect 29783 7772 29828 7800
rect 27764 7760 27770 7772
rect 29822 7760 29828 7772
rect 29880 7760 29886 7812
rect 32033 7803 32091 7809
rect 32033 7769 32045 7803
rect 32079 7769 32091 7803
rect 32033 7763 32091 7769
rect 25516 7704 26924 7732
rect 25409 7695 25467 7701
rect 28718 7692 28724 7744
rect 28776 7732 28782 7744
rect 28813 7735 28871 7741
rect 28813 7732 28825 7735
rect 28776 7704 28825 7732
rect 28776 7692 28782 7704
rect 28813 7701 28825 7704
rect 28859 7701 28871 7735
rect 28813 7695 28871 7701
rect 28902 7692 28908 7744
rect 28960 7732 28966 7744
rect 29840 7732 29868 7760
rect 32048 7732 32076 7763
rect 33502 7760 33508 7812
rect 33560 7800 33566 7812
rect 34514 7800 34520 7812
rect 33560 7772 34520 7800
rect 33560 7760 33566 7772
rect 34514 7760 34520 7772
rect 34572 7760 34578 7812
rect 35161 7803 35219 7809
rect 35161 7769 35173 7803
rect 35207 7769 35219 7803
rect 35161 7763 35219 7769
rect 28960 7704 29005 7732
rect 29840 7704 32076 7732
rect 35176 7732 35204 7763
rect 35618 7760 35624 7812
rect 35676 7760 35682 7812
rect 37458 7760 37464 7812
rect 37516 7800 37522 7812
rect 38289 7803 38347 7809
rect 38289 7800 38301 7803
rect 37516 7772 38301 7800
rect 37516 7760 37522 7772
rect 38289 7769 38301 7772
rect 38335 7769 38347 7803
rect 40052 7800 40080 7828
rect 38289 7763 38347 7769
rect 38626 7772 40080 7800
rect 36538 7732 36544 7744
rect 35176 7704 36544 7732
rect 28960 7692 28966 7704
rect 36538 7692 36544 7704
rect 36596 7692 36602 7744
rect 36630 7692 36636 7744
rect 36688 7732 36694 7744
rect 37737 7735 37795 7741
rect 37737 7732 37749 7735
rect 36688 7704 37749 7732
rect 36688 7692 36694 7704
rect 37737 7701 37749 7704
rect 37783 7732 37795 7735
rect 38626 7732 38654 7772
rect 40954 7760 40960 7812
rect 41012 7800 41018 7812
rect 41417 7803 41475 7809
rect 41417 7800 41429 7803
rect 41012 7772 41429 7800
rect 41012 7760 41018 7772
rect 41417 7769 41429 7772
rect 41463 7769 41475 7803
rect 42705 7803 42763 7809
rect 42705 7800 42717 7803
rect 41417 7763 41475 7769
rect 41708 7772 42717 7800
rect 37783 7704 38654 7732
rect 38933 7735 38991 7741
rect 37783 7701 37795 7704
rect 37737 7695 37795 7701
rect 38933 7701 38945 7735
rect 38979 7732 38991 7735
rect 39114 7732 39120 7744
rect 38979 7704 39120 7732
rect 38979 7701 38991 7704
rect 38933 7695 38991 7701
rect 39114 7692 39120 7704
rect 39172 7692 39178 7744
rect 41322 7692 41328 7744
rect 41380 7732 41386 7744
rect 41708 7732 41736 7772
rect 42705 7769 42717 7772
rect 42751 7769 42763 7803
rect 42812 7800 42840 7908
rect 42886 7896 42892 7948
rect 42944 7936 42950 7948
rect 45370 7936 45376 7948
rect 42944 7908 45376 7936
rect 42944 7896 42950 7908
rect 45370 7896 45376 7908
rect 45428 7896 45434 7948
rect 45756 7945 45784 7976
rect 46937 7973 46949 7976
rect 46983 7973 46995 8007
rect 46937 7967 46995 7973
rect 47026 7964 47032 8016
rect 47084 8004 47090 8016
rect 47084 7976 47129 8004
rect 47084 7964 47090 7976
rect 47394 7964 47400 8016
rect 47452 8004 47458 8016
rect 49712 8004 49740 8032
rect 53374 8004 53380 8016
rect 47452 7976 49740 8004
rect 50172 7976 53380 8004
rect 47452 7964 47458 7976
rect 45741 7939 45799 7945
rect 45741 7905 45753 7939
rect 45787 7905 45799 7939
rect 45741 7899 45799 7905
rect 45830 7896 45836 7948
rect 45888 7936 45894 7948
rect 46845 7939 46903 7945
rect 46845 7936 46857 7939
rect 45888 7908 46857 7936
rect 45888 7896 45894 7908
rect 46845 7905 46857 7908
rect 46891 7936 46903 7939
rect 47210 7936 47216 7948
rect 46891 7908 47216 7936
rect 46891 7905 46903 7908
rect 46845 7899 46903 7905
rect 47210 7896 47216 7908
rect 47268 7896 47274 7948
rect 49326 7936 49332 7948
rect 47320 7908 49332 7936
rect 42978 7828 42984 7880
rect 43036 7868 43042 7880
rect 43806 7868 43812 7880
rect 43036 7840 43812 7868
rect 43036 7828 43042 7840
rect 43806 7828 43812 7840
rect 43864 7828 43870 7880
rect 45646 7868 45652 7880
rect 45607 7840 45652 7868
rect 45646 7828 45652 7840
rect 45704 7828 45710 7880
rect 47026 7828 47032 7880
rect 47084 7868 47090 7880
rect 47121 7871 47179 7877
rect 47121 7868 47133 7871
rect 47084 7840 47133 7868
rect 47084 7828 47090 7840
rect 47121 7837 47133 7840
rect 47167 7868 47179 7871
rect 47320 7868 47348 7908
rect 49326 7896 49332 7908
rect 49384 7896 49390 7948
rect 49694 7896 49700 7948
rect 49752 7936 49758 7948
rect 50172 7936 50200 7976
rect 53374 7964 53380 7976
rect 53432 8004 53438 8016
rect 54021 8007 54079 8013
rect 54021 8004 54033 8007
rect 53432 7976 54033 8004
rect 53432 7964 53438 7976
rect 54021 7973 54033 7976
rect 54067 7973 54079 8007
rect 54021 7967 54079 7973
rect 57698 7964 57704 8016
rect 57756 8004 57762 8016
rect 59832 8004 59860 8044
rect 61010 8032 61016 8044
rect 61068 8032 61074 8084
rect 61102 8032 61108 8084
rect 61160 8072 61166 8084
rect 62393 8075 62451 8081
rect 62393 8072 62405 8075
rect 61160 8044 62405 8072
rect 61160 8032 61166 8044
rect 62393 8041 62405 8044
rect 62439 8041 62451 8075
rect 62393 8035 62451 8041
rect 66349 8075 66407 8081
rect 66349 8041 66361 8075
rect 66395 8072 66407 8075
rect 66395 8044 72188 8072
rect 66395 8041 66407 8044
rect 66349 8035 66407 8041
rect 57756 7976 59860 8004
rect 59909 8007 59967 8013
rect 57756 7964 57762 7976
rect 59909 7973 59921 8007
rect 59955 8004 59967 8007
rect 60090 8004 60096 8016
rect 59955 7976 60096 8004
rect 59955 7973 59967 7976
rect 59909 7967 59967 7973
rect 60090 7964 60096 7976
rect 60148 7964 60154 8016
rect 66254 8004 66260 8016
rect 63328 7976 66260 8004
rect 52638 7936 52644 7948
rect 49752 7908 50200 7936
rect 50264 7908 52644 7936
rect 49752 7896 49758 7908
rect 48222 7868 48228 7880
rect 47167 7840 47348 7868
rect 48183 7840 48228 7868
rect 47167 7837 47179 7840
rect 47121 7831 47179 7837
rect 48222 7828 48228 7840
rect 48280 7828 48286 7880
rect 48314 7828 48320 7880
rect 48372 7868 48378 7880
rect 48372 7840 48417 7868
rect 48372 7828 48378 7840
rect 46842 7800 46848 7812
rect 42812 7772 46848 7800
rect 42705 7763 42763 7769
rect 41380 7704 41736 7732
rect 41785 7735 41843 7741
rect 41380 7692 41386 7704
rect 41785 7701 41797 7735
rect 41831 7732 41843 7735
rect 42886 7732 42892 7744
rect 41831 7704 42892 7732
rect 41831 7701 41843 7704
rect 41785 7695 41843 7701
rect 42886 7692 42892 7704
rect 42944 7692 42950 7744
rect 43180 7741 43208 7772
rect 46842 7760 46848 7772
rect 46900 7760 46906 7812
rect 47210 7760 47216 7812
rect 47268 7800 47274 7812
rect 50264 7800 50292 7908
rect 52638 7896 52644 7908
rect 52696 7896 52702 7948
rect 52730 7896 52736 7948
rect 52788 7936 52794 7948
rect 53469 7939 53527 7945
rect 53469 7936 53481 7939
rect 52788 7908 53481 7936
rect 52788 7896 52794 7908
rect 53469 7905 53481 7908
rect 53515 7905 53527 7939
rect 53469 7899 53527 7905
rect 55306 7896 55312 7948
rect 55364 7936 55370 7948
rect 56321 7939 56379 7945
rect 56321 7936 56333 7939
rect 55364 7908 56333 7936
rect 55364 7896 55370 7908
rect 56321 7905 56333 7908
rect 56367 7905 56379 7939
rect 56321 7899 56379 7905
rect 56597 7939 56655 7945
rect 56597 7905 56609 7939
rect 56643 7936 56655 7939
rect 57146 7936 57152 7948
rect 56643 7908 57152 7936
rect 56643 7905 56655 7908
rect 56597 7899 56655 7905
rect 57146 7896 57152 7908
rect 57204 7896 57210 7948
rect 57330 7896 57336 7948
rect 57388 7936 57394 7948
rect 57388 7908 58940 7936
rect 57388 7896 57394 7908
rect 51166 7828 51172 7880
rect 51224 7877 51230 7880
rect 51224 7871 51246 7877
rect 51234 7837 51246 7871
rect 51224 7831 51246 7837
rect 51224 7828 51230 7831
rect 51442 7828 51448 7880
rect 51500 7868 51506 7880
rect 53009 7871 53067 7877
rect 51500 7840 52132 7868
rect 51500 7828 51506 7840
rect 50430 7800 50436 7812
rect 47268 7772 50292 7800
rect 50343 7772 50436 7800
rect 47268 7760 47274 7772
rect 50430 7760 50436 7772
rect 50488 7800 50494 7812
rect 50982 7800 50988 7812
rect 50488 7772 50988 7800
rect 50488 7760 50494 7772
rect 50982 7760 50988 7772
rect 51040 7760 51046 7812
rect 51350 7800 51356 7812
rect 51311 7772 51356 7800
rect 51350 7760 51356 7772
rect 51408 7760 51414 7812
rect 51810 7760 51816 7812
rect 51868 7800 51874 7812
rect 51997 7803 52055 7809
rect 51997 7800 52009 7803
rect 51868 7772 52009 7800
rect 51868 7760 51874 7772
rect 51997 7769 52009 7772
rect 52043 7769 52055 7803
rect 52104 7800 52132 7840
rect 53009 7837 53021 7871
rect 53055 7868 53067 7871
rect 53190 7868 53196 7880
rect 53055 7840 53196 7868
rect 53055 7837 53067 7840
rect 53009 7831 53067 7837
rect 53190 7828 53196 7840
rect 53248 7868 53254 7880
rect 54846 7868 54852 7880
rect 53248 7840 54852 7868
rect 53248 7828 53254 7840
rect 54846 7828 54852 7840
rect 54904 7828 54910 7880
rect 54941 7871 54999 7877
rect 54941 7837 54953 7871
rect 54987 7837 54999 7871
rect 54941 7831 54999 7837
rect 53926 7800 53932 7812
rect 52104 7772 53932 7800
rect 51997 7763 52055 7769
rect 53926 7760 53932 7772
rect 53984 7760 53990 7812
rect 54956 7800 54984 7831
rect 55674 7828 55680 7880
rect 55732 7868 55738 7880
rect 55861 7871 55919 7877
rect 55861 7868 55873 7871
rect 55732 7840 55873 7868
rect 55732 7828 55738 7840
rect 55861 7837 55873 7840
rect 55907 7868 55919 7871
rect 55907 7840 56364 7868
rect 55907 7837 55919 7840
rect 55861 7831 55919 7837
rect 55950 7800 55956 7812
rect 54956 7772 55956 7800
rect 55950 7760 55956 7772
rect 56008 7760 56014 7812
rect 43165 7735 43223 7741
rect 43165 7701 43177 7735
rect 43211 7701 43223 7735
rect 44082 7732 44088 7744
rect 44043 7704 44088 7732
rect 43165 7695 43223 7701
rect 44082 7692 44088 7704
rect 44140 7692 44146 7744
rect 44174 7692 44180 7744
rect 44232 7732 44238 7744
rect 44637 7735 44695 7741
rect 44637 7732 44649 7735
rect 44232 7704 44649 7732
rect 44232 7692 44238 7704
rect 44637 7701 44649 7704
rect 44683 7732 44695 7735
rect 46385 7735 46443 7741
rect 46385 7732 46397 7735
rect 44683 7704 46397 7732
rect 44683 7701 44695 7704
rect 44637 7695 44695 7701
rect 46385 7701 46397 7704
rect 46431 7732 46443 7735
rect 48866 7732 48872 7744
rect 46431 7704 48872 7732
rect 46431 7701 46443 7704
rect 46385 7695 46443 7701
rect 48866 7692 48872 7704
rect 48924 7732 48930 7744
rect 51902 7732 51908 7744
rect 48924 7704 51908 7732
rect 48924 7692 48930 7704
rect 51902 7692 51908 7704
rect 51960 7692 51966 7744
rect 52086 7692 52092 7744
rect 52144 7732 52150 7744
rect 52197 7735 52255 7741
rect 52197 7732 52209 7735
rect 52144 7704 52209 7732
rect 52144 7692 52150 7704
rect 52197 7701 52209 7704
rect 52243 7701 52255 7735
rect 52914 7732 52920 7744
rect 52875 7704 52920 7732
rect 52197 7695 52255 7701
rect 52914 7692 52920 7704
rect 52972 7692 52978 7744
rect 55769 7735 55827 7741
rect 55769 7701 55781 7735
rect 55815 7732 55827 7735
rect 55858 7732 55864 7744
rect 55815 7704 55864 7732
rect 55815 7701 55827 7704
rect 55769 7695 55827 7701
rect 55858 7692 55864 7704
rect 55916 7692 55922 7744
rect 56336 7732 56364 7840
rect 58802 7800 58808 7812
rect 57822 7772 58808 7800
rect 58802 7760 58808 7772
rect 58860 7760 58866 7812
rect 58912 7800 58940 7908
rect 59170 7896 59176 7948
rect 59228 7936 59234 7948
rect 59449 7939 59507 7945
rect 59449 7936 59461 7939
rect 59228 7908 59461 7936
rect 59228 7896 59234 7908
rect 59449 7905 59461 7908
rect 59495 7905 59507 7939
rect 60918 7936 60924 7948
rect 60879 7908 60924 7936
rect 59449 7899 59507 7905
rect 60918 7896 60924 7908
rect 60976 7896 60982 7948
rect 61010 7896 61016 7948
rect 61068 7936 61074 7948
rect 63328 7945 63356 7976
rect 66254 7964 66260 7976
rect 66312 7964 66318 8016
rect 69106 8004 69112 8016
rect 69067 7976 69112 8004
rect 69106 7964 69112 7976
rect 69164 7964 69170 8016
rect 71317 8007 71375 8013
rect 71317 7973 71329 8007
rect 71363 8004 71375 8007
rect 71866 8004 71872 8016
rect 71363 7976 71872 8004
rect 71363 7973 71375 7976
rect 71317 7967 71375 7973
rect 71866 7964 71872 7976
rect 71924 7964 71930 8016
rect 63313 7939 63371 7945
rect 63313 7936 63325 7939
rect 61068 7908 63325 7936
rect 61068 7896 61074 7908
rect 63313 7905 63325 7908
rect 63359 7905 63371 7939
rect 66070 7936 66076 7948
rect 63313 7899 63371 7905
rect 63604 7908 65380 7936
rect 66031 7908 66076 7936
rect 59541 7871 59599 7877
rect 59541 7837 59553 7871
rect 59587 7868 59599 7871
rect 60182 7868 60188 7880
rect 59587 7840 60188 7868
rect 59587 7837 59599 7840
rect 59541 7831 59599 7837
rect 60182 7828 60188 7840
rect 60240 7828 60246 7880
rect 60642 7868 60648 7880
rect 60603 7840 60648 7868
rect 60642 7828 60648 7840
rect 60700 7828 60706 7880
rect 62206 7828 62212 7880
rect 62264 7868 62270 7880
rect 63604 7868 63632 7908
rect 62264 7840 63632 7868
rect 62264 7828 62270 7840
rect 65150 7828 65156 7880
rect 65208 7868 65214 7880
rect 65352 7868 65380 7908
rect 66070 7896 66076 7908
rect 66128 7896 66134 7948
rect 66346 7896 66352 7948
rect 66404 7936 66410 7948
rect 67266 7936 67272 7948
rect 66404 7908 67272 7936
rect 66404 7896 66410 7908
rect 67266 7896 67272 7908
rect 67324 7936 67330 7948
rect 67361 7939 67419 7945
rect 67361 7936 67373 7939
rect 67324 7908 67373 7936
rect 67324 7896 67330 7908
rect 67361 7905 67373 7908
rect 67407 7905 67419 7939
rect 67361 7899 67419 7905
rect 67637 7939 67695 7945
rect 67637 7905 67649 7939
rect 67683 7936 67695 7939
rect 69661 7939 69719 7945
rect 69661 7936 69673 7939
rect 67683 7908 69673 7936
rect 67683 7905 67695 7908
rect 67637 7899 67695 7905
rect 69661 7905 69673 7908
rect 69707 7905 69719 7939
rect 69661 7899 69719 7905
rect 65981 7871 66039 7877
rect 65981 7868 65993 7871
rect 65208 7840 65253 7868
rect 65352 7840 65993 7868
rect 65208 7828 65214 7840
rect 65981 7837 65993 7840
rect 66027 7837 66039 7871
rect 69750 7868 69756 7880
rect 69711 7840 69756 7868
rect 65981 7831 66039 7837
rect 69750 7828 69756 7840
rect 69808 7828 69814 7880
rect 70397 7871 70455 7877
rect 70397 7837 70409 7871
rect 70443 7868 70455 7871
rect 70578 7868 70584 7880
rect 70443 7840 70584 7868
rect 70443 7837 70455 7840
rect 70397 7831 70455 7837
rect 70578 7828 70584 7840
rect 70636 7828 70642 7880
rect 71498 7868 71504 7880
rect 71459 7840 71504 7868
rect 71498 7828 71504 7840
rect 71556 7828 71562 7880
rect 71866 7828 71872 7880
rect 71924 7868 71930 7880
rect 72160 7877 72188 8044
rect 73154 8032 73160 8084
rect 73212 8072 73218 8084
rect 73212 8044 76236 8072
rect 73212 8032 73218 8044
rect 72970 7964 72976 8016
rect 73028 8004 73034 8016
rect 75365 8007 75423 8013
rect 75365 8004 75377 8007
rect 73028 7976 75377 8004
rect 73028 7964 73034 7976
rect 75365 7973 75377 7976
rect 75411 7973 75423 8007
rect 75365 7967 75423 7973
rect 76208 8004 76236 8044
rect 76466 8032 76472 8084
rect 76524 8072 76530 8084
rect 79042 8072 79048 8084
rect 76524 8044 79048 8072
rect 76524 8032 76530 8044
rect 79042 8032 79048 8044
rect 79100 8032 79106 8084
rect 79137 8075 79195 8081
rect 79137 8041 79149 8075
rect 79183 8072 79195 8075
rect 79183 8044 84424 8072
rect 79183 8041 79195 8044
rect 79137 8035 79195 8041
rect 78858 8004 78864 8016
rect 76208 7976 78864 8004
rect 74718 7936 74724 7948
rect 74679 7908 74724 7936
rect 74718 7896 74724 7908
rect 74776 7896 74782 7948
rect 76208 7945 76236 7976
rect 78858 7964 78864 7976
rect 78916 7964 78922 8016
rect 79965 8007 80023 8013
rect 79965 7973 79977 8007
rect 80011 8004 80023 8007
rect 80517 8007 80575 8013
rect 80517 8004 80529 8007
rect 80011 7976 80529 8004
rect 80011 7973 80023 7976
rect 79965 7967 80023 7973
rect 80517 7973 80529 7976
rect 80563 7973 80575 8007
rect 80517 7967 80575 7973
rect 81710 7964 81716 8016
rect 81768 8004 81774 8016
rect 81768 7976 84148 8004
rect 81768 7964 81774 7976
rect 84120 7948 84148 7976
rect 76193 7939 76251 7945
rect 76193 7905 76205 7939
rect 76239 7905 76251 7939
rect 76193 7899 76251 7905
rect 76282 7896 76288 7948
rect 76340 7936 76346 7948
rect 78033 7939 78091 7945
rect 78033 7936 78045 7939
rect 76340 7908 78045 7936
rect 76340 7896 76346 7908
rect 78033 7905 78045 7908
rect 78079 7905 78091 7939
rect 78033 7899 78091 7905
rect 78122 7896 78128 7948
rect 78180 7936 78186 7948
rect 78769 7939 78827 7945
rect 78769 7936 78781 7939
rect 78180 7908 78781 7936
rect 78180 7896 78186 7908
rect 78769 7905 78781 7908
rect 78815 7905 78827 7939
rect 80701 7939 80759 7945
rect 80701 7936 80713 7939
rect 78769 7899 78827 7905
rect 80532 7908 80713 7936
rect 80532 7880 80560 7908
rect 80701 7905 80713 7908
rect 80747 7905 80759 7939
rect 81434 7936 81440 7948
rect 81395 7908 81440 7936
rect 80701 7899 80759 7905
rect 81434 7896 81440 7908
rect 81492 7896 81498 7948
rect 83826 7936 83832 7948
rect 83787 7908 83832 7936
rect 83826 7896 83832 7908
rect 83884 7896 83890 7948
rect 84102 7936 84108 7948
rect 84015 7908 84108 7936
rect 84102 7896 84108 7908
rect 84160 7896 84166 7948
rect 84396 7936 84424 8044
rect 84838 8032 84844 8084
rect 84896 8072 84902 8084
rect 92842 8072 92848 8084
rect 84896 8044 92848 8072
rect 84896 8032 84902 8044
rect 86678 8004 86684 8016
rect 86639 7976 86684 8004
rect 86678 7964 86684 7976
rect 86736 7964 86742 8016
rect 88996 7945 89024 8044
rect 92842 8032 92848 8044
rect 92900 8032 92906 8084
rect 93578 8081 93584 8084
rect 93535 8075 93584 8081
rect 93535 8041 93547 8075
rect 93581 8041 93584 8075
rect 93535 8035 93584 8041
rect 93578 8032 93584 8035
rect 93636 8032 93642 8084
rect 88705 7939 88763 7945
rect 88705 7936 88717 7939
rect 84396 7908 88717 7936
rect 88705 7905 88717 7908
rect 88751 7905 88763 7939
rect 88705 7899 88763 7905
rect 88981 7939 89039 7945
rect 88981 7905 88993 7939
rect 89027 7905 89039 7939
rect 89438 7936 89444 7948
rect 89399 7908 89444 7936
rect 88981 7899 89039 7905
rect 89438 7896 89444 7908
rect 89496 7896 89502 7948
rect 91186 7896 91192 7948
rect 91244 7936 91250 7948
rect 92109 7939 92167 7945
rect 92109 7936 92121 7939
rect 91244 7908 92121 7936
rect 91244 7896 91250 7908
rect 92109 7905 92121 7908
rect 92155 7905 92167 7939
rect 92474 7936 92480 7948
rect 92109 7899 92167 7905
rect 92216 7908 92480 7936
rect 72053 7871 72111 7877
rect 71924 7862 72004 7868
rect 72053 7862 72065 7871
rect 71924 7840 72065 7862
rect 71924 7828 71930 7840
rect 71976 7837 72065 7840
rect 72099 7837 72111 7871
rect 71976 7834 72111 7837
rect 72053 7831 72111 7834
rect 72159 7871 72217 7877
rect 72159 7837 72171 7871
rect 72205 7837 72217 7871
rect 72159 7831 72217 7837
rect 72329 7871 72387 7877
rect 72329 7837 72341 7871
rect 72375 7837 72387 7871
rect 72329 7831 72387 7837
rect 58912 7772 60734 7800
rect 58342 7732 58348 7744
rect 56336 7704 58348 7732
rect 58342 7692 58348 7704
rect 58400 7732 58406 7744
rect 58529 7735 58587 7741
rect 58529 7732 58541 7735
rect 58400 7704 58541 7732
rect 58400 7692 58406 7704
rect 58529 7701 58541 7704
rect 58575 7732 58587 7735
rect 59170 7732 59176 7744
rect 58575 7704 59176 7732
rect 58575 7701 58587 7704
rect 58529 7695 58587 7701
rect 59170 7692 59176 7704
rect 59228 7692 59234 7744
rect 60706 7732 60734 7772
rect 61930 7760 61936 7812
rect 61988 7760 61994 7812
rect 62666 7760 62672 7812
rect 62724 7800 62730 7812
rect 64969 7803 65027 7809
rect 62724 7772 64920 7800
rect 62724 7760 62730 7772
rect 64782 7732 64788 7744
rect 60706 7704 64788 7732
rect 64782 7692 64788 7704
rect 64840 7692 64846 7744
rect 64892 7732 64920 7772
rect 64969 7769 64981 7803
rect 65015 7800 65027 7803
rect 67634 7800 67640 7812
rect 65015 7772 67640 7800
rect 65015 7769 65027 7772
rect 64969 7763 65027 7769
rect 67634 7760 67640 7772
rect 67692 7760 67698 7812
rect 70305 7803 70363 7809
rect 70305 7800 70317 7803
rect 68862 7772 70317 7800
rect 70305 7769 70317 7772
rect 70351 7769 70363 7803
rect 70305 7763 70363 7769
rect 66901 7735 66959 7741
rect 66901 7732 66913 7735
rect 64892 7704 66913 7732
rect 66901 7701 66913 7704
rect 66947 7732 66959 7735
rect 67726 7732 67732 7744
rect 66947 7704 67732 7732
rect 66947 7701 66959 7704
rect 66901 7695 66959 7701
rect 67726 7692 67732 7704
rect 67784 7692 67790 7744
rect 67910 7692 67916 7744
rect 67968 7732 67974 7744
rect 72344 7732 72372 7831
rect 72418 7828 72424 7880
rect 72476 7868 72482 7880
rect 73065 7871 73123 7877
rect 72476 7840 72521 7868
rect 72476 7828 72482 7840
rect 73065 7837 73077 7871
rect 73111 7868 73123 7871
rect 73154 7868 73160 7880
rect 73111 7840 73160 7868
rect 73111 7837 73123 7840
rect 73065 7831 73123 7837
rect 73154 7828 73160 7840
rect 73212 7828 73218 7880
rect 74902 7828 74908 7880
rect 74960 7868 74966 7880
rect 74960 7840 75005 7868
rect 74960 7828 74966 7840
rect 78674 7828 78680 7880
rect 78732 7868 78738 7880
rect 78861 7871 78919 7877
rect 78861 7868 78873 7871
rect 78732 7840 78873 7868
rect 78732 7828 78738 7840
rect 78861 7837 78873 7840
rect 78907 7868 78919 7871
rect 79781 7871 79839 7877
rect 79781 7868 79793 7871
rect 78907 7840 79793 7868
rect 78907 7837 78919 7840
rect 78861 7831 78919 7837
rect 79781 7837 79793 7840
rect 79827 7868 79839 7871
rect 79870 7868 79876 7880
rect 79827 7840 79876 7868
rect 79827 7837 79839 7840
rect 79781 7831 79839 7837
rect 79870 7828 79876 7840
rect 79928 7828 79934 7880
rect 79965 7871 80023 7877
rect 79965 7837 79977 7871
rect 80011 7837 80023 7871
rect 79965 7831 80023 7837
rect 76466 7800 76472 7812
rect 72436 7772 76472 7800
rect 72436 7744 72464 7772
rect 76466 7760 76472 7772
rect 76524 7760 76530 7812
rect 77849 7803 77907 7809
rect 77849 7769 77861 7803
rect 77895 7800 77907 7803
rect 78582 7800 78588 7812
rect 77895 7772 78588 7800
rect 77895 7769 77907 7772
rect 77849 7763 77907 7769
rect 78582 7760 78588 7772
rect 78640 7760 78646 7812
rect 79980 7800 80008 7831
rect 80054 7828 80060 7880
rect 80112 7868 80118 7880
rect 80425 7871 80483 7877
rect 80425 7868 80437 7871
rect 80112 7840 80437 7868
rect 80112 7828 80118 7840
rect 80425 7837 80437 7840
rect 80471 7837 80483 7871
rect 80425 7831 80483 7837
rect 80514 7828 80520 7880
rect 80572 7828 80578 7880
rect 82630 7868 82636 7880
rect 82591 7840 82636 7868
rect 82630 7828 82636 7840
rect 82688 7828 82694 7880
rect 82814 7828 82820 7880
rect 82872 7868 82878 7880
rect 82909 7871 82967 7877
rect 82909 7868 82921 7871
rect 82872 7840 82921 7868
rect 82872 7828 82878 7840
rect 82909 7837 82921 7840
rect 82955 7837 82967 7871
rect 83642 7868 83648 7880
rect 83603 7840 83648 7868
rect 82909 7831 82967 7837
rect 83642 7828 83648 7840
rect 83700 7828 83706 7880
rect 86126 7828 86132 7880
rect 86184 7868 86190 7880
rect 86497 7871 86555 7877
rect 86497 7868 86509 7871
rect 86184 7840 86509 7868
rect 86184 7828 86190 7840
rect 86497 7837 86509 7840
rect 86543 7837 86555 7871
rect 86497 7831 86555 7837
rect 89714 7828 89720 7880
rect 89772 7868 89778 7880
rect 90450 7868 90456 7880
rect 89772 7840 89817 7868
rect 90411 7840 90456 7868
rect 89772 7828 89778 7840
rect 90450 7828 90456 7840
rect 90508 7828 90514 7880
rect 91741 7871 91799 7877
rect 91741 7837 91753 7871
rect 91787 7868 91799 7871
rect 92216 7868 92244 7908
rect 92474 7896 92480 7908
rect 92532 7896 92538 7948
rect 91787 7840 92244 7868
rect 91787 7837 91799 7840
rect 91741 7831 91799 7837
rect 79980 7772 80928 7800
rect 67968 7704 72372 7732
rect 67968 7692 67974 7704
rect 72418 7692 72424 7744
rect 72476 7692 72482 7744
rect 72605 7735 72663 7741
rect 72605 7701 72617 7735
rect 72651 7732 72663 7735
rect 74626 7732 74632 7744
rect 72651 7704 74632 7732
rect 72651 7701 72663 7704
rect 72605 7695 72663 7701
rect 74626 7692 74632 7704
rect 74684 7692 74690 7744
rect 77662 7692 77668 7744
rect 77720 7732 77726 7744
rect 80026 7732 80054 7772
rect 77720 7704 80054 7732
rect 77720 7692 77726 7704
rect 80422 7692 80428 7744
rect 80480 7732 80486 7744
rect 80701 7735 80759 7741
rect 80701 7732 80713 7735
rect 80480 7704 80713 7732
rect 80480 7692 80486 7704
rect 80701 7701 80713 7704
rect 80747 7701 80759 7735
rect 80900 7732 80928 7772
rect 82170 7760 82176 7812
rect 82228 7800 82234 7812
rect 84838 7800 84844 7812
rect 82228 7772 84844 7800
rect 82228 7760 82234 7772
rect 84838 7760 84844 7772
rect 84896 7760 84902 7812
rect 88426 7800 88432 7812
rect 88274 7772 88432 7800
rect 88426 7760 88432 7772
rect 88484 7800 88490 7812
rect 89254 7800 89260 7812
rect 88484 7772 89260 7800
rect 88484 7760 88490 7772
rect 89254 7760 89260 7772
rect 89312 7800 89318 7812
rect 89622 7800 89628 7812
rect 89312 7772 89628 7800
rect 89312 7760 89318 7772
rect 89622 7760 89628 7772
rect 89680 7800 89686 7812
rect 90468 7800 90496 7828
rect 89680 7772 90496 7800
rect 89680 7760 89686 7772
rect 90818 7760 90824 7812
rect 90876 7800 90882 7812
rect 91756 7800 91784 7831
rect 93394 7828 93400 7880
rect 93452 7868 93458 7880
rect 94041 7871 94099 7877
rect 94041 7868 94053 7871
rect 93452 7840 94053 7868
rect 93452 7828 93458 7840
rect 94041 7837 94053 7840
rect 94087 7837 94099 7871
rect 94041 7831 94099 7837
rect 90876 7772 91784 7800
rect 90876 7760 90882 7772
rect 93026 7760 93032 7812
rect 93084 7760 93090 7812
rect 84378 7732 84384 7744
rect 80900 7704 84384 7732
rect 80701 7695 80759 7701
rect 84378 7692 84384 7704
rect 84436 7692 84442 7744
rect 87230 7732 87236 7744
rect 87191 7704 87236 7732
rect 87230 7692 87236 7704
rect 87288 7692 87294 7744
rect 90637 7735 90695 7741
rect 90637 7701 90649 7735
rect 90683 7732 90695 7735
rect 90726 7732 90732 7744
rect 90683 7704 90732 7732
rect 90683 7701 90695 7704
rect 90637 7695 90695 7701
rect 90726 7692 90732 7704
rect 90784 7692 90790 7744
rect 94225 7735 94283 7741
rect 94225 7701 94237 7735
rect 94271 7732 94283 7735
rect 95142 7732 95148 7744
rect 94271 7704 95148 7732
rect 94271 7701 94283 7704
rect 94225 7695 94283 7701
rect 95142 7692 95148 7704
rect 95200 7692 95206 7744
rect 1104 7642 95011 7664
rect 1104 7590 24386 7642
rect 24438 7590 24450 7642
rect 24502 7590 24514 7642
rect 24566 7590 24578 7642
rect 24630 7590 24642 7642
rect 24694 7590 47823 7642
rect 47875 7590 47887 7642
rect 47939 7590 47951 7642
rect 48003 7590 48015 7642
rect 48067 7590 48079 7642
rect 48131 7590 71260 7642
rect 71312 7590 71324 7642
rect 71376 7590 71388 7642
rect 71440 7590 71452 7642
rect 71504 7590 71516 7642
rect 71568 7590 94697 7642
rect 94749 7590 94761 7642
rect 94813 7590 94825 7642
rect 94877 7590 94889 7642
rect 94941 7590 94953 7642
rect 95005 7590 95011 7642
rect 1104 7568 95011 7590
rect 5718 7528 5724 7540
rect 1964 7500 5724 7528
rect 1964 7401 1992 7500
rect 2222 7460 2228 7472
rect 2183 7432 2228 7460
rect 2222 7420 2228 7432
rect 2280 7420 2286 7472
rect 4062 7460 4068 7472
rect 3450 7432 4068 7460
rect 4062 7420 4068 7432
rect 4120 7420 4126 7472
rect 4430 7460 4436 7472
rect 4391 7432 4436 7460
rect 4430 7420 4436 7432
rect 4488 7420 4494 7472
rect 4816 7460 4844 7500
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 5905 7531 5963 7537
rect 5905 7497 5917 7531
rect 5951 7528 5963 7531
rect 8202 7528 8208 7540
rect 5951 7500 8208 7528
rect 5951 7497 5963 7500
rect 5905 7491 5963 7497
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 18322 7528 18328 7540
rect 14476 7500 18184 7528
rect 18283 7500 18328 7528
rect 9582 7460 9588 7472
rect 4816 7432 4922 7460
rect 9495 7432 9588 7460
rect 9582 7420 9588 7432
rect 9640 7460 9646 7472
rect 12986 7460 12992 7472
rect 9640 7432 12992 7460
rect 9640 7420 9646 7432
rect 12986 7420 12992 7432
rect 13044 7460 13050 7472
rect 13722 7460 13728 7472
rect 13044 7432 13728 7460
rect 13044 7420 13050 7432
rect 13722 7420 13728 7432
rect 13780 7420 13786 7472
rect 14476 7469 14504 7500
rect 14461 7463 14519 7469
rect 14461 7429 14473 7463
rect 14507 7429 14519 7463
rect 14461 7423 14519 7429
rect 16298 7420 16304 7472
rect 16356 7460 16362 7472
rect 16853 7463 16911 7469
rect 16853 7460 16865 7463
rect 16356 7432 16865 7460
rect 16356 7420 16362 7432
rect 16853 7429 16865 7432
rect 16899 7429 16911 7463
rect 16853 7423 16911 7429
rect 17310 7420 17316 7472
rect 17368 7460 17374 7472
rect 17681 7463 17739 7469
rect 17681 7460 17693 7463
rect 17368 7432 17693 7460
rect 17368 7420 17374 7432
rect 17681 7429 17693 7432
rect 17727 7429 17739 7463
rect 18156 7460 18184 7500
rect 18322 7488 18328 7500
rect 18380 7488 18386 7540
rect 18690 7488 18696 7540
rect 18748 7528 18754 7540
rect 18969 7531 19027 7537
rect 18969 7528 18981 7531
rect 18748 7500 18981 7528
rect 18748 7488 18754 7500
rect 18969 7497 18981 7500
rect 19015 7497 19027 7531
rect 18969 7491 19027 7497
rect 21818 7488 21824 7540
rect 21876 7528 21882 7540
rect 24673 7531 24731 7537
rect 24673 7528 24685 7531
rect 21876 7500 24685 7528
rect 21876 7488 21882 7500
rect 24673 7497 24685 7500
rect 24719 7497 24731 7531
rect 27522 7528 27528 7540
rect 27483 7500 27528 7528
rect 24673 7491 24731 7497
rect 27522 7488 27528 7500
rect 27580 7488 27586 7540
rect 28442 7528 28448 7540
rect 28000 7500 28448 7528
rect 18874 7460 18880 7472
rect 18156 7432 18880 7460
rect 17681 7423 17739 7429
rect 18874 7420 18880 7432
rect 18932 7420 18938 7472
rect 20070 7460 20076 7472
rect 19076 7432 20076 7460
rect 1949 7395 2007 7401
rect 1949 7361 1961 7395
rect 1995 7361 2007 7395
rect 1949 7355 2007 7361
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7392 6699 7395
rect 6822 7392 6828 7404
rect 6687 7364 6828 7392
rect 6687 7361 6699 7364
rect 6641 7355 6699 7361
rect 3694 7324 3700 7336
rect 3655 7296 3700 7324
rect 3694 7284 3700 7296
rect 3752 7284 3758 7336
rect 3970 7284 3976 7336
rect 4028 7324 4034 7336
rect 4157 7327 4215 7333
rect 4157 7324 4169 7327
rect 4028 7296 4169 7324
rect 4028 7284 4034 7296
rect 4157 7293 4169 7296
rect 4203 7324 4215 7327
rect 6656 7324 6684 7355
rect 6822 7352 6828 7364
rect 6880 7392 6886 7404
rect 7193 7395 7251 7401
rect 7193 7392 7205 7395
rect 6880 7364 7205 7392
rect 6880 7352 6886 7364
rect 7193 7361 7205 7364
rect 7239 7392 7251 7395
rect 9490 7392 9496 7404
rect 7239 7364 9496 7392
rect 7239 7361 7251 7364
rect 7193 7355 7251 7361
rect 9490 7352 9496 7364
rect 9548 7352 9554 7404
rect 10042 7392 10048 7404
rect 9955 7364 10048 7392
rect 10042 7352 10048 7364
rect 10100 7392 10106 7404
rect 10686 7392 10692 7404
rect 10100 7364 10692 7392
rect 10100 7352 10106 7364
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 11977 7395 12035 7401
rect 11977 7392 11989 7395
rect 11072 7364 11989 7392
rect 4203 7296 6684 7324
rect 4203 7293 4215 7296
rect 4157 7287 4215 7293
rect 8294 7188 8300 7200
rect 8255 7160 8300 7188
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 10229 7191 10287 7197
rect 10229 7188 10241 7191
rect 9732 7160 10241 7188
rect 9732 7148 9738 7160
rect 10229 7157 10241 7160
rect 10275 7188 10287 7191
rect 10778 7188 10784 7200
rect 10275 7160 10784 7188
rect 10275 7157 10287 7160
rect 10229 7151 10287 7157
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 10962 7148 10968 7200
rect 11020 7188 11026 7200
rect 11072 7197 11100 7364
rect 11977 7361 11989 7364
rect 12023 7361 12035 7395
rect 18230 7392 18236 7404
rect 11977 7355 12035 7361
rect 13722 7284 13728 7336
rect 13780 7324 13786 7336
rect 14185 7327 14243 7333
rect 14185 7324 14197 7327
rect 13780 7296 14197 7324
rect 13780 7284 13786 7296
rect 14185 7293 14197 7296
rect 14231 7293 14243 7327
rect 14185 7287 14243 7293
rect 15580 7256 15608 7378
rect 18191 7364 18236 7392
rect 18230 7352 18236 7364
rect 18288 7352 18294 7404
rect 18417 7395 18475 7401
rect 18417 7361 18429 7395
rect 18463 7392 18475 7395
rect 18598 7392 18604 7404
rect 18463 7364 18604 7392
rect 18463 7361 18475 7364
rect 18417 7355 18475 7361
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 19076 7401 19104 7432
rect 20070 7420 20076 7432
rect 20128 7420 20134 7472
rect 20990 7420 20996 7472
rect 21048 7420 21054 7472
rect 22278 7460 22284 7472
rect 21192 7432 22284 7460
rect 19061 7395 19119 7401
rect 19061 7361 19073 7395
rect 19107 7361 19119 7395
rect 19061 7355 19119 7361
rect 19613 7395 19671 7401
rect 19613 7361 19625 7395
rect 19659 7392 19671 7395
rect 20254 7392 20260 7404
rect 19659 7364 20260 7392
rect 19659 7361 19671 7364
rect 19613 7355 19671 7361
rect 16209 7327 16267 7333
rect 16209 7293 16221 7327
rect 16255 7324 16267 7327
rect 19628 7324 19656 7355
rect 20254 7352 20260 7364
rect 20312 7352 20318 7404
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7392 20499 7395
rect 21192 7392 21220 7432
rect 22278 7420 22284 7432
rect 22336 7460 22342 7472
rect 26142 7460 26148 7472
rect 22336 7432 22600 7460
rect 26103 7432 26148 7460
rect 22336 7420 22342 7432
rect 20487 7364 21220 7392
rect 20487 7361 20499 7364
rect 20441 7355 20499 7361
rect 21266 7352 21272 7404
rect 21324 7392 21330 7404
rect 22097 7395 22155 7401
rect 22097 7392 22109 7395
rect 21324 7364 22109 7392
rect 21324 7352 21330 7364
rect 22097 7361 22109 7364
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 22462 7324 22468 7336
rect 16255 7296 19656 7324
rect 21100 7296 22468 7324
rect 16255 7293 16267 7296
rect 16209 7287 16267 7293
rect 21100 7256 21128 7296
rect 22462 7284 22468 7296
rect 22520 7284 22526 7336
rect 22572 7324 22600 7432
rect 26142 7420 26148 7432
rect 26200 7420 26206 7472
rect 26234 7420 26240 7472
rect 26292 7460 26298 7472
rect 28000 7469 28028 7500
rect 28442 7488 28448 7500
rect 28500 7488 28506 7540
rect 30742 7488 30748 7540
rect 30800 7528 30806 7540
rect 35437 7531 35495 7537
rect 35437 7528 35449 7531
rect 30800 7500 35449 7528
rect 30800 7488 30806 7500
rect 35437 7497 35449 7500
rect 35483 7497 35495 7531
rect 35437 7491 35495 7497
rect 36538 7488 36544 7540
rect 36596 7528 36602 7540
rect 39761 7531 39819 7537
rect 39761 7528 39773 7531
rect 36596 7500 39773 7528
rect 36596 7488 36602 7500
rect 39761 7497 39773 7500
rect 39807 7497 39819 7531
rect 39761 7491 39819 7497
rect 39850 7488 39856 7540
rect 39908 7528 39914 7540
rect 41598 7528 41604 7540
rect 39908 7500 41604 7528
rect 39908 7488 39914 7500
rect 41598 7488 41604 7500
rect 41656 7488 41662 7540
rect 42426 7488 42432 7540
rect 42484 7528 42490 7540
rect 42613 7531 42671 7537
rect 42613 7528 42625 7531
rect 42484 7500 42625 7528
rect 42484 7488 42490 7500
rect 42613 7497 42625 7500
rect 42659 7497 42671 7531
rect 42978 7528 42984 7540
rect 42939 7500 42984 7528
rect 42613 7491 42671 7497
rect 42978 7488 42984 7500
rect 43036 7488 43042 7540
rect 44177 7531 44235 7537
rect 44177 7497 44189 7531
rect 44223 7528 44235 7531
rect 44358 7528 44364 7540
rect 44223 7500 44364 7528
rect 44223 7497 44235 7500
rect 44177 7491 44235 7497
rect 44358 7488 44364 7500
rect 44416 7528 44422 7540
rect 44910 7528 44916 7540
rect 44416 7500 44916 7528
rect 44416 7488 44422 7500
rect 44910 7488 44916 7500
rect 44968 7488 44974 7540
rect 45462 7528 45468 7540
rect 45423 7500 45468 7528
rect 45462 7488 45468 7500
rect 45520 7488 45526 7540
rect 46566 7528 46572 7540
rect 46527 7500 46572 7528
rect 46566 7488 46572 7500
rect 46624 7488 46630 7540
rect 47213 7531 47271 7537
rect 47213 7497 47225 7531
rect 47259 7528 47271 7531
rect 47302 7528 47308 7540
rect 47259 7500 47308 7528
rect 47259 7497 47271 7500
rect 47213 7491 47271 7497
rect 47302 7488 47308 7500
rect 47360 7488 47366 7540
rect 49237 7531 49295 7537
rect 49237 7497 49249 7531
rect 49283 7528 49295 7531
rect 50338 7528 50344 7540
rect 49283 7500 50344 7528
rect 49283 7497 49295 7500
rect 49237 7491 49295 7497
rect 50338 7488 50344 7500
rect 50396 7488 50402 7540
rect 51350 7488 51356 7540
rect 51408 7528 51414 7540
rect 52181 7531 52239 7537
rect 52181 7528 52193 7531
rect 51408 7500 52193 7528
rect 51408 7488 51414 7500
rect 52181 7497 52193 7500
rect 52227 7497 52239 7531
rect 52181 7491 52239 7497
rect 52270 7488 52276 7540
rect 52328 7528 52334 7540
rect 57698 7528 57704 7540
rect 52328 7500 57704 7528
rect 52328 7488 52334 7500
rect 57698 7488 57704 7500
rect 57756 7488 57762 7540
rect 58618 7488 58624 7540
rect 58676 7528 58682 7540
rect 60550 7528 60556 7540
rect 58676 7500 59676 7528
rect 60511 7500 60556 7528
rect 58676 7488 58682 7500
rect 27985 7463 28043 7469
rect 26292 7432 27844 7460
rect 26292 7420 26298 7432
rect 23658 7392 23664 7404
rect 22770 7378 23664 7392
rect 22756 7364 23664 7378
rect 22756 7324 22784 7364
rect 23658 7352 23664 7364
rect 23716 7352 23722 7404
rect 25130 7392 25136 7404
rect 25070 7378 25136 7392
rect 25056 7364 25136 7378
rect 23106 7324 23112 7336
rect 22572 7296 22784 7324
rect 23067 7296 23112 7324
rect 23106 7284 23112 7296
rect 23164 7284 23170 7336
rect 23382 7284 23388 7336
rect 23440 7324 23446 7336
rect 25056 7324 25084 7364
rect 25130 7352 25136 7364
rect 25188 7352 25194 7404
rect 27706 7392 27712 7404
rect 27667 7364 27712 7392
rect 27706 7352 27712 7364
rect 27764 7352 27770 7404
rect 27816 7392 27844 7432
rect 27985 7429 27997 7463
rect 28031 7429 28043 7463
rect 27985 7423 28043 7429
rect 29638 7420 29644 7472
rect 29696 7460 29702 7472
rect 29917 7463 29975 7469
rect 29917 7460 29929 7463
rect 29696 7432 29929 7460
rect 29696 7420 29702 7432
rect 29917 7429 29929 7432
rect 29963 7429 29975 7463
rect 29917 7423 29975 7429
rect 31754 7420 31760 7472
rect 31812 7460 31818 7472
rect 32398 7460 32404 7472
rect 31812 7432 32404 7460
rect 31812 7420 31818 7432
rect 32398 7420 32404 7432
rect 32456 7420 32462 7472
rect 33134 7460 33140 7472
rect 33095 7432 33140 7460
rect 33134 7420 33140 7432
rect 33192 7420 33198 7472
rect 33594 7420 33600 7472
rect 33652 7420 33658 7472
rect 34885 7463 34943 7469
rect 34885 7429 34897 7463
rect 34931 7460 34943 7463
rect 41506 7460 41512 7472
rect 34931 7432 36400 7460
rect 34931 7429 34943 7432
rect 34885 7423 34943 7429
rect 35802 7392 35808 7404
rect 27816 7364 28842 7392
rect 35763 7364 35808 7392
rect 35802 7352 35808 7364
rect 35860 7352 35866 7404
rect 35894 7352 35900 7404
rect 35952 7352 35958 7404
rect 36372 7392 36400 7432
rect 36648 7432 41512 7460
rect 36648 7392 36676 7432
rect 41506 7420 41512 7432
rect 41564 7420 41570 7472
rect 42996 7460 43024 7488
rect 41616 7432 43024 7460
rect 36372 7364 36676 7392
rect 36722 7352 36728 7404
rect 36780 7392 36786 7404
rect 36817 7395 36875 7401
rect 36817 7392 36829 7395
rect 36780 7364 36829 7392
rect 36780 7352 36786 7364
rect 36817 7361 36829 7364
rect 36863 7361 36875 7395
rect 36817 7355 36875 7361
rect 26421 7327 26479 7333
rect 23440 7296 25084 7324
rect 25148 7296 26372 7324
rect 23440 7284 23446 7296
rect 25148 7256 25176 7296
rect 15580 7228 21128 7256
rect 21192 7228 25176 7256
rect 26344 7256 26372 7296
rect 26421 7293 26433 7327
rect 26467 7324 26479 7327
rect 26602 7324 26608 7336
rect 26467 7296 26608 7324
rect 26467 7293 26479 7296
rect 26421 7287 26479 7293
rect 26602 7284 26608 7296
rect 26660 7324 26666 7336
rect 27154 7324 27160 7336
rect 26660 7296 27160 7324
rect 26660 7284 26666 7296
rect 27154 7284 27160 7296
rect 27212 7284 27218 7336
rect 27893 7327 27951 7333
rect 27893 7293 27905 7327
rect 27939 7324 27951 7327
rect 28718 7324 28724 7336
rect 27939 7296 28724 7324
rect 27939 7293 27951 7296
rect 27893 7287 27951 7293
rect 28718 7284 28724 7296
rect 28776 7284 28782 7336
rect 30190 7324 30196 7336
rect 30151 7296 30196 7324
rect 30190 7284 30196 7296
rect 30248 7284 30254 7336
rect 32858 7324 32864 7336
rect 32819 7296 32864 7324
rect 32858 7284 32864 7296
rect 32916 7284 32922 7336
rect 35713 7327 35771 7333
rect 32968 7296 35664 7324
rect 28626 7256 28632 7268
rect 26344 7228 28632 7256
rect 11057 7191 11115 7197
rect 11057 7188 11069 7191
rect 11020 7160 11069 7188
rect 11020 7148 11026 7160
rect 11057 7157 11069 7160
rect 11103 7157 11115 7191
rect 11057 7151 11115 7157
rect 19334 7148 19340 7200
rect 19392 7188 19398 7200
rect 21192 7188 21220 7228
rect 28626 7216 28632 7228
rect 28684 7216 28690 7268
rect 31662 7216 31668 7268
rect 31720 7256 31726 7268
rect 32968 7256 32996 7296
rect 31720 7228 32996 7256
rect 35636 7256 35664 7296
rect 35713 7293 35725 7327
rect 35759 7324 35771 7327
rect 35912 7324 35940 7352
rect 36630 7324 36636 7336
rect 35759 7296 35940 7324
rect 36464 7296 36636 7324
rect 35759 7293 35771 7296
rect 35713 7287 35771 7293
rect 36464 7256 36492 7296
rect 36630 7284 36636 7296
rect 36688 7284 36694 7336
rect 36832 7324 36860 7355
rect 38102 7352 38108 7404
rect 38160 7392 38166 7404
rect 38197 7395 38255 7401
rect 38197 7392 38209 7395
rect 38160 7364 38209 7392
rect 38160 7352 38166 7364
rect 38197 7361 38209 7364
rect 38243 7392 38255 7395
rect 38838 7392 38844 7404
rect 38243 7364 38844 7392
rect 38243 7361 38255 7364
rect 38197 7355 38255 7361
rect 38838 7352 38844 7364
rect 38896 7352 38902 7404
rect 39117 7395 39175 7401
rect 39117 7361 39129 7395
rect 39163 7392 39175 7395
rect 40126 7392 40132 7404
rect 39163 7364 39988 7392
rect 40087 7364 40132 7392
rect 39163 7361 39175 7364
rect 39117 7355 39175 7361
rect 39022 7324 39028 7336
rect 36832 7296 38884 7324
rect 38983 7296 39028 7324
rect 35636 7228 36492 7256
rect 31720 7216 31726 7228
rect 36538 7216 36544 7268
rect 36596 7256 36602 7268
rect 38749 7259 38807 7265
rect 38749 7256 38761 7259
rect 36596 7228 38761 7256
rect 36596 7216 36602 7228
rect 38749 7225 38761 7228
rect 38795 7225 38807 7259
rect 38856 7256 38884 7296
rect 39022 7284 39028 7296
rect 39080 7284 39086 7336
rect 39390 7256 39396 7268
rect 38856 7228 39396 7256
rect 38749 7219 38807 7225
rect 39390 7216 39396 7228
rect 39448 7216 39454 7268
rect 39960 7256 39988 7364
rect 40126 7352 40132 7364
rect 40184 7352 40190 7404
rect 41049 7395 41107 7401
rect 41049 7392 41061 7395
rect 40696 7364 41061 7392
rect 40221 7327 40279 7333
rect 40221 7293 40233 7327
rect 40267 7324 40279 7327
rect 40586 7324 40592 7336
rect 40267 7296 40592 7324
rect 40267 7293 40279 7296
rect 40221 7287 40279 7293
rect 40586 7284 40592 7296
rect 40644 7284 40650 7336
rect 40126 7256 40132 7268
rect 39960 7228 40132 7256
rect 40126 7216 40132 7228
rect 40184 7256 40190 7268
rect 40696 7256 40724 7364
rect 41049 7361 41061 7364
rect 41095 7392 41107 7395
rect 41616 7392 41644 7432
rect 43070 7420 43076 7472
rect 43128 7420 43134 7472
rect 44082 7420 44088 7472
rect 44140 7460 44146 7472
rect 49694 7460 49700 7472
rect 44140 7432 49700 7460
rect 44140 7420 44146 7432
rect 49694 7420 49700 7432
rect 49752 7420 49758 7472
rect 49973 7463 50031 7469
rect 49973 7429 49985 7463
rect 50019 7460 50031 7463
rect 52917 7463 52975 7469
rect 52917 7460 52929 7463
rect 50019 7432 52929 7460
rect 50019 7429 50031 7432
rect 49973 7423 50031 7429
rect 52917 7429 52929 7432
rect 52963 7429 52975 7463
rect 52917 7423 52975 7429
rect 55858 7420 55864 7472
rect 55916 7420 55922 7472
rect 57517 7463 57575 7469
rect 57517 7429 57529 7463
rect 57563 7460 57575 7463
rect 58345 7463 58403 7469
rect 58345 7460 58357 7463
rect 57563 7432 58357 7460
rect 57563 7429 57575 7432
rect 57517 7423 57575 7429
rect 58345 7429 58357 7432
rect 58391 7429 58403 7463
rect 58345 7423 58403 7429
rect 59354 7420 59360 7472
rect 59412 7420 59418 7472
rect 59648 7460 59676 7500
rect 60550 7488 60556 7500
rect 60608 7488 60614 7540
rect 60826 7528 60832 7540
rect 60739 7500 60832 7528
rect 60826 7488 60832 7500
rect 60884 7528 60890 7540
rect 61562 7528 61568 7540
rect 60884 7500 61568 7528
rect 60884 7488 60890 7500
rect 61562 7488 61568 7500
rect 61620 7488 61626 7540
rect 63034 7488 63040 7540
rect 63092 7528 63098 7540
rect 64785 7531 64843 7537
rect 64785 7528 64797 7531
rect 63092 7500 64797 7528
rect 63092 7488 63098 7500
rect 64785 7497 64797 7500
rect 64831 7528 64843 7531
rect 66809 7531 66867 7537
rect 64831 7500 65564 7528
rect 64831 7497 64843 7500
rect 64785 7491 64843 7497
rect 62577 7463 62635 7469
rect 62577 7460 62589 7463
rect 59648 7432 62589 7460
rect 62577 7429 62589 7432
rect 62623 7429 62635 7463
rect 63494 7460 63500 7472
rect 63455 7432 63500 7460
rect 62577 7423 62635 7429
rect 63494 7420 63500 7432
rect 63552 7420 63558 7472
rect 65536 7460 65564 7500
rect 66809 7497 66821 7531
rect 66855 7528 66867 7531
rect 67542 7528 67548 7540
rect 66855 7500 67548 7528
rect 66855 7497 66867 7500
rect 66809 7491 66867 7497
rect 67542 7488 67548 7500
rect 67600 7488 67606 7540
rect 67634 7488 67640 7540
rect 67692 7528 67698 7540
rect 67821 7531 67879 7537
rect 67821 7528 67833 7531
rect 67692 7500 67833 7528
rect 67692 7488 67698 7500
rect 67821 7497 67833 7500
rect 67867 7497 67879 7531
rect 67821 7491 67879 7497
rect 68002 7488 68008 7540
rect 68060 7528 68066 7540
rect 74350 7528 74356 7540
rect 68060 7500 69704 7528
rect 68060 7488 68066 7500
rect 69676 7460 69704 7500
rect 71424 7500 74356 7528
rect 70489 7463 70547 7469
rect 70489 7460 70501 7463
rect 63880 7432 65472 7460
rect 41095 7364 41644 7392
rect 42061 7395 42119 7401
rect 41095 7361 41107 7364
rect 41049 7355 41107 7361
rect 42061 7361 42073 7395
rect 42107 7392 42119 7395
rect 42426 7392 42432 7404
rect 42107 7364 42432 7392
rect 42107 7361 42119 7364
rect 42061 7355 42119 7361
rect 42426 7352 42432 7364
rect 42484 7352 42490 7404
rect 42797 7395 42855 7401
rect 42797 7361 42809 7395
rect 42843 7361 42855 7395
rect 42797 7355 42855 7361
rect 42889 7395 42947 7401
rect 42889 7361 42901 7395
rect 42935 7392 42947 7395
rect 43088 7392 43116 7420
rect 63880 7404 63908 7432
rect 42935 7364 43116 7392
rect 42935 7361 42947 7364
rect 42889 7355 42947 7361
rect 40862 7324 40868 7336
rect 40823 7296 40868 7324
rect 40862 7284 40868 7296
rect 40920 7284 40926 7336
rect 40954 7284 40960 7336
rect 41012 7324 41018 7336
rect 41141 7327 41199 7333
rect 41012 7296 41057 7324
rect 41012 7284 41018 7296
rect 41141 7293 41153 7327
rect 41187 7324 41199 7327
rect 41230 7324 41236 7336
rect 41187 7296 41236 7324
rect 41187 7293 41199 7296
rect 41141 7287 41199 7293
rect 41230 7284 41236 7296
rect 41288 7284 41294 7336
rect 41598 7284 41604 7336
rect 41656 7316 41662 7336
rect 41781 7327 41839 7333
rect 41781 7316 41793 7327
rect 41656 7293 41793 7316
rect 41827 7293 41839 7327
rect 42812 7324 42840 7355
rect 46566 7352 46572 7404
rect 46624 7392 46630 7404
rect 49142 7392 49148 7404
rect 46624 7364 49148 7392
rect 46624 7352 46630 7364
rect 49142 7352 49148 7364
rect 49200 7352 49206 7404
rect 49510 7352 49516 7404
rect 49568 7392 49574 7404
rect 49789 7395 49847 7401
rect 49789 7392 49801 7395
rect 49568 7364 49801 7392
rect 49568 7352 49574 7364
rect 49789 7361 49801 7364
rect 49835 7361 49847 7395
rect 52086 7392 52092 7404
rect 49789 7355 49847 7361
rect 51552 7364 52092 7392
rect 43070 7324 43076 7336
rect 42812 7296 43076 7324
rect 41656 7288 41839 7293
rect 41656 7284 41662 7288
rect 41781 7287 41839 7288
rect 43070 7284 43076 7296
rect 43128 7284 43134 7336
rect 43438 7284 43444 7336
rect 43496 7324 43502 7336
rect 46109 7327 46167 7333
rect 46109 7324 46121 7327
rect 43496 7296 46121 7324
rect 43496 7284 43502 7296
rect 46109 7293 46121 7296
rect 46155 7324 46167 7327
rect 47302 7324 47308 7336
rect 46155 7296 47308 7324
rect 46155 7293 46167 7296
rect 46109 7287 46167 7293
rect 47302 7284 47308 7296
rect 47360 7284 47366 7336
rect 49326 7284 49332 7336
rect 49384 7324 49390 7336
rect 51552 7324 51580 7364
rect 52086 7352 52092 7364
rect 52144 7352 52150 7404
rect 52273 7395 52331 7401
rect 52273 7361 52285 7395
rect 52319 7361 52331 7395
rect 53558 7392 53564 7404
rect 53519 7364 53564 7392
rect 52273 7355 52331 7361
rect 49384 7296 51580 7324
rect 49384 7284 49390 7296
rect 51626 7284 51632 7336
rect 51684 7324 51690 7336
rect 52178 7324 52184 7336
rect 51684 7296 52184 7324
rect 51684 7284 51690 7296
rect 52178 7284 52184 7296
rect 52236 7284 52242 7336
rect 41874 7256 41880 7268
rect 40184 7228 40724 7256
rect 41835 7228 41880 7256
rect 40184 7216 40190 7228
rect 41874 7216 41880 7228
rect 41932 7216 41938 7268
rect 42058 7216 42064 7268
rect 42116 7256 42122 7268
rect 43165 7259 43223 7265
rect 43165 7256 43177 7259
rect 42116 7228 43177 7256
rect 42116 7216 42122 7228
rect 43165 7225 43177 7228
rect 43211 7256 43223 7259
rect 45554 7256 45560 7268
rect 43211 7228 45560 7256
rect 43211 7225 43223 7228
rect 43165 7219 43223 7225
rect 45554 7216 45560 7228
rect 45612 7216 45618 7268
rect 47857 7259 47915 7265
rect 47857 7256 47869 7259
rect 45664 7228 47869 7256
rect 19392 7160 21220 7188
rect 19392 7148 19398 7160
rect 22462 7148 22468 7200
rect 22520 7188 22526 7200
rect 23382 7188 23388 7200
rect 22520 7160 23388 7188
rect 22520 7148 22526 7160
rect 23382 7148 23388 7160
rect 23440 7148 23446 7200
rect 23658 7188 23664 7200
rect 23619 7160 23664 7188
rect 23658 7148 23664 7160
rect 23716 7148 23722 7200
rect 24210 7188 24216 7200
rect 24171 7160 24216 7188
rect 24210 7148 24216 7160
rect 24268 7148 24274 7200
rect 25130 7148 25136 7200
rect 25188 7188 25194 7200
rect 27246 7188 27252 7200
rect 25188 7160 27252 7188
rect 25188 7148 25194 7160
rect 27246 7148 27252 7160
rect 27304 7148 27310 7200
rect 27985 7191 28043 7197
rect 27985 7157 27997 7191
rect 28031 7188 28043 7191
rect 28074 7188 28080 7200
rect 28031 7160 28080 7188
rect 28031 7157 28043 7160
rect 27985 7151 28043 7157
rect 28074 7148 28080 7160
rect 28132 7188 28138 7200
rect 28902 7188 28908 7200
rect 28132 7160 28908 7188
rect 28132 7148 28138 7160
rect 28902 7148 28908 7160
rect 28960 7188 28966 7200
rect 30653 7191 30711 7197
rect 30653 7188 30665 7191
rect 28960 7160 30665 7188
rect 28960 7148 28966 7160
rect 30653 7157 30665 7160
rect 30699 7188 30711 7191
rect 32766 7188 32772 7200
rect 30699 7160 32772 7188
rect 30699 7157 30711 7160
rect 30653 7151 30711 7157
rect 32766 7148 32772 7160
rect 32824 7188 32830 7200
rect 33778 7188 33784 7200
rect 32824 7160 33784 7188
rect 32824 7148 32830 7160
rect 33778 7148 33784 7160
rect 33836 7148 33842 7200
rect 33870 7148 33876 7200
rect 33928 7188 33934 7200
rect 35802 7188 35808 7200
rect 33928 7160 35808 7188
rect 33928 7148 33934 7160
rect 35802 7148 35808 7160
rect 35860 7188 35866 7200
rect 37642 7188 37648 7200
rect 35860 7160 37648 7188
rect 35860 7148 35866 7160
rect 37642 7148 37648 7160
rect 37700 7148 37706 7200
rect 37737 7191 37795 7197
rect 37737 7157 37749 7191
rect 37783 7188 37795 7191
rect 37826 7188 37832 7200
rect 37783 7160 37832 7188
rect 37783 7157 37795 7160
rect 37737 7151 37795 7157
rect 37826 7148 37832 7160
rect 37884 7188 37890 7200
rect 38286 7188 38292 7200
rect 37884 7160 38292 7188
rect 37884 7148 37890 7160
rect 38286 7148 38292 7160
rect 38344 7148 38350 7200
rect 38838 7148 38844 7200
rect 38896 7188 38902 7200
rect 39850 7188 39856 7200
rect 38896 7160 39856 7188
rect 38896 7148 38902 7160
rect 39850 7148 39856 7160
rect 39908 7148 39914 7200
rect 41138 7148 41144 7200
rect 41196 7188 41202 7200
rect 41325 7191 41383 7197
rect 41325 7188 41337 7191
rect 41196 7160 41337 7188
rect 41196 7148 41202 7160
rect 41325 7157 41337 7160
rect 41371 7157 41383 7191
rect 41966 7188 41972 7200
rect 41927 7160 41972 7188
rect 41325 7151 41383 7157
rect 41966 7148 41972 7160
rect 42024 7148 42030 7200
rect 44910 7188 44916 7200
rect 44871 7160 44916 7188
rect 44910 7148 44916 7160
rect 44968 7148 44974 7200
rect 45462 7148 45468 7200
rect 45520 7188 45526 7200
rect 45664 7188 45692 7228
rect 47857 7225 47869 7228
rect 47903 7256 47915 7259
rect 48222 7256 48228 7268
rect 47903 7228 48228 7256
rect 47903 7225 47915 7228
rect 47857 7219 47915 7225
rect 48222 7216 48228 7228
rect 48280 7216 48286 7268
rect 48501 7259 48559 7265
rect 48501 7225 48513 7259
rect 48547 7256 48559 7259
rect 48682 7256 48688 7268
rect 48547 7228 48688 7256
rect 48547 7225 48559 7228
rect 48501 7219 48559 7225
rect 45520 7160 45692 7188
rect 45520 7148 45526 7160
rect 45738 7148 45744 7200
rect 45796 7188 45802 7200
rect 48516 7188 48544 7219
rect 48682 7216 48688 7228
rect 48740 7256 48746 7268
rect 51810 7256 51816 7268
rect 48740 7228 51816 7256
rect 48740 7216 48746 7228
rect 51810 7216 51816 7228
rect 51868 7256 51874 7268
rect 52086 7256 52092 7268
rect 51868 7228 52092 7256
rect 51868 7216 51874 7228
rect 52086 7216 52092 7228
rect 52144 7256 52150 7268
rect 52288 7256 52316 7355
rect 53558 7352 53564 7364
rect 53616 7352 53622 7404
rect 57238 7392 57244 7404
rect 57199 7364 57244 7392
rect 57238 7352 57244 7364
rect 57296 7352 57302 7404
rect 58066 7392 58072 7404
rect 58027 7364 58072 7392
rect 58066 7352 58072 7364
rect 58124 7352 58130 7404
rect 60737 7395 60795 7401
rect 60737 7392 60749 7395
rect 60568 7364 60749 7392
rect 53745 7327 53803 7333
rect 53745 7293 53757 7327
rect 53791 7324 53803 7327
rect 53791 7296 53880 7324
rect 53791 7293 53803 7296
rect 53745 7287 53803 7293
rect 52144 7228 52316 7256
rect 52144 7216 52150 7228
rect 45796 7160 48544 7188
rect 45796 7148 45802 7160
rect 53650 7148 53656 7200
rect 53708 7188 53714 7200
rect 53852 7188 53880 7296
rect 54202 7284 54208 7336
rect 54260 7324 54266 7336
rect 54573 7327 54631 7333
rect 54573 7324 54585 7327
rect 54260 7296 54585 7324
rect 54260 7284 54266 7296
rect 54573 7293 54585 7296
rect 54619 7293 54631 7327
rect 54846 7324 54852 7336
rect 54807 7296 54852 7324
rect 54573 7287 54631 7293
rect 54846 7284 54852 7296
rect 54904 7284 54910 7336
rect 54938 7284 54944 7336
rect 54996 7324 55002 7336
rect 60458 7324 60464 7336
rect 54996 7296 60464 7324
rect 54996 7284 55002 7296
rect 60458 7284 60464 7296
rect 60516 7284 60522 7336
rect 55950 7216 55956 7268
rect 56008 7256 56014 7268
rect 56008 7228 56456 7256
rect 56008 7216 56014 7228
rect 56428 7200 56456 7228
rect 59354 7216 59360 7268
rect 59412 7256 59418 7268
rect 60568 7256 60596 7364
rect 60737 7361 60749 7364
rect 60783 7361 60795 7395
rect 60737 7355 60795 7361
rect 60921 7395 60979 7401
rect 60921 7361 60933 7395
rect 60967 7392 60979 7395
rect 61930 7392 61936 7404
rect 60967 7364 61936 7392
rect 60967 7361 60979 7364
rect 60921 7355 60979 7361
rect 61930 7352 61936 7364
rect 61988 7352 61994 7404
rect 62666 7392 62672 7404
rect 62627 7364 62672 7392
rect 62666 7352 62672 7364
rect 62724 7352 62730 7404
rect 63862 7392 63868 7404
rect 63823 7364 63868 7392
rect 63862 7352 63868 7364
rect 63920 7352 63926 7404
rect 64325 7395 64383 7401
rect 64325 7361 64337 7395
rect 64371 7392 64383 7395
rect 64506 7392 64512 7404
rect 64371 7364 64512 7392
rect 64371 7361 64383 7364
rect 64325 7355 64383 7361
rect 64506 7352 64512 7364
rect 64564 7352 64570 7404
rect 64601 7395 64659 7401
rect 64601 7361 64613 7395
rect 64647 7392 64659 7395
rect 64690 7392 64696 7404
rect 64647 7364 64696 7392
rect 64647 7361 64659 7364
rect 64601 7355 64659 7361
rect 64690 7352 64696 7364
rect 64748 7352 64754 7404
rect 61562 7324 61568 7336
rect 61475 7296 61568 7324
rect 61562 7284 61568 7296
rect 61620 7324 61626 7336
rect 61620 7296 62988 7324
rect 61620 7284 61626 7296
rect 60918 7256 60924 7268
rect 59412 7228 60924 7256
rect 59412 7216 59418 7228
rect 60918 7216 60924 7228
rect 60976 7216 60982 7268
rect 61102 7256 61108 7268
rect 61063 7228 61108 7256
rect 61102 7216 61108 7228
rect 61160 7216 61166 7268
rect 61933 7259 61991 7265
rect 61933 7225 61945 7259
rect 61979 7256 61991 7259
rect 62114 7256 62120 7268
rect 61979 7228 62120 7256
rect 61979 7225 61991 7228
rect 61933 7219 61991 7225
rect 62114 7216 62120 7228
rect 62172 7216 62178 7268
rect 62960 7256 62988 7296
rect 64138 7284 64144 7336
rect 64196 7324 64202 7336
rect 64417 7327 64475 7333
rect 64417 7324 64429 7327
rect 64196 7296 64429 7324
rect 64196 7284 64202 7296
rect 64417 7293 64429 7296
rect 64463 7324 64475 7327
rect 65334 7324 65340 7336
rect 64463 7296 65340 7324
rect 64463 7293 64475 7296
rect 64417 7287 64475 7293
rect 65334 7284 65340 7296
rect 65392 7284 65398 7336
rect 65444 7324 65472 7432
rect 65536 7432 66484 7460
rect 69676 7432 70501 7460
rect 65536 7401 65564 7432
rect 65521 7395 65579 7401
rect 65521 7361 65533 7395
rect 65567 7361 65579 7395
rect 65521 7355 65579 7361
rect 65610 7352 65616 7404
rect 65668 7392 65674 7404
rect 65797 7395 65855 7401
rect 65668 7364 65713 7392
rect 65668 7352 65674 7364
rect 65797 7361 65809 7395
rect 65843 7392 65855 7395
rect 66346 7392 66352 7404
rect 65843 7364 66352 7392
rect 65843 7361 65855 7364
rect 65797 7355 65855 7361
rect 65812 7324 65840 7355
rect 66346 7352 66352 7364
rect 66404 7352 66410 7404
rect 66456 7401 66484 7432
rect 70489 7429 70501 7432
rect 70535 7460 70547 7463
rect 71424 7460 71452 7500
rect 74350 7488 74356 7500
rect 74408 7488 74414 7540
rect 74810 7528 74816 7540
rect 74460 7500 74816 7528
rect 70535 7432 71452 7460
rect 70535 7429 70547 7432
rect 70489 7423 70547 7429
rect 71958 7420 71964 7472
rect 72016 7420 72022 7472
rect 72418 7420 72424 7472
rect 72476 7460 72482 7472
rect 72476 7432 73016 7460
rect 72476 7420 72482 7432
rect 66441 7395 66499 7401
rect 66441 7361 66453 7395
rect 66487 7361 66499 7395
rect 66441 7355 66499 7361
rect 66625 7395 66683 7401
rect 66625 7361 66637 7395
rect 66671 7392 66683 7395
rect 66714 7392 66720 7404
rect 66671 7364 66720 7392
rect 66671 7361 66683 7364
rect 66625 7355 66683 7361
rect 66714 7352 66720 7364
rect 66772 7352 66778 7404
rect 67450 7352 67456 7404
rect 67508 7401 67514 7404
rect 67508 7395 67557 7401
rect 67508 7361 67511 7395
rect 67545 7361 67557 7395
rect 67508 7355 67557 7361
rect 67508 7352 67514 7355
rect 68094 7352 68100 7404
rect 68152 7392 68158 7404
rect 68741 7395 68799 7401
rect 68741 7392 68753 7395
rect 68152 7364 68753 7392
rect 68152 7352 68158 7364
rect 68741 7361 68753 7364
rect 68787 7361 68799 7395
rect 69566 7392 69572 7404
rect 69479 7364 69572 7392
rect 68741 7355 68799 7361
rect 69566 7352 69572 7364
rect 69624 7352 69630 7404
rect 72988 7401 73016 7432
rect 72973 7395 73031 7401
rect 72973 7361 72985 7395
rect 73019 7392 73031 7395
rect 74460 7392 74488 7500
rect 74810 7488 74816 7500
rect 74868 7488 74874 7540
rect 75089 7531 75147 7537
rect 75089 7497 75101 7531
rect 75135 7528 75147 7531
rect 76098 7528 76104 7540
rect 75135 7500 76104 7528
rect 75135 7497 75147 7500
rect 75089 7491 75147 7497
rect 76098 7488 76104 7500
rect 76156 7488 76162 7540
rect 76469 7531 76527 7537
rect 76469 7497 76481 7531
rect 76515 7497 76527 7531
rect 76469 7491 76527 7497
rect 76374 7460 76380 7472
rect 74736 7432 76380 7460
rect 74736 7401 74764 7432
rect 76374 7420 76380 7432
rect 76432 7420 76438 7472
rect 73019 7364 74488 7392
rect 74721 7395 74779 7401
rect 73019 7361 73031 7364
rect 72973 7355 73031 7361
rect 74721 7361 74733 7395
rect 74767 7361 74779 7395
rect 76006 7392 76012 7404
rect 75967 7364 76012 7392
rect 74721 7355 74779 7361
rect 76006 7352 76012 7364
rect 76064 7352 76070 7404
rect 76282 7392 76288 7404
rect 76243 7364 76288 7392
rect 76282 7352 76288 7364
rect 76340 7352 76346 7404
rect 76484 7392 76512 7491
rect 76650 7488 76656 7540
rect 76708 7528 76714 7540
rect 76929 7531 76987 7537
rect 76929 7528 76941 7531
rect 76708 7500 76941 7528
rect 76708 7488 76714 7500
rect 76929 7497 76941 7500
rect 76975 7497 76987 7531
rect 78122 7528 78128 7540
rect 78083 7500 78128 7528
rect 76929 7491 76987 7497
rect 78122 7488 78128 7500
rect 78180 7488 78186 7540
rect 78674 7488 78680 7540
rect 78732 7528 78738 7540
rect 78732 7500 80560 7528
rect 78732 7488 78738 7500
rect 79704 7469 79732 7500
rect 77757 7463 77815 7469
rect 77757 7429 77769 7463
rect 77803 7460 77815 7463
rect 78769 7463 78827 7469
rect 78769 7460 78781 7463
rect 77803 7432 78781 7460
rect 77803 7429 77815 7432
rect 77757 7423 77815 7429
rect 78769 7429 78781 7432
rect 78815 7429 78827 7463
rect 78769 7423 78827 7429
rect 79689 7463 79747 7469
rect 79689 7429 79701 7463
rect 79735 7429 79747 7463
rect 79689 7423 79747 7429
rect 79919 7429 79977 7435
rect 79919 7426 79931 7429
rect 77662 7392 77668 7404
rect 76484 7364 77668 7392
rect 77662 7352 77668 7364
rect 77720 7352 77726 7404
rect 77938 7392 77944 7404
rect 77899 7364 77944 7392
rect 77938 7352 77944 7364
rect 77996 7352 78002 7404
rect 78674 7392 78680 7404
rect 78635 7364 78680 7392
rect 78674 7352 78680 7364
rect 78732 7352 78738 7404
rect 78858 7392 78864 7404
rect 78819 7364 78864 7392
rect 78858 7352 78864 7364
rect 78916 7392 78922 7404
rect 79904 7395 79931 7426
rect 79965 7395 79977 7429
rect 79904 7392 79977 7395
rect 80330 7392 80336 7404
rect 78916 7390 79640 7392
rect 79704 7390 80336 7392
rect 78916 7364 80336 7390
rect 78916 7352 78922 7364
rect 79612 7362 79732 7364
rect 80330 7352 80336 7364
rect 80388 7352 80394 7404
rect 65444 7296 65840 7324
rect 67358 7284 67364 7336
rect 67416 7324 67422 7336
rect 68646 7324 68652 7336
rect 67416 7296 67461 7324
rect 68607 7296 68652 7324
rect 67416 7284 67422 7296
rect 68646 7284 68652 7296
rect 68704 7284 68710 7336
rect 68830 7284 68836 7336
rect 68888 7324 68894 7336
rect 69477 7327 69535 7333
rect 69477 7324 69489 7327
rect 68888 7296 69489 7324
rect 68888 7284 68894 7296
rect 69477 7293 69489 7296
rect 69523 7293 69535 7327
rect 69477 7287 69535 7293
rect 65981 7259 66039 7265
rect 62960 7228 64644 7256
rect 56321 7191 56379 7197
rect 56321 7188 56333 7191
rect 53708 7160 56333 7188
rect 53708 7148 53714 7160
rect 56321 7157 56333 7160
rect 56367 7157 56379 7191
rect 56321 7151 56379 7157
rect 56410 7148 56416 7200
rect 56468 7188 56474 7200
rect 59817 7191 59875 7197
rect 59817 7188 59829 7191
rect 56468 7160 59829 7188
rect 56468 7148 56474 7160
rect 59817 7157 59829 7160
rect 59863 7157 59875 7191
rect 59817 7151 59875 7157
rect 62025 7191 62083 7197
rect 62025 7157 62037 7191
rect 62071 7188 62083 7191
rect 62482 7188 62488 7200
rect 62071 7160 62488 7188
rect 62071 7157 62083 7160
rect 62025 7151 62083 7157
rect 62482 7148 62488 7160
rect 62540 7148 62546 7200
rect 64616 7197 64644 7228
rect 65981 7225 65993 7259
rect 66027 7256 66039 7259
rect 67082 7256 67088 7268
rect 66027 7228 67088 7256
rect 66027 7225 66039 7228
rect 65981 7219 66039 7225
rect 67082 7216 67088 7228
rect 67140 7216 67146 7268
rect 64601 7191 64659 7197
rect 64601 7157 64613 7191
rect 64647 7188 64659 7191
rect 65150 7188 65156 7200
rect 64647 7160 65156 7188
rect 64647 7157 64659 7160
rect 64601 7151 64659 7157
rect 65150 7148 65156 7160
rect 65208 7148 65214 7200
rect 66622 7188 66628 7200
rect 66583 7160 66628 7188
rect 66622 7148 66628 7160
rect 66680 7148 66686 7200
rect 67266 7148 67272 7200
rect 67324 7188 67330 7200
rect 68278 7188 68284 7200
rect 67324 7160 68284 7188
rect 67324 7148 67330 7160
rect 68278 7148 68284 7160
rect 68336 7148 68342 7200
rect 68462 7188 68468 7200
rect 68423 7160 68468 7188
rect 68462 7148 68468 7160
rect 68520 7148 68526 7200
rect 69584 7188 69612 7352
rect 72697 7327 72755 7333
rect 72697 7324 72709 7327
rect 69952 7296 72709 7324
rect 69952 7265 69980 7296
rect 72697 7293 72709 7296
rect 72743 7293 72755 7327
rect 73522 7324 73528 7336
rect 73483 7296 73528 7324
rect 72697 7287 72755 7293
rect 73522 7284 73528 7296
rect 73580 7284 73586 7336
rect 74626 7324 74632 7336
rect 74587 7296 74632 7324
rect 74626 7284 74632 7296
rect 74684 7284 74690 7336
rect 76101 7327 76159 7333
rect 76101 7293 76113 7327
rect 76147 7324 76159 7327
rect 78692 7324 78720 7352
rect 80532 7333 80560 7500
rect 82630 7488 82636 7540
rect 82688 7528 82694 7540
rect 83274 7528 83280 7540
rect 82688 7500 83280 7528
rect 82688 7488 82694 7500
rect 83274 7488 83280 7500
rect 83332 7528 83338 7540
rect 85301 7531 85359 7537
rect 83332 7500 84608 7528
rect 83332 7488 83338 7500
rect 80698 7460 80704 7472
rect 80659 7432 80704 7460
rect 80698 7420 80704 7432
rect 80756 7420 80762 7472
rect 81342 7420 81348 7472
rect 81400 7460 81406 7472
rect 83185 7463 83243 7469
rect 81400 7432 83044 7460
rect 81400 7420 81406 7432
rect 83016 7401 83044 7432
rect 83185 7429 83197 7463
rect 83231 7460 83243 7463
rect 83231 7432 84516 7460
rect 83231 7429 83243 7432
rect 83185 7423 83243 7429
rect 84488 7404 84516 7432
rect 83001 7395 83059 7401
rect 83001 7361 83013 7395
rect 83047 7361 83059 7395
rect 83001 7355 83059 7361
rect 83274 7352 83280 7404
rect 83332 7392 83338 7404
rect 84197 7395 84255 7401
rect 83332 7364 83377 7392
rect 83332 7352 83338 7364
rect 84197 7361 84209 7395
rect 84243 7361 84255 7395
rect 84197 7355 84255 7361
rect 84289 7395 84347 7401
rect 84289 7361 84301 7395
rect 84335 7361 84347 7395
rect 84470 7392 84476 7404
rect 84383 7364 84476 7392
rect 84289 7355 84347 7361
rect 76147 7296 78720 7324
rect 80517 7327 80575 7333
rect 76147 7293 76159 7296
rect 76101 7287 76159 7293
rect 80517 7293 80529 7327
rect 80563 7324 80575 7327
rect 81618 7324 81624 7336
rect 80563 7296 81624 7324
rect 80563 7293 80575 7296
rect 80517 7287 80575 7293
rect 69937 7259 69995 7265
rect 69937 7225 69949 7259
rect 69983 7225 69995 7259
rect 69937 7219 69995 7225
rect 74534 7216 74540 7268
rect 74592 7256 74598 7268
rect 76116 7256 76144 7287
rect 81618 7284 81624 7296
rect 81676 7284 81682 7336
rect 81710 7284 81716 7336
rect 81768 7324 81774 7336
rect 81768 7296 81813 7324
rect 81768 7284 81774 7296
rect 84212 7268 84240 7355
rect 84194 7256 84200 7268
rect 74592 7228 76144 7256
rect 76208 7228 84200 7256
rect 74592 7216 74598 7228
rect 71225 7191 71283 7197
rect 71225 7188 71237 7191
rect 69584 7160 71237 7188
rect 71225 7157 71237 7160
rect 71271 7157 71283 7191
rect 71225 7151 71283 7157
rect 71958 7148 71964 7200
rect 72016 7188 72022 7200
rect 76208 7188 76236 7228
rect 84194 7216 84200 7228
rect 84252 7216 84258 7268
rect 84304 7256 84332 7355
rect 84470 7352 84476 7364
rect 84528 7352 84534 7404
rect 84580 7401 84608 7500
rect 85301 7497 85313 7531
rect 85347 7528 85359 7531
rect 85482 7528 85488 7540
rect 85347 7500 85488 7528
rect 85347 7497 85359 7500
rect 85301 7491 85359 7497
rect 85482 7488 85488 7500
rect 85540 7488 85546 7540
rect 85942 7488 85948 7540
rect 86000 7528 86006 7540
rect 86037 7531 86095 7537
rect 86037 7528 86049 7531
rect 86000 7500 86049 7528
rect 86000 7488 86006 7500
rect 86037 7497 86049 7500
rect 86083 7497 86095 7531
rect 86586 7528 86592 7540
rect 86547 7500 86592 7528
rect 86037 7491 86095 7497
rect 86586 7488 86592 7500
rect 86644 7488 86650 7540
rect 92842 7488 92848 7540
rect 92900 7528 92906 7540
rect 93121 7531 93179 7537
rect 93121 7528 93133 7531
rect 92900 7500 93133 7528
rect 92900 7488 92906 7500
rect 93121 7497 93133 7500
rect 93167 7497 93179 7531
rect 93121 7491 93179 7497
rect 84749 7463 84807 7469
rect 84749 7429 84761 7463
rect 84795 7460 84807 7463
rect 88334 7460 88340 7472
rect 84795 7432 88340 7460
rect 84795 7429 84807 7432
rect 84749 7423 84807 7429
rect 88334 7420 88340 7432
rect 88392 7420 88398 7472
rect 89162 7460 89168 7472
rect 89123 7432 89168 7460
rect 89162 7420 89168 7432
rect 89220 7420 89226 7472
rect 90450 7420 90456 7472
rect 90508 7460 90514 7472
rect 93026 7460 93032 7472
rect 90508 7432 93032 7460
rect 90508 7420 90514 7432
rect 84565 7395 84623 7401
rect 84565 7361 84577 7395
rect 84611 7361 84623 7395
rect 84565 7355 84623 7361
rect 85945 7395 86003 7401
rect 85945 7361 85957 7395
rect 85991 7392 86003 7395
rect 86034 7392 86040 7404
rect 85991 7364 86040 7392
rect 85991 7361 86003 7364
rect 85945 7355 86003 7361
rect 86034 7352 86040 7364
rect 86092 7352 86098 7404
rect 87509 7395 87567 7401
rect 87509 7392 87521 7395
rect 87064 7364 87521 7392
rect 85022 7284 85028 7336
rect 85080 7324 85086 7336
rect 87064 7324 87092 7364
rect 87509 7361 87521 7364
rect 87555 7392 87567 7395
rect 88245 7395 88303 7401
rect 87555 7364 88196 7392
rect 87555 7361 87567 7364
rect 87509 7355 87567 7361
rect 85080 7296 87092 7324
rect 85080 7284 85086 7296
rect 87138 7284 87144 7336
rect 87196 7324 87202 7336
rect 87233 7327 87291 7333
rect 87233 7324 87245 7327
rect 87196 7296 87245 7324
rect 87196 7284 87202 7296
rect 87233 7293 87245 7296
rect 87279 7293 87291 7327
rect 87233 7287 87291 7293
rect 84654 7256 84660 7268
rect 84304 7228 84660 7256
rect 84654 7216 84660 7228
rect 84712 7216 84718 7268
rect 88168 7256 88196 7364
rect 88245 7361 88257 7395
rect 88291 7392 88303 7395
rect 88426 7392 88432 7404
rect 88291 7364 88432 7392
rect 88291 7361 88303 7364
rect 88245 7355 88303 7361
rect 88426 7352 88432 7364
rect 88484 7352 88490 7404
rect 91002 7352 91008 7404
rect 91060 7392 91066 7404
rect 92308 7401 92336 7432
rect 93026 7420 93032 7432
rect 93084 7420 93090 7472
rect 91557 7395 91615 7401
rect 91557 7392 91569 7395
rect 91060 7364 91569 7392
rect 91060 7352 91066 7364
rect 91557 7361 91569 7364
rect 91603 7392 91615 7395
rect 92293 7395 92351 7401
rect 91603 7364 91968 7392
rect 91603 7361 91615 7364
rect 91557 7355 91615 7361
rect 88886 7284 88892 7336
rect 88944 7324 88950 7336
rect 88981 7327 89039 7333
rect 88981 7324 88993 7327
rect 88944 7296 88993 7324
rect 88944 7284 88950 7296
rect 88981 7293 88993 7296
rect 89027 7293 89039 7327
rect 88981 7287 89039 7293
rect 89441 7327 89499 7333
rect 89441 7293 89453 7327
rect 89487 7293 89499 7327
rect 89441 7287 89499 7293
rect 89070 7256 89076 7268
rect 88168 7228 89076 7256
rect 89070 7216 89076 7228
rect 89128 7256 89134 7268
rect 89456 7256 89484 7287
rect 90174 7284 90180 7336
rect 90232 7324 90238 7336
rect 91281 7327 91339 7333
rect 91281 7324 91293 7327
rect 90232 7296 91293 7324
rect 90232 7284 90238 7296
rect 91281 7293 91293 7296
rect 91327 7293 91339 7327
rect 91940 7324 91968 7364
rect 92293 7361 92305 7395
rect 92339 7361 92351 7395
rect 92934 7392 92940 7404
rect 92895 7364 92940 7392
rect 92293 7355 92351 7361
rect 92934 7352 92940 7364
rect 92992 7352 92998 7404
rect 94133 7327 94191 7333
rect 94133 7324 94145 7327
rect 91940 7296 94145 7324
rect 91281 7287 91339 7293
rect 94133 7293 94145 7296
rect 94179 7293 94191 7327
rect 94133 7287 94191 7293
rect 89714 7256 89720 7268
rect 89128 7228 89720 7256
rect 89128 7216 89134 7228
rect 89714 7216 89720 7228
rect 89772 7216 89778 7268
rect 72016 7160 76236 7188
rect 76285 7191 76343 7197
rect 72016 7148 72022 7160
rect 76285 7157 76297 7191
rect 76331 7188 76343 7191
rect 76466 7188 76472 7200
rect 76331 7160 76472 7188
rect 76331 7157 76343 7160
rect 76285 7151 76343 7157
rect 76466 7148 76472 7160
rect 76524 7148 76530 7200
rect 79870 7188 79876 7200
rect 79831 7160 79876 7188
rect 79870 7148 79876 7160
rect 79928 7148 79934 7200
rect 80054 7148 80060 7200
rect 80112 7188 80118 7200
rect 82814 7188 82820 7200
rect 80112 7160 80157 7188
rect 82775 7160 82820 7188
rect 80112 7148 80118 7160
rect 82814 7148 82820 7160
rect 82872 7148 82878 7200
rect 88429 7191 88487 7197
rect 88429 7157 88441 7191
rect 88475 7188 88487 7191
rect 89806 7188 89812 7200
rect 88475 7160 89812 7188
rect 88475 7157 88487 7160
rect 88429 7151 88487 7157
rect 89806 7148 89812 7160
rect 89864 7148 89870 7200
rect 92477 7191 92535 7197
rect 92477 7157 92489 7191
rect 92523 7188 92535 7191
rect 92750 7188 92756 7200
rect 92523 7160 92756 7188
rect 92523 7157 92535 7160
rect 92477 7151 92535 7157
rect 92750 7148 92756 7160
rect 92808 7148 92814 7200
rect 1104 7098 94852 7120
rect 1104 7046 12668 7098
rect 12720 7046 12732 7098
rect 12784 7046 12796 7098
rect 12848 7046 12860 7098
rect 12912 7046 12924 7098
rect 12976 7046 36105 7098
rect 36157 7046 36169 7098
rect 36221 7046 36233 7098
rect 36285 7046 36297 7098
rect 36349 7046 36361 7098
rect 36413 7046 59542 7098
rect 59594 7046 59606 7098
rect 59658 7046 59670 7098
rect 59722 7046 59734 7098
rect 59786 7046 59798 7098
rect 59850 7046 82979 7098
rect 83031 7046 83043 7098
rect 83095 7046 83107 7098
rect 83159 7046 83171 7098
rect 83223 7046 83235 7098
rect 83287 7046 94852 7098
rect 1104 7024 94852 7046
rect 12342 6984 12348 6996
rect 10060 6956 12348 6984
rect 4246 6848 4252 6860
rect 4159 6820 4252 6848
rect 4246 6808 4252 6820
rect 4304 6848 4310 6860
rect 5166 6848 5172 6860
rect 4304 6820 5172 6848
rect 4304 6808 4310 6820
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 9674 6848 9680 6860
rect 8128 6820 9680 6848
rect 8128 6792 8156 6820
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 9858 6808 9864 6860
rect 9916 6848 9922 6860
rect 10060 6857 10088 6956
rect 12342 6944 12348 6956
rect 12400 6984 12406 6996
rect 13722 6984 13728 6996
rect 12400 6956 13728 6984
rect 12400 6944 12406 6956
rect 10686 6876 10692 6928
rect 10744 6876 10750 6928
rect 10045 6851 10103 6857
rect 10045 6848 10057 6851
rect 9916 6820 10057 6848
rect 9916 6808 9922 6820
rect 10045 6817 10057 6820
rect 10091 6817 10103 6851
rect 10704 6848 10732 6876
rect 12912 6857 12940 6956
rect 13722 6944 13728 6956
rect 13780 6944 13786 6996
rect 20898 6944 20904 6996
rect 20956 6984 20962 6996
rect 21453 6987 21511 6993
rect 21453 6984 21465 6987
rect 20956 6956 21465 6984
rect 20956 6944 20962 6956
rect 21453 6953 21465 6956
rect 21499 6953 21511 6987
rect 21453 6947 21511 6953
rect 22097 6987 22155 6993
rect 22097 6953 22109 6987
rect 22143 6984 22155 6987
rect 22278 6984 22284 6996
rect 22143 6956 22284 6984
rect 22143 6953 22155 6956
rect 22097 6947 22155 6953
rect 22278 6944 22284 6956
rect 22336 6944 22342 6996
rect 25130 6984 25136 6996
rect 22388 6956 25136 6984
rect 16669 6919 16727 6925
rect 14476 6888 14688 6916
rect 12894 6851 12952 6857
rect 10704 6820 11928 6848
rect 10045 6811 10103 6817
rect 3053 6783 3111 6789
rect 3053 6749 3065 6783
rect 3099 6749 3111 6783
rect 4154 6780 4160 6792
rect 4115 6752 4160 6780
rect 3053 6743 3111 6749
rect 3068 6712 3096 6743
rect 4154 6740 4160 6752
rect 4212 6740 4218 6792
rect 6914 6780 6920 6792
rect 4264 6752 6920 6780
rect 4264 6712 4292 6752
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 7193 6783 7251 6789
rect 7193 6749 7205 6783
rect 7239 6749 7251 6783
rect 7193 6743 7251 6749
rect 7469 6783 7527 6789
rect 7469 6749 7481 6783
rect 7515 6780 7527 6783
rect 7558 6780 7564 6792
rect 7515 6752 7564 6780
rect 7515 6749 7527 6752
rect 7469 6743 7527 6749
rect 6730 6712 6736 6724
rect 3068 6684 4292 6712
rect 4540 6684 6736 6712
rect 3237 6647 3295 6653
rect 3237 6613 3249 6647
rect 3283 6644 3295 6647
rect 4154 6644 4160 6656
rect 3283 6616 4160 6644
rect 3283 6613 3295 6616
rect 3237 6607 3295 6613
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4540 6653 4568 6684
rect 6730 6672 6736 6684
rect 6788 6672 6794 6724
rect 7208 6712 7236 6743
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 8110 6780 8116 6792
rect 8023 6752 8116 6780
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 10321 6783 10379 6789
rect 10321 6776 10333 6783
rect 10244 6749 10333 6776
rect 10367 6749 10379 6783
rect 10244 6748 10379 6749
rect 8294 6712 8300 6724
rect 7208 6684 8300 6712
rect 8294 6672 8300 6684
rect 8352 6672 8358 6724
rect 8389 6715 8447 6721
rect 8389 6681 8401 6715
rect 8435 6712 8447 6715
rect 8570 6712 8576 6724
rect 8435 6684 8576 6712
rect 8435 6681 8447 6684
rect 8389 6675 8447 6681
rect 8570 6672 8576 6684
rect 8628 6672 8634 6724
rect 4525 6647 4583 6653
rect 4525 6613 4537 6647
rect 4571 6613 4583 6647
rect 5074 6644 5080 6656
rect 5035 6616 5080 6644
rect 4525 6607 4583 6613
rect 5074 6604 5080 6616
rect 5132 6604 5138 6656
rect 6638 6644 6644 6656
rect 6599 6616 6644 6644
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 9585 6647 9643 6653
rect 9585 6613 9597 6647
rect 9631 6644 9643 6647
rect 10134 6644 10140 6656
rect 9631 6616 10140 6644
rect 9631 6613 9643 6616
rect 9585 6607 9643 6613
rect 10134 6604 10140 6616
rect 10192 6644 10198 6656
rect 10244 6644 10272 6748
rect 10321 6743 10379 6748
rect 10778 6740 10784 6792
rect 10836 6780 10842 6792
rect 11900 6789 11928 6820
rect 12894 6817 12906 6851
rect 12940 6817 12952 6851
rect 12894 6811 12952 6817
rect 13449 6851 13507 6857
rect 13449 6817 13461 6851
rect 13495 6848 13507 6851
rect 14476 6848 14504 6888
rect 13495 6820 14504 6848
rect 14553 6851 14611 6857
rect 13495 6817 13507 6820
rect 13449 6811 13507 6817
rect 14553 6817 14565 6851
rect 14599 6817 14611 6851
rect 14660 6848 14688 6888
rect 16669 6885 16681 6919
rect 16715 6916 16727 6919
rect 16942 6916 16948 6928
rect 16715 6888 16948 6916
rect 16715 6885 16727 6888
rect 16669 6879 16727 6885
rect 16942 6876 16948 6888
rect 17000 6916 17006 6928
rect 17954 6916 17960 6928
rect 17000 6888 17960 6916
rect 17000 6876 17006 6888
rect 17954 6876 17960 6888
rect 18012 6876 18018 6928
rect 18230 6876 18236 6928
rect 18288 6916 18294 6928
rect 18288 6888 20208 6916
rect 18288 6876 18294 6888
rect 20180 6857 20208 6888
rect 22186 6876 22192 6928
rect 22244 6916 22250 6928
rect 22388 6916 22416 6956
rect 25130 6944 25136 6956
rect 25188 6944 25194 6996
rect 28074 6984 28080 6996
rect 25240 6956 26648 6984
rect 28035 6956 28080 6984
rect 22244 6888 22416 6916
rect 22925 6919 22983 6925
rect 22244 6876 22250 6888
rect 22925 6885 22937 6919
rect 22971 6916 22983 6919
rect 22971 6888 23704 6916
rect 22971 6885 22983 6888
rect 22925 6879 22983 6885
rect 20165 6851 20223 6857
rect 14660 6820 20116 6848
rect 14553 6811 14611 6817
rect 10965 6783 11023 6789
rect 10965 6780 10977 6783
rect 10836 6752 10977 6780
rect 10836 6740 10842 6752
rect 10965 6749 10977 6752
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6749 11943 6783
rect 12618 6780 12624 6792
rect 12531 6752 12624 6780
rect 11885 6743 11943 6749
rect 12618 6740 12624 6752
rect 12676 6780 12682 6792
rect 13464 6780 13492 6811
rect 12676 6752 13492 6780
rect 12676 6740 12682 6752
rect 10502 6672 10508 6724
rect 10560 6712 10566 6724
rect 14568 6712 14596 6811
rect 14645 6783 14703 6789
rect 14645 6749 14657 6783
rect 14691 6780 14703 6783
rect 15010 6780 15016 6792
rect 14691 6752 15016 6780
rect 14691 6749 14703 6752
rect 14645 6743 14703 6749
rect 15010 6740 15016 6752
rect 15068 6740 15074 6792
rect 15286 6780 15292 6792
rect 15247 6752 15292 6780
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 17310 6740 17316 6792
rect 17368 6780 17374 6792
rect 18785 6783 18843 6789
rect 18785 6780 18797 6783
rect 17368 6752 18797 6780
rect 17368 6740 17374 6752
rect 18785 6749 18797 6752
rect 18831 6749 18843 6783
rect 19981 6783 20039 6789
rect 19981 6780 19993 6783
rect 18785 6743 18843 6749
rect 19444 6752 19993 6780
rect 10560 6684 14596 6712
rect 10560 6672 10566 6684
rect 10192 6616 10272 6644
rect 10192 6604 10198 6616
rect 10410 6604 10416 6656
rect 10468 6644 10474 6656
rect 11241 6647 11299 6653
rect 11241 6644 11253 6647
rect 10468 6616 11253 6644
rect 10468 6604 10474 6616
rect 11241 6613 11253 6616
rect 11287 6644 11299 6647
rect 11701 6647 11759 6653
rect 11701 6644 11713 6647
rect 11287 6616 11713 6644
rect 11287 6613 11299 6616
rect 11241 6607 11299 6613
rect 11701 6613 11713 6616
rect 11747 6613 11759 6647
rect 11701 6607 11759 6613
rect 13630 6604 13636 6656
rect 13688 6644 13694 6656
rect 14277 6647 14335 6653
rect 14277 6644 14289 6647
rect 13688 6616 14289 6644
rect 13688 6604 13694 6616
rect 14277 6613 14289 6616
rect 14323 6613 14335 6647
rect 15304 6644 15332 6740
rect 17954 6672 17960 6724
rect 18012 6712 18018 6724
rect 19444 6721 19472 6752
rect 19981 6749 19993 6752
rect 20027 6749 20039 6783
rect 20088 6780 20116 6820
rect 20165 6817 20177 6851
rect 20211 6848 20223 6851
rect 20438 6848 20444 6860
rect 20211 6820 20444 6848
rect 20211 6817 20223 6820
rect 20165 6811 20223 6817
rect 20438 6808 20444 6820
rect 20496 6808 20502 6860
rect 20530 6808 20536 6860
rect 20588 6848 20594 6860
rect 23569 6851 23627 6857
rect 23569 6848 23581 6851
rect 20588 6820 23581 6848
rect 20588 6808 20594 6820
rect 23569 6817 23581 6820
rect 23615 6817 23627 6851
rect 23569 6811 23627 6817
rect 23014 6780 23020 6792
rect 20088 6752 22876 6780
rect 22975 6752 23020 6780
rect 19981 6743 20039 6749
rect 19429 6715 19487 6721
rect 19429 6712 19441 6715
rect 18012 6684 19441 6712
rect 18012 6672 18018 6684
rect 19429 6681 19441 6684
rect 19475 6681 19487 6715
rect 19996 6712 20024 6743
rect 20993 6715 21051 6721
rect 20993 6712 21005 6715
rect 19996 6684 21005 6712
rect 19429 6675 19487 6681
rect 20993 6681 21005 6684
rect 21039 6712 21051 6715
rect 22094 6712 22100 6724
rect 21039 6684 22100 6712
rect 21039 6681 21051 6684
rect 20993 6675 21051 6681
rect 22066 6672 22100 6684
rect 22152 6672 22158 6724
rect 22738 6712 22744 6724
rect 22699 6684 22744 6712
rect 22738 6672 22744 6684
rect 22796 6672 22802 6724
rect 22848 6712 22876 6752
rect 23014 6740 23020 6752
rect 23072 6740 23078 6792
rect 23676 6789 23704 6888
rect 24854 6848 24860 6860
rect 24815 6820 24860 6848
rect 24854 6808 24860 6820
rect 24912 6808 24918 6860
rect 23661 6783 23719 6789
rect 23661 6749 23673 6783
rect 23707 6780 23719 6783
rect 23750 6780 23756 6792
rect 23707 6752 23756 6780
rect 23707 6749 23719 6752
rect 23661 6743 23719 6749
rect 23750 6740 23756 6752
rect 23808 6780 23814 6792
rect 25240 6780 25268 6956
rect 25317 6851 25375 6857
rect 25317 6817 25329 6851
rect 25363 6848 25375 6851
rect 26326 6848 26332 6860
rect 25363 6820 26332 6848
rect 25363 6817 25375 6820
rect 25317 6811 25375 6817
rect 26326 6808 26332 6820
rect 26384 6808 26390 6860
rect 26620 6848 26648 6956
rect 28074 6944 28080 6956
rect 28132 6944 28138 6996
rect 28442 6944 28448 6996
rect 28500 6984 28506 6996
rect 28721 6987 28779 6993
rect 28721 6984 28733 6987
rect 28500 6956 28733 6984
rect 28500 6944 28506 6956
rect 28721 6953 28733 6956
rect 28767 6953 28779 6987
rect 28721 6947 28779 6953
rect 32235 6987 32293 6993
rect 32235 6953 32247 6987
rect 32281 6984 32293 6987
rect 34054 6984 34060 6996
rect 32281 6956 34060 6984
rect 32281 6953 32293 6956
rect 32235 6947 32293 6953
rect 34054 6944 34060 6956
rect 34112 6944 34118 6996
rect 35158 6993 35164 6996
rect 35148 6987 35164 6993
rect 35148 6953 35160 6987
rect 35148 6947 35164 6953
rect 35158 6944 35164 6947
rect 35216 6944 35222 6996
rect 35250 6944 35256 6996
rect 35308 6984 35314 6996
rect 36998 6984 37004 6996
rect 35308 6956 37004 6984
rect 35308 6944 35314 6956
rect 36998 6944 37004 6956
rect 37056 6944 37062 6996
rect 37826 6984 37832 6996
rect 37787 6956 37832 6984
rect 37826 6944 37832 6956
rect 37884 6944 37890 6996
rect 38933 6987 38991 6993
rect 38933 6953 38945 6987
rect 38979 6984 38991 6987
rect 39022 6984 39028 6996
rect 38979 6956 39028 6984
rect 38979 6953 38991 6956
rect 38933 6947 38991 6953
rect 39022 6944 39028 6956
rect 39080 6944 39086 6996
rect 40770 6944 40776 6996
rect 40828 6984 40834 6996
rect 41049 6987 41107 6993
rect 41049 6984 41061 6987
rect 40828 6956 41061 6984
rect 40828 6944 40834 6956
rect 41049 6953 41061 6956
rect 41095 6953 41107 6987
rect 41049 6947 41107 6953
rect 41506 6944 41512 6996
rect 41564 6984 41570 6996
rect 45738 6984 45744 6996
rect 41564 6956 45744 6984
rect 41564 6944 41570 6956
rect 45738 6944 45744 6956
rect 45796 6944 45802 6996
rect 49237 6987 49295 6993
rect 49237 6984 49249 6987
rect 48332 6956 49249 6984
rect 26694 6876 26700 6928
rect 26752 6916 26758 6928
rect 31202 6916 31208 6928
rect 26752 6888 31208 6916
rect 26752 6876 26758 6888
rect 31202 6876 31208 6888
rect 31260 6876 31266 6928
rect 32858 6916 32864 6928
rect 32508 6888 32864 6916
rect 28442 6848 28448 6860
rect 26620 6820 28448 6848
rect 28442 6808 28448 6820
rect 28500 6808 28506 6860
rect 29454 6808 29460 6860
rect 29512 6848 29518 6860
rect 29917 6851 29975 6857
rect 29917 6848 29929 6851
rect 29512 6820 29929 6848
rect 29512 6808 29518 6820
rect 29917 6817 29929 6820
rect 29963 6817 29975 6851
rect 29917 6811 29975 6817
rect 30190 6808 30196 6860
rect 30248 6848 30254 6860
rect 32508 6857 32536 6888
rect 32858 6876 32864 6888
rect 32916 6916 32922 6928
rect 32916 6888 33548 6916
rect 32916 6876 32922 6888
rect 32493 6851 32551 6857
rect 32493 6848 32505 6851
rect 30248 6820 32505 6848
rect 30248 6808 30254 6820
rect 32493 6817 32505 6820
rect 32539 6817 32551 6851
rect 32493 6811 32551 6817
rect 32953 6851 33011 6857
rect 32953 6817 32965 6851
rect 32999 6848 33011 6851
rect 33134 6848 33140 6860
rect 32999 6820 33140 6848
rect 32999 6817 33011 6820
rect 32953 6811 33011 6817
rect 33134 6808 33140 6820
rect 33192 6808 33198 6860
rect 33410 6848 33416 6860
rect 33371 6820 33416 6848
rect 33410 6808 33416 6820
rect 33468 6808 33474 6860
rect 33520 6848 33548 6888
rect 34146 6876 34152 6928
rect 34204 6916 34210 6928
rect 34204 6888 34249 6916
rect 34204 6876 34210 6888
rect 36170 6876 36176 6928
rect 36228 6916 36234 6928
rect 37366 6916 37372 6928
rect 36228 6888 37372 6916
rect 36228 6876 36234 6888
rect 37366 6876 37372 6888
rect 37424 6876 37430 6928
rect 38010 6876 38016 6928
rect 38068 6916 38074 6928
rect 38068 6888 39252 6916
rect 38068 6876 38074 6888
rect 34882 6848 34888 6860
rect 33520 6820 34888 6848
rect 34882 6808 34888 6820
rect 34940 6808 34946 6860
rect 35802 6808 35808 6860
rect 35860 6848 35866 6860
rect 36633 6851 36691 6857
rect 36633 6848 36645 6851
rect 35860 6820 36645 6848
rect 35860 6808 35866 6820
rect 36633 6817 36645 6820
rect 36679 6817 36691 6851
rect 37274 6848 37280 6860
rect 37235 6820 37280 6848
rect 36633 6811 36691 6817
rect 23808 6752 25268 6780
rect 27341 6783 27399 6789
rect 23808 6740 23814 6752
rect 27341 6749 27353 6783
rect 27387 6780 27399 6783
rect 30098 6780 30104 6792
rect 27387 6752 30104 6780
rect 27387 6749 27399 6752
rect 27341 6743 27399 6749
rect 30098 6740 30104 6752
rect 30156 6740 30162 6792
rect 33318 6780 33324 6792
rect 33279 6752 33324 6780
rect 33318 6740 33324 6752
rect 33376 6740 33382 6792
rect 33778 6740 33784 6792
rect 33836 6780 33842 6792
rect 34698 6780 34704 6792
rect 33836 6752 34284 6780
rect 34348 6767 34704 6780
rect 33836 6740 33842 6752
rect 34256 6724 34284 6752
rect 34331 6761 34704 6767
rect 34331 6727 34343 6761
rect 34377 6752 34704 6761
rect 34377 6727 34389 6752
rect 34698 6740 34704 6752
rect 34756 6740 34762 6792
rect 36648 6780 36676 6811
rect 37274 6808 37280 6820
rect 37332 6808 37338 6860
rect 38470 6848 38476 6860
rect 38431 6820 38476 6848
rect 38470 6808 38476 6820
rect 38528 6808 38534 6860
rect 38838 6808 38844 6860
rect 38896 6848 38902 6860
rect 39224 6848 39252 6888
rect 40218 6876 40224 6928
rect 40276 6916 40282 6928
rect 40405 6919 40463 6925
rect 40405 6916 40417 6919
rect 40276 6888 40417 6916
rect 40276 6876 40282 6888
rect 40405 6885 40417 6888
rect 40451 6916 40463 6919
rect 40862 6916 40868 6928
rect 40451 6888 40868 6916
rect 40451 6885 40463 6888
rect 40405 6879 40463 6885
rect 40862 6876 40868 6888
rect 40920 6876 40926 6928
rect 41230 6876 41236 6928
rect 41288 6916 41294 6928
rect 43070 6916 43076 6928
rect 41288 6888 43076 6916
rect 41288 6876 41294 6888
rect 43070 6876 43076 6888
rect 43128 6876 43134 6928
rect 40034 6848 40040 6860
rect 38896 6820 39160 6848
rect 39224 6820 39620 6848
rect 39995 6820 40040 6848
rect 38896 6808 38902 6820
rect 39022 6780 39028 6792
rect 36648 6752 39028 6780
rect 39022 6740 39028 6752
rect 39080 6740 39086 6792
rect 39132 6789 39160 6820
rect 39117 6783 39175 6789
rect 39117 6749 39129 6783
rect 39163 6749 39175 6783
rect 39117 6743 39175 6749
rect 39393 6783 39451 6789
rect 39393 6749 39405 6783
rect 39439 6780 39451 6783
rect 39592 6780 39620 6820
rect 40034 6808 40040 6820
rect 40092 6808 40098 6860
rect 40497 6851 40555 6857
rect 40497 6817 40509 6851
rect 40543 6848 40555 6851
rect 41966 6848 41972 6860
rect 40543 6820 41972 6848
rect 40543 6817 40555 6820
rect 40497 6811 40555 6817
rect 41966 6808 41972 6820
rect 42024 6808 42030 6860
rect 42886 6848 42892 6860
rect 42847 6820 42892 6848
rect 42886 6808 42892 6820
rect 42944 6808 42950 6860
rect 43438 6848 43444 6860
rect 42996 6820 43444 6848
rect 40770 6780 40776 6792
rect 39439 6752 39528 6780
rect 39592 6752 40776 6780
rect 39439 6749 39451 6752
rect 39393 6743 39451 6749
rect 25590 6712 25596 6724
rect 22848 6684 24900 6712
rect 25551 6684 25596 6712
rect 18230 6644 18236 6656
rect 15304 6616 18236 6644
rect 14277 6607 14335 6613
rect 18230 6604 18236 6616
rect 18288 6604 18294 6656
rect 22066 6644 22094 6672
rect 22922 6644 22928 6656
rect 22066 6616 22928 6644
rect 22922 6604 22928 6616
rect 22980 6604 22986 6656
rect 23017 6647 23075 6653
rect 23017 6613 23029 6647
rect 23063 6644 23075 6647
rect 23382 6644 23388 6656
rect 23063 6616 23388 6644
rect 23063 6613 23075 6616
rect 23017 6607 23075 6613
rect 23382 6604 23388 6616
rect 23440 6604 23446 6656
rect 24029 6647 24087 6653
rect 24029 6613 24041 6647
rect 24075 6644 24087 6647
rect 24118 6644 24124 6656
rect 24075 6616 24124 6644
rect 24075 6613 24087 6616
rect 24029 6607 24087 6613
rect 24118 6604 24124 6616
rect 24176 6604 24182 6656
rect 24872 6644 24900 6684
rect 25590 6672 25596 6684
rect 25648 6672 25654 6724
rect 26234 6672 26240 6724
rect 26292 6672 26298 6724
rect 26896 6684 28120 6712
rect 26896 6644 26924 6684
rect 24872 6616 26924 6644
rect 28092 6644 28120 6684
rect 28166 6672 28172 6724
rect 28224 6712 28230 6724
rect 28537 6715 28595 6721
rect 28537 6712 28549 6715
rect 28224 6684 28549 6712
rect 28224 6672 28230 6684
rect 28537 6681 28549 6684
rect 28583 6681 28595 6715
rect 30466 6712 30472 6724
rect 28537 6675 28595 6681
rect 28644 6684 30052 6712
rect 30427 6684 30472 6712
rect 28644 6644 28672 6684
rect 28092 6616 28672 6644
rect 28718 6604 28724 6656
rect 28776 6653 28782 6656
rect 28776 6647 28795 6653
rect 28783 6613 28795 6647
rect 28776 6607 28795 6613
rect 28905 6647 28963 6653
rect 28905 6613 28917 6647
rect 28951 6644 28963 6647
rect 29730 6644 29736 6656
rect 28951 6616 29736 6644
rect 28951 6613 28963 6616
rect 28905 6607 28963 6613
rect 28776 6604 28782 6607
rect 29730 6604 29736 6616
rect 29788 6604 29794 6656
rect 30024 6644 30052 6684
rect 30466 6672 30472 6684
rect 30524 6672 30530 6724
rect 31662 6672 31668 6724
rect 31720 6672 31726 6724
rect 33042 6712 33048 6724
rect 32232 6684 33048 6712
rect 32232 6644 32260 6684
rect 33042 6672 33048 6684
rect 33100 6672 33106 6724
rect 33870 6672 33876 6724
rect 33928 6712 33934 6724
rect 34057 6715 34115 6721
rect 34057 6712 34069 6715
rect 33928 6684 34069 6712
rect 33928 6672 33934 6684
rect 34057 6681 34069 6684
rect 34103 6681 34115 6715
rect 34238 6712 34244 6724
rect 34151 6684 34244 6712
rect 34057 6675 34115 6681
rect 34238 6672 34244 6684
rect 34296 6672 34302 6724
rect 34331 6721 34389 6727
rect 34514 6672 34520 6724
rect 34572 6712 34578 6724
rect 35618 6712 35624 6724
rect 34572 6684 35624 6712
rect 34572 6672 34578 6684
rect 35618 6672 35624 6684
rect 35676 6672 35682 6724
rect 39500 6712 39528 6752
rect 40770 6740 40776 6752
rect 40828 6780 40834 6792
rect 40957 6783 41015 6789
rect 40957 6780 40969 6783
rect 40828 6752 40969 6780
rect 40828 6740 40834 6752
rect 40957 6749 40969 6752
rect 41003 6749 41015 6783
rect 41138 6780 41144 6792
rect 41099 6752 41144 6780
rect 40957 6743 41015 6749
rect 41138 6740 41144 6752
rect 41196 6740 41202 6792
rect 42797 6783 42855 6789
rect 42797 6780 42809 6783
rect 41386 6752 42809 6780
rect 40310 6712 40316 6724
rect 36464 6684 39436 6712
rect 39500 6684 40316 6712
rect 30024 6616 32260 6644
rect 33410 6604 33416 6656
rect 33468 6644 33474 6656
rect 34882 6644 34888 6656
rect 33468 6616 34888 6644
rect 33468 6604 33474 6616
rect 34882 6604 34888 6616
rect 34940 6644 34946 6656
rect 36464 6644 36492 6684
rect 34940 6616 36492 6644
rect 34940 6604 34946 6616
rect 36722 6604 36728 6656
rect 36780 6644 36786 6656
rect 38930 6644 38936 6656
rect 36780 6616 38936 6644
rect 36780 6604 36786 6616
rect 38930 6604 38936 6616
rect 38988 6604 38994 6656
rect 39298 6644 39304 6656
rect 39259 6616 39304 6644
rect 39298 6604 39304 6616
rect 39356 6604 39362 6656
rect 39408 6644 39436 6684
rect 40310 6672 40316 6684
rect 40368 6672 40374 6724
rect 40862 6672 40868 6724
rect 40920 6712 40926 6724
rect 41386 6712 41414 6752
rect 42797 6749 42809 6752
rect 42843 6780 42855 6783
rect 42996 6780 43024 6820
rect 43438 6808 43444 6820
rect 43496 6808 43502 6860
rect 44634 6848 44640 6860
rect 44595 6820 44640 6848
rect 44634 6808 44640 6820
rect 44692 6808 44698 6860
rect 44910 6808 44916 6860
rect 44968 6848 44974 6860
rect 45465 6851 45523 6857
rect 45465 6848 45477 6851
rect 44968 6820 45477 6848
rect 44968 6808 44974 6820
rect 45465 6817 45477 6820
rect 45511 6848 45523 6851
rect 45830 6848 45836 6860
rect 45511 6820 45836 6848
rect 45511 6817 45523 6820
rect 45465 6811 45523 6817
rect 45830 6808 45836 6820
rect 45888 6808 45894 6860
rect 48332 6848 48360 6956
rect 49237 6953 49249 6956
rect 49283 6984 49295 6987
rect 49602 6984 49608 6996
rect 49283 6956 49608 6984
rect 49283 6953 49295 6956
rect 49237 6947 49295 6953
rect 49602 6944 49608 6956
rect 49660 6944 49666 6996
rect 50604 6987 50662 6993
rect 50604 6953 50616 6987
rect 50650 6984 50662 6987
rect 52641 6987 52699 6993
rect 52641 6984 52653 6987
rect 50650 6956 52653 6984
rect 50650 6953 50662 6956
rect 50604 6947 50662 6953
rect 52641 6953 52653 6956
rect 52687 6953 52699 6987
rect 52641 6947 52699 6953
rect 53282 6944 53288 6996
rect 53340 6984 53346 6996
rect 53745 6987 53803 6993
rect 53745 6984 53757 6987
rect 53340 6956 53757 6984
rect 53340 6944 53346 6956
rect 53745 6953 53757 6956
rect 53791 6953 53803 6987
rect 53745 6947 53803 6953
rect 54573 6987 54631 6993
rect 54573 6953 54585 6987
rect 54619 6984 54631 6987
rect 54846 6984 54852 6996
rect 54619 6956 54852 6984
rect 54619 6953 54631 6956
rect 54573 6947 54631 6953
rect 54846 6944 54852 6956
rect 54904 6944 54910 6996
rect 58526 6984 58532 6996
rect 58487 6956 58532 6984
rect 58526 6944 58532 6956
rect 58584 6944 58590 6996
rect 61102 6944 61108 6996
rect 61160 6984 61166 6996
rect 61160 6956 64828 6984
rect 61160 6944 61166 6956
rect 51902 6876 51908 6928
rect 51960 6916 51966 6928
rect 56778 6916 56784 6928
rect 51960 6888 56784 6916
rect 51960 6876 51966 6888
rect 56778 6876 56784 6888
rect 56836 6876 56842 6928
rect 48774 6848 48780 6860
rect 46032 6820 48360 6848
rect 48735 6820 48780 6848
rect 42843 6752 43024 6780
rect 42843 6749 42855 6752
rect 42797 6743 42855 6749
rect 43070 6740 43076 6792
rect 43128 6780 43134 6792
rect 45189 6783 45247 6789
rect 45189 6780 45201 6783
rect 43128 6752 45201 6780
rect 43128 6740 43134 6752
rect 45189 6749 45201 6752
rect 45235 6749 45247 6783
rect 45189 6743 45247 6749
rect 45278 6740 45284 6792
rect 45336 6780 45342 6792
rect 46032 6789 46060 6820
rect 48774 6808 48780 6820
rect 48832 6808 48838 6860
rect 49421 6851 49479 6857
rect 49421 6817 49433 6851
rect 49467 6848 49479 6851
rect 50062 6848 50068 6860
rect 49467 6820 50068 6848
rect 49467 6817 49479 6820
rect 49421 6811 49479 6817
rect 50062 6808 50068 6820
rect 50120 6808 50126 6860
rect 50338 6848 50344 6860
rect 50299 6820 50344 6848
rect 50338 6808 50344 6820
rect 50396 6808 50402 6860
rect 50982 6808 50988 6860
rect 51040 6848 51046 6860
rect 53193 6851 53251 6857
rect 53193 6848 53205 6851
rect 51040 6820 53205 6848
rect 51040 6808 51046 6820
rect 53193 6817 53205 6820
rect 53239 6817 53251 6851
rect 53193 6811 53251 6817
rect 53466 6808 53472 6860
rect 53524 6848 53530 6860
rect 56410 6848 56416 6860
rect 53524 6820 54524 6848
rect 56371 6820 56416 6848
rect 53524 6808 53530 6820
rect 46017 6783 46075 6789
rect 45336 6752 45381 6780
rect 45336 6740 45342 6752
rect 46017 6749 46029 6783
rect 46063 6749 46075 6783
rect 46017 6743 46075 6749
rect 47857 6783 47915 6789
rect 47857 6749 47869 6783
rect 47903 6780 47915 6783
rect 47903 6752 49464 6780
rect 47903 6749 47915 6752
rect 47857 6743 47915 6749
rect 40920 6684 41414 6712
rect 41969 6715 42027 6721
rect 40920 6672 40926 6684
rect 41969 6681 41981 6715
rect 42015 6712 42027 6715
rect 43162 6712 43168 6724
rect 42015 6684 43168 6712
rect 42015 6681 42027 6684
rect 41969 6675 42027 6681
rect 41984 6644 42012 6675
rect 43162 6672 43168 6684
rect 43220 6672 43226 6724
rect 43346 6672 43352 6724
rect 43404 6712 43410 6724
rect 43533 6715 43591 6721
rect 43533 6712 43545 6715
rect 43404 6684 43545 6712
rect 43404 6672 43410 6684
rect 43533 6681 43545 6684
rect 43579 6681 43591 6715
rect 43533 6675 43591 6681
rect 44634 6672 44640 6724
rect 44692 6712 44698 6724
rect 46032 6712 46060 6743
rect 44692 6684 46060 6712
rect 46201 6715 46259 6721
rect 44692 6672 44698 6684
rect 46201 6681 46213 6715
rect 46247 6712 46259 6715
rect 46247 6684 47348 6712
rect 46247 6681 46259 6684
rect 46201 6675 46259 6681
rect 47320 6656 47348 6684
rect 49142 6672 49148 6724
rect 49200 6712 49206 6724
rect 49237 6715 49295 6721
rect 49237 6712 49249 6715
rect 49200 6684 49249 6712
rect 49200 6672 49206 6684
rect 49237 6681 49249 6684
rect 49283 6681 49295 6715
rect 49436 6712 49464 6752
rect 49510 6740 49516 6792
rect 49568 6780 49574 6792
rect 52733 6783 52791 6789
rect 49568 6752 49613 6780
rect 49568 6740 49574 6752
rect 52733 6749 52745 6783
rect 52779 6780 52791 6783
rect 53650 6780 53656 6792
rect 52779 6752 53656 6780
rect 52779 6749 52791 6752
rect 52733 6743 52791 6749
rect 53650 6740 53656 6752
rect 53708 6740 53714 6792
rect 54389 6783 54447 6789
rect 54389 6749 54401 6783
rect 54435 6749 54447 6783
rect 54389 6743 54447 6749
rect 52914 6712 52920 6724
rect 49436 6684 49832 6712
rect 51842 6684 52920 6712
rect 49237 6675 49295 6681
rect 42426 6644 42432 6656
rect 39408 6616 42012 6644
rect 42387 6616 42432 6644
rect 42426 6604 42432 6616
rect 42484 6604 42490 6656
rect 42886 6604 42892 6656
rect 42944 6644 42950 6656
rect 43625 6647 43683 6653
rect 43625 6644 43637 6647
rect 42944 6616 43637 6644
rect 42944 6604 42950 6616
rect 43625 6613 43637 6616
rect 43671 6644 43683 6647
rect 44910 6644 44916 6656
rect 43671 6616 44916 6644
rect 43671 6613 43683 6616
rect 43625 6607 43683 6613
rect 44910 6604 44916 6616
rect 44968 6604 44974 6656
rect 45462 6644 45468 6656
rect 45423 6616 45468 6644
rect 45462 6604 45468 6616
rect 45520 6604 45526 6656
rect 47302 6604 47308 6656
rect 47360 6604 47366 6656
rect 49694 6644 49700 6656
rect 49655 6616 49700 6644
rect 49694 6604 49700 6616
rect 49752 6604 49758 6656
rect 49804 6644 49832 6684
rect 52914 6672 52920 6684
rect 52972 6672 52978 6724
rect 54404 6712 54432 6743
rect 53576 6684 54432 6712
rect 53576 6656 53604 6684
rect 51626 6644 51632 6656
rect 49804 6616 51632 6644
rect 51626 6604 51632 6616
rect 51684 6604 51690 6656
rect 52089 6647 52147 6653
rect 52089 6613 52101 6647
rect 52135 6644 52147 6647
rect 53558 6644 53564 6656
rect 52135 6616 53564 6644
rect 52135 6613 52147 6616
rect 52089 6607 52147 6613
rect 53558 6604 53564 6616
rect 53616 6604 53622 6656
rect 54496 6644 54524 6820
rect 56410 6808 56416 6820
rect 56468 6808 56474 6860
rect 56502 6808 56508 6860
rect 56560 6848 56566 6860
rect 57977 6851 58035 6857
rect 57977 6848 57989 6851
rect 56560 6820 57989 6848
rect 56560 6808 56566 6820
rect 57977 6817 57989 6820
rect 58023 6817 58035 6851
rect 57977 6811 58035 6817
rect 60642 6808 60648 6860
rect 60700 6848 60706 6860
rect 60737 6851 60795 6857
rect 60737 6848 60749 6851
rect 60700 6820 60749 6848
rect 60700 6808 60706 6820
rect 60737 6817 60749 6820
rect 60783 6817 60795 6851
rect 60737 6811 60795 6817
rect 60918 6808 60924 6860
rect 60976 6848 60982 6860
rect 62040 6857 62068 6956
rect 64800 6916 64828 6956
rect 65150 6944 65156 6996
rect 65208 6984 65214 6996
rect 65245 6987 65303 6993
rect 65245 6984 65257 6987
rect 65208 6956 65257 6984
rect 65208 6944 65214 6956
rect 65245 6953 65257 6956
rect 65291 6953 65303 6987
rect 67818 6984 67824 6996
rect 65245 6947 65303 6953
rect 65352 6956 67824 6984
rect 65352 6916 65380 6956
rect 67818 6944 67824 6956
rect 67876 6944 67882 6996
rect 67931 6987 67989 6993
rect 67931 6953 67943 6987
rect 67977 6984 67989 6987
rect 68462 6984 68468 6996
rect 67977 6956 68468 6984
rect 67977 6953 67989 6956
rect 67931 6947 67989 6953
rect 68462 6944 68468 6956
rect 68520 6944 68526 6996
rect 68738 6944 68744 6996
rect 68796 6984 68802 6996
rect 72970 6984 72976 6996
rect 68796 6956 72976 6984
rect 68796 6944 68802 6956
rect 72970 6944 72976 6956
rect 73028 6944 73034 6996
rect 77938 6944 77944 6996
rect 77996 6984 78002 6996
rect 79962 6984 79968 6996
rect 77996 6956 79968 6984
rect 77996 6944 78002 6956
rect 79962 6944 79968 6956
rect 80020 6944 80026 6996
rect 80330 6944 80336 6996
rect 80388 6984 80394 6996
rect 81529 6987 81587 6993
rect 80388 6956 80652 6984
rect 80388 6944 80394 6956
rect 64800 6888 65380 6916
rect 68278 6876 68284 6928
rect 68336 6916 68342 6928
rect 69198 6916 69204 6928
rect 68336 6888 69204 6916
rect 68336 6876 68342 6888
rect 69198 6876 69204 6888
rect 69256 6876 69262 6928
rect 74169 6919 74227 6925
rect 74169 6885 74181 6919
rect 74215 6885 74227 6919
rect 77956 6916 77984 6944
rect 74169 6879 74227 6885
rect 74552 6888 74764 6916
rect 61841 6851 61899 6857
rect 61841 6848 61853 6851
rect 60976 6820 61853 6848
rect 60976 6808 60982 6820
rect 61841 6817 61853 6820
rect 61887 6817 61899 6851
rect 61841 6811 61899 6817
rect 62025 6851 62083 6857
rect 62025 6817 62037 6851
rect 62071 6817 62083 6851
rect 62025 6811 62083 6817
rect 62482 6808 62488 6860
rect 62540 6848 62546 6860
rect 62761 6851 62819 6857
rect 62761 6848 62773 6851
rect 62540 6820 62773 6848
rect 62540 6808 62546 6820
rect 62761 6817 62773 6820
rect 62807 6817 62819 6851
rect 62942 6848 62948 6860
rect 62903 6820 62948 6848
rect 62761 6811 62819 6817
rect 62942 6808 62948 6820
rect 63000 6808 63006 6860
rect 63218 6848 63224 6860
rect 63052 6820 63224 6848
rect 56321 6783 56379 6789
rect 56321 6749 56333 6783
rect 56367 6780 56379 6783
rect 57238 6780 57244 6792
rect 56367 6752 57244 6780
rect 56367 6749 56379 6752
rect 56321 6743 56379 6749
rect 57238 6740 57244 6752
rect 57296 6740 57302 6792
rect 59446 6740 59452 6792
rect 59504 6780 59510 6792
rect 59541 6783 59599 6789
rect 59541 6780 59553 6783
rect 59504 6752 59553 6780
rect 59504 6740 59510 6752
rect 59541 6749 59553 6752
rect 59587 6749 59599 6783
rect 59541 6743 59599 6749
rect 59817 6783 59875 6789
rect 59817 6749 59829 6783
rect 59863 6780 59875 6783
rect 59906 6780 59912 6792
rect 59863 6752 59912 6780
rect 59863 6749 59875 6752
rect 59817 6743 59875 6749
rect 59906 6740 59912 6752
rect 59964 6740 59970 6792
rect 59998 6740 60004 6792
rect 60056 6780 60062 6792
rect 60274 6780 60280 6792
rect 60056 6752 60280 6780
rect 60056 6740 60062 6752
rect 60274 6740 60280 6752
rect 60332 6740 60338 6792
rect 60826 6780 60832 6792
rect 60787 6752 60832 6780
rect 60826 6740 60832 6752
rect 60884 6740 60890 6792
rect 61010 6740 61016 6792
rect 61068 6780 61074 6792
rect 61654 6780 61660 6792
rect 61068 6752 61660 6780
rect 61068 6740 61074 6752
rect 61654 6740 61660 6752
rect 61712 6740 61718 6792
rect 61930 6780 61936 6792
rect 61891 6752 61936 6780
rect 61930 6740 61936 6752
rect 61988 6740 61994 6792
rect 62114 6740 62120 6792
rect 62172 6780 62178 6792
rect 62669 6783 62727 6789
rect 62172 6752 62217 6780
rect 62172 6740 62178 6752
rect 62669 6749 62681 6783
rect 62715 6780 62727 6783
rect 63052 6780 63080 6820
rect 63218 6808 63224 6820
rect 63276 6848 63282 6860
rect 65150 6848 65156 6860
rect 63276 6820 65156 6848
rect 63276 6808 63282 6820
rect 65150 6808 65156 6820
rect 65208 6808 65214 6860
rect 65426 6808 65432 6860
rect 65484 6848 65490 6860
rect 68646 6848 68652 6860
rect 65484 6820 68652 6848
rect 65484 6808 65490 6820
rect 68646 6808 68652 6820
rect 68704 6808 68710 6860
rect 69290 6848 69296 6860
rect 69251 6820 69296 6848
rect 69290 6808 69296 6820
rect 69348 6808 69354 6860
rect 71593 6851 71651 6857
rect 71593 6817 71605 6851
rect 71639 6848 71651 6851
rect 74184 6848 74212 6879
rect 71639 6820 74212 6848
rect 71639 6817 71651 6820
rect 71593 6811 71651 6817
rect 74350 6808 74356 6860
rect 74408 6848 74414 6860
rect 74552 6848 74580 6888
rect 74408 6820 74580 6848
rect 74629 6851 74687 6857
rect 74408 6808 74414 6820
rect 74629 6817 74641 6851
rect 74675 6817 74687 6851
rect 74736 6848 74764 6888
rect 75196 6888 75408 6916
rect 75196 6848 75224 6888
rect 74736 6820 75224 6848
rect 75273 6851 75331 6857
rect 74629 6811 74687 6817
rect 75273 6817 75285 6851
rect 75319 6817 75331 6851
rect 75380 6848 75408 6888
rect 76116 6888 77984 6916
rect 76116 6848 76144 6888
rect 78030 6876 78036 6928
rect 78088 6916 78094 6928
rect 80514 6916 80520 6928
rect 78088 6888 80520 6916
rect 78088 6876 78094 6888
rect 80514 6876 80520 6888
rect 80572 6876 80578 6928
rect 78858 6848 78864 6860
rect 75380 6820 76144 6848
rect 76208 6820 78864 6848
rect 75273 6811 75331 6817
rect 63494 6780 63500 6792
rect 62715 6752 63080 6780
rect 63455 6752 63500 6780
rect 62715 6749 62727 6752
rect 62669 6743 62727 6749
rect 63494 6740 63500 6752
rect 63552 6740 63558 6792
rect 64874 6740 64880 6792
rect 64932 6780 64938 6792
rect 66806 6780 66812 6792
rect 64932 6752 65564 6780
rect 64932 6740 64938 6752
rect 56962 6712 56968 6724
rect 56923 6684 56968 6712
rect 56962 6672 56968 6684
rect 57020 6672 57026 6724
rect 61102 6712 61108 6724
rect 57946 6684 61108 6712
rect 57425 6647 57483 6653
rect 57425 6644 57437 6647
rect 54496 6616 57437 6644
rect 57425 6613 57437 6616
rect 57471 6644 57483 6647
rect 57946 6644 57974 6684
rect 61102 6672 61108 6684
rect 61160 6672 61166 6724
rect 63773 6715 63831 6721
rect 63773 6712 63785 6715
rect 61212 6684 63785 6712
rect 57471 6616 57974 6644
rect 57471 6613 57483 6616
rect 57425 6607 57483 6613
rect 59538 6604 59544 6656
rect 59596 6644 59602 6656
rect 59633 6647 59691 6653
rect 59633 6644 59645 6647
rect 59596 6616 59645 6644
rect 59596 6604 59602 6616
rect 59633 6613 59645 6616
rect 59679 6613 59691 6647
rect 59998 6644 60004 6656
rect 59959 6616 60004 6644
rect 59633 6607 59691 6613
rect 59998 6604 60004 6616
rect 60056 6604 60062 6656
rect 61212 6653 61240 6684
rect 63773 6681 63785 6684
rect 63819 6681 63831 6715
rect 65426 6712 65432 6724
rect 63773 6675 63831 6681
rect 65168 6684 65432 6712
rect 61197 6647 61255 6653
rect 61197 6613 61209 6647
rect 61243 6613 61255 6647
rect 61654 6644 61660 6656
rect 61615 6616 61660 6644
rect 61197 6607 61255 6613
rect 61654 6604 61660 6616
rect 61712 6604 61718 6656
rect 62945 6647 63003 6653
rect 62945 6613 62957 6647
rect 62991 6644 63003 6647
rect 65168 6644 65196 6684
rect 65426 6672 65432 6684
rect 65484 6672 65490 6724
rect 65536 6712 65564 6752
rect 65812 6752 66812 6780
rect 65812 6712 65840 6752
rect 66806 6740 66812 6752
rect 66864 6740 66870 6792
rect 68186 6740 68192 6792
rect 68244 6780 68250 6792
rect 70302 6780 70308 6792
rect 68244 6752 70308 6780
rect 68244 6740 68250 6752
rect 70302 6740 70308 6752
rect 70360 6740 70366 6792
rect 71130 6740 71136 6792
rect 71188 6780 71194 6792
rect 71317 6783 71375 6789
rect 71317 6780 71329 6783
rect 71188 6752 71329 6780
rect 71188 6740 71194 6752
rect 71317 6749 71329 6752
rect 71363 6749 71375 6783
rect 74534 6780 74540 6792
rect 74447 6752 74540 6780
rect 71317 6743 71375 6749
rect 74534 6740 74540 6752
rect 74592 6740 74598 6792
rect 65536 6684 65840 6712
rect 66070 6672 66076 6724
rect 66128 6712 66134 6724
rect 66165 6715 66223 6721
rect 66165 6712 66177 6715
rect 66128 6684 66177 6712
rect 66128 6672 66134 6684
rect 66165 6681 66177 6684
rect 66211 6681 66223 6715
rect 69753 6715 69811 6721
rect 69753 6712 69765 6715
rect 66165 6675 66223 6681
rect 67560 6684 69765 6712
rect 62991 6616 65196 6644
rect 62991 6613 63003 6616
rect 62945 6607 63003 6613
rect 65242 6604 65248 6656
rect 65300 6644 65306 6656
rect 67560 6644 67588 6684
rect 69753 6681 69765 6684
rect 69799 6681 69811 6715
rect 71866 6712 71872 6724
rect 69753 6675 69811 6681
rect 69860 6684 71872 6712
rect 65300 6616 67588 6644
rect 65300 6604 65306 6616
rect 67634 6604 67640 6656
rect 67692 6644 67698 6656
rect 68741 6647 68799 6653
rect 68741 6644 68753 6647
rect 67692 6616 68753 6644
rect 67692 6604 67698 6616
rect 68741 6613 68753 6616
rect 68787 6644 68799 6647
rect 69860 6644 69888 6684
rect 71866 6672 71872 6684
rect 71924 6672 71930 6724
rect 72050 6672 72056 6724
rect 72108 6672 72114 6724
rect 73154 6672 73160 6724
rect 73212 6712 73218 6724
rect 73617 6715 73675 6721
rect 73617 6712 73629 6715
rect 73212 6684 73629 6712
rect 73212 6672 73218 6684
rect 73617 6681 73629 6684
rect 73663 6681 73675 6715
rect 73617 6675 73675 6681
rect 68787 6616 69888 6644
rect 68787 6613 68799 6616
rect 68741 6607 68799 6613
rect 70394 6604 70400 6656
rect 70452 6644 70458 6656
rect 70670 6644 70676 6656
rect 70452 6616 70676 6644
rect 70452 6604 70458 6616
rect 70670 6604 70676 6616
rect 70728 6604 70734 6656
rect 70762 6604 70768 6656
rect 70820 6644 70826 6656
rect 72418 6644 72424 6656
rect 70820 6616 72424 6644
rect 70820 6604 70826 6616
rect 72418 6604 72424 6616
rect 72476 6604 72482 6656
rect 73065 6647 73123 6653
rect 73065 6613 73077 6647
rect 73111 6644 73123 6647
rect 74552 6644 74580 6740
rect 74644 6712 74672 6811
rect 75178 6740 75184 6792
rect 75236 6780 75242 6792
rect 75288 6780 75316 6811
rect 75454 6780 75460 6792
rect 75236 6752 75316 6780
rect 75415 6752 75460 6780
rect 75236 6740 75242 6752
rect 75454 6740 75460 6752
rect 75512 6740 75518 6792
rect 76208 6789 76236 6820
rect 78858 6808 78864 6820
rect 78916 6808 78922 6860
rect 80422 6848 80428 6860
rect 80383 6820 80428 6848
rect 80422 6808 80428 6820
rect 80480 6808 80486 6860
rect 80624 6848 80652 6956
rect 81176 6956 81480 6984
rect 80701 6919 80759 6925
rect 80701 6885 80713 6919
rect 80747 6916 80759 6919
rect 81176 6916 81204 6956
rect 80747 6888 81204 6916
rect 80747 6885 80759 6888
rect 80701 6879 80759 6885
rect 81452 6848 81480 6956
rect 81529 6953 81541 6987
rect 81575 6984 81587 6987
rect 82630 6984 82636 6996
rect 81575 6956 82636 6984
rect 81575 6953 81587 6956
rect 81529 6947 81587 6953
rect 82630 6944 82636 6956
rect 82688 6944 82694 6996
rect 83642 6944 83648 6996
rect 83700 6984 83706 6996
rect 84010 6984 84016 6996
rect 83700 6956 84016 6984
rect 83700 6944 83706 6956
rect 84010 6944 84016 6956
rect 84068 6984 84074 6996
rect 84381 6987 84439 6993
rect 84381 6984 84393 6987
rect 84068 6956 84393 6984
rect 84068 6944 84074 6956
rect 84381 6953 84393 6956
rect 84427 6953 84439 6987
rect 84381 6947 84439 6953
rect 84470 6944 84476 6996
rect 84528 6984 84534 6996
rect 84749 6987 84807 6993
rect 84749 6984 84761 6987
rect 84528 6956 84761 6984
rect 84528 6944 84534 6956
rect 84749 6953 84761 6956
rect 84795 6953 84807 6987
rect 84749 6947 84807 6953
rect 88153 6987 88211 6993
rect 88153 6953 88165 6987
rect 88199 6984 88211 6987
rect 88426 6984 88432 6996
rect 88199 6956 88432 6984
rect 88199 6953 88211 6956
rect 88153 6947 88211 6953
rect 88426 6944 88432 6956
rect 88484 6944 88490 6996
rect 89714 6984 89720 6996
rect 88720 6956 89720 6984
rect 84102 6876 84108 6928
rect 84160 6916 84166 6928
rect 85022 6916 85028 6928
rect 84160 6888 85028 6916
rect 84160 6876 84166 6888
rect 85022 6876 85028 6888
rect 85080 6876 85086 6928
rect 87049 6919 87107 6925
rect 87049 6885 87061 6919
rect 87095 6916 87107 6919
rect 87138 6916 87144 6928
rect 87095 6888 87144 6916
rect 87095 6885 87107 6888
rect 87049 6879 87107 6885
rect 87138 6876 87144 6888
rect 87196 6916 87202 6928
rect 87966 6916 87972 6928
rect 87196 6888 87972 6916
rect 87196 6876 87202 6888
rect 87966 6876 87972 6888
rect 88024 6916 88030 6928
rect 88720 6916 88748 6956
rect 89714 6944 89720 6956
rect 89772 6984 89778 6996
rect 90174 6984 90180 6996
rect 89772 6956 90180 6984
rect 89772 6944 89778 6956
rect 90174 6944 90180 6956
rect 90232 6944 90238 6996
rect 92842 6944 92848 6996
rect 92900 6984 92906 6996
rect 93397 6987 93455 6993
rect 93397 6984 93409 6987
rect 92900 6956 93409 6984
rect 92900 6944 92906 6956
rect 93397 6953 93409 6956
rect 93443 6984 93455 6987
rect 93762 6984 93768 6996
rect 93443 6956 93768 6984
rect 93443 6953 93455 6956
rect 93397 6947 93455 6953
rect 93762 6944 93768 6956
rect 93820 6944 93826 6996
rect 88024 6888 88748 6916
rect 88024 6876 88030 6888
rect 82449 6851 82507 6857
rect 82449 6848 82461 6851
rect 80624 6820 81204 6848
rect 81452 6820 82461 6848
rect 81176 6814 81204 6820
rect 82449 6817 82461 6820
rect 82495 6817 82507 6851
rect 81176 6799 81296 6814
rect 82449 6811 82507 6817
rect 82538 6808 82544 6860
rect 82596 6848 82602 6860
rect 84473 6851 84531 6857
rect 84473 6848 84485 6851
rect 82596 6820 84485 6848
rect 82596 6808 82602 6820
rect 84473 6817 84485 6820
rect 84519 6848 84531 6851
rect 87230 6848 87236 6860
rect 84519 6820 87236 6848
rect 84519 6817 84531 6820
rect 84473 6811 84531 6817
rect 87230 6808 87236 6820
rect 87288 6808 87294 6860
rect 88242 6848 88248 6860
rect 87340 6820 88248 6848
rect 81176 6793 81311 6799
rect 75549 6783 75607 6789
rect 75549 6749 75561 6783
rect 75595 6780 75607 6783
rect 76193 6783 76251 6789
rect 76193 6780 76205 6783
rect 75595 6752 76205 6780
rect 75595 6749 75607 6752
rect 75549 6743 75607 6749
rect 76193 6749 76205 6752
rect 76239 6749 76251 6783
rect 76193 6743 76251 6749
rect 76377 6783 76435 6789
rect 76377 6749 76389 6783
rect 76423 6780 76435 6783
rect 76926 6780 76932 6792
rect 76423 6752 76932 6780
rect 76423 6749 76435 6752
rect 76377 6743 76435 6749
rect 75273 6715 75331 6721
rect 75273 6712 75285 6715
rect 74644 6684 75285 6712
rect 75273 6681 75285 6684
rect 75319 6681 75331 6715
rect 75273 6675 75331 6681
rect 75638 6672 75644 6724
rect 75696 6712 75702 6724
rect 76392 6712 76420 6743
rect 76926 6740 76932 6752
rect 76984 6740 76990 6792
rect 77294 6780 77300 6792
rect 77255 6752 77300 6780
rect 77294 6740 77300 6752
rect 77352 6740 77358 6792
rect 77754 6740 77760 6792
rect 77812 6780 77818 6792
rect 78309 6783 78367 6789
rect 78309 6780 78321 6783
rect 77812 6752 78321 6780
rect 77812 6740 77818 6752
rect 78309 6749 78321 6752
rect 78355 6749 78367 6783
rect 78309 6743 78367 6749
rect 78950 6740 78956 6792
rect 79008 6780 79014 6792
rect 79413 6783 79471 6789
rect 79413 6780 79425 6783
rect 79008 6752 79425 6780
rect 79008 6740 79014 6752
rect 79413 6749 79425 6752
rect 79459 6780 79471 6783
rect 79778 6780 79784 6792
rect 79459 6752 79784 6780
rect 79459 6749 79471 6752
rect 79413 6743 79471 6749
rect 79778 6740 79784 6752
rect 79836 6740 79842 6792
rect 80330 6780 80336 6792
rect 80291 6752 80336 6780
rect 80330 6740 80336 6752
rect 80388 6740 80394 6792
rect 81176 6786 81265 6793
rect 81253 6759 81265 6786
rect 81299 6759 81311 6793
rect 81618 6780 81624 6792
rect 81253 6753 81311 6759
rect 81579 6752 81624 6780
rect 81618 6740 81624 6752
rect 81676 6740 81682 6792
rect 82170 6780 82176 6792
rect 82131 6752 82176 6780
rect 82170 6740 82176 6752
rect 82228 6740 82234 6792
rect 84378 6780 84384 6792
rect 84339 6752 84384 6780
rect 84378 6740 84384 6752
rect 84436 6740 84442 6792
rect 84562 6740 84568 6792
rect 84620 6780 84626 6792
rect 85209 6783 85267 6789
rect 85209 6780 85221 6783
rect 84620 6752 85221 6780
rect 84620 6740 84626 6752
rect 85209 6749 85221 6752
rect 85255 6749 85267 6783
rect 85209 6743 85267 6749
rect 86678 6740 86684 6792
rect 86736 6780 86742 6792
rect 86865 6783 86923 6789
rect 86865 6780 86877 6783
rect 86736 6752 86877 6780
rect 86736 6740 86742 6752
rect 86865 6749 86877 6752
rect 86911 6749 86923 6783
rect 86865 6743 86923 6749
rect 86954 6740 86960 6792
rect 87012 6780 87018 6792
rect 87340 6780 87368 6820
rect 88242 6808 88248 6820
rect 88300 6808 88306 6860
rect 88720 6857 88748 6888
rect 89806 6876 89812 6928
rect 89864 6916 89870 6928
rect 89901 6919 89959 6925
rect 89901 6916 89913 6919
rect 89864 6888 89913 6916
rect 89864 6876 89870 6888
rect 89901 6885 89913 6888
rect 89947 6916 89959 6919
rect 90726 6916 90732 6928
rect 89947 6888 90732 6916
rect 89947 6885 89959 6888
rect 89901 6879 89959 6885
rect 90726 6876 90732 6888
rect 90784 6876 90790 6928
rect 88705 6851 88763 6857
rect 88705 6817 88717 6851
rect 88751 6817 88763 6851
rect 88705 6811 88763 6817
rect 89438 6808 89444 6860
rect 89496 6848 89502 6860
rect 90913 6851 90971 6857
rect 90913 6848 90925 6851
rect 89496 6820 90925 6848
rect 89496 6808 89502 6820
rect 90913 6817 90925 6820
rect 90959 6817 90971 6851
rect 92382 6848 92388 6860
rect 92343 6820 92388 6848
rect 90913 6811 90971 6817
rect 92382 6808 92388 6820
rect 92440 6808 92446 6860
rect 94038 6848 94044 6860
rect 92584 6820 94044 6848
rect 87012 6752 87368 6780
rect 87012 6740 87018 6752
rect 87414 6740 87420 6792
rect 87472 6780 87478 6792
rect 87969 6783 88027 6789
rect 87969 6780 87981 6783
rect 87472 6752 87981 6780
rect 87472 6740 87478 6752
rect 87969 6749 87981 6752
rect 88015 6749 88027 6783
rect 87969 6743 88027 6749
rect 88981 6783 89039 6789
rect 88981 6749 88993 6783
rect 89027 6780 89039 6783
rect 89070 6780 89076 6792
rect 89027 6752 89076 6780
rect 89027 6749 89039 6752
rect 88981 6743 89039 6749
rect 89070 6740 89076 6752
rect 89128 6740 89134 6792
rect 89622 6780 89628 6792
rect 89583 6752 89628 6780
rect 89622 6740 89628 6752
rect 89680 6740 89686 6792
rect 89898 6740 89904 6792
rect 89956 6780 89962 6792
rect 90453 6783 90511 6789
rect 90453 6780 90465 6783
rect 89956 6752 90465 6780
rect 89956 6740 89962 6752
rect 90453 6749 90465 6752
rect 90499 6780 90511 6783
rect 92584 6780 92612 6820
rect 94038 6808 94044 6820
rect 94096 6808 94102 6860
rect 90499 6752 92612 6780
rect 92661 6783 92719 6789
rect 90499 6749 90511 6752
rect 90453 6743 90511 6749
rect 92661 6749 92673 6783
rect 92707 6780 92719 6783
rect 93854 6780 93860 6792
rect 92707 6752 93860 6780
rect 92707 6749 92719 6752
rect 92661 6743 92719 6749
rect 93854 6740 93860 6752
rect 93912 6740 93918 6792
rect 76742 6712 76748 6724
rect 75696 6684 76420 6712
rect 76703 6684 76748 6712
rect 75696 6672 75702 6684
rect 76742 6672 76748 6684
rect 76800 6672 76806 6724
rect 78490 6672 78496 6724
rect 78548 6712 78554 6724
rect 78861 6715 78919 6721
rect 78861 6712 78873 6715
rect 78548 6684 78873 6712
rect 78548 6672 78554 6684
rect 78861 6681 78873 6684
rect 78907 6681 78919 6715
rect 78861 6675 78919 6681
rect 81345 6715 81403 6721
rect 81345 6681 81357 6715
rect 81391 6712 81403 6715
rect 81710 6712 81716 6724
rect 81391 6684 81716 6712
rect 81391 6681 81403 6684
rect 81345 6675 81403 6681
rect 81710 6672 81716 6684
rect 81768 6712 81774 6724
rect 83826 6712 83832 6724
rect 81768 6684 82768 6712
rect 83674 6684 83832 6712
rect 81768 6672 81774 6684
rect 73111 6616 74580 6644
rect 73111 6613 73123 6616
rect 73065 6607 73123 6613
rect 74626 6604 74632 6656
rect 74684 6644 74690 6656
rect 76466 6644 76472 6656
rect 74684 6616 76472 6644
rect 74684 6604 74690 6616
rect 76466 6604 76472 6616
rect 76524 6604 76530 6656
rect 76558 6604 76564 6656
rect 76616 6644 76622 6656
rect 76616 6616 76661 6644
rect 76616 6604 76622 6616
rect 76834 6604 76840 6656
rect 76892 6644 76898 6656
rect 77757 6647 77815 6653
rect 77757 6644 77769 6647
rect 76892 6616 77769 6644
rect 76892 6604 76898 6616
rect 77757 6613 77769 6616
rect 77803 6613 77815 6647
rect 77757 6607 77815 6613
rect 79870 6604 79876 6656
rect 79928 6644 79934 6656
rect 81437 6647 81495 6653
rect 81437 6644 81449 6647
rect 79928 6616 81449 6644
rect 79928 6604 79934 6616
rect 81437 6613 81449 6616
rect 81483 6644 81495 6647
rect 82538 6644 82544 6656
rect 81483 6616 82544 6644
rect 81483 6613 81495 6616
rect 81437 6607 81495 6613
rect 82538 6604 82544 6616
rect 82596 6604 82602 6656
rect 82740 6644 82768 6684
rect 83826 6672 83832 6684
rect 83884 6672 83890 6724
rect 84102 6672 84108 6724
rect 84160 6712 84166 6724
rect 88886 6712 88892 6724
rect 84160 6684 88892 6712
rect 84160 6672 84166 6684
rect 88886 6672 88892 6684
rect 88944 6672 88950 6724
rect 91833 6715 91891 6721
rect 91833 6712 91845 6715
rect 89824 6684 91845 6712
rect 83921 6647 83979 6653
rect 83921 6644 83933 6647
rect 82740 6616 83933 6644
rect 83921 6613 83933 6616
rect 83967 6644 83979 6647
rect 84010 6644 84016 6656
rect 83967 6616 84016 6644
rect 83967 6613 83979 6616
rect 83921 6607 83979 6613
rect 84010 6604 84016 6616
rect 84068 6604 84074 6656
rect 85853 6647 85911 6653
rect 85853 6613 85865 6647
rect 85899 6644 85911 6647
rect 86954 6644 86960 6656
rect 85899 6616 86960 6644
rect 85899 6613 85911 6616
rect 85853 6607 85911 6613
rect 86954 6604 86960 6616
rect 87012 6604 87018 6656
rect 87046 6604 87052 6656
rect 87104 6644 87110 6656
rect 89824 6644 89852 6684
rect 91833 6681 91845 6684
rect 91879 6681 91891 6715
rect 91833 6675 91891 6681
rect 93118 6672 93124 6724
rect 93176 6712 93182 6724
rect 93949 6715 94007 6721
rect 93949 6712 93961 6715
rect 93176 6684 93961 6712
rect 93176 6672 93182 6684
rect 93949 6681 93961 6684
rect 93995 6681 94007 6715
rect 93949 6675 94007 6681
rect 87104 6616 89852 6644
rect 87104 6604 87110 6616
rect 90726 6604 90732 6656
rect 90784 6644 90790 6656
rect 92750 6644 92756 6656
rect 90784 6616 92756 6644
rect 90784 6604 90790 6616
rect 92750 6604 92756 6616
rect 92808 6604 92814 6656
rect 1104 6554 95011 6576
rect 1104 6502 24386 6554
rect 24438 6502 24450 6554
rect 24502 6502 24514 6554
rect 24566 6502 24578 6554
rect 24630 6502 24642 6554
rect 24694 6502 47823 6554
rect 47875 6502 47887 6554
rect 47939 6502 47951 6554
rect 48003 6502 48015 6554
rect 48067 6502 48079 6554
rect 48131 6502 71260 6554
rect 71312 6502 71324 6554
rect 71376 6502 71388 6554
rect 71440 6502 71452 6554
rect 71504 6502 71516 6554
rect 71568 6502 94697 6554
rect 94749 6502 94761 6554
rect 94813 6502 94825 6554
rect 94877 6502 94889 6554
rect 94941 6502 94953 6554
rect 95005 6502 95011 6554
rect 1104 6480 95011 6502
rect 4246 6400 4252 6452
rect 4304 6440 4310 6452
rect 4709 6443 4767 6449
rect 4709 6440 4721 6443
rect 4304 6412 4721 6440
rect 4304 6400 4310 6412
rect 4709 6409 4721 6412
rect 4755 6440 4767 6443
rect 5074 6440 5080 6452
rect 4755 6412 5080 6440
rect 4755 6409 4767 6412
rect 4709 6403 4767 6409
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 5166 6400 5172 6452
rect 5224 6440 5230 6452
rect 10502 6440 10508 6452
rect 5224 6412 10508 6440
rect 5224 6400 5230 6412
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 15010 6440 15016 6452
rect 14971 6412 15016 6440
rect 15010 6400 15016 6412
rect 15068 6400 15074 6452
rect 17954 6440 17960 6452
rect 17915 6412 17960 6440
rect 17954 6400 17960 6412
rect 18012 6400 18018 6452
rect 19426 6440 19432 6452
rect 18708 6412 19432 6440
rect 5997 6375 6055 6381
rect 5997 6341 6009 6375
rect 6043 6372 6055 6375
rect 6638 6372 6644 6384
rect 6043 6344 6644 6372
rect 6043 6341 6055 6344
rect 5997 6335 6055 6341
rect 6638 6332 6644 6344
rect 6696 6372 6702 6384
rect 7558 6372 7564 6384
rect 6696 6344 7564 6372
rect 6696 6332 6702 6344
rect 6840 6313 6868 6344
rect 7558 6332 7564 6344
rect 7616 6372 7622 6384
rect 7616 6344 9996 6372
rect 7616 6332 7622 6344
rect 6825 6307 6883 6313
rect 6825 6273 6837 6307
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6304 7527 6307
rect 8110 6304 8116 6316
rect 7515 6276 8116 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 8386 6304 8392 6316
rect 8251 6276 8392 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 8386 6264 8392 6276
rect 8444 6264 8450 6316
rect 8496 6313 8524 6344
rect 8481 6307 8539 6313
rect 8481 6273 8493 6307
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6304 9275 6307
rect 9674 6304 9680 6316
rect 9263 6276 9680 6304
rect 9263 6273 9275 6276
rect 9217 6267 9275 6273
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 9858 6304 9864 6316
rect 9819 6276 9864 6304
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 9968 6304 9996 6344
rect 10134 6304 10140 6316
rect 9968 6276 10140 6304
rect 10134 6264 10140 6276
rect 10192 6304 10198 6316
rect 10192 6276 10548 6304
rect 10192 6264 10198 6276
rect 5718 6196 5724 6248
rect 5776 6236 5782 6248
rect 6549 6239 6607 6245
rect 6549 6236 6561 6239
rect 5776 6208 6561 6236
rect 5776 6196 5782 6208
rect 6549 6205 6561 6208
rect 6595 6205 6607 6239
rect 6549 6199 6607 6205
rect 10520 6168 10548 6276
rect 10594 6264 10600 6316
rect 10652 6304 10658 6316
rect 10778 6304 10784 6316
rect 10652 6276 10784 6304
rect 10652 6264 10658 6276
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 14277 6307 14335 6313
rect 14277 6273 14289 6307
rect 14323 6304 14335 6307
rect 14826 6304 14832 6316
rect 14323 6276 14832 6304
rect 14323 6273 14335 6276
rect 14277 6267 14335 6273
rect 14826 6264 14832 6276
rect 14884 6264 14890 6316
rect 18708 6313 18736 6412
rect 19426 6400 19432 6412
rect 19484 6400 19490 6452
rect 20530 6440 20536 6452
rect 20491 6412 20536 6440
rect 20530 6400 20536 6412
rect 20588 6400 20594 6452
rect 22186 6440 22192 6452
rect 21008 6412 22192 6440
rect 19242 6332 19248 6384
rect 19300 6372 19306 6384
rect 20898 6372 20904 6384
rect 19300 6344 20904 6372
rect 19300 6332 19306 6344
rect 20898 6332 20904 6344
rect 20956 6332 20962 6384
rect 18693 6307 18751 6313
rect 18693 6273 18705 6307
rect 18739 6273 18751 6307
rect 19521 6307 19579 6313
rect 19521 6304 19533 6307
rect 18693 6267 18751 6273
rect 19260 6276 19533 6304
rect 10686 6196 10692 6248
rect 10744 6236 10750 6248
rect 10744 6208 14412 6236
rect 10744 6196 10750 6208
rect 10778 6168 10784 6180
rect 10520 6140 10784 6168
rect 10778 6128 10784 6140
rect 10836 6168 10842 6180
rect 11701 6171 11759 6177
rect 11701 6168 11713 6171
rect 10836 6140 11713 6168
rect 10836 6128 10842 6140
rect 11701 6137 11713 6140
rect 11747 6168 11759 6171
rect 12618 6168 12624 6180
rect 11747 6140 12624 6168
rect 11747 6137 11759 6140
rect 11701 6131 11759 6137
rect 12618 6128 12624 6140
rect 12676 6128 12682 6180
rect 14384 6177 14412 6208
rect 17954 6196 17960 6248
rect 18012 6236 18018 6248
rect 18417 6239 18475 6245
rect 18417 6236 18429 6239
rect 18012 6208 18429 6236
rect 18012 6196 18018 6208
rect 18417 6205 18429 6208
rect 18463 6205 18475 6239
rect 18417 6199 18475 6205
rect 18601 6239 18659 6245
rect 18601 6205 18613 6239
rect 18647 6236 18659 6239
rect 19260 6236 19288 6276
rect 19521 6273 19533 6276
rect 19567 6304 19579 6307
rect 19702 6304 19708 6316
rect 19567 6276 19708 6304
rect 19567 6273 19579 6276
rect 19521 6267 19579 6273
rect 19702 6264 19708 6276
rect 19760 6264 19766 6316
rect 20349 6307 20407 6313
rect 20349 6304 20361 6307
rect 19904 6276 20361 6304
rect 18647 6208 19288 6236
rect 19337 6239 19395 6245
rect 18647 6205 18659 6208
rect 18601 6199 18659 6205
rect 19337 6205 19349 6239
rect 19383 6205 19395 6239
rect 19337 6199 19395 6205
rect 14369 6171 14427 6177
rect 14369 6137 14381 6171
rect 14415 6168 14427 6171
rect 19242 6168 19248 6180
rect 14415 6140 19248 6168
rect 14415 6137 14427 6140
rect 14369 6131 14427 6137
rect 19242 6128 19248 6140
rect 19300 6128 19306 6180
rect 19352 6168 19380 6199
rect 19904 6177 19932 6276
rect 20349 6273 20361 6276
rect 20395 6273 20407 6307
rect 20349 6267 20407 6273
rect 20438 6264 20444 6316
rect 20496 6304 20502 6316
rect 21008 6313 21036 6412
rect 22186 6400 22192 6412
rect 22244 6400 22250 6452
rect 22738 6400 22744 6452
rect 22796 6440 22802 6452
rect 26605 6443 26663 6449
rect 26605 6440 26617 6443
rect 22796 6412 26617 6440
rect 22796 6400 22802 6412
rect 22646 6332 22652 6384
rect 22704 6372 22710 6384
rect 22925 6375 22983 6381
rect 22925 6372 22937 6375
rect 22704 6344 22937 6372
rect 22704 6332 22710 6344
rect 22925 6341 22937 6344
rect 22971 6341 22983 6375
rect 22925 6335 22983 6341
rect 20533 6307 20591 6313
rect 20533 6304 20545 6307
rect 20496 6276 20545 6304
rect 20496 6264 20502 6276
rect 20533 6273 20545 6276
rect 20579 6304 20591 6307
rect 20993 6307 21051 6313
rect 20993 6304 21005 6307
rect 20579 6276 21005 6304
rect 20579 6273 20591 6276
rect 20533 6267 20591 6273
rect 20993 6273 21005 6276
rect 21039 6273 21051 6307
rect 20993 6267 21051 6273
rect 21174 6264 21180 6316
rect 21232 6304 21238 6316
rect 23198 6304 23204 6316
rect 21232 6276 23204 6304
rect 21232 6264 21238 6276
rect 23198 6264 23204 6276
rect 23256 6264 23262 6316
rect 23768 6313 23796 6412
rect 26605 6409 26617 6412
rect 26651 6440 26663 6443
rect 28166 6440 28172 6452
rect 26651 6412 28172 6440
rect 26651 6409 26663 6412
rect 26605 6403 26663 6409
rect 28166 6400 28172 6412
rect 28224 6400 28230 6452
rect 32306 6440 32312 6452
rect 28276 6412 32312 6440
rect 25222 6332 25228 6384
rect 25280 6372 25286 6384
rect 25590 6372 25596 6384
rect 25280 6344 25596 6372
rect 25280 6332 25286 6344
rect 25590 6332 25596 6344
rect 25648 6332 25654 6384
rect 26418 6332 26424 6384
rect 26476 6372 26482 6384
rect 28276 6372 28304 6412
rect 32306 6400 32312 6412
rect 32364 6400 32370 6452
rect 32401 6443 32459 6449
rect 32401 6409 32413 6443
rect 32447 6440 32459 6443
rect 33318 6440 33324 6452
rect 32447 6412 33324 6440
rect 32447 6409 32459 6412
rect 32401 6403 32459 6409
rect 33318 6400 33324 6412
rect 33376 6440 33382 6452
rect 39298 6440 39304 6452
rect 33376 6412 36308 6440
rect 39259 6412 39304 6440
rect 33376 6400 33382 6412
rect 26476 6344 28304 6372
rect 26476 6332 26482 6344
rect 29730 6332 29736 6384
rect 29788 6372 29794 6384
rect 33134 6372 33140 6384
rect 29788 6344 31754 6372
rect 33095 6344 33140 6372
rect 29788 6332 29794 6344
rect 23477 6307 23535 6313
rect 23477 6273 23489 6307
rect 23523 6273 23535 6307
rect 23477 6267 23535 6273
rect 23753 6307 23811 6313
rect 23753 6273 23765 6307
rect 23799 6273 23811 6307
rect 23753 6267 23811 6273
rect 23014 6196 23020 6248
rect 23072 6236 23078 6248
rect 23492 6236 23520 6267
rect 26510 6264 26516 6316
rect 26568 6304 26574 6316
rect 27525 6307 27583 6313
rect 27525 6304 27537 6307
rect 26568 6276 27537 6304
rect 26568 6264 26574 6276
rect 27525 6273 27537 6276
rect 27571 6273 27583 6307
rect 30101 6307 30159 6313
rect 27525 6267 27583 6273
rect 23072 6208 23520 6236
rect 23661 6239 23719 6245
rect 23072 6196 23078 6208
rect 23661 6205 23673 6239
rect 23707 6236 23719 6239
rect 24210 6236 24216 6248
rect 23707 6208 24216 6236
rect 23707 6205 23719 6208
rect 23661 6199 23719 6205
rect 24210 6196 24216 6208
rect 24268 6236 24274 6248
rect 24762 6236 24768 6248
rect 24268 6208 24768 6236
rect 24268 6196 24274 6208
rect 24762 6196 24768 6208
rect 24820 6196 24826 6248
rect 24857 6239 24915 6245
rect 24857 6205 24869 6239
rect 24903 6205 24915 6239
rect 25130 6236 25136 6248
rect 25091 6208 25136 6236
rect 24857 6199 24915 6205
rect 19889 6171 19947 6177
rect 19352 6140 19472 6168
rect 7745 6103 7803 6109
rect 7745 6069 7757 6103
rect 7791 6100 7803 6103
rect 8570 6100 8576 6112
rect 7791 6072 8576 6100
rect 7791 6069 7803 6072
rect 7745 6063 7803 6069
rect 8570 6060 8576 6072
rect 8628 6100 8634 6112
rect 9401 6103 9459 6109
rect 9401 6100 9413 6103
rect 8628 6072 9413 6100
rect 8628 6060 8634 6072
rect 9401 6069 9413 6072
rect 9447 6100 9459 6103
rect 10410 6100 10416 6112
rect 9447 6072 10416 6100
rect 9447 6069 9459 6072
rect 9401 6063 9459 6069
rect 10410 6060 10416 6072
rect 10468 6100 10474 6112
rect 11057 6103 11115 6109
rect 11057 6100 11069 6103
rect 10468 6072 11069 6100
rect 10468 6060 10474 6072
rect 11057 6069 11069 6072
rect 11103 6069 11115 6103
rect 18506 6100 18512 6112
rect 18467 6072 18512 6100
rect 11057 6063 11115 6069
rect 18506 6060 18512 6072
rect 18564 6060 18570 6112
rect 19444 6100 19472 6140
rect 19889 6137 19901 6171
rect 19935 6137 19947 6171
rect 22738 6168 22744 6180
rect 19889 6131 19947 6137
rect 19996 6140 22744 6168
rect 19610 6100 19616 6112
rect 19444 6072 19616 6100
rect 19610 6060 19616 6072
rect 19668 6100 19674 6112
rect 19996 6100 20024 6140
rect 22738 6128 22744 6140
rect 22796 6128 22802 6180
rect 19668 6072 20024 6100
rect 22465 6103 22523 6109
rect 19668 6060 19674 6072
rect 22465 6069 22477 6103
rect 22511 6100 22523 6103
rect 22830 6100 22836 6112
rect 22511 6072 22836 6100
rect 22511 6069 22523 6072
rect 22465 6063 22523 6069
rect 22830 6060 22836 6072
rect 22888 6060 22894 6112
rect 23750 6100 23756 6112
rect 23711 6072 23756 6100
rect 23750 6060 23756 6072
rect 23808 6060 23814 6112
rect 23937 6103 23995 6109
rect 23937 6069 23949 6103
rect 23983 6100 23995 6103
rect 24302 6100 24308 6112
rect 23983 6072 24308 6100
rect 23983 6069 23995 6072
rect 23937 6063 23995 6069
rect 24302 6060 24308 6072
rect 24360 6060 24366 6112
rect 24872 6100 24900 6199
rect 25130 6196 25136 6208
rect 25188 6196 25194 6248
rect 25866 6196 25872 6248
rect 25924 6236 25930 6248
rect 27433 6239 27491 6245
rect 27433 6236 27445 6239
rect 25924 6208 27445 6236
rect 25924 6196 25930 6208
rect 27433 6205 27445 6208
rect 27479 6205 27491 6239
rect 27433 6199 27491 6205
rect 26234 6128 26240 6180
rect 26292 6168 26298 6180
rect 27157 6171 27215 6177
rect 27157 6168 27169 6171
rect 26292 6140 27169 6168
rect 26292 6128 26298 6140
rect 27157 6137 27169 6140
rect 27203 6137 27215 6171
rect 28736 6168 28764 6290
rect 30101 6273 30113 6307
rect 30147 6304 30159 6307
rect 30190 6304 30196 6316
rect 30147 6276 30196 6304
rect 30147 6273 30159 6276
rect 30101 6267 30159 6273
rect 30190 6264 30196 6276
rect 30248 6264 30254 6316
rect 29825 6239 29883 6245
rect 29825 6205 29837 6239
rect 29871 6236 29883 6239
rect 30742 6236 30748 6248
rect 29871 6208 30748 6236
rect 29871 6205 29883 6208
rect 29825 6199 29883 6205
rect 30742 6196 30748 6208
rect 30800 6196 30806 6248
rect 31726 6236 31754 6344
rect 33134 6332 33140 6344
rect 33192 6332 33198 6384
rect 33226 6332 33232 6384
rect 33284 6372 33290 6384
rect 33594 6372 33600 6384
rect 33284 6344 33600 6372
rect 33284 6332 33290 6344
rect 33594 6332 33600 6344
rect 33652 6332 33658 6384
rect 34882 6372 34888 6384
rect 34843 6344 34888 6372
rect 34882 6332 34888 6344
rect 34940 6332 34946 6384
rect 32490 6264 32496 6316
rect 32548 6304 32554 6316
rect 32858 6304 32864 6316
rect 32548 6276 32864 6304
rect 32548 6264 32554 6276
rect 32858 6264 32864 6276
rect 32916 6264 32922 6316
rect 34698 6264 34704 6316
rect 34756 6304 34762 6316
rect 34756 6276 35756 6304
rect 34756 6264 34762 6276
rect 35618 6236 35624 6248
rect 31726 6208 35624 6236
rect 35618 6196 35624 6208
rect 35676 6196 35682 6248
rect 35728 6236 35756 6276
rect 35894 6264 35900 6316
rect 35952 6304 35958 6316
rect 36280 6313 36308 6412
rect 39298 6400 39304 6412
rect 39356 6400 39362 6452
rect 40218 6440 40224 6452
rect 40179 6412 40224 6440
rect 40218 6400 40224 6412
rect 40276 6400 40282 6452
rect 41230 6440 41236 6452
rect 40328 6412 41236 6440
rect 40328 6372 40356 6412
rect 41230 6400 41236 6412
rect 41288 6400 41294 6452
rect 43717 6443 43775 6449
rect 43717 6409 43729 6443
rect 43763 6440 43775 6443
rect 44726 6440 44732 6452
rect 43763 6412 44732 6440
rect 43763 6409 43775 6412
rect 43717 6403 43775 6409
rect 44726 6400 44732 6412
rect 44784 6400 44790 6452
rect 45186 6440 45192 6452
rect 45147 6412 45192 6440
rect 45186 6400 45192 6412
rect 45244 6400 45250 6452
rect 46382 6400 46388 6452
rect 46440 6440 46446 6452
rect 46937 6443 46995 6449
rect 46937 6440 46949 6443
rect 46440 6412 46949 6440
rect 46440 6400 46446 6412
rect 46937 6409 46949 6412
rect 46983 6440 46995 6443
rect 48130 6440 48136 6452
rect 46983 6412 48136 6440
rect 46983 6409 46995 6412
rect 46937 6403 46995 6409
rect 48130 6400 48136 6412
rect 48188 6400 48194 6452
rect 48682 6440 48688 6452
rect 48240 6412 48688 6440
rect 48038 6372 48044 6384
rect 39132 6344 40356 6372
rect 40880 6344 48044 6372
rect 35989 6307 36047 6313
rect 35989 6304 36001 6307
rect 35952 6276 36001 6304
rect 35952 6264 35958 6276
rect 35989 6273 36001 6276
rect 36035 6273 36047 6307
rect 35989 6267 36047 6273
rect 36265 6307 36323 6313
rect 36265 6273 36277 6307
rect 36311 6304 36323 6307
rect 38010 6304 38016 6316
rect 36311 6276 38016 6304
rect 36311 6273 36323 6276
rect 36265 6267 36323 6273
rect 38010 6264 38016 6276
rect 38068 6264 38074 6316
rect 38562 6264 38568 6316
rect 38620 6304 38626 6316
rect 39132 6313 39160 6344
rect 39117 6307 39175 6313
rect 39117 6304 39129 6307
rect 38620 6276 39129 6304
rect 38620 6264 38626 6276
rect 39117 6273 39129 6276
rect 39163 6273 39175 6307
rect 39117 6267 39175 6273
rect 39301 6307 39359 6313
rect 39301 6273 39313 6307
rect 39347 6273 39359 6307
rect 40126 6304 40132 6316
rect 40087 6276 40132 6304
rect 39301 6267 39359 6273
rect 37918 6236 37924 6248
rect 35728 6208 37924 6236
rect 37918 6196 37924 6208
rect 37976 6196 37982 6248
rect 39022 6196 39028 6248
rect 39080 6236 39086 6248
rect 39316 6236 39344 6267
rect 40126 6264 40132 6276
rect 40184 6264 40190 6316
rect 40310 6304 40316 6316
rect 40271 6276 40316 6304
rect 40310 6264 40316 6276
rect 40368 6264 40374 6316
rect 40880 6245 40908 6344
rect 48038 6332 48044 6344
rect 48096 6332 48102 6384
rect 40957 6307 41015 6313
rect 40957 6273 40969 6307
rect 41003 6273 41015 6307
rect 40957 6267 41015 6273
rect 42061 6307 42119 6313
rect 42061 6273 42073 6307
rect 42107 6304 42119 6307
rect 44174 6304 44180 6316
rect 42107 6276 44180 6304
rect 42107 6273 42119 6276
rect 42061 6267 42119 6273
rect 39080 6208 39344 6236
rect 39080 6196 39086 6208
rect 27157 6131 27215 6137
rect 27448 6140 28764 6168
rect 27448 6112 27476 6140
rect 30098 6128 30104 6180
rect 30156 6168 30162 6180
rect 32674 6168 32680 6180
rect 30156 6140 32680 6168
rect 30156 6128 30162 6140
rect 32674 6128 32680 6140
rect 32732 6128 32738 6180
rect 34238 6128 34244 6180
rect 34296 6168 34302 6180
rect 35342 6168 35348 6180
rect 34296 6140 35348 6168
rect 34296 6128 34302 6140
rect 35342 6128 35348 6140
rect 35400 6128 35406 6180
rect 39316 6168 39344 6208
rect 40865 6239 40923 6245
rect 40865 6205 40877 6239
rect 40911 6205 40923 6239
rect 40972 6236 41000 6267
rect 44174 6264 44180 6276
rect 44232 6264 44238 6316
rect 44542 6304 44548 6316
rect 44503 6276 44548 6304
rect 44542 6264 44548 6276
rect 44600 6264 44606 6316
rect 45554 6304 45560 6316
rect 45515 6276 45560 6304
rect 45554 6264 45560 6276
rect 45612 6264 45618 6316
rect 46198 6304 46204 6316
rect 46159 6276 46204 6304
rect 46198 6264 46204 6276
rect 46256 6264 46262 6316
rect 46385 6307 46443 6313
rect 46385 6273 46397 6307
rect 46431 6304 46443 6307
rect 48133 6307 48191 6313
rect 46431 6276 47992 6304
rect 46431 6273 46443 6276
rect 46385 6267 46443 6273
rect 43165 6239 43223 6245
rect 40972 6208 43116 6236
rect 40865 6199 40923 6205
rect 40954 6168 40960 6180
rect 39316 6140 40960 6168
rect 40954 6128 40960 6140
rect 41012 6128 41018 6180
rect 41325 6171 41383 6177
rect 41325 6137 41337 6171
rect 41371 6168 41383 6171
rect 42702 6168 42708 6180
rect 41371 6140 42708 6168
rect 41371 6137 41383 6140
rect 41325 6131 41383 6137
rect 42702 6128 42708 6140
rect 42760 6128 42766 6180
rect 43088 6168 43116 6208
rect 43165 6205 43177 6239
rect 43211 6236 43223 6239
rect 44082 6236 44088 6248
rect 43211 6208 44088 6236
rect 43211 6205 43223 6208
rect 43165 6199 43223 6205
rect 44082 6196 44088 6208
rect 44140 6196 44146 6248
rect 44637 6239 44695 6245
rect 44637 6205 44649 6239
rect 44683 6205 44695 6239
rect 45462 6236 45468 6248
rect 45423 6208 45468 6236
rect 44637 6199 44695 6205
rect 44652 6168 44680 6199
rect 45462 6196 45468 6208
rect 45520 6196 45526 6248
rect 46216 6236 46244 6264
rect 46934 6236 46940 6248
rect 46216 6208 46940 6236
rect 46934 6196 46940 6208
rect 46992 6196 46998 6248
rect 47964 6245 47992 6276
rect 48133 6273 48145 6307
rect 48179 6304 48191 6307
rect 48240 6304 48268 6412
rect 48682 6400 48688 6412
rect 48740 6400 48746 6452
rect 49510 6440 49516 6452
rect 48976 6412 49516 6440
rect 48314 6332 48320 6384
rect 48372 6372 48378 6384
rect 48976 6372 49004 6412
rect 49510 6400 49516 6412
rect 49568 6440 49574 6452
rect 49789 6443 49847 6449
rect 49789 6440 49801 6443
rect 49568 6412 49801 6440
rect 49568 6400 49574 6412
rect 49789 6409 49801 6412
rect 49835 6409 49847 6443
rect 49789 6403 49847 6409
rect 49973 6443 50031 6449
rect 49973 6409 49985 6443
rect 50019 6440 50031 6443
rect 50154 6440 50160 6452
rect 50019 6412 50160 6440
rect 50019 6409 50031 6412
rect 49973 6403 50031 6409
rect 50154 6400 50160 6412
rect 50212 6400 50218 6452
rect 52089 6443 52147 6449
rect 52089 6409 52101 6443
rect 52135 6440 52147 6443
rect 56134 6440 56140 6452
rect 52135 6412 54156 6440
rect 52135 6409 52147 6412
rect 52089 6403 52147 6409
rect 49878 6372 49884 6384
rect 48372 6344 49004 6372
rect 49839 6344 49884 6372
rect 48372 6332 48378 6344
rect 48179 6276 48268 6304
rect 48402 6307 48460 6313
rect 48179 6273 48191 6276
rect 48133 6267 48191 6273
rect 48402 6273 48414 6307
rect 48448 6304 48460 6307
rect 48516 6304 48636 6310
rect 48774 6304 48780 6316
rect 48448 6282 48780 6304
rect 48448 6276 48544 6282
rect 48608 6276 48780 6282
rect 48448 6273 48460 6276
rect 48402 6267 48460 6273
rect 48774 6264 48780 6276
rect 48832 6264 48838 6316
rect 48976 6313 49004 6344
rect 49878 6332 49884 6344
rect 49936 6372 49942 6384
rect 50617 6375 50675 6381
rect 50617 6372 50629 6375
rect 49936 6344 50629 6372
rect 49936 6332 49942 6344
rect 50617 6341 50629 6344
rect 50663 6341 50675 6375
rect 53834 6372 53840 6384
rect 53795 6344 53840 6372
rect 50617 6335 50675 6341
rect 53834 6332 53840 6344
rect 53892 6332 53898 6384
rect 49142 6313 49148 6316
rect 48961 6307 49019 6313
rect 48961 6273 48973 6307
rect 49007 6273 49019 6307
rect 48961 6267 49019 6273
rect 49139 6267 49148 6313
rect 49200 6304 49206 6316
rect 49200 6276 49239 6304
rect 49142 6264 49148 6267
rect 49200 6264 49206 6276
rect 50062 6264 50068 6316
rect 50120 6304 50126 6316
rect 51721 6307 51779 6313
rect 51721 6304 51733 6307
rect 50120 6276 51733 6304
rect 50120 6264 50126 6276
rect 51721 6273 51733 6276
rect 51767 6304 51779 6307
rect 52270 6304 52276 6316
rect 51767 6276 52276 6304
rect 51767 6273 51779 6276
rect 51721 6267 51779 6273
rect 52270 6264 52276 6276
rect 52328 6264 52334 6316
rect 47949 6239 48007 6245
rect 47949 6205 47961 6239
rect 47995 6205 48007 6239
rect 48222 6236 48228 6248
rect 48183 6208 48228 6236
rect 47949 6199 48007 6205
rect 48222 6196 48228 6208
rect 48280 6196 48286 6248
rect 48318 6239 48376 6245
rect 48318 6205 48330 6239
rect 48364 6224 48376 6239
rect 48364 6205 48445 6224
rect 48318 6199 48445 6205
rect 48332 6196 48445 6199
rect 51442 6196 51448 6248
rect 51500 6236 51506 6248
rect 51629 6239 51687 6245
rect 51629 6236 51641 6239
rect 51500 6208 51641 6236
rect 51500 6196 51506 6208
rect 51629 6205 51641 6208
rect 51675 6205 51687 6239
rect 53650 6236 53656 6248
rect 53611 6208 53656 6236
rect 51629 6199 51687 6205
rect 53650 6196 53656 6208
rect 53708 6196 53714 6248
rect 53926 6236 53932 6248
rect 53887 6208 53932 6236
rect 53926 6196 53932 6208
rect 53984 6196 53990 6248
rect 54128 6236 54156 6412
rect 54496 6412 56140 6440
rect 54496 6313 54524 6412
rect 56134 6400 56140 6412
rect 56192 6400 56198 6452
rect 58161 6443 58219 6449
rect 58161 6409 58173 6443
rect 58207 6440 58219 6443
rect 58250 6440 58256 6452
rect 58207 6412 58256 6440
rect 58207 6409 58219 6412
rect 58161 6403 58219 6409
rect 58250 6400 58256 6412
rect 58308 6440 58314 6452
rect 58986 6440 58992 6452
rect 58308 6412 58992 6440
rect 58308 6400 58314 6412
rect 58986 6400 58992 6412
rect 59044 6400 59050 6452
rect 59538 6440 59544 6452
rect 59499 6412 59544 6440
rect 59538 6400 59544 6412
rect 59596 6400 59602 6452
rect 60642 6440 60648 6452
rect 60603 6412 60648 6440
rect 60642 6400 60648 6412
rect 60700 6400 60706 6452
rect 62114 6400 62120 6452
rect 62172 6440 62178 6452
rect 64601 6443 64659 6449
rect 64601 6440 64613 6443
rect 62172 6412 64613 6440
rect 62172 6400 62178 6412
rect 64601 6409 64613 6412
rect 64647 6409 64659 6443
rect 64601 6403 64659 6409
rect 65337 6443 65395 6449
rect 65337 6409 65349 6443
rect 65383 6440 65395 6443
rect 65610 6440 65616 6452
rect 65383 6412 65616 6440
rect 65383 6409 65395 6412
rect 65337 6403 65395 6409
rect 65610 6400 65616 6412
rect 65668 6400 65674 6452
rect 65702 6400 65708 6452
rect 65760 6440 65766 6452
rect 67361 6443 67419 6449
rect 67361 6440 67373 6443
rect 65760 6412 67373 6440
rect 65760 6400 65766 6412
rect 67361 6409 67373 6412
rect 67407 6440 67419 6443
rect 67634 6440 67640 6452
rect 67407 6412 67640 6440
rect 67407 6409 67419 6412
rect 67361 6403 67419 6409
rect 67634 6400 67640 6412
rect 67692 6400 67698 6452
rect 68554 6440 68560 6452
rect 68515 6412 68560 6440
rect 68554 6400 68560 6412
rect 68612 6440 68618 6452
rect 71498 6440 71504 6452
rect 68612 6412 71504 6440
rect 68612 6400 68618 6412
rect 71498 6400 71504 6412
rect 71556 6400 71562 6452
rect 71593 6443 71651 6449
rect 71593 6409 71605 6443
rect 71639 6440 71651 6443
rect 72050 6440 72056 6452
rect 71639 6412 72056 6440
rect 71639 6409 71651 6412
rect 71593 6403 71651 6409
rect 72050 6400 72056 6412
rect 72108 6400 72114 6452
rect 72145 6443 72203 6449
rect 72145 6409 72157 6443
rect 72191 6409 72203 6443
rect 72145 6403 72203 6409
rect 74721 6443 74779 6449
rect 74721 6409 74733 6443
rect 74767 6440 74779 6443
rect 75362 6440 75368 6452
rect 74767 6412 75368 6440
rect 74767 6409 74779 6412
rect 74721 6403 74779 6409
rect 55030 6332 55036 6384
rect 55088 6372 55094 6384
rect 56505 6375 56563 6381
rect 55088 6344 55246 6372
rect 55088 6332 55094 6344
rect 56505 6341 56517 6375
rect 56551 6372 56563 6375
rect 58710 6372 58716 6384
rect 56551 6344 58020 6372
rect 58671 6344 58716 6372
rect 56551 6341 56563 6344
rect 56505 6335 56563 6341
rect 54481 6307 54539 6313
rect 54481 6273 54493 6307
rect 54527 6273 54539 6307
rect 54481 6267 54539 6273
rect 54757 6239 54815 6245
rect 54757 6236 54769 6239
rect 54128 6208 54769 6236
rect 54757 6205 54769 6208
rect 54803 6205 54815 6239
rect 54757 6199 54815 6205
rect 54846 6196 54852 6248
rect 54904 6236 54910 6248
rect 56520 6236 56548 6335
rect 56965 6307 57023 6313
rect 56965 6273 56977 6307
rect 57011 6273 57023 6307
rect 56965 6267 57023 6273
rect 57149 6307 57207 6313
rect 57149 6273 57161 6307
rect 57195 6304 57207 6307
rect 57882 6304 57888 6316
rect 57195 6276 57888 6304
rect 57195 6273 57207 6276
rect 57149 6267 57207 6273
rect 54904 6208 56548 6236
rect 56980 6236 57008 6267
rect 57882 6264 57888 6276
rect 57940 6264 57946 6316
rect 57698 6236 57704 6248
rect 56980 6208 57704 6236
rect 54904 6196 54910 6208
rect 57698 6196 57704 6208
rect 57756 6196 57762 6248
rect 57992 6236 58020 6344
rect 58710 6332 58716 6344
rect 58768 6332 58774 6384
rect 59170 6332 59176 6384
rect 59228 6372 59234 6384
rect 67450 6372 67456 6384
rect 59228 6344 67456 6372
rect 59228 6332 59234 6344
rect 67450 6332 67456 6344
rect 67508 6332 67514 6384
rect 67726 6332 67732 6384
rect 67784 6372 67790 6384
rect 70029 6375 70087 6381
rect 67784 6344 68862 6372
rect 67784 6332 67790 6344
rect 70029 6341 70041 6375
rect 70075 6372 70087 6375
rect 72160 6372 72188 6403
rect 75362 6400 75368 6412
rect 75420 6400 75426 6452
rect 75454 6400 75460 6452
rect 75512 6440 75518 6452
rect 76285 6443 76343 6449
rect 76285 6440 76297 6443
rect 75512 6412 76297 6440
rect 75512 6400 75518 6412
rect 76285 6409 76297 6412
rect 76331 6409 76343 6443
rect 76285 6403 76343 6409
rect 76374 6400 76380 6452
rect 76432 6440 76438 6452
rect 76432 6412 77340 6440
rect 76432 6400 76438 6412
rect 74626 6372 74632 6384
rect 70075 6344 72188 6372
rect 72528 6344 74632 6372
rect 70075 6341 70087 6344
rect 70029 6335 70087 6341
rect 58894 6264 58900 6316
rect 58952 6304 58958 6316
rect 59354 6304 59360 6316
rect 58952 6276 59360 6304
rect 58952 6264 58958 6276
rect 59354 6264 59360 6276
rect 59412 6264 59418 6316
rect 59541 6307 59599 6313
rect 59541 6273 59553 6307
rect 59587 6273 59599 6307
rect 60553 6307 60611 6313
rect 60553 6304 60565 6307
rect 59541 6267 59599 6273
rect 59924 6276 60565 6304
rect 59262 6236 59268 6248
rect 57992 6208 59268 6236
rect 59262 6196 59268 6208
rect 59320 6236 59326 6248
rect 59556 6236 59584 6267
rect 59320 6208 59584 6236
rect 59320 6196 59326 6208
rect 46293 6171 46351 6177
rect 46293 6168 46305 6171
rect 43088 6140 44588 6168
rect 44652 6140 46305 6168
rect 26694 6100 26700 6112
rect 24872 6072 26700 6100
rect 26694 6060 26700 6072
rect 26752 6060 26758 6112
rect 27430 6060 27436 6112
rect 27488 6060 27494 6112
rect 28353 6103 28411 6109
rect 28353 6069 28365 6103
rect 28399 6100 28411 6103
rect 28810 6100 28816 6112
rect 28399 6072 28816 6100
rect 28399 6069 28411 6072
rect 28353 6063 28411 6069
rect 28810 6060 28816 6072
rect 28868 6100 28874 6112
rect 33870 6100 33876 6112
rect 28868 6072 33876 6100
rect 28868 6060 28874 6072
rect 33870 6060 33876 6072
rect 33928 6060 33934 6112
rect 34146 6060 34152 6112
rect 34204 6100 34210 6112
rect 37645 6103 37703 6109
rect 37645 6100 37657 6103
rect 34204 6072 37657 6100
rect 34204 6060 34210 6072
rect 37645 6069 37657 6072
rect 37691 6069 37703 6103
rect 44266 6100 44272 6112
rect 44227 6072 44272 6100
rect 37645 6063 37703 6069
rect 44266 6060 44272 6072
rect 44324 6060 44330 6112
rect 44560 6100 44588 6140
rect 46293 6137 46305 6140
rect 46339 6137 46351 6171
rect 48417 6168 48445 6196
rect 49602 6168 49608 6180
rect 48417 6140 49608 6168
rect 46293 6131 46351 6137
rect 49602 6128 49608 6140
rect 49660 6128 49666 6180
rect 50893 6171 50951 6177
rect 50893 6168 50905 6171
rect 49712 6140 50905 6168
rect 45738 6100 45744 6112
rect 44560 6072 45744 6100
rect 45738 6060 45744 6072
rect 45796 6060 45802 6112
rect 46934 6060 46940 6112
rect 46992 6100 46998 6112
rect 48314 6100 48320 6112
rect 46992 6072 48320 6100
rect 46992 6060 46998 6072
rect 48314 6060 48320 6072
rect 48372 6060 48378 6112
rect 48774 6060 48780 6112
rect 48832 6100 48838 6112
rect 49145 6103 49203 6109
rect 49145 6100 49157 6103
rect 48832 6072 49157 6100
rect 48832 6060 48838 6072
rect 49145 6069 49157 6072
rect 49191 6100 49203 6103
rect 49712 6100 49740 6140
rect 50893 6137 50905 6140
rect 50939 6137 50951 6171
rect 50893 6131 50951 6137
rect 49191 6072 49740 6100
rect 50157 6103 50215 6109
rect 49191 6069 49203 6072
rect 49145 6063 49203 6069
rect 50157 6069 50169 6103
rect 50203 6100 50215 6103
rect 50706 6100 50712 6112
rect 50203 6072 50712 6100
rect 50203 6069 50215 6072
rect 50157 6063 50215 6069
rect 50706 6060 50712 6072
rect 50764 6060 50770 6112
rect 51077 6103 51135 6109
rect 51077 6069 51089 6103
rect 51123 6100 51135 6103
rect 51350 6100 51356 6112
rect 51123 6072 51356 6100
rect 51123 6069 51135 6072
rect 51077 6063 51135 6069
rect 51350 6060 51356 6072
rect 51408 6060 51414 6112
rect 56962 6060 56968 6112
rect 57020 6100 57026 6112
rect 57057 6103 57115 6109
rect 57057 6100 57069 6103
rect 57020 6072 57069 6100
rect 57020 6060 57026 6072
rect 57057 6069 57069 6072
rect 57103 6069 57115 6103
rect 57057 6063 57115 6069
rect 57146 6060 57152 6112
rect 57204 6100 57210 6112
rect 59924 6100 59952 6276
rect 60553 6273 60565 6276
rect 60599 6273 60611 6307
rect 60553 6267 60611 6273
rect 60737 6307 60795 6313
rect 60737 6273 60749 6307
rect 60783 6304 60795 6307
rect 61654 6304 61660 6316
rect 60783 6276 61660 6304
rect 60783 6273 60795 6276
rect 60737 6267 60795 6273
rect 61654 6264 61660 6276
rect 61712 6264 61718 6316
rect 61841 6307 61899 6313
rect 61841 6273 61853 6307
rect 61887 6304 61899 6307
rect 61930 6304 61936 6316
rect 61887 6276 61936 6304
rect 61887 6273 61899 6276
rect 61841 6267 61899 6273
rect 61930 6264 61936 6276
rect 61988 6304 61994 6316
rect 63586 6304 63592 6316
rect 61988 6276 63592 6304
rect 61988 6264 61994 6276
rect 63586 6264 63592 6276
rect 63644 6264 63650 6316
rect 63770 6304 63776 6316
rect 63731 6276 63776 6304
rect 63770 6264 63776 6276
rect 63828 6264 63834 6316
rect 64506 6304 64512 6316
rect 64467 6276 64512 6304
rect 64506 6264 64512 6276
rect 64564 6264 64570 6316
rect 64690 6304 64696 6316
rect 64651 6276 64696 6304
rect 64690 6264 64696 6276
rect 64748 6264 64754 6316
rect 65150 6304 65156 6316
rect 65111 6276 65156 6304
rect 65150 6264 65156 6276
rect 65208 6264 65214 6316
rect 65334 6304 65340 6316
rect 65295 6276 65340 6304
rect 65334 6264 65340 6276
rect 65392 6304 65398 6316
rect 66070 6304 66076 6316
rect 65392 6276 66076 6304
rect 65392 6264 65398 6276
rect 66070 6264 66076 6276
rect 66128 6304 66134 6316
rect 66717 6307 66775 6313
rect 66128 6276 66576 6304
rect 66128 6264 66134 6276
rect 59998 6196 60004 6248
rect 60056 6236 60062 6248
rect 61749 6239 61807 6245
rect 61749 6236 61761 6239
rect 60056 6208 61761 6236
rect 60056 6196 60062 6208
rect 61749 6205 61761 6208
rect 61795 6205 61807 6239
rect 66162 6236 66168 6248
rect 61749 6199 61807 6205
rect 61856 6208 66168 6236
rect 60093 6171 60151 6177
rect 60093 6137 60105 6171
rect 60139 6168 60151 6171
rect 61010 6168 61016 6180
rect 60139 6140 61016 6168
rect 60139 6137 60151 6140
rect 60093 6131 60151 6137
rect 61010 6128 61016 6140
rect 61068 6128 61074 6180
rect 61102 6128 61108 6180
rect 61160 6168 61166 6180
rect 61856 6168 61884 6208
rect 66162 6196 66168 6208
rect 66220 6196 66226 6248
rect 64598 6168 64604 6180
rect 61160 6140 61884 6168
rect 61948 6140 64604 6168
rect 61160 6128 61166 6140
rect 61948 6100 61976 6140
rect 64598 6128 64604 6140
rect 64656 6128 64662 6180
rect 62114 6100 62120 6112
rect 57204 6072 61976 6100
rect 62075 6072 62120 6100
rect 57204 6060 57210 6072
rect 62114 6060 62120 6072
rect 62172 6060 62178 6112
rect 63310 6100 63316 6112
rect 63271 6072 63316 6100
rect 63310 6060 63316 6072
rect 63368 6060 63374 6112
rect 63494 6060 63500 6112
rect 63552 6100 63558 6112
rect 63957 6103 64015 6109
rect 63957 6100 63969 6103
rect 63552 6072 63969 6100
rect 63552 6060 63558 6072
rect 63957 6069 63969 6072
rect 64003 6100 64015 6103
rect 65242 6100 65248 6112
rect 64003 6072 65248 6100
rect 64003 6069 64015 6072
rect 63957 6063 64015 6069
rect 65242 6060 65248 6072
rect 65300 6060 65306 6112
rect 65886 6100 65892 6112
rect 65847 6072 65892 6100
rect 65886 6060 65892 6072
rect 65944 6060 65950 6112
rect 66070 6060 66076 6112
rect 66128 6100 66134 6112
rect 66441 6103 66499 6109
rect 66441 6100 66453 6103
rect 66128 6072 66453 6100
rect 66128 6060 66134 6072
rect 66441 6069 66453 6072
rect 66487 6069 66499 6103
rect 66548 6100 66576 6276
rect 66717 6273 66729 6307
rect 66763 6304 66775 6307
rect 67542 6304 67548 6316
rect 66763 6276 67548 6304
rect 66763 6273 66775 6276
rect 66717 6267 66775 6273
rect 67542 6264 67548 6276
rect 67600 6264 67606 6316
rect 70302 6264 70308 6316
rect 70360 6304 70366 6316
rect 70762 6304 70768 6316
rect 70360 6276 70768 6304
rect 70360 6264 70366 6276
rect 70762 6264 70768 6276
rect 70820 6264 70826 6316
rect 71406 6304 71412 6316
rect 71367 6276 71412 6304
rect 71406 6264 71412 6276
rect 71464 6264 71470 6316
rect 71682 6304 71688 6316
rect 71643 6276 71688 6304
rect 71682 6264 71688 6276
rect 71740 6264 71746 6316
rect 72528 6313 72556 6344
rect 74626 6332 74632 6344
rect 74684 6332 74690 6384
rect 76006 6372 76012 6384
rect 74828 6344 76012 6372
rect 72513 6307 72571 6313
rect 72513 6273 72525 6307
rect 72559 6273 72571 6307
rect 73522 6304 73528 6316
rect 73483 6276 73528 6304
rect 72513 6267 72571 6273
rect 66809 6239 66867 6245
rect 66809 6205 66821 6239
rect 66855 6236 66867 6239
rect 66855 6208 70256 6236
rect 66855 6205 66867 6208
rect 66809 6199 66867 6205
rect 66622 6128 66628 6180
rect 66680 6168 66686 6180
rect 70228 6168 70256 6208
rect 71498 6196 71504 6248
rect 71556 6236 71562 6248
rect 72528 6236 72556 6267
rect 73522 6264 73528 6276
rect 73580 6264 73586 6316
rect 73709 6307 73767 6313
rect 73709 6273 73721 6307
rect 73755 6273 73767 6307
rect 73709 6267 73767 6273
rect 71556 6208 72556 6236
rect 72605 6239 72663 6245
rect 71556 6196 71562 6208
rect 72605 6205 72617 6239
rect 72651 6236 72663 6239
rect 73617 6239 73675 6245
rect 73617 6236 73629 6239
rect 72651 6208 73629 6236
rect 72651 6205 72663 6208
rect 72605 6199 72663 6205
rect 73617 6205 73629 6208
rect 73663 6205 73675 6239
rect 73724 6236 73752 6267
rect 74350 6264 74356 6316
rect 74408 6304 74414 6316
rect 74828 6313 74856 6344
rect 76006 6332 76012 6344
rect 76064 6372 76070 6384
rect 77312 6372 77340 6412
rect 77386 6400 77392 6452
rect 77444 6440 77450 6452
rect 83182 6440 83188 6452
rect 77444 6412 83188 6440
rect 77444 6400 77450 6412
rect 83182 6400 83188 6412
rect 83240 6400 83246 6452
rect 83277 6443 83335 6449
rect 83277 6409 83289 6443
rect 83323 6440 83335 6443
rect 94130 6440 94136 6452
rect 83323 6412 90588 6440
rect 94091 6412 94136 6440
rect 83323 6409 83335 6412
rect 83277 6403 83335 6409
rect 78766 6372 78772 6384
rect 76064 6344 77248 6372
rect 77312 6344 77524 6372
rect 78727 6344 78772 6372
rect 76064 6332 76070 6344
rect 74537 6307 74595 6313
rect 74537 6304 74549 6307
rect 74408 6276 74549 6304
rect 74408 6264 74414 6276
rect 74537 6273 74549 6276
rect 74583 6273 74595 6307
rect 74537 6267 74595 6273
rect 74813 6307 74871 6313
rect 74813 6273 74825 6307
rect 74859 6273 74871 6307
rect 74813 6267 74871 6273
rect 74994 6264 75000 6316
rect 75052 6304 75058 6316
rect 77220 6313 77248 6344
rect 75549 6307 75607 6313
rect 75549 6304 75561 6307
rect 75052 6276 75561 6304
rect 75052 6264 75058 6276
rect 75549 6273 75561 6276
rect 75595 6273 75607 6307
rect 75549 6267 75607 6273
rect 77205 6307 77263 6313
rect 77205 6273 77217 6307
rect 77251 6273 77263 6307
rect 77205 6267 77263 6273
rect 77389 6307 77447 6313
rect 77389 6273 77401 6307
rect 77435 6273 77447 6307
rect 77496 6304 77524 6344
rect 78766 6332 78772 6344
rect 78824 6332 78830 6384
rect 79226 6372 79232 6384
rect 79187 6344 79232 6372
rect 79226 6332 79232 6344
rect 79284 6332 79290 6384
rect 79686 6332 79692 6384
rect 79744 6372 79750 6384
rect 80698 6372 80704 6384
rect 79744 6344 80704 6372
rect 79744 6332 79750 6344
rect 80698 6332 80704 6344
rect 80756 6332 80762 6384
rect 84102 6372 84108 6384
rect 83384 6344 84108 6372
rect 83384 6316 83412 6344
rect 84102 6332 84108 6344
rect 84160 6332 84166 6384
rect 87046 6372 87052 6384
rect 84672 6344 87052 6372
rect 79965 6307 80023 6313
rect 79965 6304 79977 6307
rect 77496 6276 79977 6304
rect 77389 6267 77447 6273
rect 79965 6273 79977 6276
rect 80011 6273 80023 6307
rect 79965 6267 80023 6273
rect 82909 6307 82967 6313
rect 82909 6273 82921 6307
rect 82955 6304 82967 6307
rect 83366 6304 83372 6316
rect 82955 6276 83372 6304
rect 82955 6273 82967 6276
rect 82909 6267 82967 6273
rect 75273 6239 75331 6245
rect 75273 6236 75285 6239
rect 73724 6208 75285 6236
rect 73617 6199 73675 6205
rect 75273 6205 75285 6208
rect 75319 6205 75331 6239
rect 75454 6236 75460 6248
rect 75415 6208 75460 6236
rect 75273 6199 75331 6205
rect 75454 6196 75460 6208
rect 75512 6196 75518 6248
rect 75632 6239 75690 6245
rect 75632 6236 75644 6239
rect 75564 6208 75644 6236
rect 74353 6171 74411 6177
rect 74353 6168 74365 6171
rect 66680 6140 68232 6168
rect 70228 6140 74365 6168
rect 66680 6128 66686 6140
rect 68094 6100 68100 6112
rect 66548 6072 68100 6100
rect 66441 6063 66499 6069
rect 68094 6060 68100 6072
rect 68152 6060 68158 6112
rect 68204 6100 68232 6140
rect 74353 6137 74365 6140
rect 74399 6137 74411 6171
rect 74353 6131 74411 6137
rect 70394 6100 70400 6112
rect 68204 6072 70400 6100
rect 70394 6060 70400 6072
rect 70452 6060 70458 6112
rect 71225 6103 71283 6109
rect 71225 6069 71237 6103
rect 71271 6100 71283 6103
rect 72142 6100 72148 6112
rect 71271 6072 72148 6100
rect 71271 6069 71283 6072
rect 71225 6063 71283 6069
rect 72142 6060 72148 6072
rect 72200 6060 72206 6112
rect 73522 6060 73528 6112
rect 73580 6100 73586 6112
rect 73982 6100 73988 6112
rect 73580 6072 73988 6100
rect 73580 6060 73586 6072
rect 73982 6060 73988 6072
rect 74040 6060 74046 6112
rect 75454 6060 75460 6112
rect 75512 6100 75518 6112
rect 75564 6100 75592 6208
rect 75632 6205 75644 6208
rect 75678 6205 75690 6239
rect 75632 6199 75690 6205
rect 75733 6239 75791 6245
rect 75733 6205 75745 6239
rect 75779 6236 75791 6239
rect 75779 6208 76420 6236
rect 75779 6205 75791 6208
rect 75733 6199 75791 6205
rect 76392 6177 76420 6208
rect 76558 6196 76564 6248
rect 76616 6236 76622 6248
rect 76745 6239 76803 6245
rect 76745 6236 76757 6239
rect 76616 6208 76757 6236
rect 76616 6196 76622 6208
rect 76745 6205 76757 6208
rect 76791 6205 76803 6239
rect 76745 6199 76803 6205
rect 76377 6171 76435 6177
rect 76377 6137 76389 6171
rect 76423 6168 76435 6171
rect 77205 6171 77263 6177
rect 77205 6168 77217 6171
rect 76423 6140 77217 6168
rect 76423 6137 76435 6140
rect 76377 6131 76435 6137
rect 77205 6137 77217 6140
rect 77251 6137 77263 6171
rect 77205 6131 77263 6137
rect 75512 6072 75592 6100
rect 75512 6060 75518 6072
rect 76650 6060 76656 6112
rect 76708 6100 76714 6112
rect 77404 6100 77432 6267
rect 83366 6264 83372 6276
rect 83424 6264 83430 6316
rect 83734 6264 83740 6316
rect 83792 6304 83798 6316
rect 83921 6307 83979 6313
rect 83921 6304 83933 6307
rect 83792 6276 83933 6304
rect 83792 6264 83798 6276
rect 83921 6273 83933 6276
rect 83967 6273 83979 6307
rect 83921 6267 83979 6273
rect 80238 6236 80244 6248
rect 80199 6208 80244 6236
rect 80238 6196 80244 6208
rect 80296 6196 80302 6248
rect 81250 6196 81256 6248
rect 81308 6236 81314 6248
rect 81618 6236 81624 6248
rect 81308 6208 81624 6236
rect 81308 6196 81314 6208
rect 81618 6196 81624 6208
rect 81676 6196 81682 6248
rect 81986 6236 81992 6248
rect 81947 6208 81992 6236
rect 81986 6196 81992 6208
rect 82044 6196 82050 6248
rect 82814 6236 82820 6248
rect 82775 6208 82820 6236
rect 82814 6196 82820 6208
rect 82872 6196 82878 6248
rect 78582 6128 78588 6180
rect 78640 6168 78646 6180
rect 84672 6168 84700 6344
rect 87046 6332 87052 6344
rect 87104 6332 87110 6384
rect 90560 6381 90588 6412
rect 94130 6400 94136 6412
rect 94188 6400 94194 6452
rect 90545 6375 90603 6381
rect 90545 6341 90557 6375
rect 90591 6341 90603 6375
rect 90545 6335 90603 6341
rect 91830 6332 91836 6384
rect 91888 6372 91894 6384
rect 91888 6344 92428 6372
rect 91888 6332 91894 6344
rect 84746 6264 84752 6316
rect 84804 6304 84810 6316
rect 85022 6304 85028 6316
rect 84804 6276 84849 6304
rect 84983 6276 85028 6304
rect 84804 6264 84810 6276
rect 85022 6264 85028 6276
rect 85080 6304 85086 6316
rect 85482 6304 85488 6316
rect 85080 6276 85488 6304
rect 85080 6264 85086 6276
rect 85482 6264 85488 6276
rect 85540 6304 85546 6316
rect 85758 6304 85764 6316
rect 85540 6276 85620 6304
rect 85719 6276 85764 6304
rect 85540 6264 85546 6276
rect 85592 6236 85620 6276
rect 85758 6264 85764 6276
rect 85816 6264 85822 6316
rect 86512 6304 86632 6314
rect 86668 6307 86726 6313
rect 86668 6304 86680 6307
rect 86052 6286 86680 6304
rect 86052 6276 86540 6286
rect 86604 6276 86680 6286
rect 86052 6236 86080 6276
rect 86668 6273 86680 6276
rect 86714 6273 86726 6307
rect 86668 6267 86726 6273
rect 86862 6264 86868 6316
rect 86920 6304 86926 6316
rect 87414 6304 87420 6316
rect 86920 6276 87420 6304
rect 86920 6264 86926 6276
rect 87414 6264 87420 6276
rect 87472 6264 87478 6316
rect 88337 6307 88395 6313
rect 88337 6273 88349 6307
rect 88383 6304 88395 6307
rect 88426 6304 88432 6316
rect 88383 6276 88432 6304
rect 88383 6273 88395 6276
rect 88337 6267 88395 6273
rect 88426 6264 88432 6276
rect 88484 6264 88490 6316
rect 85592 6208 86080 6236
rect 86126 6196 86132 6248
rect 86184 6236 86190 6248
rect 86405 6239 86463 6245
rect 86405 6236 86417 6239
rect 86184 6208 86417 6236
rect 86184 6196 86190 6208
rect 86405 6205 86417 6208
rect 86451 6205 86463 6239
rect 86405 6199 86463 6205
rect 88886 6196 88892 6248
rect 88944 6236 88950 6248
rect 89073 6239 89131 6245
rect 89073 6236 89085 6239
rect 88944 6208 89085 6236
rect 88944 6196 88950 6208
rect 89073 6205 89085 6208
rect 89119 6205 89131 6239
rect 89073 6199 89131 6205
rect 89456 6236 89484 6290
rect 90818 6264 90824 6316
rect 90876 6304 90882 6316
rect 90876 6276 90921 6304
rect 90876 6264 90882 6276
rect 91278 6264 91284 6316
rect 91336 6304 91342 6316
rect 92400 6313 92428 6344
rect 92109 6307 92167 6313
rect 92109 6304 92121 6307
rect 91336 6276 92121 6304
rect 91336 6264 91342 6276
rect 92109 6273 92121 6276
rect 92155 6273 92167 6307
rect 92109 6267 92167 6273
rect 92385 6307 92443 6313
rect 92385 6273 92397 6307
rect 92431 6273 92443 6307
rect 93026 6304 93032 6316
rect 92987 6276 93032 6304
rect 92385 6267 92443 6273
rect 93026 6264 93032 6276
rect 93084 6264 93090 6316
rect 89898 6236 89904 6248
rect 89456 6208 89904 6236
rect 89456 6168 89484 6208
rect 89898 6196 89904 6208
rect 89956 6196 89962 6248
rect 78640 6140 80054 6168
rect 78640 6128 78646 6140
rect 77846 6100 77852 6112
rect 76708 6072 77432 6100
rect 77807 6072 77852 6100
rect 76708 6060 76714 6072
rect 77846 6060 77852 6072
rect 77904 6060 77910 6112
rect 80026 6100 80054 6140
rect 81268 6140 84700 6168
rect 88168 6140 89484 6168
rect 81268 6100 81296 6140
rect 80026 6072 81296 6100
rect 81526 6060 81532 6112
rect 81584 6100 81590 6112
rect 83458 6100 83464 6112
rect 81584 6072 83464 6100
rect 81584 6060 81590 6072
rect 83458 6060 83464 6072
rect 83516 6060 83522 6112
rect 83826 6060 83832 6112
rect 83884 6100 83890 6112
rect 84013 6103 84071 6109
rect 84013 6100 84025 6103
rect 83884 6072 84025 6100
rect 83884 6060 83890 6072
rect 84013 6069 84025 6072
rect 84059 6100 84071 6103
rect 84378 6100 84384 6112
rect 84059 6072 84384 6100
rect 84059 6069 84071 6072
rect 84013 6063 84071 6069
rect 84378 6060 84384 6072
rect 84436 6100 84442 6112
rect 85758 6100 85764 6112
rect 84436 6072 85764 6100
rect 84436 6060 84442 6072
rect 85758 6060 85764 6072
rect 85816 6060 85822 6112
rect 85945 6103 86003 6109
rect 85945 6069 85957 6103
rect 85991 6100 86003 6103
rect 87598 6100 87604 6112
rect 85991 6072 87604 6100
rect 85991 6069 86003 6072
rect 85945 6063 86003 6069
rect 87598 6060 87604 6072
rect 87656 6060 87662 6112
rect 87690 6060 87696 6112
rect 87748 6100 87754 6112
rect 88168 6109 88196 6140
rect 88153 6103 88211 6109
rect 88153 6100 88165 6103
rect 87748 6072 88165 6100
rect 87748 6060 87754 6072
rect 88153 6069 88165 6072
rect 88199 6069 88211 6103
rect 88153 6063 88211 6069
rect 91002 6060 91008 6112
rect 91060 6100 91066 6112
rect 91373 6103 91431 6109
rect 91373 6100 91385 6103
rect 91060 6072 91385 6100
rect 91060 6060 91066 6072
rect 91373 6069 91385 6072
rect 91419 6100 91431 6103
rect 91830 6100 91836 6112
rect 91419 6072 91836 6100
rect 91419 6069 91431 6072
rect 91373 6063 91431 6069
rect 91830 6060 91836 6072
rect 91888 6060 91894 6112
rect 92750 6060 92756 6112
rect 92808 6100 92814 6112
rect 93305 6103 93363 6109
rect 93305 6100 93317 6103
rect 92808 6072 93317 6100
rect 92808 6060 92814 6072
rect 93305 6069 93317 6072
rect 93351 6069 93363 6103
rect 93305 6063 93363 6069
rect 1104 6010 94852 6032
rect 1104 5958 12668 6010
rect 12720 5958 12732 6010
rect 12784 5958 12796 6010
rect 12848 5958 12860 6010
rect 12912 5958 12924 6010
rect 12976 5958 36105 6010
rect 36157 5958 36169 6010
rect 36221 5958 36233 6010
rect 36285 5958 36297 6010
rect 36349 5958 36361 6010
rect 36413 5958 59542 6010
rect 59594 5958 59606 6010
rect 59658 5958 59670 6010
rect 59722 5958 59734 6010
rect 59786 5958 59798 6010
rect 59850 5958 82979 6010
rect 83031 5958 83043 6010
rect 83095 5958 83107 6010
rect 83159 5958 83171 6010
rect 83223 5958 83235 6010
rect 83287 5958 94852 6010
rect 1104 5936 94852 5958
rect 9490 5856 9496 5908
rect 9548 5896 9554 5908
rect 10321 5899 10379 5905
rect 10321 5896 10333 5899
rect 9548 5868 10333 5896
rect 9548 5856 9554 5868
rect 10321 5865 10333 5868
rect 10367 5896 10379 5899
rect 10686 5896 10692 5908
rect 10367 5868 10692 5896
rect 10367 5865 10379 5868
rect 10321 5859 10379 5865
rect 10686 5856 10692 5868
rect 10744 5856 10750 5908
rect 19886 5896 19892 5908
rect 19847 5868 19892 5896
rect 19886 5856 19892 5868
rect 19944 5856 19950 5908
rect 20548 5868 22784 5896
rect 8573 5831 8631 5837
rect 8573 5797 8585 5831
rect 8619 5828 8631 5831
rect 20548 5828 20576 5868
rect 22649 5831 22707 5837
rect 22649 5828 22661 5831
rect 8619 5800 12434 5828
rect 8619 5797 8631 5800
rect 8573 5791 8631 5797
rect 3970 5760 3976 5772
rect 3931 5732 3976 5760
rect 3970 5720 3976 5732
rect 4028 5720 4034 5772
rect 6365 5763 6423 5769
rect 6365 5729 6377 5763
rect 6411 5760 6423 5763
rect 6822 5760 6828 5772
rect 6411 5732 6828 5760
rect 6411 5729 6423 5732
rect 6365 5723 6423 5729
rect 6822 5720 6828 5732
rect 6880 5720 6886 5772
rect 7101 5763 7159 5769
rect 7101 5729 7113 5763
rect 7147 5760 7159 5763
rect 9217 5763 9275 5769
rect 9217 5760 9229 5763
rect 7147 5732 9229 5760
rect 7147 5729 7159 5732
rect 7101 5723 7159 5729
rect 9217 5729 9229 5732
rect 9263 5729 9275 5763
rect 9217 5723 9275 5729
rect 5718 5692 5724 5704
rect 5382 5664 5724 5692
rect 5718 5652 5724 5664
rect 5776 5652 5782 5704
rect 9309 5695 9367 5701
rect 9309 5661 9321 5695
rect 9355 5661 9367 5695
rect 12406 5692 12434 5800
rect 16316 5800 20576 5828
rect 20640 5800 22661 5828
rect 16316 5769 16344 5800
rect 16301 5763 16359 5769
rect 14292 5732 15516 5760
rect 14292 5701 14320 5732
rect 15488 5701 15516 5732
rect 16301 5729 16313 5763
rect 16347 5729 16359 5763
rect 16301 5723 16359 5729
rect 18506 5720 18512 5772
rect 18564 5760 18570 5772
rect 19521 5763 19579 5769
rect 19521 5760 19533 5763
rect 18564 5732 19533 5760
rect 18564 5720 18570 5732
rect 19521 5729 19533 5732
rect 19567 5729 19579 5763
rect 19521 5723 19579 5729
rect 19702 5720 19708 5772
rect 19760 5760 19766 5772
rect 20533 5763 20591 5769
rect 20533 5760 20545 5763
rect 19760 5732 20545 5760
rect 19760 5720 19766 5732
rect 20533 5729 20545 5732
rect 20579 5729 20591 5763
rect 20533 5723 20591 5729
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 12406 5664 14289 5692
rect 9309 5655 9367 5661
rect 14277 5661 14289 5664
rect 14323 5661 14335 5695
rect 15289 5695 15347 5701
rect 15289 5692 15301 5695
rect 14277 5655 14335 5661
rect 14384 5664 15301 5692
rect 4246 5624 4252 5636
rect 4207 5596 4252 5624
rect 4246 5584 4252 5596
rect 4304 5584 4310 5636
rect 5736 5624 5764 5652
rect 9324 5624 9352 5655
rect 13078 5624 13084 5636
rect 5736 5596 7590 5624
rect 9324 5596 13084 5624
rect 5718 5556 5724 5568
rect 5679 5528 5724 5556
rect 5718 5516 5724 5528
rect 5776 5516 5782 5568
rect 7484 5556 7512 5596
rect 13078 5584 13084 5596
rect 13136 5624 13142 5636
rect 14384 5624 14412 5664
rect 15289 5661 15301 5664
rect 15335 5661 15347 5695
rect 15289 5655 15347 5661
rect 15473 5695 15531 5701
rect 15473 5661 15485 5695
rect 15519 5661 15531 5695
rect 19610 5692 19616 5704
rect 19571 5664 19616 5692
rect 15473 5655 15531 5661
rect 19610 5652 19616 5664
rect 19668 5652 19674 5704
rect 20640 5701 20668 5800
rect 22649 5797 22661 5800
rect 22695 5797 22707 5831
rect 22756 5828 22784 5868
rect 22830 5856 22836 5908
rect 22888 5896 22894 5908
rect 23109 5899 23167 5905
rect 23109 5896 23121 5899
rect 22888 5868 23121 5896
rect 22888 5856 22894 5868
rect 23109 5865 23121 5868
rect 23155 5896 23167 5899
rect 23566 5896 23572 5908
rect 23155 5868 23572 5896
rect 23155 5865 23167 5868
rect 23109 5859 23167 5865
rect 23566 5856 23572 5868
rect 23624 5856 23630 5908
rect 25682 5896 25688 5908
rect 24688 5868 25688 5896
rect 23750 5828 23756 5840
rect 22756 5800 23756 5828
rect 22649 5791 22707 5797
rect 22664 5760 22692 5791
rect 23750 5788 23756 5800
rect 23808 5788 23814 5840
rect 24688 5828 24716 5868
rect 25682 5856 25688 5868
rect 25740 5856 25746 5908
rect 25866 5896 25872 5908
rect 25827 5868 25872 5896
rect 25866 5856 25872 5868
rect 25924 5856 25930 5908
rect 28718 5896 28724 5908
rect 25976 5868 28724 5896
rect 24044 5800 24716 5828
rect 23017 5763 23075 5769
rect 21652 5732 22600 5760
rect 22664 5732 22968 5760
rect 20625 5695 20683 5701
rect 20625 5661 20637 5695
rect 20671 5661 20683 5695
rect 20625 5655 20683 5661
rect 14550 5624 14556 5636
rect 13136 5596 14412 5624
rect 14511 5596 14556 5624
rect 13136 5584 13142 5596
rect 14550 5584 14556 5596
rect 14608 5584 14614 5636
rect 19426 5584 19432 5636
rect 19484 5624 19490 5636
rect 21652 5633 21680 5732
rect 21821 5695 21879 5701
rect 21821 5661 21833 5695
rect 21867 5692 21879 5695
rect 22572 5692 22600 5732
rect 22646 5692 22652 5704
rect 21867 5664 22508 5692
rect 22572 5664 22652 5692
rect 21867 5661 21879 5664
rect 21821 5655 21879 5661
rect 21637 5627 21695 5633
rect 21637 5624 21649 5627
rect 19484 5596 21649 5624
rect 19484 5584 19490 5596
rect 21637 5593 21649 5596
rect 21683 5593 21695 5627
rect 21637 5587 21695 5593
rect 21913 5627 21971 5633
rect 21913 5593 21925 5627
rect 21959 5624 21971 5627
rect 22094 5624 22100 5636
rect 21959 5596 22100 5624
rect 21959 5593 21971 5596
rect 21913 5587 21971 5593
rect 22094 5584 22100 5596
rect 22152 5584 22158 5636
rect 22189 5627 22247 5633
rect 22189 5593 22201 5627
rect 22235 5624 22247 5627
rect 22370 5624 22376 5636
rect 22235 5596 22376 5624
rect 22235 5593 22247 5596
rect 22189 5587 22247 5593
rect 22370 5584 22376 5596
rect 22428 5584 22434 5636
rect 8386 5556 8392 5568
rect 7484 5528 8392 5556
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 9858 5556 9864 5568
rect 9819 5528 9864 5556
rect 9858 5516 9864 5528
rect 9916 5556 9922 5568
rect 10778 5556 10784 5568
rect 9916 5528 10784 5556
rect 9916 5516 9922 5528
rect 10778 5516 10784 5528
rect 10836 5556 10842 5568
rect 11149 5559 11207 5565
rect 11149 5556 11161 5559
rect 10836 5528 11161 5556
rect 10836 5516 10842 5528
rect 11149 5525 11161 5528
rect 11195 5525 11207 5559
rect 22002 5556 22008 5568
rect 21963 5528 22008 5556
rect 11149 5519 11207 5525
rect 22002 5516 22008 5528
rect 22060 5516 22066 5568
rect 22480 5556 22508 5664
rect 22646 5652 22652 5664
rect 22704 5652 22710 5704
rect 22830 5692 22836 5704
rect 22791 5664 22836 5692
rect 22830 5652 22836 5664
rect 22888 5652 22894 5704
rect 22940 5694 22968 5732
rect 23017 5729 23029 5763
rect 23063 5760 23075 5763
rect 23290 5760 23296 5772
rect 23063 5732 23296 5760
rect 23063 5729 23075 5732
rect 23017 5723 23075 5729
rect 23290 5720 23296 5732
rect 23348 5720 23354 5772
rect 24044 5701 24072 5800
rect 24946 5788 24952 5840
rect 25004 5828 25010 5840
rect 25976 5828 26004 5868
rect 28718 5856 28724 5868
rect 28776 5856 28782 5908
rect 34241 5899 34299 5905
rect 34241 5865 34253 5899
rect 34287 5896 34299 5899
rect 40126 5896 40132 5908
rect 34287 5868 40132 5896
rect 34287 5865 34299 5868
rect 34241 5859 34299 5865
rect 40126 5856 40132 5868
rect 40184 5856 40190 5908
rect 40773 5899 40831 5905
rect 40773 5865 40785 5899
rect 40819 5896 40831 5899
rect 41598 5896 41604 5908
rect 40819 5868 41604 5896
rect 40819 5865 40831 5868
rect 40773 5859 40831 5865
rect 41598 5856 41604 5868
rect 41656 5896 41662 5908
rect 42886 5896 42892 5908
rect 41656 5868 42892 5896
rect 41656 5856 41662 5868
rect 42886 5856 42892 5868
rect 42944 5856 42950 5908
rect 42981 5899 43039 5905
rect 42981 5865 42993 5899
rect 43027 5896 43039 5899
rect 44542 5896 44548 5908
rect 43027 5868 44548 5896
rect 43027 5865 43039 5868
rect 42981 5859 43039 5865
rect 44542 5856 44548 5868
rect 44600 5856 44606 5908
rect 46658 5856 46664 5908
rect 46716 5896 46722 5908
rect 47765 5899 47823 5905
rect 47765 5896 47777 5899
rect 46716 5868 47777 5896
rect 46716 5856 46722 5868
rect 47765 5865 47777 5868
rect 47811 5865 47823 5899
rect 47765 5859 47823 5865
rect 48038 5856 48044 5908
rect 48096 5896 48102 5908
rect 49510 5896 49516 5908
rect 48096 5868 49516 5896
rect 48096 5856 48102 5868
rect 49510 5856 49516 5868
rect 49568 5856 49574 5908
rect 49786 5896 49792 5908
rect 49747 5868 49792 5896
rect 49786 5856 49792 5868
rect 49844 5856 49850 5908
rect 50798 5896 50804 5908
rect 50759 5868 50804 5896
rect 50798 5856 50804 5868
rect 50856 5856 50862 5908
rect 51442 5896 51448 5908
rect 51403 5868 51448 5896
rect 51442 5856 51448 5868
rect 51500 5856 51506 5908
rect 51718 5856 51724 5908
rect 51776 5896 51782 5908
rect 51997 5899 52055 5905
rect 51997 5896 52009 5899
rect 51776 5868 52009 5896
rect 51776 5856 51782 5868
rect 51997 5865 52009 5868
rect 52043 5865 52055 5899
rect 51997 5859 52055 5865
rect 52546 5856 52552 5908
rect 52604 5896 52610 5908
rect 52825 5899 52883 5905
rect 52825 5896 52837 5899
rect 52604 5868 52837 5896
rect 52604 5856 52610 5868
rect 52825 5865 52837 5868
rect 52871 5865 52883 5899
rect 52825 5859 52883 5865
rect 53282 5856 53288 5908
rect 53340 5896 53346 5908
rect 53377 5899 53435 5905
rect 53377 5896 53389 5899
rect 53340 5868 53389 5896
rect 53340 5856 53346 5868
rect 53377 5865 53389 5868
rect 53423 5865 53435 5899
rect 53377 5859 53435 5865
rect 53742 5856 53748 5908
rect 53800 5896 53806 5908
rect 53929 5899 53987 5905
rect 53929 5896 53941 5899
rect 53800 5868 53941 5896
rect 53800 5856 53806 5868
rect 53929 5865 53941 5868
rect 53975 5865 53987 5899
rect 54478 5896 54484 5908
rect 54439 5868 54484 5896
rect 53929 5859 53987 5865
rect 54478 5856 54484 5868
rect 54536 5856 54542 5908
rect 59446 5896 59452 5908
rect 55048 5868 59452 5896
rect 28442 5828 28448 5840
rect 25004 5800 26004 5828
rect 28403 5800 28448 5828
rect 25004 5788 25010 5800
rect 28442 5788 28448 5800
rect 28500 5788 28506 5840
rect 28966 5800 32628 5828
rect 24118 5720 24124 5772
rect 24176 5760 24182 5772
rect 26973 5763 27031 5769
rect 26973 5760 26985 5763
rect 24176 5732 26985 5760
rect 24176 5720 24182 5732
rect 26973 5729 26985 5732
rect 27019 5729 27031 5763
rect 26973 5723 27031 5729
rect 27062 5720 27068 5772
rect 27120 5760 27126 5772
rect 28966 5760 28994 5800
rect 27120 5732 28994 5760
rect 27120 5720 27126 5732
rect 31754 5720 31760 5772
rect 31812 5760 31818 5772
rect 32033 5763 32091 5769
rect 32033 5760 32045 5763
rect 31812 5732 32045 5760
rect 31812 5720 31818 5732
rect 32033 5729 32045 5732
rect 32079 5760 32091 5763
rect 32490 5760 32496 5772
rect 32079 5732 32496 5760
rect 32079 5729 32091 5732
rect 32033 5723 32091 5729
rect 32490 5720 32496 5732
rect 32548 5720 32554 5772
rect 32600 5760 32628 5800
rect 35526 5788 35532 5840
rect 35584 5828 35590 5840
rect 36817 5831 36875 5837
rect 36817 5828 36829 5831
rect 35584 5800 36829 5828
rect 35584 5788 35590 5800
rect 36817 5797 36829 5800
rect 36863 5797 36875 5831
rect 38102 5828 38108 5840
rect 38063 5800 38108 5828
rect 36817 5791 36875 5797
rect 38102 5788 38108 5800
rect 38160 5788 38166 5840
rect 38838 5828 38844 5840
rect 38799 5800 38844 5828
rect 38838 5788 38844 5800
rect 38896 5788 38902 5840
rect 39022 5788 39028 5840
rect 39080 5828 39086 5840
rect 39393 5831 39451 5837
rect 39393 5828 39405 5831
rect 39080 5800 39405 5828
rect 39080 5788 39086 5800
rect 39393 5797 39405 5800
rect 39439 5797 39451 5831
rect 39393 5791 39451 5797
rect 40310 5788 40316 5840
rect 40368 5828 40374 5840
rect 41230 5828 41236 5840
rect 40368 5800 41236 5828
rect 40368 5788 40374 5800
rect 41230 5788 41236 5800
rect 41288 5788 41294 5840
rect 43993 5831 44051 5837
rect 43993 5797 44005 5831
rect 44039 5828 44051 5831
rect 44358 5828 44364 5840
rect 44039 5800 44364 5828
rect 44039 5797 44051 5800
rect 43993 5791 44051 5797
rect 44358 5788 44364 5800
rect 44416 5788 44422 5840
rect 45278 5788 45284 5840
rect 45336 5828 45342 5840
rect 46569 5831 46627 5837
rect 46569 5828 46581 5831
rect 45336 5800 46581 5828
rect 45336 5788 45342 5800
rect 46569 5797 46581 5800
rect 46615 5797 46627 5831
rect 46569 5791 46627 5797
rect 49694 5788 49700 5840
rect 49752 5828 49758 5840
rect 51350 5828 51356 5840
rect 49752 5800 51074 5828
rect 51311 5800 51356 5828
rect 49752 5788 49758 5800
rect 35066 5760 35072 5772
rect 32600 5732 35072 5760
rect 35066 5720 35072 5732
rect 35124 5760 35130 5772
rect 35437 5763 35495 5769
rect 35437 5760 35449 5763
rect 35124 5732 35449 5760
rect 35124 5720 35130 5732
rect 35437 5729 35449 5732
rect 35483 5760 35495 5763
rect 35894 5760 35900 5772
rect 35483 5732 35900 5760
rect 35483 5729 35495 5732
rect 35437 5723 35495 5729
rect 35894 5720 35900 5732
rect 35952 5720 35958 5772
rect 35989 5763 36047 5769
rect 35989 5729 36001 5763
rect 36035 5760 36047 5763
rect 36446 5760 36452 5772
rect 36035 5732 36452 5760
rect 36035 5729 36047 5732
rect 35989 5723 36047 5729
rect 36446 5720 36452 5732
rect 36504 5720 36510 5772
rect 37458 5720 37464 5772
rect 37516 5760 37522 5772
rect 40129 5763 40187 5769
rect 40129 5760 40141 5763
rect 37516 5732 40141 5760
rect 37516 5720 37522 5732
rect 40129 5729 40141 5732
rect 40175 5760 40187 5763
rect 40862 5760 40868 5772
rect 40175 5732 40868 5760
rect 40175 5729 40187 5732
rect 40129 5723 40187 5729
rect 40862 5720 40868 5732
rect 40920 5720 40926 5772
rect 41509 5763 41567 5769
rect 41509 5729 41521 5763
rect 41555 5760 41567 5763
rect 44266 5760 44272 5772
rect 41555 5732 44272 5760
rect 41555 5729 41567 5732
rect 41509 5723 41567 5729
rect 44266 5720 44272 5732
rect 44324 5720 44330 5772
rect 45189 5763 45247 5769
rect 45189 5729 45201 5763
rect 45235 5760 45247 5763
rect 45646 5760 45652 5772
rect 45235 5732 45652 5760
rect 45235 5729 45247 5732
rect 45189 5723 45247 5729
rect 45646 5720 45652 5732
rect 45704 5720 45710 5772
rect 45738 5720 45744 5772
rect 45796 5760 45802 5772
rect 48222 5760 48228 5772
rect 45796 5732 48228 5760
rect 45796 5720 45802 5732
rect 48222 5720 48228 5732
rect 48280 5720 48286 5772
rect 48777 5763 48835 5769
rect 48777 5729 48789 5763
rect 48823 5760 48835 5763
rect 51046 5760 51074 5800
rect 51350 5788 51356 5800
rect 51408 5788 51414 5840
rect 55048 5828 55076 5868
rect 59446 5856 59452 5868
rect 59504 5856 59510 5908
rect 60090 5896 60096 5908
rect 60051 5868 60096 5896
rect 60090 5856 60096 5868
rect 60148 5856 60154 5908
rect 62114 5905 62120 5908
rect 62104 5899 62120 5905
rect 62104 5865 62116 5899
rect 62104 5859 62120 5865
rect 62114 5856 62120 5859
rect 62172 5856 62178 5908
rect 62298 5856 62304 5908
rect 62356 5896 62362 5908
rect 63402 5896 63408 5908
rect 62356 5868 63408 5896
rect 62356 5856 62362 5868
rect 63402 5856 63408 5868
rect 63460 5856 63466 5908
rect 65061 5899 65119 5905
rect 65061 5865 65073 5899
rect 65107 5896 65119 5899
rect 67358 5896 67364 5908
rect 65107 5868 67364 5896
rect 65107 5865 65119 5868
rect 65061 5859 65119 5865
rect 67358 5856 67364 5868
rect 67416 5856 67422 5908
rect 68094 5896 68100 5908
rect 68055 5868 68100 5896
rect 68094 5856 68100 5868
rect 68152 5896 68158 5908
rect 68649 5899 68707 5905
rect 68649 5896 68661 5899
rect 68152 5868 68661 5896
rect 68152 5856 68158 5868
rect 68649 5865 68661 5868
rect 68695 5865 68707 5899
rect 69198 5896 69204 5908
rect 69159 5868 69204 5896
rect 68649 5859 68707 5865
rect 69198 5856 69204 5868
rect 69256 5856 69262 5908
rect 69290 5856 69296 5908
rect 69348 5896 69354 5908
rect 70118 5896 70124 5908
rect 69348 5868 70124 5896
rect 69348 5856 69354 5868
rect 70118 5856 70124 5868
rect 70176 5856 70182 5908
rect 70397 5899 70455 5905
rect 70397 5865 70409 5899
rect 70443 5896 70455 5899
rect 70578 5896 70584 5908
rect 70443 5868 70584 5896
rect 70443 5865 70455 5868
rect 70397 5859 70455 5865
rect 70578 5856 70584 5868
rect 70636 5856 70642 5908
rect 70946 5896 70952 5908
rect 70907 5868 70952 5896
rect 70946 5856 70952 5868
rect 71004 5856 71010 5908
rect 71406 5856 71412 5908
rect 71464 5896 71470 5908
rect 74350 5896 74356 5908
rect 71464 5868 74356 5896
rect 71464 5856 71470 5868
rect 74350 5856 74356 5868
rect 74408 5856 74414 5908
rect 74902 5856 74908 5908
rect 74960 5896 74966 5908
rect 75273 5899 75331 5905
rect 75273 5896 75285 5899
rect 74960 5868 75285 5896
rect 74960 5856 74966 5868
rect 75273 5865 75285 5868
rect 75319 5896 75331 5899
rect 75319 5868 76236 5896
rect 75319 5865 75331 5868
rect 75273 5859 75331 5865
rect 58894 5828 58900 5840
rect 51460 5800 55076 5828
rect 55140 5800 58900 5828
rect 51460 5760 51488 5800
rect 48823 5732 50476 5760
rect 51046 5732 51488 5760
rect 48823 5729 48835 5732
rect 48777 5723 48835 5729
rect 24029 5695 24087 5701
rect 22940 5666 23060 5694
rect 23032 5636 23060 5666
rect 24029 5661 24041 5695
rect 24075 5661 24087 5695
rect 24029 5655 24087 5661
rect 24210 5652 24216 5704
rect 24268 5692 24274 5704
rect 24765 5695 24823 5701
rect 24765 5692 24777 5695
rect 24268 5664 24777 5692
rect 24268 5652 24274 5664
rect 24765 5661 24777 5664
rect 24811 5661 24823 5695
rect 24765 5655 24823 5661
rect 24854 5652 24860 5704
rect 24912 5692 24918 5704
rect 24949 5695 25007 5701
rect 24949 5692 24961 5695
rect 24912 5664 24961 5692
rect 24912 5652 24918 5664
rect 24949 5661 24961 5664
rect 24995 5692 25007 5695
rect 25222 5692 25228 5704
rect 24995 5664 25228 5692
rect 24995 5661 25007 5664
rect 24949 5655 25007 5661
rect 25222 5652 25228 5664
rect 25280 5652 25286 5704
rect 25406 5692 25412 5704
rect 25367 5664 25412 5692
rect 25406 5652 25412 5664
rect 25464 5652 25470 5704
rect 25682 5692 25688 5704
rect 25595 5664 25688 5692
rect 25682 5652 25688 5664
rect 25740 5692 25746 5704
rect 26142 5692 26148 5704
rect 25740 5664 26148 5692
rect 25740 5652 25746 5664
rect 26142 5652 26148 5664
rect 26200 5652 26206 5704
rect 26694 5692 26700 5704
rect 26655 5664 26700 5692
rect 26694 5652 26700 5664
rect 26752 5652 26758 5704
rect 38010 5652 38016 5704
rect 38068 5652 38074 5704
rect 41230 5692 41236 5704
rect 41191 5664 41236 5692
rect 41230 5652 41236 5664
rect 41288 5652 41294 5704
rect 44450 5692 44456 5704
rect 44100 5664 44456 5692
rect 23014 5584 23020 5636
rect 23072 5584 23078 5636
rect 23106 5584 23112 5636
rect 23164 5624 23170 5636
rect 23164 5596 23209 5624
rect 23164 5584 23170 5596
rect 23474 5584 23480 5636
rect 23532 5624 23538 5636
rect 25501 5627 25559 5633
rect 25501 5624 25513 5627
rect 23532 5596 25513 5624
rect 23532 5584 23538 5596
rect 25501 5593 25513 5596
rect 25547 5593 25559 5627
rect 25501 5587 25559 5593
rect 25590 5584 25596 5636
rect 25648 5624 25654 5636
rect 27430 5624 27436 5636
rect 25648 5596 27436 5624
rect 25648 5584 25654 5596
rect 27430 5584 27436 5596
rect 27488 5584 27494 5636
rect 29822 5584 29828 5636
rect 29880 5624 29886 5636
rect 30285 5627 30343 5633
rect 30285 5624 30297 5627
rect 29880 5596 30297 5624
rect 29880 5584 29886 5596
rect 30285 5593 30297 5596
rect 30331 5593 30343 5627
rect 32766 5624 32772 5636
rect 32727 5596 32772 5624
rect 30285 5587 30343 5593
rect 32766 5584 32772 5596
rect 32824 5584 32830 5636
rect 33226 5584 33232 5636
rect 33284 5584 33290 5636
rect 37458 5624 37464 5636
rect 35268 5596 37464 5624
rect 23124 5556 23152 5584
rect 22480 5528 23152 5556
rect 24026 5516 24032 5568
rect 24084 5556 24090 5568
rect 24854 5556 24860 5568
rect 24084 5528 24860 5556
rect 24084 5516 24090 5528
rect 24854 5516 24860 5528
rect 24912 5516 24918 5568
rect 24949 5559 25007 5565
rect 24949 5525 24961 5559
rect 24995 5556 25007 5559
rect 25130 5556 25136 5568
rect 24995 5528 25136 5556
rect 24995 5525 25007 5528
rect 24949 5519 25007 5525
rect 25130 5516 25136 5528
rect 25188 5516 25194 5568
rect 25222 5516 25228 5568
rect 25280 5556 25286 5568
rect 32582 5556 32588 5568
rect 25280 5528 32588 5556
rect 25280 5516 25286 5528
rect 32582 5516 32588 5528
rect 32640 5516 32646 5568
rect 32674 5516 32680 5568
rect 32732 5556 32738 5568
rect 35268 5556 35296 5596
rect 37458 5584 37464 5596
rect 37516 5584 37522 5636
rect 37553 5627 37611 5633
rect 37553 5593 37565 5627
rect 37599 5624 37611 5627
rect 38028 5624 38056 5652
rect 37599 5596 38654 5624
rect 37599 5593 37611 5596
rect 37553 5587 37611 5593
rect 32732 5528 35296 5556
rect 38626 5556 38654 5596
rect 42518 5584 42524 5636
rect 42576 5584 42582 5636
rect 44100 5556 44128 5664
rect 44450 5652 44456 5664
rect 44508 5652 44514 5704
rect 44637 5695 44695 5701
rect 44637 5661 44649 5695
rect 44683 5692 44695 5695
rect 47670 5692 47676 5704
rect 44683 5664 47676 5692
rect 44683 5661 44695 5664
rect 44637 5655 44695 5661
rect 47670 5652 47676 5664
rect 47728 5652 47734 5704
rect 48682 5692 48688 5704
rect 48643 5664 48688 5692
rect 48682 5652 48688 5664
rect 48740 5652 48746 5704
rect 48869 5695 48927 5701
rect 48869 5661 48881 5695
rect 48915 5661 48927 5695
rect 49510 5692 49516 5704
rect 49471 5664 49516 5692
rect 48869 5655 48927 5661
rect 44468 5624 44496 5652
rect 46017 5627 46075 5633
rect 46017 5624 46029 5627
rect 44468 5596 46029 5624
rect 46017 5593 46029 5596
rect 46063 5624 46075 5627
rect 46198 5624 46204 5636
rect 46063 5596 46204 5624
rect 46063 5593 46075 5596
rect 46017 5587 46075 5593
rect 46198 5584 46204 5596
rect 46256 5584 46262 5636
rect 47302 5624 47308 5636
rect 47263 5596 47308 5624
rect 47302 5584 47308 5596
rect 47360 5584 47366 5636
rect 48884 5624 48912 5655
rect 49510 5652 49516 5664
rect 49568 5652 49574 5704
rect 49602 5652 49608 5704
rect 49660 5692 49666 5704
rect 50246 5692 50252 5704
rect 49660 5664 50252 5692
rect 49660 5652 49666 5664
rect 50246 5652 50252 5664
rect 50304 5652 50310 5704
rect 50448 5701 50476 5732
rect 51534 5720 51540 5772
rect 51592 5760 51598 5772
rect 51592 5732 51637 5760
rect 51592 5720 51598 5732
rect 50341 5695 50399 5701
rect 50341 5661 50353 5695
rect 50387 5661 50399 5695
rect 50341 5655 50399 5661
rect 50433 5695 50491 5701
rect 50433 5661 50445 5695
rect 50479 5661 50491 5695
rect 50614 5692 50620 5704
rect 50575 5664 50620 5692
rect 50433 5655 50491 5661
rect 49620 5624 49648 5652
rect 48884 5596 49648 5624
rect 49789 5627 49847 5633
rect 49789 5593 49801 5627
rect 49835 5624 49847 5627
rect 50062 5624 50068 5636
rect 49835 5596 50068 5624
rect 49835 5593 49847 5596
rect 49789 5587 49847 5593
rect 50062 5584 50068 5596
rect 50120 5584 50126 5636
rect 50356 5624 50384 5655
rect 50614 5652 50620 5664
rect 50672 5652 50678 5704
rect 50706 5652 50712 5704
rect 50764 5692 50770 5704
rect 51261 5695 51319 5701
rect 51261 5692 51273 5695
rect 50764 5664 51273 5692
rect 50764 5652 50770 5664
rect 51261 5661 51273 5664
rect 51307 5692 51319 5695
rect 51736 5692 51856 5694
rect 55140 5692 55168 5800
rect 58894 5788 58900 5800
rect 58952 5788 58958 5840
rect 60274 5788 60280 5840
rect 60332 5828 60338 5840
rect 60332 5800 61884 5828
rect 60332 5788 60338 5800
rect 55214 5720 55220 5772
rect 55272 5760 55278 5772
rect 55585 5763 55643 5769
rect 55585 5760 55597 5763
rect 55272 5732 55597 5760
rect 55272 5720 55278 5732
rect 55585 5729 55597 5732
rect 55631 5729 55643 5763
rect 55585 5723 55643 5729
rect 56597 5763 56655 5769
rect 56597 5729 56609 5763
rect 56643 5760 56655 5763
rect 58802 5760 58808 5772
rect 56643 5732 58808 5760
rect 56643 5729 56655 5732
rect 56597 5723 56655 5729
rect 58802 5720 58808 5732
rect 58860 5720 58866 5772
rect 60734 5760 60740 5772
rect 60695 5732 60740 5760
rect 60734 5720 60740 5732
rect 60792 5720 60798 5772
rect 61856 5769 61884 5800
rect 63586 5788 63592 5840
rect 63644 5828 63650 5840
rect 64690 5828 64696 5840
rect 63644 5800 64696 5828
rect 63644 5788 63650 5800
rect 61841 5763 61899 5769
rect 61841 5729 61853 5763
rect 61887 5760 61899 5763
rect 63494 5760 63500 5772
rect 61887 5732 63500 5760
rect 61887 5729 61899 5732
rect 61841 5723 61899 5729
rect 63494 5720 63500 5732
rect 63552 5720 63558 5772
rect 63880 5769 63908 5800
rect 64690 5788 64696 5800
rect 64748 5828 64754 5840
rect 65702 5828 65708 5840
rect 64748 5800 65708 5828
rect 64748 5788 64754 5800
rect 65702 5788 65708 5800
rect 65760 5788 65766 5840
rect 67542 5828 67548 5840
rect 67455 5800 67548 5828
rect 67542 5788 67548 5800
rect 67600 5828 67606 5840
rect 74994 5828 75000 5840
rect 67600 5800 75000 5828
rect 67600 5788 67606 5800
rect 74994 5788 75000 5800
rect 75052 5788 75058 5840
rect 75089 5831 75147 5837
rect 75089 5797 75101 5831
rect 75135 5828 75147 5831
rect 76006 5828 76012 5840
rect 75135 5800 76012 5828
rect 75135 5797 75147 5800
rect 75089 5791 75147 5797
rect 76006 5788 76012 5800
rect 76064 5788 76070 5840
rect 63865 5763 63923 5769
rect 63865 5729 63877 5763
rect 63911 5729 63923 5763
rect 64598 5760 64604 5772
rect 64559 5732 64604 5760
rect 63865 5723 63923 5729
rect 64598 5720 64604 5732
rect 64656 5720 64662 5772
rect 66070 5760 66076 5772
rect 66031 5732 66076 5760
rect 66070 5720 66076 5732
rect 66128 5720 66134 5772
rect 66162 5720 66168 5772
rect 66220 5760 66226 5772
rect 71958 5760 71964 5772
rect 66220 5732 69980 5760
rect 71919 5732 71964 5760
rect 66220 5720 66226 5732
rect 51307 5666 55168 5692
rect 51307 5664 51764 5666
rect 51828 5664 55168 5666
rect 55677 5695 55735 5701
rect 51307 5661 51319 5664
rect 51261 5655 51319 5661
rect 55677 5661 55689 5695
rect 55723 5661 55735 5695
rect 55677 5655 55735 5661
rect 54386 5624 54392 5636
rect 50172 5596 50384 5624
rect 50448 5596 54392 5624
rect 38626 5528 44128 5556
rect 32732 5516 32738 5528
rect 44174 5516 44180 5568
rect 44232 5556 44238 5568
rect 44453 5559 44511 5565
rect 44453 5556 44465 5559
rect 44232 5528 44465 5556
rect 44232 5516 44238 5528
rect 44453 5525 44465 5528
rect 44499 5525 44511 5559
rect 44453 5519 44511 5525
rect 49142 5516 49148 5568
rect 49200 5556 49206 5568
rect 49329 5559 49387 5565
rect 49329 5556 49341 5559
rect 49200 5528 49341 5556
rect 49200 5516 49206 5528
rect 49329 5525 49341 5528
rect 49375 5556 49387 5559
rect 50172 5556 50200 5596
rect 49375 5528 50200 5556
rect 49375 5525 49387 5528
rect 49329 5519 49387 5525
rect 50246 5516 50252 5568
rect 50304 5556 50310 5568
rect 50448 5556 50476 5596
rect 54386 5584 54392 5596
rect 54444 5624 54450 5636
rect 55692 5624 55720 5655
rect 56686 5652 56692 5704
rect 56744 5692 56750 5704
rect 56781 5695 56839 5701
rect 56781 5692 56793 5695
rect 56744 5664 56793 5692
rect 56744 5652 56750 5664
rect 56781 5661 56793 5664
rect 56827 5661 56839 5695
rect 56962 5692 56968 5704
rect 56923 5664 56968 5692
rect 56781 5655 56839 5661
rect 56962 5652 56968 5664
rect 57020 5652 57026 5704
rect 57057 5695 57115 5701
rect 57057 5661 57069 5695
rect 57103 5692 57115 5695
rect 57238 5692 57244 5704
rect 57103 5664 57244 5692
rect 57103 5661 57115 5664
rect 57057 5655 57115 5661
rect 57238 5652 57244 5664
rect 57296 5692 57302 5704
rect 57517 5695 57575 5701
rect 57517 5692 57529 5695
rect 57296 5664 57529 5692
rect 57296 5652 57302 5664
rect 57517 5661 57529 5664
rect 57563 5661 57575 5695
rect 57517 5655 57575 5661
rect 57624 5664 58020 5692
rect 54444 5596 55720 5624
rect 54444 5584 54450 5596
rect 56134 5584 56140 5636
rect 56192 5624 56198 5636
rect 57624 5624 57652 5664
rect 56192 5596 57652 5624
rect 56192 5584 56198 5596
rect 57698 5584 57704 5636
rect 57756 5624 57762 5636
rect 57882 5624 57888 5636
rect 57756 5596 57801 5624
rect 57843 5596 57888 5624
rect 57756 5584 57762 5596
rect 57882 5584 57888 5596
rect 57940 5584 57946 5636
rect 57992 5624 58020 5664
rect 58434 5652 58440 5704
rect 58492 5692 58498 5704
rect 58897 5695 58955 5701
rect 58897 5692 58909 5695
rect 58492 5664 58909 5692
rect 58492 5652 58498 5664
rect 58897 5661 58909 5664
rect 58943 5661 58955 5695
rect 58897 5655 58955 5661
rect 59446 5652 59452 5704
rect 59504 5692 59510 5704
rect 60826 5692 60832 5704
rect 59504 5664 60734 5692
rect 60787 5664 60832 5692
rect 59504 5652 59510 5664
rect 59354 5624 59360 5636
rect 57992 5596 58480 5624
rect 50304 5528 50476 5556
rect 50304 5516 50310 5528
rect 52270 5516 52276 5568
rect 52328 5556 52334 5568
rect 54846 5556 54852 5568
rect 52328 5528 54852 5556
rect 52328 5516 52334 5528
rect 54846 5516 54852 5528
rect 54904 5516 54910 5568
rect 55858 5516 55864 5568
rect 55916 5556 55922 5568
rect 56045 5559 56103 5565
rect 56045 5556 56057 5559
rect 55916 5528 56057 5556
rect 55916 5516 55922 5528
rect 56045 5525 56057 5528
rect 56091 5525 56103 5559
rect 56045 5519 56103 5525
rect 56778 5516 56784 5568
rect 56836 5556 56842 5568
rect 58345 5559 58403 5565
rect 58345 5556 58357 5559
rect 56836 5528 58357 5556
rect 56836 5516 56842 5528
rect 58345 5525 58357 5528
rect 58391 5525 58403 5559
rect 58452 5556 58480 5596
rect 59096 5596 59360 5624
rect 59096 5556 59124 5596
rect 59354 5584 59360 5596
rect 59412 5624 59418 5636
rect 60274 5624 60280 5636
rect 59412 5596 60280 5624
rect 59412 5584 59418 5596
rect 60274 5584 60280 5596
rect 60332 5584 60338 5636
rect 60706 5624 60734 5664
rect 60826 5652 60832 5664
rect 60884 5652 60890 5704
rect 63678 5652 63684 5704
rect 63736 5692 63742 5704
rect 64693 5695 64751 5701
rect 64693 5692 64705 5695
rect 63736 5664 64705 5692
rect 63736 5652 63742 5664
rect 64693 5661 64705 5664
rect 64739 5661 64751 5695
rect 64693 5655 64751 5661
rect 65797 5695 65855 5701
rect 65797 5661 65809 5695
rect 65843 5661 65855 5695
rect 67726 5692 67732 5704
rect 67206 5664 67732 5692
rect 65797 5655 65855 5661
rect 63402 5624 63408 5636
rect 60706 5596 62528 5624
rect 63315 5596 63408 5624
rect 58452 5528 59124 5556
rect 58345 5519 58403 5525
rect 59170 5516 59176 5568
rect 59228 5556 59234 5568
rect 59449 5559 59507 5565
rect 59449 5556 59461 5559
rect 59228 5528 59461 5556
rect 59228 5516 59234 5528
rect 59449 5525 59461 5528
rect 59495 5525 59507 5559
rect 59449 5519 59507 5525
rect 59814 5516 59820 5568
rect 59872 5556 59878 5568
rect 60366 5556 60372 5568
rect 59872 5528 60372 5556
rect 59872 5516 59878 5528
rect 60366 5516 60372 5528
rect 60424 5516 60430 5568
rect 61197 5559 61255 5565
rect 61197 5525 61209 5559
rect 61243 5556 61255 5559
rect 62390 5556 62396 5568
rect 61243 5528 62396 5556
rect 61243 5525 61255 5528
rect 61197 5519 61255 5525
rect 62390 5516 62396 5528
rect 62448 5516 62454 5568
rect 62500 5556 62528 5596
rect 63402 5584 63408 5596
rect 63460 5624 63466 5636
rect 64874 5624 64880 5636
rect 63460 5596 64880 5624
rect 63460 5584 63466 5596
rect 64874 5584 64880 5596
rect 64932 5584 64938 5636
rect 64506 5556 64512 5568
rect 62500 5528 64512 5556
rect 64506 5516 64512 5528
rect 64564 5516 64570 5568
rect 65812 5556 65840 5655
rect 67726 5652 67732 5664
rect 67784 5652 67790 5704
rect 69842 5692 69848 5704
rect 69803 5664 69848 5692
rect 69842 5652 69848 5664
rect 69900 5652 69906 5704
rect 67450 5584 67456 5636
rect 67508 5624 67514 5636
rect 69952 5624 69980 5732
rect 71958 5720 71964 5732
rect 72016 5720 72022 5772
rect 73154 5760 73160 5772
rect 73115 5732 73160 5760
rect 73154 5720 73160 5732
rect 73212 5720 73218 5772
rect 73246 5720 73252 5772
rect 73304 5760 73310 5772
rect 73304 5732 75592 5760
rect 73304 5720 73310 5732
rect 75564 5704 75592 5732
rect 70118 5652 70124 5704
rect 70176 5692 70182 5704
rect 71406 5692 71412 5704
rect 70176 5664 71412 5692
rect 70176 5652 70182 5664
rect 71406 5652 71412 5664
rect 71464 5652 71470 5704
rect 71774 5692 71780 5704
rect 71735 5664 71780 5692
rect 71774 5652 71780 5664
rect 71832 5652 71838 5704
rect 73338 5652 73344 5704
rect 73396 5692 73402 5704
rect 74902 5692 74908 5704
rect 73396 5664 74908 5692
rect 73396 5652 73402 5664
rect 74902 5652 74908 5664
rect 74960 5652 74966 5704
rect 75270 5692 75276 5704
rect 75231 5664 75276 5692
rect 75270 5652 75276 5664
rect 75328 5652 75334 5704
rect 75365 5695 75423 5701
rect 75365 5661 75377 5695
rect 75411 5661 75423 5695
rect 75546 5692 75552 5704
rect 75459 5664 75552 5692
rect 75365 5655 75423 5661
rect 75178 5624 75184 5636
rect 67508 5596 69888 5624
rect 69952 5596 75184 5624
rect 67508 5584 67514 5596
rect 67634 5556 67640 5568
rect 65812 5528 67640 5556
rect 67634 5516 67640 5528
rect 67692 5556 67698 5568
rect 68186 5556 68192 5568
rect 67692 5528 68192 5556
rect 67692 5516 67698 5528
rect 68186 5516 68192 5528
rect 68244 5516 68250 5568
rect 69860 5556 69888 5596
rect 75178 5584 75184 5596
rect 75236 5584 75242 5636
rect 75380 5624 75408 5655
rect 75546 5652 75552 5664
rect 75604 5652 75610 5704
rect 76208 5692 76236 5868
rect 76282 5856 76288 5908
rect 76340 5896 76346 5908
rect 77846 5896 77852 5908
rect 76340 5868 77852 5896
rect 76340 5856 76346 5868
rect 77846 5856 77852 5868
rect 77904 5856 77910 5908
rect 79045 5899 79103 5905
rect 79045 5865 79057 5899
rect 79091 5896 79103 5899
rect 80974 5896 80980 5908
rect 79091 5868 80980 5896
rect 79091 5865 79103 5868
rect 79045 5859 79103 5865
rect 80974 5856 80980 5868
rect 81032 5856 81038 5908
rect 82814 5856 82820 5908
rect 82872 5896 82878 5908
rect 82909 5899 82967 5905
rect 82909 5896 82921 5899
rect 82872 5868 82921 5896
rect 82872 5856 82878 5868
rect 82909 5865 82921 5868
rect 82955 5865 82967 5899
rect 83458 5896 83464 5908
rect 83419 5868 83464 5896
rect 82909 5859 82967 5865
rect 83458 5856 83464 5868
rect 83516 5856 83522 5908
rect 84746 5856 84752 5908
rect 84804 5896 84810 5908
rect 85853 5899 85911 5905
rect 84804 5868 85252 5896
rect 84804 5856 84810 5868
rect 76742 5788 76748 5840
rect 76800 5828 76806 5840
rect 77389 5831 77447 5837
rect 77389 5828 77401 5831
rect 76800 5800 77401 5828
rect 76800 5788 76806 5800
rect 77389 5797 77401 5800
rect 77435 5797 77447 5831
rect 77389 5791 77447 5797
rect 80790 5788 80796 5840
rect 80848 5828 80854 5840
rect 81253 5831 81311 5837
rect 81253 5828 81265 5831
rect 80848 5800 81265 5828
rect 80848 5788 80854 5800
rect 81253 5797 81265 5800
rect 81299 5797 81311 5831
rect 81253 5791 81311 5797
rect 82722 5788 82728 5840
rect 82780 5828 82786 5840
rect 84286 5828 84292 5840
rect 82780 5800 84292 5828
rect 82780 5788 82786 5800
rect 84286 5788 84292 5800
rect 84344 5828 84350 5840
rect 85117 5831 85175 5837
rect 85117 5828 85129 5831
rect 84344 5800 85129 5828
rect 84344 5788 84350 5800
rect 85117 5797 85129 5800
rect 85163 5797 85175 5831
rect 85224 5828 85252 5868
rect 85853 5865 85865 5899
rect 85899 5896 85911 5899
rect 86402 5896 86408 5908
rect 85899 5868 86408 5896
rect 85899 5865 85911 5868
rect 85853 5859 85911 5865
rect 86402 5856 86408 5868
rect 86460 5856 86466 5908
rect 87598 5856 87604 5908
rect 87656 5896 87662 5908
rect 88429 5899 88487 5905
rect 88429 5896 88441 5899
rect 87656 5868 88441 5896
rect 87656 5856 87662 5868
rect 88429 5865 88441 5868
rect 88475 5896 88487 5899
rect 89806 5896 89812 5908
rect 88475 5868 89812 5896
rect 88475 5865 88487 5868
rect 88429 5859 88487 5865
rect 89806 5856 89812 5868
rect 89864 5856 89870 5908
rect 93118 5896 93124 5908
rect 91204 5868 93124 5896
rect 86126 5828 86132 5840
rect 85224 5800 86132 5828
rect 85117 5791 85175 5797
rect 86126 5788 86132 5800
rect 86184 5828 86190 5840
rect 87230 5828 87236 5840
rect 86184 5800 87236 5828
rect 86184 5788 86190 5800
rect 87230 5788 87236 5800
rect 87288 5788 87294 5840
rect 78769 5763 78827 5769
rect 78769 5729 78781 5763
rect 78815 5760 78827 5763
rect 78815 5732 80100 5760
rect 78815 5729 78827 5732
rect 78769 5723 78827 5729
rect 76377 5695 76435 5701
rect 76377 5692 76389 5695
rect 76208 5664 76389 5692
rect 76377 5661 76389 5664
rect 76423 5692 76435 5695
rect 77113 5695 77171 5701
rect 77113 5692 77125 5695
rect 76423 5664 77125 5692
rect 76423 5661 76435 5664
rect 76377 5655 76435 5661
rect 77113 5661 77125 5664
rect 77159 5661 77171 5695
rect 77113 5655 77171 5661
rect 78677 5695 78735 5701
rect 78677 5661 78689 5695
rect 78723 5692 78735 5695
rect 78723 5664 78812 5692
rect 78723 5661 78735 5664
rect 78677 5655 78735 5661
rect 78784 5636 78812 5664
rect 79042 5652 79048 5704
rect 79100 5692 79106 5704
rect 79686 5692 79692 5704
rect 79100 5664 79692 5692
rect 79100 5652 79106 5664
rect 79686 5652 79692 5664
rect 79744 5652 79750 5704
rect 80072 5682 80100 5732
rect 80698 5720 80704 5772
rect 80756 5760 80762 5772
rect 81526 5760 81532 5772
rect 80756 5732 80801 5760
rect 81268 5732 81532 5760
rect 80756 5720 80762 5732
rect 80425 5695 80483 5701
rect 80072 5654 80192 5682
rect 80425 5661 80437 5695
rect 80471 5692 80483 5695
rect 81268 5692 81296 5732
rect 81526 5720 81532 5732
rect 81584 5720 81590 5772
rect 81618 5720 81624 5772
rect 81676 5760 81682 5772
rect 84013 5763 84071 5769
rect 84013 5760 84025 5763
rect 81676 5732 84025 5760
rect 81676 5720 81682 5732
rect 84013 5729 84025 5732
rect 84059 5729 84071 5763
rect 84013 5723 84071 5729
rect 86586 5720 86592 5772
rect 86644 5760 86650 5772
rect 86644 5732 87092 5760
rect 86644 5720 86650 5732
rect 80471 5664 81296 5692
rect 80471 5661 80483 5664
rect 80425 5655 80483 5661
rect 75454 5624 75460 5636
rect 75380 5596 75460 5624
rect 75454 5584 75460 5596
rect 75512 5624 75518 5636
rect 75822 5624 75828 5636
rect 75512 5596 75828 5624
rect 75512 5584 75518 5596
rect 75822 5584 75828 5596
rect 75880 5584 75886 5636
rect 75914 5584 75920 5636
rect 75972 5624 75978 5636
rect 76101 5627 76159 5633
rect 76101 5624 76113 5627
rect 75972 5596 76113 5624
rect 75972 5584 75978 5596
rect 76101 5593 76113 5596
rect 76147 5593 76159 5627
rect 76101 5587 76159 5593
rect 78766 5584 78772 5636
rect 78824 5584 78830 5636
rect 74074 5556 74080 5568
rect 69860 5528 74080 5556
rect 74074 5516 74080 5528
rect 74132 5516 74138 5568
rect 75270 5516 75276 5568
rect 75328 5556 75334 5568
rect 76282 5556 76288 5568
rect 75328 5528 76288 5556
rect 75328 5516 75334 5528
rect 76282 5516 76288 5528
rect 76340 5516 76346 5568
rect 76466 5556 76472 5568
rect 76427 5528 76472 5556
rect 76466 5516 76472 5528
rect 76524 5516 76530 5568
rect 76653 5559 76711 5565
rect 76653 5525 76665 5559
rect 76699 5556 76711 5559
rect 76926 5556 76932 5568
rect 76699 5528 76932 5556
rect 76699 5525 76711 5528
rect 76653 5519 76711 5525
rect 76926 5516 76932 5528
rect 76984 5516 76990 5568
rect 77573 5559 77631 5565
rect 77573 5525 77585 5559
rect 77619 5556 77631 5559
rect 77662 5556 77668 5568
rect 77619 5528 77668 5556
rect 77619 5525 77631 5528
rect 77573 5519 77631 5525
rect 77662 5516 77668 5528
rect 77720 5516 77726 5568
rect 79505 5559 79563 5565
rect 79505 5525 79517 5559
rect 79551 5556 79563 5559
rect 79870 5556 79876 5568
rect 79551 5528 79876 5556
rect 79551 5525 79563 5528
rect 79505 5519 79563 5525
rect 79870 5516 79876 5528
rect 79928 5516 79934 5568
rect 79962 5516 79968 5568
rect 80020 5556 80026 5568
rect 80054 5556 80060 5568
rect 80020 5528 80060 5556
rect 80020 5516 80026 5528
rect 80054 5516 80060 5528
rect 80112 5516 80118 5568
rect 80164 5556 80192 5654
rect 81342 5652 81348 5704
rect 81400 5652 81406 5704
rect 81986 5652 81992 5704
rect 82044 5692 82050 5704
rect 86954 5692 86960 5704
rect 82044 5664 84700 5692
rect 86915 5664 86960 5692
rect 82044 5652 82050 5664
rect 80330 5584 80336 5636
rect 80388 5624 80394 5636
rect 81360 5624 81388 5652
rect 81805 5627 81863 5633
rect 81805 5624 81817 5627
rect 80388 5596 81817 5624
rect 80388 5584 80394 5596
rect 81805 5593 81817 5596
rect 81851 5624 81863 5627
rect 84565 5627 84623 5633
rect 84565 5624 84577 5627
rect 81851 5596 84577 5624
rect 81851 5593 81863 5596
rect 81805 5587 81863 5593
rect 84565 5593 84577 5596
rect 84611 5593 84623 5627
rect 84672 5624 84700 5664
rect 86954 5652 86960 5664
rect 87012 5652 87018 5704
rect 87064 5692 87092 5732
rect 87966 5720 87972 5772
rect 88024 5760 88030 5772
rect 89625 5763 89683 5769
rect 88024 5732 88069 5760
rect 88024 5720 88030 5732
rect 89625 5729 89637 5763
rect 89671 5760 89683 5763
rect 89714 5760 89720 5772
rect 89671 5732 89720 5760
rect 89671 5729 89683 5732
rect 89625 5723 89683 5729
rect 89714 5720 89720 5732
rect 89772 5720 89778 5772
rect 87693 5695 87751 5701
rect 87693 5692 87705 5695
rect 87064 5664 87705 5692
rect 87693 5661 87705 5664
rect 87739 5661 87751 5695
rect 87693 5655 87751 5661
rect 87782 5652 87788 5704
rect 87840 5692 87846 5704
rect 88613 5695 88671 5701
rect 88613 5692 88625 5695
rect 87840 5664 88625 5692
rect 87840 5652 87846 5664
rect 88613 5661 88625 5664
rect 88659 5661 88671 5695
rect 89346 5692 89352 5704
rect 89307 5664 89352 5692
rect 88613 5655 88671 5661
rect 89346 5652 89352 5664
rect 89404 5652 89410 5704
rect 91204 5692 91232 5868
rect 93118 5856 93124 5868
rect 93176 5856 93182 5908
rect 93394 5896 93400 5908
rect 93355 5868 93400 5896
rect 93394 5856 93400 5868
rect 93452 5856 93458 5908
rect 93762 5856 93768 5908
rect 93820 5896 93826 5908
rect 93857 5899 93915 5905
rect 93857 5896 93869 5899
rect 93820 5868 93869 5896
rect 93820 5856 93826 5868
rect 93857 5865 93869 5868
rect 93903 5865 93915 5899
rect 93857 5859 93915 5865
rect 92750 5828 92756 5840
rect 92711 5800 92756 5828
rect 92750 5788 92756 5800
rect 92808 5788 92814 5840
rect 91278 5720 91284 5772
rect 91336 5760 91342 5772
rect 91557 5763 91615 5769
rect 91557 5760 91569 5763
rect 91336 5732 91569 5760
rect 91336 5720 91342 5732
rect 91557 5729 91569 5732
rect 91603 5729 91615 5763
rect 91557 5723 91615 5729
rect 91830 5692 91836 5704
rect 89686 5664 91232 5692
rect 91791 5664 91836 5692
rect 89686 5624 89714 5664
rect 91830 5652 91836 5664
rect 91888 5652 91894 5704
rect 92477 5695 92535 5701
rect 92477 5661 92489 5695
rect 92523 5661 92535 5695
rect 93210 5692 93216 5704
rect 93171 5664 93216 5692
rect 92477 5655 92535 5661
rect 84672 5596 89714 5624
rect 84565 5587 84623 5593
rect 89898 5584 89904 5636
rect 89956 5624 89962 5636
rect 92492 5624 92520 5655
rect 93210 5652 93216 5664
rect 93268 5652 93274 5704
rect 89956 5596 92520 5624
rect 89956 5584 89962 5596
rect 81434 5556 81440 5568
rect 80164 5528 81440 5556
rect 81434 5516 81440 5528
rect 81492 5516 81498 5568
rect 81618 5516 81624 5568
rect 81676 5556 81682 5568
rect 82449 5559 82507 5565
rect 82449 5556 82461 5559
rect 81676 5528 82461 5556
rect 81676 5516 81682 5528
rect 82449 5525 82461 5528
rect 82495 5556 82507 5559
rect 86034 5556 86040 5568
rect 82495 5528 86040 5556
rect 82495 5525 82507 5528
rect 82449 5519 82507 5525
rect 86034 5516 86040 5528
rect 86092 5516 86098 5568
rect 86773 5559 86831 5565
rect 86773 5525 86785 5559
rect 86819 5556 86831 5559
rect 87138 5556 87144 5568
rect 86819 5528 87144 5556
rect 86819 5525 86831 5528
rect 86773 5519 86831 5525
rect 87138 5516 87144 5528
rect 87196 5516 87202 5568
rect 87230 5516 87236 5568
rect 87288 5556 87294 5568
rect 90177 5559 90235 5565
rect 90177 5556 90189 5559
rect 87288 5528 90189 5556
rect 87288 5516 87294 5528
rect 90177 5525 90189 5528
rect 90223 5556 90235 5559
rect 90637 5559 90695 5565
rect 90637 5556 90649 5559
rect 90223 5528 90649 5556
rect 90223 5525 90235 5528
rect 90177 5519 90235 5525
rect 90637 5525 90649 5528
rect 90683 5525 90695 5559
rect 90637 5519 90695 5525
rect 1104 5466 95011 5488
rect 1104 5414 24386 5466
rect 24438 5414 24450 5466
rect 24502 5414 24514 5466
rect 24566 5414 24578 5466
rect 24630 5414 24642 5466
rect 24694 5414 47823 5466
rect 47875 5414 47887 5466
rect 47939 5414 47951 5466
rect 48003 5414 48015 5466
rect 48067 5414 48079 5466
rect 48131 5414 71260 5466
rect 71312 5414 71324 5466
rect 71376 5414 71388 5466
rect 71440 5414 71452 5466
rect 71504 5414 71516 5466
rect 71568 5414 94697 5466
rect 94749 5414 94761 5466
rect 94813 5414 94825 5466
rect 94877 5414 94889 5466
rect 94941 5414 94953 5466
rect 95005 5414 95011 5466
rect 1104 5392 95011 5414
rect 4246 5352 4252 5364
rect 4207 5324 4252 5352
rect 4246 5312 4252 5324
rect 4304 5312 4310 5364
rect 8297 5355 8355 5361
rect 8297 5321 8309 5355
rect 8343 5352 8355 5355
rect 8386 5352 8392 5364
rect 8343 5324 8392 5352
rect 8343 5321 8355 5324
rect 8297 5315 8355 5321
rect 8386 5312 8392 5324
rect 8444 5312 8450 5364
rect 22097 5355 22155 5361
rect 22097 5321 22109 5355
rect 22143 5352 22155 5355
rect 22370 5352 22376 5364
rect 22143 5324 22376 5352
rect 22143 5321 22155 5324
rect 22097 5315 22155 5321
rect 22370 5312 22376 5324
rect 22428 5312 22434 5364
rect 22833 5355 22891 5361
rect 22833 5321 22845 5355
rect 22879 5352 22891 5355
rect 23474 5352 23480 5364
rect 22879 5324 23480 5352
rect 22879 5321 22891 5324
rect 22833 5315 22891 5321
rect 23474 5312 23480 5324
rect 23532 5312 23538 5364
rect 23750 5312 23756 5364
rect 23808 5352 23814 5364
rect 24762 5352 24768 5364
rect 23808 5324 24768 5352
rect 23808 5312 23814 5324
rect 24762 5312 24768 5324
rect 24820 5312 24826 5364
rect 24872 5324 33548 5352
rect 9582 5284 9588 5296
rect 9543 5256 9588 5284
rect 9582 5244 9588 5256
rect 9640 5244 9646 5296
rect 12986 5284 12992 5296
rect 12947 5256 12992 5284
rect 12986 5244 12992 5256
rect 13044 5244 13050 5296
rect 22002 5244 22008 5296
rect 22060 5284 22066 5296
rect 23293 5287 23351 5293
rect 23293 5284 23305 5287
rect 22060 5256 23305 5284
rect 22060 5244 22066 5256
rect 4338 5216 4344 5228
rect 4299 5188 4344 5216
rect 4338 5176 4344 5188
rect 4396 5176 4402 5228
rect 5718 5176 5724 5228
rect 5776 5216 5782 5228
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 5776 5188 6837 5216
rect 5776 5176 5782 5188
rect 6825 5185 6837 5188
rect 6871 5216 6883 5219
rect 14458 5216 14464 5228
rect 6871 5188 14464 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 14458 5176 14464 5188
rect 14516 5176 14522 5228
rect 22094 5176 22100 5228
rect 22152 5216 22158 5228
rect 22554 5216 22560 5228
rect 22152 5188 22560 5216
rect 22152 5176 22158 5188
rect 22554 5176 22560 5188
rect 22612 5176 22618 5228
rect 22756 5225 22784 5256
rect 23293 5253 23305 5256
rect 23339 5284 23351 5287
rect 23566 5284 23572 5296
rect 23339 5256 23572 5284
rect 23339 5253 23351 5256
rect 23293 5247 23351 5253
rect 23566 5244 23572 5256
rect 23624 5284 23630 5296
rect 24210 5284 24216 5296
rect 23624 5256 24216 5284
rect 23624 5244 23630 5256
rect 24210 5244 24216 5256
rect 24268 5244 24274 5296
rect 24394 5244 24400 5296
rect 24452 5284 24458 5296
rect 24872 5284 24900 5324
rect 24452 5256 24900 5284
rect 26145 5287 26203 5293
rect 24452 5244 24458 5256
rect 26145 5253 26157 5287
rect 26191 5284 26203 5287
rect 26234 5284 26240 5296
rect 26191 5256 26240 5284
rect 26191 5253 26203 5256
rect 26145 5247 26203 5253
rect 26234 5244 26240 5256
rect 26292 5244 26298 5296
rect 27341 5287 27399 5293
rect 27341 5284 27353 5287
rect 26620 5256 27353 5284
rect 22741 5219 22799 5225
rect 22741 5185 22753 5219
rect 22787 5185 22799 5219
rect 22741 5179 22799 5185
rect 22830 5176 22836 5228
rect 22888 5216 22894 5228
rect 23477 5219 23535 5225
rect 23477 5216 23489 5219
rect 22888 5188 23489 5216
rect 22888 5176 22894 5188
rect 23477 5185 23489 5188
rect 23523 5216 23535 5219
rect 24026 5216 24032 5228
rect 23523 5188 24032 5216
rect 23523 5185 23535 5188
rect 23477 5179 23535 5185
rect 24026 5176 24032 5188
rect 24084 5176 24090 5228
rect 25038 5176 25044 5228
rect 25096 5176 25102 5228
rect 13722 5108 13728 5160
rect 13780 5148 13786 5160
rect 14737 5151 14795 5157
rect 14737 5148 14749 5151
rect 13780 5120 14749 5148
rect 13780 5108 13786 5120
rect 14737 5117 14749 5120
rect 14783 5148 14795 5151
rect 15470 5148 15476 5160
rect 14783 5120 15476 5148
rect 14783 5117 14795 5120
rect 14737 5111 14795 5117
rect 15470 5108 15476 5120
rect 15528 5108 15534 5160
rect 15930 5108 15936 5160
rect 15988 5148 15994 5160
rect 24854 5148 24860 5160
rect 15988 5120 24860 5148
rect 15988 5108 15994 5120
rect 24854 5108 24860 5120
rect 24912 5108 24918 5160
rect 26421 5151 26479 5157
rect 26421 5117 26433 5151
rect 26467 5148 26479 5151
rect 26510 5148 26516 5160
rect 26467 5120 26516 5148
rect 26467 5117 26479 5120
rect 26421 5111 26479 5117
rect 26510 5108 26516 5120
rect 26568 5108 26574 5160
rect 8478 5040 8484 5092
rect 8536 5080 8542 5092
rect 24394 5080 24400 5092
rect 8536 5052 24400 5080
rect 8536 5040 8542 5052
rect 24394 5040 24400 5052
rect 24452 5040 24458 5092
rect 6917 5015 6975 5021
rect 6917 4981 6929 5015
rect 6963 5012 6975 5015
rect 7006 5012 7012 5024
rect 6963 4984 7012 5012
rect 6963 4981 6975 4984
rect 6917 4975 6975 4981
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 23658 5012 23664 5024
rect 23619 4984 23664 5012
rect 23658 4972 23664 4984
rect 23716 4972 23722 5024
rect 24210 5012 24216 5024
rect 24171 4984 24216 5012
rect 24210 4972 24216 4984
rect 24268 4972 24274 5024
rect 24670 5012 24676 5024
rect 24631 4984 24676 5012
rect 24670 4972 24676 4984
rect 24728 4972 24734 5024
rect 24762 4972 24768 5024
rect 24820 5012 24826 5024
rect 26620 5012 26648 5256
rect 27341 5253 27353 5256
rect 27387 5253 27399 5287
rect 28258 5284 28264 5296
rect 28219 5256 28264 5284
rect 27341 5247 27399 5253
rect 28258 5244 28264 5256
rect 28316 5244 28322 5296
rect 33226 5284 33232 5296
rect 31050 5256 33232 5284
rect 33226 5244 33232 5256
rect 33284 5244 33290 5296
rect 28721 5219 28779 5225
rect 28721 5185 28733 5219
rect 28767 5185 28779 5219
rect 28721 5179 28779 5185
rect 27246 5148 27252 5160
rect 27207 5120 27252 5148
rect 27246 5108 27252 5120
rect 27304 5108 27310 5160
rect 26694 5040 26700 5092
rect 26752 5080 26758 5092
rect 28736 5080 28764 5179
rect 31754 5176 31760 5228
rect 31812 5216 31818 5228
rect 32674 5216 32680 5228
rect 31812 5188 31857 5216
rect 32635 5188 32680 5216
rect 31812 5176 31818 5188
rect 32674 5176 32680 5188
rect 32732 5176 32738 5228
rect 31481 5151 31539 5157
rect 31481 5117 31493 5151
rect 31527 5148 31539 5151
rect 32585 5151 32643 5157
rect 31527 5120 31754 5148
rect 31527 5117 31539 5120
rect 31481 5111 31539 5117
rect 26752 5052 28764 5080
rect 31726 5080 31754 5120
rect 32585 5117 32597 5151
rect 32631 5117 32643 5151
rect 33520 5148 33548 5324
rect 34238 5312 34244 5364
rect 34296 5352 34302 5364
rect 34425 5355 34483 5361
rect 34425 5352 34437 5355
rect 34296 5324 34437 5352
rect 34296 5312 34302 5324
rect 34425 5321 34437 5324
rect 34471 5321 34483 5355
rect 37918 5352 37924 5364
rect 37879 5324 37924 5352
rect 34425 5315 34483 5321
rect 37918 5312 37924 5324
rect 37976 5312 37982 5364
rect 39669 5355 39727 5361
rect 39669 5321 39681 5355
rect 39715 5352 39727 5355
rect 40034 5352 40040 5364
rect 39715 5324 40040 5352
rect 39715 5321 39727 5324
rect 39669 5315 39727 5321
rect 40034 5312 40040 5324
rect 40092 5352 40098 5364
rect 40129 5355 40187 5361
rect 40129 5352 40141 5355
rect 40092 5324 40141 5352
rect 40092 5312 40098 5324
rect 40129 5321 40141 5324
rect 40175 5321 40187 5355
rect 40862 5352 40868 5364
rect 40823 5324 40868 5352
rect 40129 5315 40187 5321
rect 40862 5312 40868 5324
rect 40920 5312 40926 5364
rect 80054 5352 80060 5364
rect 41386 5324 80060 5352
rect 33594 5244 33600 5296
rect 33652 5284 33658 5296
rect 41386 5284 41414 5324
rect 80054 5312 80060 5324
rect 80112 5312 80118 5364
rect 81986 5352 81992 5364
rect 80164 5324 81992 5352
rect 33652 5256 41414 5284
rect 41509 5287 41567 5293
rect 33652 5244 33658 5256
rect 41509 5253 41521 5287
rect 41555 5284 41567 5287
rect 42058 5284 42064 5296
rect 41555 5256 42064 5284
rect 41555 5253 41567 5256
rect 41509 5247 41567 5253
rect 42058 5244 42064 5256
rect 42116 5244 42122 5296
rect 42702 5244 42708 5296
rect 42760 5284 42766 5296
rect 44269 5287 44327 5293
rect 44269 5284 44281 5287
rect 42760 5256 44281 5284
rect 42760 5244 42766 5256
rect 44269 5253 44281 5256
rect 44315 5253 44327 5287
rect 44269 5247 44327 5253
rect 45554 5244 45560 5296
rect 45612 5284 45618 5296
rect 46293 5287 46351 5293
rect 46293 5284 46305 5287
rect 45612 5256 46305 5284
rect 45612 5244 45618 5256
rect 46293 5253 46305 5256
rect 46339 5253 46351 5287
rect 46293 5247 46351 5253
rect 47762 5244 47768 5296
rect 47820 5284 47826 5296
rect 48225 5287 48283 5293
rect 48225 5284 48237 5287
rect 47820 5256 48237 5284
rect 47820 5244 47826 5256
rect 48225 5253 48237 5256
rect 48271 5284 48283 5287
rect 49405 5287 49463 5293
rect 49405 5284 49417 5287
rect 48271 5256 49417 5284
rect 48271 5253 48283 5256
rect 48225 5247 48283 5253
rect 49405 5253 49417 5256
rect 49451 5284 49463 5287
rect 49602 5284 49608 5296
rect 49451 5253 49464 5284
rect 49563 5256 49608 5284
rect 49405 5247 49464 5253
rect 36357 5219 36415 5225
rect 36357 5185 36369 5219
rect 36403 5216 36415 5219
rect 36446 5216 36452 5228
rect 36403 5188 36452 5216
rect 36403 5185 36415 5188
rect 36357 5179 36415 5185
rect 36446 5176 36452 5188
rect 36504 5176 36510 5228
rect 36722 5176 36728 5228
rect 36780 5216 36786 5228
rect 37645 5219 37703 5225
rect 37645 5216 37657 5219
rect 36780 5188 37657 5216
rect 36780 5176 36786 5188
rect 37645 5185 37657 5188
rect 37691 5185 37703 5219
rect 37645 5179 37703 5185
rect 38010 5176 38016 5228
rect 38068 5216 38074 5228
rect 42978 5216 42984 5228
rect 38068 5188 42748 5216
rect 42939 5188 42984 5216
rect 38068 5176 38074 5188
rect 36906 5148 36912 5160
rect 33520 5120 36584 5148
rect 36819 5120 36912 5148
rect 32585 5111 32643 5117
rect 32309 5083 32367 5089
rect 32309 5080 32321 5083
rect 31726 5052 32321 5080
rect 26752 5040 26758 5052
rect 32309 5049 32321 5052
rect 32355 5049 32367 5083
rect 32309 5043 32367 5049
rect 24820 4984 26648 5012
rect 24820 4972 24826 4984
rect 28442 4972 28448 5024
rect 28500 5012 28506 5024
rect 28905 5015 28963 5021
rect 28905 5012 28917 5015
rect 28500 4984 28917 5012
rect 28500 4972 28506 4984
rect 28905 4981 28917 4984
rect 28951 4981 28963 5015
rect 30006 5012 30012 5024
rect 29967 4984 30012 5012
rect 28905 4975 28963 4981
rect 30006 4972 30012 4984
rect 30064 4972 30070 5024
rect 30098 4972 30104 5024
rect 30156 5012 30162 5024
rect 32600 5012 32628 5111
rect 32766 5040 32772 5092
rect 32824 5080 32830 5092
rect 33410 5080 33416 5092
rect 32824 5052 33416 5080
rect 32824 5040 32830 5052
rect 33410 5040 33416 5052
rect 33468 5080 33474 5092
rect 33781 5083 33839 5089
rect 33781 5080 33793 5083
rect 33468 5052 33793 5080
rect 33468 5040 33474 5052
rect 33781 5049 33793 5052
rect 33827 5049 33839 5083
rect 36556 5080 36584 5120
rect 36906 5108 36912 5120
rect 36964 5148 36970 5160
rect 41230 5148 41236 5160
rect 36964 5120 41236 5148
rect 36964 5108 36970 5120
rect 41230 5108 41236 5120
rect 41288 5108 41294 5160
rect 41322 5108 41328 5160
rect 41380 5148 41386 5160
rect 41969 5151 42027 5157
rect 41969 5148 41981 5151
rect 41380 5120 41981 5148
rect 41380 5108 41386 5120
rect 41969 5117 41981 5120
rect 42015 5117 42027 5151
rect 41969 5111 42027 5117
rect 41782 5080 41788 5092
rect 36556 5052 41788 5080
rect 33781 5043 33839 5049
rect 41782 5040 41788 5052
rect 41840 5040 41846 5092
rect 42720 5080 42748 5188
rect 42978 5176 42984 5188
rect 43036 5176 43042 5228
rect 45922 5216 45928 5228
rect 45402 5188 45928 5216
rect 45922 5176 45928 5188
rect 45980 5176 45986 5228
rect 48130 5216 48136 5228
rect 48091 5188 48136 5216
rect 48130 5176 48136 5188
rect 48188 5176 48194 5228
rect 49436 5216 49464 5247
rect 49602 5244 49608 5256
rect 49660 5244 49666 5296
rect 49712 5256 51074 5284
rect 49712 5216 49740 5256
rect 50062 5216 50068 5228
rect 49436 5188 49740 5216
rect 50023 5188 50068 5216
rect 50062 5176 50068 5188
rect 50120 5176 50126 5228
rect 50154 5176 50160 5228
rect 50212 5216 50218 5228
rect 50893 5219 50951 5225
rect 50893 5216 50905 5219
rect 50212 5188 50905 5216
rect 50212 5176 50218 5188
rect 50893 5185 50905 5188
rect 50939 5185 50951 5219
rect 51046 5216 51074 5256
rect 51994 5244 52000 5296
rect 52052 5284 52058 5296
rect 52178 5284 52184 5296
rect 52052 5256 52184 5284
rect 52052 5244 52058 5256
rect 52178 5244 52184 5256
rect 52236 5244 52242 5296
rect 53561 5287 53619 5293
rect 53561 5253 53573 5287
rect 53607 5284 53619 5287
rect 53742 5284 53748 5296
rect 53607 5256 53748 5284
rect 53607 5253 53619 5256
rect 53561 5247 53619 5253
rect 53742 5244 53748 5256
rect 53800 5244 53806 5296
rect 55122 5244 55128 5296
rect 55180 5244 55186 5296
rect 55858 5284 55864 5296
rect 55819 5256 55864 5284
rect 55858 5244 55864 5256
rect 55916 5244 55922 5296
rect 56594 5244 56600 5296
rect 56652 5284 56658 5296
rect 57882 5284 57888 5296
rect 56652 5256 57888 5284
rect 56652 5244 56658 5256
rect 57882 5244 57888 5256
rect 57940 5284 57946 5296
rect 58161 5287 58219 5293
rect 58161 5284 58173 5287
rect 57940 5256 58173 5284
rect 57940 5244 57946 5256
rect 58161 5253 58173 5256
rect 58207 5284 58219 5287
rect 62298 5284 62304 5296
rect 58207 5256 60136 5284
rect 61962 5256 62304 5284
rect 58207 5253 58219 5256
rect 58161 5247 58219 5253
rect 53193 5219 53251 5225
rect 53193 5216 53205 5219
rect 51046 5188 53205 5216
rect 50893 5179 50951 5185
rect 53193 5185 53205 5188
rect 53239 5185 53251 5219
rect 53374 5216 53380 5228
rect 53335 5188 53380 5216
rect 53193 5179 53251 5185
rect 53374 5176 53380 5188
rect 53432 5176 53438 5228
rect 53466 5176 53472 5228
rect 53524 5216 53530 5228
rect 56778 5216 56784 5228
rect 53524 5188 53569 5216
rect 56739 5188 56784 5216
rect 53524 5176 53530 5188
rect 56778 5176 56784 5188
rect 56836 5176 56842 5228
rect 56965 5219 57023 5225
rect 56965 5185 56977 5219
rect 57011 5185 57023 5219
rect 56965 5179 57023 5185
rect 43070 5148 43076 5160
rect 43031 5120 43076 5148
rect 43070 5108 43076 5120
rect 43128 5108 43134 5160
rect 43990 5148 43996 5160
rect 43951 5120 43996 5148
rect 43990 5108 43996 5120
rect 44048 5108 44054 5160
rect 44358 5108 44364 5160
rect 44416 5148 44422 5160
rect 44416 5120 45968 5148
rect 44416 5108 44422 5120
rect 45738 5080 45744 5092
rect 42720 5052 43116 5080
rect 45699 5052 45744 5080
rect 30156 4984 32628 5012
rect 30156 4972 30162 4984
rect 34882 4972 34888 5024
rect 34940 5012 34946 5024
rect 38473 5015 38531 5021
rect 38473 5012 38485 5015
rect 34940 4984 38485 5012
rect 34940 4972 34946 4984
rect 38473 4981 38485 4984
rect 38519 5012 38531 5015
rect 39025 5015 39083 5021
rect 39025 5012 39037 5015
rect 38519 4984 39037 5012
rect 38519 4981 38531 4984
rect 38473 4975 38531 4981
rect 39025 4981 39037 4984
rect 39071 5012 39083 5015
rect 40310 5012 40316 5024
rect 39071 4984 40316 5012
rect 39071 4981 39083 4984
rect 39025 4975 39083 4981
rect 40310 4972 40316 4984
rect 40368 4972 40374 5024
rect 40954 4972 40960 5024
rect 41012 5012 41018 5024
rect 42058 5012 42064 5024
rect 41012 4984 42064 5012
rect 41012 4972 41018 4984
rect 42058 4972 42064 4984
rect 42116 4972 42122 5024
rect 42702 5012 42708 5024
rect 42663 4984 42708 5012
rect 42702 4972 42708 4984
rect 42760 4972 42766 5024
rect 43088 5012 43116 5052
rect 45738 5040 45744 5052
rect 45796 5040 45802 5092
rect 45940 5080 45968 5120
rect 47118 5108 47124 5160
rect 47176 5148 47182 5160
rect 48317 5151 48375 5157
rect 48317 5148 48329 5151
rect 47176 5120 48329 5148
rect 47176 5108 47182 5120
rect 48317 5117 48329 5120
rect 48363 5117 48375 5151
rect 48317 5111 48375 5117
rect 45940 5052 46980 5080
rect 45278 5012 45284 5024
rect 43088 4984 45284 5012
rect 45278 4972 45284 4984
rect 45336 4972 45342 5024
rect 46952 5021 46980 5052
rect 47670 5040 47676 5092
rect 47728 5080 47734 5092
rect 47765 5083 47823 5089
rect 47765 5080 47777 5083
rect 47728 5052 47777 5080
rect 47728 5040 47734 5052
rect 47765 5049 47777 5052
rect 47811 5049 47823 5083
rect 47765 5043 47823 5049
rect 46937 5015 46995 5021
rect 46937 4981 46949 5015
rect 46983 5012 46995 5015
rect 48222 5012 48228 5024
rect 46983 4984 48228 5012
rect 46983 4981 46995 4984
rect 46937 4975 46995 4981
rect 48222 4972 48228 4984
rect 48280 4972 48286 5024
rect 48332 5012 48360 5111
rect 48682 5108 48688 5160
rect 48740 5148 48746 5160
rect 50172 5148 50200 5176
rect 50338 5148 50344 5160
rect 48740 5120 50200 5148
rect 50299 5120 50344 5148
rect 48740 5108 48746 5120
rect 49252 5089 49280 5120
rect 50338 5108 50344 5120
rect 50396 5108 50402 5160
rect 51166 5148 51172 5160
rect 51127 5120 51172 5148
rect 51166 5108 51172 5120
rect 51224 5108 51230 5160
rect 55214 5148 55220 5160
rect 53668 5120 55220 5148
rect 49237 5083 49295 5089
rect 49237 5049 49249 5083
rect 49283 5049 49295 5083
rect 49602 5080 49608 5092
rect 49237 5043 49295 5049
rect 49344 5052 49608 5080
rect 49344 5012 49372 5052
rect 49602 5040 49608 5052
rect 49660 5040 49666 5092
rect 50157 5083 50215 5089
rect 50157 5049 50169 5083
rect 50203 5049 50215 5083
rect 50157 5043 50215 5049
rect 51077 5083 51135 5089
rect 51077 5049 51089 5083
rect 51123 5080 51135 5083
rect 53668 5080 53696 5120
rect 55214 5108 55220 5120
rect 55272 5108 55278 5160
rect 56134 5148 56140 5160
rect 56095 5120 56140 5148
rect 56134 5108 56140 5120
rect 56192 5108 56198 5160
rect 56980 5148 57008 5179
rect 57054 5176 57060 5228
rect 57112 5216 57118 5228
rect 57112 5188 57157 5216
rect 57112 5176 57118 5188
rect 57330 5176 57336 5228
rect 57388 5216 57394 5228
rect 57698 5216 57704 5228
rect 57388 5188 57704 5216
rect 57388 5176 57394 5188
rect 57698 5176 57704 5188
rect 57756 5216 57762 5228
rect 58069 5219 58127 5225
rect 58069 5216 58081 5219
rect 57756 5188 58081 5216
rect 57756 5176 57762 5188
rect 58069 5185 58081 5188
rect 58115 5216 58127 5219
rect 58115 5188 58204 5216
rect 58115 5185 58127 5188
rect 58069 5179 58127 5185
rect 58176 5148 58204 5188
rect 58342 5176 58348 5228
rect 58400 5216 58406 5228
rect 58400 5188 60044 5216
rect 58400 5176 58406 5188
rect 59446 5148 59452 5160
rect 56980 5120 58112 5148
rect 58176 5120 59452 5148
rect 51123 5052 53696 5080
rect 53745 5083 53803 5089
rect 51123 5049 51135 5052
rect 51077 5043 51135 5049
rect 53745 5049 53757 5083
rect 53791 5049 53803 5083
rect 54386 5080 54392 5092
rect 54347 5052 54392 5080
rect 53745 5043 53803 5049
rect 48332 4984 49372 5012
rect 49418 4972 49424 5024
rect 49476 5012 49482 5024
rect 49786 5012 49792 5024
rect 49476 4984 49792 5012
rect 49476 4972 49482 4984
rect 49786 4972 49792 4984
rect 49844 5012 49850 5024
rect 50172 5012 50200 5043
rect 49844 4984 50200 5012
rect 50249 5015 50307 5021
rect 49844 4972 49850 4984
rect 50249 4981 50261 5015
rect 50295 5012 50307 5015
rect 50985 5015 51043 5021
rect 50985 5012 50997 5015
rect 50295 4984 50997 5012
rect 50295 4981 50307 4984
rect 50249 4975 50307 4981
rect 50985 4981 50997 4984
rect 51031 4981 51043 5015
rect 50985 4975 51043 4981
rect 51721 5015 51779 5021
rect 51721 4981 51733 5015
rect 51767 5012 51779 5015
rect 51994 5012 52000 5024
rect 51767 4984 52000 5012
rect 51767 4981 51779 4984
rect 51721 4975 51779 4981
rect 51994 4972 52000 4984
rect 52052 4972 52058 5024
rect 53466 4972 53472 5024
rect 53524 5012 53530 5024
rect 53760 5012 53788 5043
rect 54386 5040 54392 5052
rect 54444 5040 54450 5092
rect 57330 5080 57336 5092
rect 56060 5052 57336 5080
rect 56060 5012 56088 5052
rect 57330 5040 57336 5052
rect 57388 5040 57394 5092
rect 58084 5089 58112 5120
rect 59446 5108 59452 5120
rect 59504 5108 59510 5160
rect 58069 5083 58127 5089
rect 58069 5049 58081 5083
rect 58115 5049 58127 5083
rect 58802 5080 58808 5092
rect 58763 5052 58808 5080
rect 58069 5043 58127 5049
rect 58802 5040 58808 5052
rect 58860 5040 58866 5092
rect 58986 5040 58992 5092
rect 59044 5080 59050 5092
rect 59909 5083 59967 5089
rect 59909 5080 59921 5083
rect 59044 5052 59921 5080
rect 59044 5040 59050 5052
rect 59909 5049 59921 5052
rect 59955 5049 59967 5083
rect 59909 5043 59967 5049
rect 53524 4984 56088 5012
rect 53524 4972 53530 4984
rect 56134 4972 56140 5024
rect 56192 5012 56198 5024
rect 56597 5015 56655 5021
rect 56597 5012 56609 5015
rect 56192 4984 56609 5012
rect 56192 4972 56198 4984
rect 56597 4981 56609 4984
rect 56643 4981 56655 5015
rect 56597 4975 56655 4981
rect 56686 4972 56692 5024
rect 56744 5012 56750 5024
rect 59078 5012 59084 5024
rect 56744 4984 59084 5012
rect 56744 4972 56750 4984
rect 59078 4972 59084 4984
rect 59136 4972 59142 5024
rect 59449 5015 59507 5021
rect 59449 4981 59461 5015
rect 59495 5012 59507 5015
rect 59814 5012 59820 5024
rect 59495 4984 59820 5012
rect 59495 4981 59507 4984
rect 59449 4975 59507 4981
rect 59814 4972 59820 4984
rect 59872 4972 59878 5024
rect 60016 5012 60044 5188
rect 60108 5080 60136 5256
rect 62298 5244 62304 5256
rect 62356 5244 62362 5296
rect 62390 5244 62396 5296
rect 62448 5284 62454 5296
rect 62448 5256 62493 5284
rect 62448 5244 62454 5256
rect 63310 5244 63316 5296
rect 63368 5284 63374 5296
rect 63773 5287 63831 5293
rect 63773 5284 63785 5287
rect 63368 5256 63785 5284
rect 63368 5244 63374 5256
rect 63773 5253 63785 5256
rect 63819 5253 63831 5287
rect 63773 5247 63831 5253
rect 64690 5244 64696 5296
rect 64748 5284 64754 5296
rect 64877 5287 64935 5293
rect 64877 5284 64889 5287
rect 64748 5256 64889 5284
rect 64748 5244 64754 5256
rect 64877 5253 64889 5256
rect 64923 5253 64935 5287
rect 64877 5247 64935 5253
rect 65886 5244 65892 5296
rect 65944 5284 65950 5296
rect 66349 5287 66407 5293
rect 66349 5284 66361 5287
rect 65944 5256 66361 5284
rect 65944 5244 65950 5256
rect 66349 5253 66361 5256
rect 66395 5253 66407 5287
rect 66349 5247 66407 5253
rect 67726 5244 67732 5296
rect 67784 5284 67790 5296
rect 68373 5287 68431 5293
rect 68373 5284 68385 5287
rect 67784 5256 68385 5284
rect 67784 5244 67790 5256
rect 68373 5253 68385 5256
rect 68419 5253 68431 5287
rect 70302 5284 70308 5296
rect 68373 5247 68431 5253
rect 69768 5256 70308 5284
rect 62669 5219 62727 5225
rect 62669 5185 62681 5219
rect 62715 5216 62727 5219
rect 63494 5216 63500 5228
rect 62715 5188 63500 5216
rect 62715 5185 62727 5188
rect 62669 5179 62727 5185
rect 63494 5176 63500 5188
rect 63552 5176 63558 5228
rect 64417 5219 64475 5225
rect 64417 5185 64429 5219
rect 64463 5216 64475 5219
rect 65334 5216 65340 5228
rect 64463 5188 65340 5216
rect 64463 5185 64475 5188
rect 64417 5179 64475 5185
rect 65334 5176 65340 5188
rect 65392 5176 65398 5228
rect 69768 5225 69796 5256
rect 70302 5244 70308 5256
rect 70360 5244 70366 5296
rect 71866 5284 71872 5296
rect 71254 5256 71872 5284
rect 71866 5244 71872 5256
rect 71924 5244 71930 5296
rect 72050 5244 72056 5296
rect 72108 5284 72114 5296
rect 73617 5287 73675 5293
rect 73617 5284 73629 5287
rect 72108 5256 73629 5284
rect 72108 5244 72114 5256
rect 73617 5253 73629 5256
rect 73663 5253 73675 5287
rect 76742 5284 76748 5296
rect 73617 5247 73675 5253
rect 75472 5256 76748 5284
rect 69753 5219 69811 5225
rect 69753 5185 69765 5219
rect 69799 5185 69811 5219
rect 69753 5179 69811 5185
rect 71774 5176 71780 5228
rect 71832 5216 71838 5228
rect 72421 5219 72479 5225
rect 72421 5216 72433 5219
rect 71832 5188 72433 5216
rect 71832 5176 71838 5188
rect 72421 5185 72433 5188
rect 72467 5185 72479 5219
rect 73709 5219 73767 5225
rect 73517 5209 73575 5215
rect 73517 5206 73529 5209
rect 72421 5179 72479 5185
rect 73448 5178 73529 5206
rect 60458 5108 60464 5160
rect 60516 5148 60522 5160
rect 60516 5120 62620 5148
rect 60516 5108 60522 5120
rect 62592 5080 62620 5120
rect 63862 5108 63868 5160
rect 63920 5148 63926 5160
rect 66901 5151 66959 5157
rect 66901 5148 66913 5151
rect 63920 5120 66913 5148
rect 63920 5108 63926 5120
rect 66901 5117 66913 5120
rect 66947 5148 66959 5151
rect 69201 5151 69259 5157
rect 69201 5148 69213 5151
rect 66947 5120 69213 5148
rect 66947 5117 66959 5120
rect 66901 5111 66959 5117
rect 69201 5117 69213 5120
rect 69247 5148 69259 5151
rect 69290 5148 69296 5160
rect 69247 5120 69296 5148
rect 69247 5117 69259 5120
rect 69201 5111 69259 5117
rect 69290 5108 69296 5120
rect 69348 5108 69354 5160
rect 70029 5151 70087 5157
rect 70029 5117 70041 5151
rect 70075 5148 70087 5151
rect 70075 5120 72096 5148
rect 70075 5117 70087 5120
rect 70029 5111 70087 5117
rect 63221 5083 63279 5089
rect 63221 5080 63233 5083
rect 60108 5052 61424 5080
rect 62592 5052 63233 5080
rect 60826 5012 60832 5024
rect 60016 4984 60832 5012
rect 60826 4972 60832 4984
rect 60884 5012 60890 5024
rect 60921 5015 60979 5021
rect 60921 5012 60933 5015
rect 60884 4984 60933 5012
rect 60884 4972 60890 4984
rect 60921 4981 60933 4984
rect 60967 4981 60979 5015
rect 61396 5012 61424 5052
rect 63221 5049 63233 5052
rect 63267 5049 63279 5083
rect 63221 5043 63279 5049
rect 64414 5040 64420 5092
rect 64472 5080 64478 5092
rect 65429 5083 65487 5089
rect 65429 5080 65441 5083
rect 64472 5052 65441 5080
rect 64472 5040 64478 5052
rect 65429 5049 65441 5052
rect 65475 5080 65487 5083
rect 71501 5083 71559 5089
rect 65475 5052 67634 5080
rect 65475 5049 65487 5052
rect 65429 5043 65487 5049
rect 63678 5012 63684 5024
rect 61396 4984 63684 5012
rect 60921 4975 60979 4981
rect 63678 4972 63684 4984
rect 63736 4972 63742 5024
rect 67606 5012 67634 5052
rect 71501 5049 71513 5083
rect 71547 5080 71559 5083
rect 71774 5080 71780 5092
rect 71547 5052 71780 5080
rect 71547 5049 71559 5052
rect 71501 5043 71559 5049
rect 71774 5040 71780 5052
rect 71832 5040 71838 5092
rect 72068 5089 72096 5120
rect 72142 5108 72148 5160
rect 72200 5148 72206 5160
rect 72329 5151 72387 5157
rect 72329 5148 72341 5151
rect 72200 5120 72341 5148
rect 72200 5108 72206 5120
rect 72329 5117 72341 5120
rect 72375 5117 72387 5151
rect 72329 5111 72387 5117
rect 72053 5083 72111 5089
rect 72053 5049 72065 5083
rect 72099 5049 72111 5083
rect 73448 5080 73476 5178
rect 73517 5175 73529 5178
rect 73563 5175 73575 5209
rect 73709 5185 73721 5219
rect 73755 5216 73767 5219
rect 73798 5216 73804 5228
rect 73755 5188 73804 5216
rect 73755 5185 73767 5188
rect 73709 5179 73767 5185
rect 73798 5176 73804 5188
rect 73856 5176 73862 5228
rect 73982 5176 73988 5228
rect 74040 5216 74046 5228
rect 74169 5219 74227 5225
rect 74169 5216 74181 5219
rect 74040 5188 74181 5216
rect 74040 5176 74046 5188
rect 74169 5185 74181 5188
rect 74215 5185 74227 5219
rect 74169 5179 74227 5185
rect 74353 5219 74411 5225
rect 74353 5185 74365 5219
rect 74399 5185 74411 5219
rect 74353 5179 74411 5185
rect 73517 5169 73575 5175
rect 74368 5148 74396 5179
rect 74442 5176 74448 5228
rect 74500 5216 74506 5228
rect 74500 5188 75224 5216
rect 74500 5176 74506 5188
rect 75196 5157 75224 5188
rect 75270 5176 75276 5228
rect 75328 5216 75334 5228
rect 75472 5225 75500 5256
rect 76742 5244 76748 5256
rect 76800 5244 76806 5296
rect 80164 5246 80192 5324
rect 81986 5312 81992 5324
rect 82044 5312 82050 5364
rect 85390 5312 85396 5364
rect 85448 5352 85454 5364
rect 86954 5352 86960 5364
rect 85448 5324 86960 5352
rect 85448 5312 85454 5324
rect 86954 5312 86960 5324
rect 87012 5352 87018 5364
rect 87690 5352 87696 5364
rect 87012 5324 87696 5352
rect 87012 5312 87018 5324
rect 87690 5312 87696 5324
rect 87748 5312 87754 5364
rect 90634 5352 90640 5364
rect 90595 5324 90640 5352
rect 90634 5312 90640 5324
rect 90692 5312 90698 5364
rect 91002 5312 91008 5364
rect 91060 5352 91066 5364
rect 91281 5355 91339 5361
rect 91281 5352 91293 5355
rect 91060 5324 91293 5352
rect 91060 5312 91066 5324
rect 91281 5321 91293 5324
rect 91327 5352 91339 5355
rect 91830 5352 91836 5364
rect 91327 5324 91836 5352
rect 91327 5321 91339 5324
rect 91281 5315 91339 5321
rect 91830 5312 91836 5324
rect 91888 5352 91894 5364
rect 93670 5352 93676 5364
rect 91888 5324 93676 5352
rect 91888 5312 91894 5324
rect 93670 5312 93676 5324
rect 93728 5312 93734 5364
rect 94038 5312 94044 5364
rect 94096 5352 94102 5364
rect 94133 5355 94191 5361
rect 94133 5352 94145 5355
rect 94096 5324 94145 5352
rect 94096 5312 94102 5324
rect 94133 5321 94145 5324
rect 94179 5321 94191 5355
rect 94133 5315 94191 5321
rect 75457 5219 75515 5225
rect 75328 5188 75373 5216
rect 75328 5176 75334 5188
rect 75457 5185 75469 5219
rect 75503 5185 75515 5219
rect 75457 5179 75515 5185
rect 75822 5176 75828 5228
rect 75880 5216 75886 5228
rect 76009 5219 76067 5225
rect 76009 5216 76021 5219
rect 75880 5188 76021 5216
rect 75880 5176 75886 5188
rect 76009 5185 76021 5188
rect 76055 5185 76067 5219
rect 76009 5179 76067 5185
rect 76193 5219 76251 5225
rect 76193 5185 76205 5219
rect 76239 5185 76251 5219
rect 76193 5179 76251 5185
rect 74997 5151 75055 5157
rect 74997 5148 75009 5151
rect 74368 5120 75009 5148
rect 74997 5117 75009 5120
rect 75043 5117 75055 5151
rect 74997 5111 75055 5117
rect 75181 5151 75239 5157
rect 75181 5117 75193 5151
rect 75227 5117 75239 5151
rect 75181 5111 75239 5117
rect 75365 5151 75423 5157
rect 75365 5117 75377 5151
rect 75411 5148 75423 5151
rect 75914 5148 75920 5160
rect 75411 5120 75920 5148
rect 75411 5117 75423 5120
rect 75365 5111 75423 5117
rect 73522 5080 73528 5092
rect 73448 5052 73528 5080
rect 72053 5043 72111 5049
rect 73522 5040 73528 5052
rect 73580 5080 73586 5092
rect 75380 5080 75408 5111
rect 75914 5108 75920 5120
rect 75972 5108 75978 5160
rect 76208 5148 76236 5179
rect 76282 5176 76288 5228
rect 76340 5216 76346 5228
rect 76653 5219 76711 5225
rect 76653 5216 76665 5219
rect 76340 5188 76665 5216
rect 76340 5176 76346 5188
rect 76653 5185 76665 5188
rect 76699 5185 76711 5219
rect 76834 5216 76840 5228
rect 76795 5188 76840 5216
rect 76653 5179 76711 5185
rect 76834 5176 76840 5188
rect 76892 5176 76898 5228
rect 76926 5176 76932 5228
rect 76984 5216 76990 5228
rect 77573 5219 77631 5225
rect 77573 5216 77585 5219
rect 76984 5188 77585 5216
rect 76984 5176 76990 5188
rect 77573 5185 77585 5188
rect 77619 5185 77631 5219
rect 77573 5179 77631 5185
rect 77662 5176 77668 5228
rect 77720 5216 77726 5228
rect 79229 5219 79287 5225
rect 77720 5188 77765 5216
rect 77720 5176 77726 5188
rect 79229 5185 79241 5219
rect 79275 5216 79287 5219
rect 80072 5218 80192 5246
rect 80606 5244 80612 5296
rect 80664 5284 80670 5296
rect 80664 5256 81466 5284
rect 80664 5244 80670 5256
rect 84010 5244 84016 5296
rect 84068 5284 84074 5296
rect 84657 5287 84715 5293
rect 84657 5284 84669 5287
rect 84068 5256 84669 5284
rect 84068 5244 84074 5256
rect 84657 5253 84669 5256
rect 84703 5284 84715 5287
rect 92014 5284 92020 5296
rect 84703 5256 92020 5284
rect 84703 5253 84715 5256
rect 84657 5247 84715 5253
rect 92014 5244 92020 5256
rect 92072 5244 92078 5296
rect 84381 5219 84439 5225
rect 80072 5216 80100 5218
rect 79275 5188 80100 5216
rect 79275 5185 79287 5188
rect 79229 5179 79287 5185
rect 84381 5185 84393 5219
rect 84427 5216 84439 5219
rect 84930 5216 84936 5228
rect 84427 5188 84936 5216
rect 84427 5185 84439 5188
rect 84381 5179 84439 5185
rect 76944 5148 76972 5176
rect 76208 5120 76972 5148
rect 77849 5151 77907 5157
rect 77849 5117 77861 5151
rect 77895 5148 77907 5151
rect 78030 5148 78036 5160
rect 77895 5120 78036 5148
rect 77895 5117 77907 5120
rect 77849 5111 77907 5117
rect 78030 5108 78036 5120
rect 78088 5108 78094 5160
rect 79137 5151 79195 5157
rect 79137 5117 79149 5151
rect 79183 5117 79195 5151
rect 79137 5111 79195 5117
rect 73580 5052 75408 5080
rect 73580 5040 73586 5052
rect 75454 5040 75460 5092
rect 75512 5080 75518 5092
rect 76101 5083 76159 5089
rect 76101 5080 76113 5083
rect 75512 5052 76113 5080
rect 75512 5040 75518 5052
rect 76101 5049 76113 5052
rect 76147 5049 76159 5083
rect 76101 5043 76159 5049
rect 77757 5083 77815 5089
rect 77757 5049 77769 5083
rect 77803 5080 77815 5083
rect 79152 5080 79180 5111
rect 77803 5052 79180 5080
rect 77803 5049 77815 5052
rect 77757 5043 77815 5049
rect 69842 5012 69848 5024
rect 67606 4984 69848 5012
rect 69842 4972 69848 4984
rect 69900 4972 69906 5024
rect 74258 5012 74264 5024
rect 74219 4984 74264 5012
rect 74258 4972 74264 4984
rect 74316 4972 74322 5024
rect 75822 4972 75828 5024
rect 75880 5012 75886 5024
rect 79244 5012 79272 5179
rect 84930 5176 84936 5188
rect 84988 5176 84994 5228
rect 85390 5176 85396 5228
rect 85448 5216 85454 5228
rect 85448 5188 85493 5216
rect 85448 5176 85454 5188
rect 85666 5176 85672 5228
rect 85724 5216 85730 5228
rect 86037 5219 86095 5225
rect 86037 5216 86049 5219
rect 85724 5188 86049 5216
rect 85724 5176 85730 5188
rect 86037 5185 86049 5188
rect 86083 5216 86095 5219
rect 86586 5216 86592 5228
rect 86083 5188 86592 5216
rect 86083 5185 86095 5188
rect 86037 5179 86095 5185
rect 86586 5176 86592 5188
rect 86644 5216 86650 5228
rect 87049 5219 87107 5225
rect 87049 5216 87061 5219
rect 86644 5188 87061 5216
rect 86644 5176 86650 5188
rect 87049 5185 87061 5188
rect 87095 5216 87107 5219
rect 87690 5216 87696 5228
rect 87095 5188 87552 5216
rect 87651 5188 87696 5216
rect 87095 5185 87107 5188
rect 87049 5179 87107 5185
rect 80238 5148 80244 5160
rect 79612 5120 80244 5148
rect 79612 5089 79640 5120
rect 80238 5108 80244 5120
rect 80296 5108 80302 5160
rect 80701 5151 80759 5157
rect 80701 5117 80713 5151
rect 80747 5117 80759 5151
rect 80974 5148 80980 5160
rect 80935 5120 80980 5148
rect 80701 5111 80759 5117
rect 79597 5083 79655 5089
rect 79597 5049 79609 5083
rect 79643 5049 79655 5083
rect 79597 5043 79655 5049
rect 75880 4984 79272 5012
rect 75880 4972 75886 4984
rect 80146 4972 80152 5024
rect 80204 5012 80210 5024
rect 80716 5012 80744 5111
rect 80974 5108 80980 5120
rect 81032 5108 81038 5160
rect 81434 5108 81440 5160
rect 81492 5148 81498 5160
rect 84562 5148 84568 5160
rect 81492 5120 82492 5148
rect 84523 5120 84568 5148
rect 81492 5108 81498 5120
rect 82464 5089 82492 5120
rect 84562 5108 84568 5120
rect 84620 5108 84626 5160
rect 86313 5151 86371 5157
rect 86313 5117 86325 5151
rect 86359 5148 86371 5151
rect 86773 5151 86831 5157
rect 86773 5148 86785 5151
rect 86359 5120 86785 5148
rect 86359 5117 86371 5120
rect 86313 5111 86371 5117
rect 86773 5117 86785 5120
rect 86819 5117 86831 5151
rect 87524 5148 87552 5188
rect 87690 5176 87696 5188
rect 87748 5176 87754 5228
rect 90177 5219 90235 5225
rect 90177 5216 90189 5219
rect 89686 5188 90189 5216
rect 89686 5148 89714 5188
rect 90177 5185 90189 5188
rect 90223 5216 90235 5219
rect 92382 5216 92388 5228
rect 90223 5188 92388 5216
rect 90223 5185 90235 5188
rect 90177 5179 90235 5185
rect 92382 5176 92388 5188
rect 92440 5176 92446 5228
rect 93026 5216 93032 5228
rect 92987 5188 93032 5216
rect 93026 5176 93032 5188
rect 93084 5176 93090 5228
rect 87524 5120 89714 5148
rect 86773 5111 86831 5117
rect 82449 5083 82507 5089
rect 82449 5049 82461 5083
rect 82495 5080 82507 5083
rect 82495 5052 84700 5080
rect 82495 5049 82507 5052
rect 82449 5043 82507 5049
rect 84672 5024 84700 5052
rect 81434 5012 81440 5024
rect 80204 4984 80249 5012
rect 80716 4984 81440 5012
rect 80204 4972 80210 4984
rect 81434 4972 81440 4984
rect 81492 5012 81498 5024
rect 82170 5012 82176 5024
rect 81492 4984 82176 5012
rect 81492 4972 81498 4984
rect 82170 4972 82176 4984
rect 82228 4972 82234 5024
rect 83093 5015 83151 5021
rect 83093 4981 83105 5015
rect 83139 5012 83151 5015
rect 83366 5012 83372 5024
rect 83139 4984 83372 5012
rect 83139 4981 83151 4984
rect 83093 4975 83151 4981
rect 83366 4972 83372 4984
rect 83424 4972 83430 5024
rect 84194 5012 84200 5024
rect 84155 4984 84200 5012
rect 84194 4972 84200 4984
rect 84252 4972 84258 5024
rect 84654 5012 84660 5024
rect 84615 4984 84660 5012
rect 84654 4972 84660 4984
rect 84712 4972 84718 5024
rect 85114 5012 85120 5024
rect 85075 4984 85120 5012
rect 85114 4972 85120 4984
rect 85172 4972 85178 5024
rect 86788 5012 86816 5111
rect 91278 5108 91284 5160
rect 91336 5148 91342 5160
rect 92109 5151 92167 5157
rect 92109 5148 92121 5151
rect 91336 5120 92121 5148
rect 91336 5108 91342 5120
rect 92109 5117 92121 5120
rect 92155 5117 92167 5151
rect 92109 5111 92167 5117
rect 88076 5052 91508 5080
rect 88076 5024 88104 5052
rect 87046 5012 87052 5024
rect 86788 4984 87052 5012
rect 87046 4972 87052 4984
rect 87104 5012 87110 5024
rect 87874 5012 87880 5024
rect 87104 4984 87880 5012
rect 87104 4972 87110 4984
rect 87874 4972 87880 4984
rect 87932 4972 87938 5024
rect 87969 5015 88027 5021
rect 87969 4981 87981 5015
rect 88015 5012 88027 5015
rect 88058 5012 88064 5024
rect 88015 4984 88064 5012
rect 88015 4981 88027 4984
rect 87969 4975 88027 4981
rect 88058 4972 88064 4984
rect 88116 4972 88122 5024
rect 88978 5012 88984 5024
rect 88939 4984 88984 5012
rect 88978 4972 88984 4984
rect 89036 5012 89042 5024
rect 89346 5012 89352 5024
rect 89036 4984 89352 5012
rect 89036 4972 89042 4984
rect 89346 4972 89352 4984
rect 89404 5012 89410 5024
rect 89533 5015 89591 5021
rect 89533 5012 89545 5015
rect 89404 4984 89545 5012
rect 89404 4972 89410 4984
rect 89533 4981 89545 4984
rect 89579 5012 89591 5015
rect 91002 5012 91008 5024
rect 89579 4984 91008 5012
rect 89579 4981 89591 4984
rect 89533 4975 89591 4981
rect 91002 4972 91008 4984
rect 91060 4972 91066 5024
rect 91480 5012 91508 5052
rect 93305 5015 93363 5021
rect 93305 5012 93317 5015
rect 91480 4984 93317 5012
rect 93305 4981 93317 4984
rect 93351 4981 93363 5015
rect 93305 4975 93363 4981
rect 1104 4922 94852 4944
rect 1104 4870 12668 4922
rect 12720 4870 12732 4922
rect 12784 4870 12796 4922
rect 12848 4870 12860 4922
rect 12912 4870 12924 4922
rect 12976 4870 36105 4922
rect 36157 4870 36169 4922
rect 36221 4870 36233 4922
rect 36285 4870 36297 4922
rect 36349 4870 36361 4922
rect 36413 4870 59542 4922
rect 59594 4870 59606 4922
rect 59658 4870 59670 4922
rect 59722 4870 59734 4922
rect 59786 4870 59798 4922
rect 59850 4870 82979 4922
rect 83031 4870 83043 4922
rect 83095 4870 83107 4922
rect 83159 4870 83171 4922
rect 83223 4870 83235 4922
rect 83287 4870 94852 4922
rect 1104 4848 94852 4870
rect 4338 4768 4344 4820
rect 4396 4808 4402 4820
rect 8481 4811 8539 4817
rect 8481 4808 8493 4811
rect 4396 4780 8493 4808
rect 4396 4768 4402 4780
rect 8481 4777 8493 4780
rect 8527 4808 8539 4811
rect 22830 4808 22836 4820
rect 8527 4780 12434 4808
rect 22791 4780 22836 4808
rect 8527 4777 8539 4780
rect 8481 4771 8539 4777
rect 6730 4672 6736 4684
rect 6691 4644 6736 4672
rect 6730 4632 6736 4644
rect 6788 4632 6794 4684
rect 7006 4672 7012 4684
rect 6967 4644 7012 4672
rect 7006 4632 7012 4644
rect 7064 4632 7070 4684
rect 8386 4604 8392 4616
rect 8142 4576 8392 4604
rect 8386 4564 8392 4576
rect 8444 4604 8450 4616
rect 9122 4604 9128 4616
rect 8444 4576 9128 4604
rect 8444 4564 8450 4576
rect 9122 4564 9128 4576
rect 9180 4564 9186 4616
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4604 9459 4607
rect 9858 4604 9864 4616
rect 9447 4576 9864 4604
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 9858 4564 9864 4576
rect 9916 4564 9922 4616
rect 10137 4607 10195 4613
rect 10137 4573 10149 4607
rect 10183 4604 10195 4607
rect 10594 4604 10600 4616
rect 10183 4576 10600 4604
rect 10183 4573 10195 4576
rect 10137 4567 10195 4573
rect 10594 4564 10600 4576
rect 10652 4564 10658 4616
rect 12406 4604 12434 4780
rect 22830 4768 22836 4780
rect 22888 4768 22894 4820
rect 23382 4768 23388 4820
rect 23440 4808 23446 4820
rect 26326 4808 26332 4820
rect 23440 4780 26332 4808
rect 23440 4768 23446 4780
rect 26326 4768 26332 4780
rect 26384 4768 26390 4820
rect 26510 4808 26516 4820
rect 26471 4780 26516 4808
rect 26510 4768 26516 4780
rect 26568 4768 26574 4820
rect 27246 4768 27252 4820
rect 27304 4808 27310 4820
rect 29733 4811 29791 4817
rect 29733 4808 29745 4811
rect 27304 4780 29745 4808
rect 27304 4768 27310 4780
rect 29733 4777 29745 4780
rect 29779 4777 29791 4811
rect 29733 4771 29791 4777
rect 31110 4768 31116 4820
rect 31168 4808 31174 4820
rect 34882 4808 34888 4820
rect 31168 4780 34888 4808
rect 31168 4768 31174 4780
rect 34882 4768 34888 4780
rect 34940 4768 34946 4820
rect 37734 4808 37740 4820
rect 34992 4780 37740 4808
rect 22373 4743 22431 4749
rect 22373 4709 22385 4743
rect 22419 4740 22431 4743
rect 23477 4743 23535 4749
rect 23477 4740 23489 4743
rect 22419 4712 23489 4740
rect 22419 4709 22431 4712
rect 22373 4703 22431 4709
rect 23477 4709 23489 4712
rect 23523 4740 23535 4743
rect 24210 4740 24216 4752
rect 23523 4712 24216 4740
rect 23523 4709 23535 4712
rect 23477 4703 23535 4709
rect 24210 4700 24216 4712
rect 24268 4700 24274 4752
rect 25501 4743 25559 4749
rect 25501 4709 25513 4743
rect 25547 4740 25559 4743
rect 30098 4740 30104 4752
rect 25547 4712 30104 4740
rect 25547 4709 25559 4712
rect 25501 4703 25559 4709
rect 30098 4700 30104 4712
rect 30156 4700 30162 4752
rect 33594 4740 33600 4752
rect 31220 4712 33600 4740
rect 23106 4632 23112 4684
rect 23164 4672 23170 4684
rect 24670 4672 24676 4684
rect 23164 4644 24676 4672
rect 23164 4632 23170 4644
rect 24670 4632 24676 4644
rect 24728 4632 24734 4684
rect 24854 4632 24860 4684
rect 24912 4672 24918 4684
rect 31220 4672 31248 4712
rect 33594 4700 33600 4712
rect 33652 4700 33658 4752
rect 34992 4749 35020 4780
rect 37734 4768 37740 4780
rect 37792 4768 37798 4820
rect 38105 4811 38163 4817
rect 38105 4777 38117 4811
rect 38151 4808 38163 4811
rect 38151 4780 41736 4808
rect 38151 4777 38163 4780
rect 38105 4771 38163 4777
rect 33689 4743 33747 4749
rect 33689 4709 33701 4743
rect 33735 4740 33747 4743
rect 34977 4743 35035 4749
rect 33735 4712 33916 4740
rect 33735 4709 33747 4712
rect 33689 4703 33747 4709
rect 24912 4644 31248 4672
rect 31297 4675 31355 4681
rect 24912 4632 24918 4644
rect 31297 4641 31309 4675
rect 31343 4672 31355 4675
rect 33410 4672 33416 4684
rect 31343 4644 33416 4672
rect 31343 4641 31355 4644
rect 31297 4635 31355 4641
rect 33410 4632 33416 4644
rect 33468 4632 33474 4684
rect 14369 4607 14427 4613
rect 14369 4604 14381 4607
rect 12406 4576 14381 4604
rect 14369 4573 14381 4576
rect 14415 4573 14427 4607
rect 14369 4567 14427 4573
rect 14458 4564 14464 4616
rect 14516 4604 14522 4616
rect 14553 4607 14611 4613
rect 14553 4604 14565 4607
rect 14516 4576 14565 4604
rect 14516 4564 14522 4576
rect 14553 4573 14565 4576
rect 14599 4573 14611 4607
rect 14553 4567 14611 4573
rect 23658 4564 23664 4616
rect 23716 4604 23722 4616
rect 25038 4604 25044 4616
rect 23716 4576 25044 4604
rect 23716 4564 23722 4576
rect 25038 4564 25044 4576
rect 25096 4564 25102 4616
rect 25130 4564 25136 4616
rect 25188 4604 25194 4616
rect 25317 4607 25375 4613
rect 25188 4576 25233 4604
rect 25188 4564 25194 4576
rect 25317 4573 25329 4607
rect 25363 4604 25375 4607
rect 25682 4604 25688 4616
rect 25363 4600 25452 4604
rect 25608 4600 25688 4604
rect 25363 4576 25688 4600
rect 25363 4573 25375 4576
rect 25317 4567 25375 4573
rect 25424 4572 25636 4576
rect 25682 4564 25688 4576
rect 25740 4564 25746 4616
rect 27801 4607 27859 4613
rect 27801 4573 27813 4607
rect 27847 4604 27859 4607
rect 29822 4604 29828 4616
rect 27847 4576 29828 4604
rect 27847 4573 27859 4576
rect 27801 4567 27859 4573
rect 29822 4564 29828 4576
rect 29880 4564 29886 4616
rect 29917 4607 29975 4613
rect 29917 4573 29929 4607
rect 29963 4604 29975 4607
rect 30834 4604 30840 4616
rect 29963 4576 30840 4604
rect 29963 4573 29975 4576
rect 29917 4567 29975 4573
rect 30834 4564 30840 4576
rect 30892 4564 30898 4616
rect 33888 4604 33916 4712
rect 34977 4709 34989 4743
rect 35023 4709 35035 4743
rect 39022 4740 39028 4752
rect 38983 4712 39028 4740
rect 34977 4703 35035 4709
rect 33965 4675 34023 4681
rect 33965 4641 33977 4675
rect 34011 4672 34023 4675
rect 34992 4672 35020 4703
rect 39022 4700 39028 4712
rect 39080 4700 39086 4752
rect 41708 4740 41736 4780
rect 41782 4768 41788 4820
rect 41840 4808 41846 4820
rect 47673 4811 47731 4817
rect 41840 4780 47624 4808
rect 41840 4768 41846 4780
rect 42978 4740 42984 4752
rect 41708 4712 42984 4740
rect 42978 4700 42984 4712
rect 43036 4700 43042 4752
rect 43346 4740 43352 4752
rect 43307 4712 43352 4740
rect 43346 4700 43352 4712
rect 43404 4700 43410 4752
rect 44361 4743 44419 4749
rect 44361 4709 44373 4743
rect 44407 4740 44419 4743
rect 44450 4740 44456 4752
rect 44407 4712 44456 4740
rect 44407 4709 44419 4712
rect 44361 4703 44419 4709
rect 44450 4700 44456 4712
rect 44508 4700 44514 4752
rect 44910 4700 44916 4752
rect 44968 4740 44974 4752
rect 45189 4743 45247 4749
rect 45189 4740 45201 4743
rect 44968 4712 45201 4740
rect 44968 4700 44974 4712
rect 45189 4709 45201 4712
rect 45235 4740 45247 4743
rect 46937 4743 46995 4749
rect 46937 4740 46949 4743
rect 45235 4712 46949 4740
rect 45235 4709 45247 4712
rect 45189 4703 45247 4709
rect 46937 4709 46949 4712
rect 46983 4740 46995 4743
rect 46983 4712 47532 4740
rect 46983 4709 46995 4712
rect 46937 4703 46995 4709
rect 34011 4644 35020 4672
rect 36633 4675 36691 4681
rect 34011 4641 34023 4644
rect 33965 4635 34023 4641
rect 36633 4641 36645 4675
rect 36679 4672 36691 4675
rect 42702 4672 42708 4684
rect 36679 4644 42708 4672
rect 36679 4641 36691 4644
rect 36633 4635 36691 4641
rect 42702 4632 42708 4644
rect 42760 4632 42766 4684
rect 45830 4632 45836 4684
rect 45888 4672 45894 4684
rect 47504 4681 47532 4712
rect 45925 4675 45983 4681
rect 45925 4672 45937 4675
rect 45888 4644 45937 4672
rect 45888 4632 45894 4644
rect 45925 4641 45937 4644
rect 45971 4641 45983 4675
rect 45925 4635 45983 4641
rect 47489 4675 47547 4681
rect 47489 4641 47501 4675
rect 47535 4641 47547 4675
rect 47596 4672 47624 4780
rect 47673 4777 47685 4811
rect 47719 4808 47731 4811
rect 48130 4808 48136 4820
rect 47719 4780 48136 4808
rect 47719 4777 47731 4780
rect 47673 4771 47731 4777
rect 48130 4768 48136 4780
rect 48188 4808 48194 4820
rect 49145 4811 49203 4817
rect 49145 4808 49157 4811
rect 48188 4780 49157 4808
rect 48188 4768 48194 4780
rect 49145 4777 49157 4780
rect 49191 4777 49203 4811
rect 49145 4771 49203 4777
rect 49602 4768 49608 4820
rect 49660 4808 49666 4820
rect 50338 4808 50344 4820
rect 49660 4780 50344 4808
rect 49660 4768 49666 4780
rect 50338 4768 50344 4780
rect 50396 4768 50402 4820
rect 50614 4768 50620 4820
rect 50672 4808 50678 4820
rect 50893 4811 50951 4817
rect 50893 4808 50905 4811
rect 50672 4780 50905 4808
rect 50672 4768 50678 4780
rect 50893 4777 50905 4780
rect 50939 4777 50951 4811
rect 50893 4771 50951 4777
rect 52362 4768 52368 4820
rect 52420 4808 52426 4820
rect 52457 4811 52515 4817
rect 52457 4808 52469 4811
rect 52420 4780 52469 4808
rect 52420 4768 52426 4780
rect 52457 4777 52469 4780
rect 52503 4777 52515 4811
rect 53742 4808 53748 4820
rect 53655 4780 53748 4808
rect 52457 4771 52515 4777
rect 53742 4768 53748 4780
rect 53800 4768 53806 4820
rect 53926 4768 53932 4820
rect 53984 4808 53990 4820
rect 54757 4811 54815 4817
rect 54757 4808 54769 4811
rect 53984 4780 54769 4808
rect 53984 4768 53990 4780
rect 54757 4777 54769 4780
rect 54803 4777 54815 4811
rect 56594 4808 56600 4820
rect 54757 4771 54815 4777
rect 54864 4780 56600 4808
rect 50062 4700 50068 4752
rect 50120 4740 50126 4752
rect 53377 4743 53435 4749
rect 53377 4740 53389 4743
rect 50120 4712 53389 4740
rect 50120 4700 50126 4712
rect 53377 4709 53389 4712
rect 53423 4709 53435 4743
rect 53377 4703 53435 4709
rect 53558 4700 53564 4752
rect 53616 4740 53622 4752
rect 53760 4740 53788 4768
rect 54864 4740 54892 4780
rect 56594 4768 56600 4780
rect 56652 4768 56658 4820
rect 56873 4811 56931 4817
rect 56873 4777 56885 4811
rect 56919 4808 56931 4811
rect 57054 4808 57060 4820
rect 56919 4780 57060 4808
rect 56919 4777 56931 4780
rect 56873 4771 56931 4777
rect 57054 4768 57060 4780
rect 57112 4768 57118 4820
rect 58158 4768 58164 4820
rect 58216 4808 58222 4820
rect 59173 4811 59231 4817
rect 59173 4808 59185 4811
rect 58216 4780 59185 4808
rect 58216 4768 58222 4780
rect 59173 4777 59185 4780
rect 59219 4777 59231 4811
rect 59173 4771 59231 4777
rect 60737 4811 60795 4817
rect 60737 4777 60749 4811
rect 60783 4808 60795 4811
rect 61286 4808 61292 4820
rect 60783 4780 61292 4808
rect 60783 4777 60795 4780
rect 60737 4771 60795 4777
rect 58069 4743 58127 4749
rect 58069 4740 58081 4743
rect 53616 4712 53696 4740
rect 53760 4712 54892 4740
rect 55784 4712 58081 4740
rect 53616 4700 53622 4712
rect 49970 4672 49976 4684
rect 47596 4644 49976 4672
rect 47489 4635 47547 4641
rect 49970 4632 49976 4644
rect 50028 4632 50034 4684
rect 36357 4607 36415 4613
rect 33888 4576 35388 4604
rect 35360 4548 35388 4576
rect 36357 4573 36369 4607
rect 36403 4573 36415 4607
rect 40402 4604 40408 4616
rect 40363 4576 40408 4604
rect 36357 4567 36415 4573
rect 22554 4496 22560 4548
rect 22612 4536 22618 4548
rect 23290 4536 23296 4548
rect 22612 4508 23296 4536
rect 22612 4496 22618 4508
rect 23290 4496 23296 4508
rect 23348 4536 23354 4548
rect 23348 4508 24072 4536
rect 23348 4496 23354 4508
rect 10318 4468 10324 4480
rect 10279 4440 10324 4468
rect 10318 4428 10324 4440
rect 10376 4428 10382 4480
rect 10686 4428 10692 4480
rect 10744 4468 10750 4480
rect 10781 4471 10839 4477
rect 10781 4468 10793 4471
rect 10744 4440 10793 4468
rect 10744 4428 10750 4440
rect 10781 4437 10793 4440
rect 10827 4437 10839 4471
rect 15378 4468 15384 4480
rect 15339 4440 15384 4468
rect 10781 4431 10839 4437
rect 15378 4428 15384 4440
rect 15436 4428 15442 4480
rect 22830 4428 22836 4480
rect 22888 4468 22894 4480
rect 23937 4471 23995 4477
rect 23937 4468 23949 4471
rect 22888 4440 23949 4468
rect 22888 4428 22894 4440
rect 23937 4437 23949 4440
rect 23983 4437 23995 4471
rect 24044 4468 24072 4508
rect 24302 4496 24308 4548
rect 24360 4536 24366 4548
rect 31110 4536 31116 4548
rect 24360 4508 31116 4536
rect 24360 4496 24366 4508
rect 31110 4496 31116 4508
rect 31168 4496 31174 4548
rect 31386 4536 31392 4548
rect 31347 4508 31392 4536
rect 31386 4496 31392 4508
rect 31444 4496 31450 4548
rect 32306 4536 32312 4548
rect 32267 4508 32312 4536
rect 32306 4496 32312 4508
rect 32364 4496 32370 4548
rect 35342 4536 35348 4548
rect 33428 4508 35020 4536
rect 35303 4508 35348 4536
rect 26142 4468 26148 4480
rect 24044 4440 26148 4468
rect 23937 4431 23995 4437
rect 26142 4428 26148 4440
rect 26200 4428 26206 4480
rect 26326 4428 26332 4480
rect 26384 4468 26390 4480
rect 33428 4468 33456 4508
rect 26384 4440 33456 4468
rect 33505 4471 33563 4477
rect 26384 4428 26390 4440
rect 33505 4437 33517 4471
rect 33551 4468 33563 4471
rect 33594 4468 33600 4480
rect 33551 4440 33600 4468
rect 33551 4437 33563 4440
rect 33505 4431 33563 4437
rect 33594 4428 33600 4440
rect 33652 4428 33658 4480
rect 34606 4428 34612 4480
rect 34664 4468 34670 4480
rect 34885 4471 34943 4477
rect 34885 4468 34897 4471
rect 34664 4440 34897 4468
rect 34664 4428 34670 4440
rect 34885 4437 34897 4440
rect 34931 4437 34943 4471
rect 34992 4468 35020 4508
rect 35342 4496 35348 4508
rect 35400 4496 35406 4548
rect 36372 4536 36400 4567
rect 40402 4564 40408 4576
rect 40460 4564 40466 4616
rect 41782 4564 41788 4616
rect 41840 4604 41846 4616
rect 42518 4604 42524 4616
rect 41840 4576 42524 4604
rect 41840 4564 41846 4576
rect 42518 4564 42524 4576
rect 42576 4564 42582 4616
rect 46017 4607 46075 4613
rect 46017 4573 46029 4607
rect 46063 4604 46075 4607
rect 47118 4604 47124 4616
rect 46063 4576 47124 4604
rect 46063 4573 46075 4576
rect 46017 4567 46075 4573
rect 47118 4564 47124 4576
rect 47176 4564 47182 4616
rect 47762 4604 47768 4616
rect 47723 4576 47768 4604
rect 47762 4564 47768 4576
rect 47820 4564 47826 4616
rect 49237 4607 49295 4613
rect 49237 4573 49249 4607
rect 49283 4604 49295 4607
rect 50080 4604 50108 4700
rect 50433 4675 50491 4681
rect 50433 4641 50445 4675
rect 50479 4672 50491 4675
rect 52270 4672 52276 4684
rect 50479 4644 52276 4672
rect 50479 4641 50491 4644
rect 50433 4635 50491 4641
rect 52270 4632 52276 4644
rect 52328 4632 52334 4684
rect 53668 4681 53696 4712
rect 53653 4675 53711 4681
rect 53653 4641 53665 4675
rect 53699 4641 53711 4675
rect 53653 4635 53711 4641
rect 51994 4604 52000 4616
rect 49283 4576 50108 4604
rect 51955 4576 52000 4604
rect 49283 4573 49295 4576
rect 49237 4567 49295 4573
rect 51994 4564 52000 4576
rect 52052 4564 52058 4616
rect 53466 4564 53472 4616
rect 53524 4604 53530 4616
rect 53561 4607 53619 4613
rect 53561 4604 53573 4607
rect 53524 4576 53573 4604
rect 53524 4564 53530 4576
rect 53561 4573 53573 4576
rect 53607 4573 53619 4607
rect 53668 4604 53696 4635
rect 54941 4607 54999 4613
rect 53668 4576 54892 4604
rect 53561 4567 53619 4573
rect 36906 4536 36912 4548
rect 36372 4508 36912 4536
rect 36906 4496 36912 4508
rect 36964 4496 36970 4548
rect 37918 4536 37924 4548
rect 37831 4508 37924 4536
rect 37918 4496 37924 4508
rect 37976 4536 37982 4548
rect 38470 4536 38476 4548
rect 37976 4508 38476 4536
rect 37976 4496 37982 4508
rect 38470 4496 38476 4508
rect 38528 4496 38534 4548
rect 40678 4536 40684 4548
rect 40639 4508 40684 4536
rect 40678 4496 40684 4508
rect 40736 4496 40742 4548
rect 42613 4539 42671 4545
rect 42613 4536 42625 4539
rect 41984 4508 42625 4536
rect 38010 4468 38016 4480
rect 34992 4440 38016 4468
rect 34885 4431 34943 4437
rect 38010 4428 38016 4440
rect 38068 4428 38074 4480
rect 40034 4428 40040 4480
rect 40092 4468 40098 4480
rect 41984 4468 42012 4508
rect 42613 4505 42625 4508
rect 42659 4505 42671 4539
rect 47394 4536 47400 4548
rect 42613 4499 42671 4505
rect 46400 4508 47400 4536
rect 42150 4468 42156 4480
rect 40092 4440 42012 4468
rect 42111 4440 42156 4468
rect 40092 4428 40098 4440
rect 42150 4428 42156 4440
rect 42208 4428 42214 4480
rect 42518 4428 42524 4480
rect 42576 4468 42582 4480
rect 43806 4468 43812 4480
rect 42576 4440 43812 4468
rect 42576 4428 42582 4440
rect 43806 4428 43812 4440
rect 43864 4468 43870 4480
rect 45922 4468 45928 4480
rect 43864 4440 45928 4468
rect 43864 4428 43870 4440
rect 45922 4428 45928 4440
rect 45980 4428 45986 4480
rect 46400 4477 46428 4508
rect 47394 4496 47400 4508
rect 47452 4496 47458 4548
rect 49786 4536 49792 4548
rect 49699 4508 49792 4536
rect 49786 4496 49792 4508
rect 49844 4536 49850 4548
rect 51534 4536 51540 4548
rect 49844 4508 51540 4536
rect 49844 4496 49850 4508
rect 51534 4496 51540 4508
rect 51592 4496 51598 4548
rect 53374 4496 53380 4548
rect 53432 4536 53438 4548
rect 53837 4539 53895 4545
rect 53837 4536 53849 4539
rect 53432 4508 53849 4536
rect 53432 4496 53438 4508
rect 53837 4505 53849 4508
rect 53883 4505 53895 4539
rect 54864 4536 54892 4576
rect 54941 4573 54953 4607
rect 54987 4604 54999 4607
rect 55784 4604 55812 4712
rect 58069 4709 58081 4712
rect 58115 4709 58127 4743
rect 60752 4740 60780 4771
rect 61286 4768 61292 4780
rect 61344 4768 61350 4820
rect 62393 4811 62451 4817
rect 62393 4777 62405 4811
rect 62439 4808 62451 4811
rect 63494 4808 63500 4820
rect 62439 4780 63500 4808
rect 62439 4777 62451 4780
rect 62393 4771 62451 4777
rect 63494 4768 63500 4780
rect 63552 4768 63558 4820
rect 63678 4768 63684 4820
rect 63736 4808 63742 4820
rect 65889 4811 65947 4817
rect 65889 4808 65901 4811
rect 63736 4780 65901 4808
rect 63736 4768 63742 4780
rect 65889 4777 65901 4780
rect 65935 4777 65947 4811
rect 65889 4771 65947 4777
rect 71682 4768 71688 4820
rect 71740 4808 71746 4820
rect 73246 4808 73252 4820
rect 71740 4780 73252 4808
rect 71740 4768 71746 4780
rect 73246 4768 73252 4780
rect 73304 4768 73310 4820
rect 73614 4808 73620 4820
rect 73575 4780 73620 4808
rect 73614 4768 73620 4780
rect 73672 4808 73678 4820
rect 74353 4811 74411 4817
rect 74353 4808 74365 4811
rect 73672 4780 74365 4808
rect 73672 4768 73678 4780
rect 74353 4777 74365 4780
rect 74399 4777 74411 4811
rect 76190 4808 76196 4820
rect 76151 4780 76196 4808
rect 74353 4771 74411 4777
rect 76190 4768 76196 4780
rect 76248 4768 76254 4820
rect 77478 4768 77484 4820
rect 77536 4808 77542 4820
rect 77941 4811 77999 4817
rect 77941 4808 77953 4811
rect 77536 4780 77953 4808
rect 77536 4768 77542 4780
rect 77941 4777 77953 4780
rect 77987 4808 77999 4811
rect 77987 4780 79548 4808
rect 77987 4777 77999 4780
rect 77941 4771 77999 4777
rect 61194 4740 61200 4752
rect 58069 4703 58127 4709
rect 58452 4712 60780 4740
rect 61155 4712 61200 4740
rect 56134 4672 56140 4684
rect 56095 4644 56140 4672
rect 56134 4632 56140 4644
rect 56192 4632 56198 4684
rect 58342 4672 58348 4684
rect 57072 4644 58348 4672
rect 54987 4576 55812 4604
rect 56018 4607 56076 4613
rect 56018 4580 56030 4607
rect 54987 4573 54999 4576
rect 54941 4567 54999 4573
rect 55968 4573 56030 4580
rect 56064 4604 56076 4607
rect 56410 4604 56416 4616
rect 56064 4576 56416 4604
rect 56064 4573 56088 4576
rect 55968 4552 56088 4573
rect 56410 4564 56416 4576
rect 56468 4564 56474 4616
rect 55858 4536 55864 4548
rect 54864 4508 55864 4536
rect 53837 4499 53895 4505
rect 46385 4471 46443 4477
rect 46385 4437 46397 4471
rect 46431 4437 46443 4471
rect 47486 4468 47492 4480
rect 47447 4440 47492 4468
rect 46385 4431 46443 4437
rect 47486 4428 47492 4440
rect 47544 4428 47550 4480
rect 47578 4428 47584 4480
rect 47636 4468 47642 4480
rect 49418 4468 49424 4480
rect 47636 4440 49424 4468
rect 47636 4428 47642 4440
rect 49418 4428 49424 4440
rect 49476 4428 49482 4480
rect 53852 4468 53880 4499
rect 55858 4496 55864 4508
rect 55916 4496 55922 4548
rect 55968 4468 55996 4552
rect 56134 4496 56140 4548
rect 56192 4536 56198 4548
rect 57072 4545 57100 4644
rect 58342 4632 58348 4644
rect 58400 4632 58406 4684
rect 57238 4604 57244 4616
rect 57199 4576 57244 4604
rect 57238 4564 57244 4576
rect 57296 4564 57302 4616
rect 57330 4564 57336 4616
rect 57388 4604 57394 4616
rect 58452 4604 58480 4712
rect 61194 4700 61200 4712
rect 61252 4700 61258 4752
rect 62945 4743 63003 4749
rect 62945 4709 62957 4743
rect 62991 4740 63003 4743
rect 64690 4740 64696 4752
rect 62991 4712 64696 4740
rect 62991 4709 63003 4712
rect 62945 4703 63003 4709
rect 64690 4700 64696 4712
rect 64748 4700 64754 4752
rect 65153 4743 65211 4749
rect 65153 4709 65165 4743
rect 65199 4740 65211 4743
rect 65334 4740 65340 4752
rect 65199 4712 65340 4740
rect 65199 4709 65211 4712
rect 65153 4703 65211 4709
rect 65334 4700 65340 4712
rect 65392 4700 65398 4752
rect 72237 4743 72295 4749
rect 72237 4740 72249 4743
rect 69400 4712 72249 4740
rect 58526 4632 58532 4684
rect 58584 4672 58590 4684
rect 59906 4672 59912 4684
rect 58584 4644 59912 4672
rect 58584 4632 58590 4644
rect 59906 4632 59912 4644
rect 59964 4672 59970 4684
rect 61749 4675 61807 4681
rect 61749 4672 61761 4675
rect 59964 4644 61761 4672
rect 59964 4632 59970 4644
rect 61749 4641 61761 4644
rect 61795 4672 61807 4675
rect 63497 4675 63555 4681
rect 61795 4644 63448 4672
rect 61795 4641 61807 4644
rect 61749 4635 61807 4641
rect 58710 4604 58716 4616
rect 57388 4576 58480 4604
rect 58671 4576 58716 4604
rect 57388 4564 57394 4576
rect 58710 4564 58716 4576
rect 58768 4564 58774 4616
rect 59078 4564 59084 4616
rect 59136 4604 59142 4616
rect 59725 4607 59783 4613
rect 59725 4604 59737 4607
rect 59136 4576 59737 4604
rect 59136 4564 59142 4576
rect 59725 4573 59737 4576
rect 59771 4604 59783 4607
rect 62942 4604 62948 4616
rect 59771 4576 62948 4604
rect 59771 4573 59783 4576
rect 59725 4567 59783 4573
rect 62942 4564 62948 4576
rect 63000 4564 63006 4616
rect 63420 4604 63448 4644
rect 63497 4641 63509 4675
rect 63543 4672 63555 4675
rect 63586 4672 63592 4684
rect 63543 4644 63592 4672
rect 63543 4641 63555 4644
rect 63497 4635 63555 4641
rect 63586 4632 63592 4644
rect 63644 4632 63650 4684
rect 64046 4672 64052 4684
rect 64007 4644 64052 4672
rect 64046 4632 64052 4644
rect 64104 4632 64110 4684
rect 64414 4632 64420 4684
rect 64472 4672 64478 4684
rect 64509 4675 64567 4681
rect 64509 4672 64521 4675
rect 64472 4644 64521 4672
rect 64472 4632 64478 4644
rect 64509 4641 64521 4644
rect 64555 4641 64567 4675
rect 67358 4672 67364 4684
rect 67319 4644 67364 4672
rect 64509 4635 64567 4641
rect 67358 4632 67364 4644
rect 67416 4632 67422 4684
rect 67634 4632 67640 4684
rect 67692 4672 67698 4684
rect 68097 4675 68155 4681
rect 68097 4672 68109 4675
rect 67692 4644 68109 4672
rect 67692 4632 67698 4644
rect 68097 4641 68109 4644
rect 68143 4641 68155 4675
rect 68097 4635 68155 4641
rect 68373 4675 68431 4681
rect 68373 4641 68385 4675
rect 68419 4672 68431 4675
rect 69400 4672 69428 4712
rect 72237 4709 72249 4712
rect 72283 4709 72295 4743
rect 72237 4703 72295 4709
rect 73798 4700 73804 4752
rect 73856 4740 73862 4752
rect 74442 4740 74448 4752
rect 73856 4712 74448 4740
rect 73856 4700 73862 4712
rect 74442 4700 74448 4712
rect 74500 4740 74506 4752
rect 74537 4743 74595 4749
rect 74537 4740 74549 4743
rect 74500 4712 74549 4740
rect 74500 4700 74506 4712
rect 74537 4709 74549 4712
rect 74583 4740 74595 4743
rect 76466 4740 76472 4752
rect 74583 4712 76472 4740
rect 74583 4709 74595 4712
rect 74537 4703 74595 4709
rect 76466 4700 76472 4712
rect 76524 4700 76530 4752
rect 77849 4743 77907 4749
rect 77849 4740 77861 4743
rect 77036 4712 77861 4740
rect 68419 4644 69428 4672
rect 69845 4675 69903 4681
rect 68419 4641 68431 4644
rect 68373 4635 68431 4641
rect 69845 4641 69857 4675
rect 69891 4672 69903 4675
rect 71685 4675 71743 4681
rect 69891 4644 71636 4672
rect 69891 4641 69903 4644
rect 69845 4635 69903 4641
rect 63862 4604 63868 4616
rect 63420 4576 63868 4604
rect 63862 4564 63868 4576
rect 63920 4564 63926 4616
rect 71515 4607 71573 4613
rect 71515 4573 71527 4607
rect 71561 4573 71573 4607
rect 71608 4604 71636 4644
rect 71685 4641 71697 4675
rect 71731 4672 71743 4675
rect 72050 4672 72056 4684
rect 71731 4644 72056 4672
rect 71731 4641 71743 4644
rect 71685 4635 71743 4641
rect 72050 4632 72056 4644
rect 72108 4632 72114 4684
rect 72697 4675 72755 4681
rect 72697 4641 72709 4675
rect 72743 4672 72755 4675
rect 74258 4672 74264 4684
rect 72743 4644 74264 4672
rect 72743 4641 72755 4644
rect 72697 4635 72755 4641
rect 74258 4632 74264 4644
rect 74316 4632 74322 4684
rect 74626 4632 74632 4684
rect 74684 4672 74690 4684
rect 75089 4675 75147 4681
rect 75089 4672 75101 4675
rect 74684 4644 75101 4672
rect 74684 4632 74690 4644
rect 75089 4641 75101 4644
rect 75135 4672 75147 4675
rect 76374 4672 76380 4684
rect 75135 4644 76380 4672
rect 75135 4641 75147 4644
rect 75089 4635 75147 4641
rect 76374 4632 76380 4644
rect 76432 4632 76438 4684
rect 77036 4681 77064 4712
rect 77849 4709 77861 4712
rect 77895 4709 77907 4743
rect 78030 4740 78036 4752
rect 77849 4703 77907 4709
rect 77956 4712 78036 4740
rect 77021 4675 77079 4681
rect 77021 4641 77033 4675
rect 77067 4641 77079 4675
rect 77021 4635 77079 4641
rect 77757 4675 77815 4681
rect 77757 4641 77769 4675
rect 77803 4672 77815 4675
rect 77956 4672 77984 4712
rect 78030 4700 78036 4712
rect 78088 4700 78094 4752
rect 77803 4644 77984 4672
rect 78048 4644 79272 4672
rect 77803 4641 77815 4644
rect 77757 4635 77815 4641
rect 72605 4607 72663 4613
rect 72605 4604 72617 4607
rect 71608 4576 72617 4604
rect 71515 4567 71573 4573
rect 72605 4573 72617 4576
rect 72651 4604 72663 4607
rect 73246 4604 73252 4616
rect 72651 4576 73252 4604
rect 72651 4573 72663 4576
rect 72605 4567 72663 4573
rect 57057 4539 57115 4545
rect 57057 4536 57069 4539
rect 56192 4508 57069 4536
rect 56192 4496 56198 4508
rect 57057 4505 57069 4508
rect 57103 4505 57115 4539
rect 57698 4536 57704 4548
rect 57659 4508 57704 4536
rect 57057 4499 57115 4505
rect 57698 4496 57704 4508
rect 57756 4496 57762 4548
rect 57882 4536 57888 4548
rect 57843 4508 57888 4536
rect 57882 4496 57888 4508
rect 57940 4536 57946 4548
rect 57940 4508 58572 4536
rect 57940 4496 57946 4508
rect 53852 4440 55996 4468
rect 56413 4471 56471 4477
rect 56413 4437 56425 4471
rect 56459 4468 56471 4471
rect 57790 4468 57796 4480
rect 56459 4440 57796 4468
rect 56459 4437 56471 4440
rect 56413 4431 56471 4437
rect 57790 4428 57796 4440
rect 57848 4428 57854 4480
rect 58544 4477 58572 4508
rect 66806 4496 66812 4548
rect 66864 4496 66870 4548
rect 67726 4496 67732 4548
rect 67784 4536 67790 4548
rect 71530 4536 71558 4567
rect 73246 4564 73252 4576
rect 73304 4564 73310 4616
rect 73430 4604 73436 4616
rect 73391 4576 73436 4604
rect 73430 4564 73436 4576
rect 73488 4564 73494 4616
rect 73522 4564 73528 4616
rect 73580 4604 73586 4616
rect 76926 4604 76932 4616
rect 73580 4576 73625 4604
rect 74184 4576 76932 4604
rect 73580 4564 73586 4576
rect 74184 4548 74212 4576
rect 76926 4564 76932 4576
rect 76984 4564 76990 4616
rect 78048 4613 78076 4644
rect 78033 4607 78091 4613
rect 78033 4604 78045 4607
rect 77220 4576 78045 4604
rect 73706 4536 73712 4548
rect 67784 4508 68862 4536
rect 71530 4508 72740 4536
rect 73667 4508 73712 4536
rect 67784 4496 67790 4508
rect 58529 4471 58587 4477
rect 58529 4437 58541 4471
rect 58575 4437 58587 4471
rect 58529 4431 58587 4437
rect 71225 4471 71283 4477
rect 71225 4437 71237 4471
rect 71271 4468 71283 4471
rect 71590 4468 71596 4480
rect 71271 4440 71596 4468
rect 71271 4437 71283 4440
rect 71225 4431 71283 4437
rect 71590 4428 71596 4440
rect 71648 4428 71654 4480
rect 72712 4468 72740 4508
rect 73706 4496 73712 4508
rect 73764 4496 73770 4548
rect 74166 4536 74172 4548
rect 74079 4508 74172 4536
rect 74166 4496 74172 4508
rect 74224 4496 74230 4548
rect 74385 4539 74443 4545
rect 74385 4505 74397 4539
rect 74431 4536 74443 4539
rect 77220 4536 77248 4576
rect 78033 4573 78045 4576
rect 78079 4573 78091 4607
rect 78033 4567 78091 4573
rect 78493 4607 78551 4613
rect 78493 4573 78505 4607
rect 78539 4573 78551 4607
rect 78493 4567 78551 4573
rect 78677 4607 78735 4613
rect 78677 4573 78689 4607
rect 78723 4604 78735 4607
rect 78723 4576 79180 4604
rect 78723 4573 78735 4576
rect 78677 4567 78735 4573
rect 78398 4536 78404 4548
rect 74431 4508 77248 4536
rect 77312 4508 78404 4536
rect 74431 4505 74443 4508
rect 74385 4499 74443 4505
rect 73522 4468 73528 4480
rect 72712 4440 73528 4468
rect 73522 4428 73528 4440
rect 73580 4428 73586 4480
rect 77312 4477 77340 4508
rect 78398 4496 78404 4508
rect 78456 4496 78462 4548
rect 78508 4536 78536 4567
rect 78766 4536 78772 4548
rect 78508 4508 78772 4536
rect 77297 4471 77355 4477
rect 77297 4437 77309 4471
rect 77343 4437 77355 4471
rect 77297 4431 77355 4437
rect 77386 4428 77392 4480
rect 77444 4468 77450 4480
rect 78508 4468 78536 4508
rect 78766 4496 78772 4508
rect 78824 4496 78830 4548
rect 77444 4440 78536 4468
rect 78585 4471 78643 4477
rect 77444 4428 77450 4440
rect 78585 4437 78597 4471
rect 78631 4468 78643 4471
rect 78674 4468 78680 4480
rect 78631 4440 78680 4468
rect 78631 4437 78643 4440
rect 78585 4431 78643 4437
rect 78674 4428 78680 4440
rect 78732 4428 78738 4480
rect 79152 4477 79180 4576
rect 79244 4536 79272 4644
rect 79520 4613 79548 4780
rect 79870 4768 79876 4820
rect 79928 4808 79934 4820
rect 82446 4808 82452 4820
rect 79928 4780 82452 4808
rect 79928 4768 79934 4780
rect 82446 4768 82452 4780
rect 82504 4768 82510 4820
rect 83200 4780 83964 4808
rect 79781 4675 79839 4681
rect 79781 4641 79793 4675
rect 79827 4672 79839 4675
rect 79962 4672 79968 4684
rect 79827 4644 79968 4672
rect 79827 4641 79839 4644
rect 79781 4635 79839 4641
rect 79962 4632 79968 4644
rect 80020 4632 80026 4684
rect 79505 4607 79563 4613
rect 79505 4573 79517 4607
rect 79551 4573 79563 4607
rect 79505 4567 79563 4573
rect 80698 4564 80704 4616
rect 80756 4604 80762 4616
rect 81253 4607 81311 4613
rect 81253 4604 81265 4607
rect 80756 4576 81265 4604
rect 80756 4564 80762 4576
rect 81253 4573 81265 4576
rect 81299 4573 81311 4607
rect 81526 4604 81532 4616
rect 81487 4576 81532 4604
rect 81253 4567 81311 4573
rect 79597 4539 79655 4545
rect 79597 4536 79609 4539
rect 79244 4508 79609 4536
rect 79597 4505 79609 4508
rect 79643 4505 79655 4539
rect 79597 4499 79655 4505
rect 79137 4471 79195 4477
rect 79137 4437 79149 4471
rect 79183 4437 79195 4471
rect 79612 4468 79640 4499
rect 79686 4496 79692 4548
rect 79744 4536 79750 4548
rect 80333 4539 80391 4545
rect 80333 4536 80345 4539
rect 79744 4508 80345 4536
rect 79744 4496 79750 4508
rect 80333 4505 80345 4508
rect 80379 4505 80391 4539
rect 81268 4536 81296 4567
rect 81526 4564 81532 4576
rect 81584 4564 81590 4616
rect 82265 4607 82323 4613
rect 82265 4573 82277 4607
rect 82311 4604 82323 4607
rect 82722 4604 82728 4616
rect 82311 4576 82728 4604
rect 82311 4573 82323 4576
rect 82265 4567 82323 4573
rect 82722 4564 82728 4576
rect 82780 4604 82786 4616
rect 83200 4604 83228 4780
rect 83936 4740 83964 4780
rect 84286 4768 84292 4820
rect 84344 4808 84350 4820
rect 85025 4811 85083 4817
rect 85025 4808 85037 4811
rect 84344 4780 85037 4808
rect 84344 4768 84350 4780
rect 85025 4777 85037 4780
rect 85071 4777 85083 4811
rect 87046 4808 87052 4820
rect 85025 4771 85083 4777
rect 86788 4780 87052 4808
rect 84378 4740 84384 4752
rect 83936 4712 84384 4740
rect 84378 4700 84384 4712
rect 84436 4700 84442 4752
rect 84930 4700 84936 4752
rect 84988 4740 84994 4752
rect 85850 4740 85856 4752
rect 84988 4712 85856 4740
rect 84988 4700 84994 4712
rect 85850 4700 85856 4712
rect 85908 4700 85914 4752
rect 86678 4672 86684 4684
rect 84028 4644 86684 4672
rect 83366 4604 83372 4616
rect 82780 4576 83228 4604
rect 83327 4576 83372 4604
rect 82780 4564 82786 4576
rect 83366 4564 83372 4576
rect 83424 4564 83430 4616
rect 83642 4604 83648 4616
rect 83603 4576 83648 4604
rect 83642 4564 83648 4576
rect 83700 4564 83706 4616
rect 83734 4564 83740 4616
rect 83792 4604 83798 4616
rect 84028 4604 84056 4644
rect 86678 4632 86684 4644
rect 86736 4632 86742 4684
rect 86788 4681 86816 4780
rect 87046 4768 87052 4780
rect 87104 4768 87110 4820
rect 87138 4768 87144 4820
rect 87196 4808 87202 4820
rect 87969 4811 88027 4817
rect 87969 4808 87981 4811
rect 87196 4780 87981 4808
rect 87196 4768 87202 4780
rect 87969 4777 87981 4780
rect 88015 4808 88027 4811
rect 88058 4808 88064 4820
rect 88015 4780 88064 4808
rect 88015 4777 88027 4780
rect 87969 4771 88027 4777
rect 88058 4768 88064 4780
rect 88116 4768 88122 4820
rect 89686 4780 89852 4808
rect 89686 4740 89714 4780
rect 87432 4712 89714 4740
rect 86773 4675 86831 4681
rect 86773 4641 86785 4675
rect 86819 4641 86831 4675
rect 86773 4635 86831 4641
rect 84378 4604 84384 4616
rect 83792 4576 84056 4604
rect 84339 4576 84384 4604
rect 83792 4564 83798 4576
rect 84378 4564 84384 4576
rect 84436 4564 84442 4616
rect 84654 4564 84660 4616
rect 84712 4604 84718 4616
rect 85669 4607 85727 4613
rect 85669 4604 85681 4607
rect 84712 4576 85681 4604
rect 84712 4564 84718 4576
rect 85669 4573 85681 4576
rect 85715 4573 85727 4607
rect 85850 4604 85856 4616
rect 85811 4576 85856 4604
rect 85669 4567 85727 4573
rect 81710 4536 81716 4548
rect 81268 4508 81716 4536
rect 80333 4499 80391 4505
rect 81710 4496 81716 4508
rect 81768 4496 81774 4548
rect 83826 4536 83832 4548
rect 82372 4508 83832 4536
rect 82372 4468 82400 4508
rect 83826 4496 83832 4508
rect 83884 4496 83890 4548
rect 85684 4536 85712 4567
rect 85850 4564 85856 4576
rect 85908 4564 85914 4616
rect 86586 4564 86592 4616
rect 86644 4604 86650 4616
rect 87049 4607 87107 4613
rect 87049 4604 87061 4607
rect 86644 4576 87061 4604
rect 86644 4564 86650 4576
rect 87049 4573 87061 4576
rect 87095 4604 87107 4607
rect 87230 4604 87236 4616
rect 87095 4576 87236 4604
rect 87095 4573 87107 4576
rect 87049 4567 87107 4573
rect 87230 4564 87236 4576
rect 87288 4564 87294 4616
rect 87432 4536 87460 4712
rect 88518 4672 88524 4684
rect 88479 4644 88524 4672
rect 88518 4632 88524 4644
rect 88576 4632 88582 4684
rect 87690 4604 87696 4616
rect 87651 4576 87696 4604
rect 87690 4564 87696 4576
rect 87748 4564 87754 4616
rect 88610 4604 88616 4616
rect 88571 4576 88616 4604
rect 88610 4564 88616 4576
rect 88668 4564 88674 4616
rect 89824 4548 89852 4780
rect 93213 4743 93271 4749
rect 93213 4740 93225 4743
rect 90560 4712 93225 4740
rect 90560 4613 90588 4712
rect 93213 4709 93225 4712
rect 93259 4709 93271 4743
rect 93213 4703 93271 4709
rect 91005 4675 91063 4681
rect 91005 4641 91017 4675
rect 91051 4672 91063 4675
rect 91925 4675 91983 4681
rect 91925 4672 91937 4675
rect 91051 4644 91937 4672
rect 91051 4641 91063 4644
rect 91005 4635 91063 4641
rect 91925 4641 91937 4644
rect 91971 4641 91983 4675
rect 91925 4635 91983 4641
rect 90545 4607 90603 4613
rect 90545 4573 90557 4607
rect 90591 4573 90603 4607
rect 90818 4604 90824 4616
rect 90779 4576 90824 4604
rect 90545 4567 90603 4573
rect 90818 4564 90824 4576
rect 90876 4564 90882 4616
rect 92014 4604 92020 4616
rect 91975 4576 92020 4604
rect 92014 4564 92020 4576
rect 92072 4564 92078 4616
rect 93029 4607 93087 4613
rect 93029 4604 93041 4607
rect 92216 4576 93041 4604
rect 85684 4508 87460 4536
rect 88886 4496 88892 4548
rect 88944 4536 88950 4548
rect 89441 4539 89499 4545
rect 89441 4536 89453 4539
rect 88944 4508 89453 4536
rect 88944 4496 88950 4508
rect 89441 4505 89453 4508
rect 89487 4505 89499 4539
rect 89622 4536 89628 4548
rect 89583 4508 89628 4536
rect 89441 4499 89499 4505
rect 79612 4440 82400 4468
rect 79137 4431 79195 4437
rect 82446 4428 82452 4480
rect 82504 4468 82510 4480
rect 84565 4471 84623 4477
rect 84565 4468 84577 4471
rect 82504 4440 84577 4468
rect 82504 4428 82510 4440
rect 84565 4437 84577 4440
rect 84611 4468 84623 4471
rect 85114 4468 85120 4480
rect 84611 4440 85120 4468
rect 84611 4437 84623 4440
rect 84565 4431 84623 4437
rect 85114 4428 85120 4440
rect 85172 4428 85178 4480
rect 85853 4471 85911 4477
rect 85853 4437 85865 4471
rect 85899 4468 85911 4471
rect 87046 4468 87052 4480
rect 85899 4440 87052 4468
rect 85899 4437 85911 4440
rect 85853 4431 85911 4437
rect 87046 4428 87052 4440
rect 87104 4428 87110 4480
rect 88981 4471 89039 4477
rect 88981 4437 88993 4471
rect 89027 4468 89039 4471
rect 89346 4468 89352 4480
rect 89027 4440 89352 4468
rect 89027 4437 89039 4440
rect 88981 4431 89039 4437
rect 89346 4428 89352 4440
rect 89404 4428 89410 4480
rect 89456 4468 89484 4499
rect 89622 4496 89628 4508
rect 89680 4496 89686 4548
rect 89806 4536 89812 4548
rect 89767 4508 89812 4536
rect 89806 4496 89812 4508
rect 89864 4496 89870 4548
rect 92106 4536 92112 4548
rect 90192 4508 92112 4536
rect 90192 4468 90220 4508
rect 92106 4496 92112 4508
rect 92164 4496 92170 4548
rect 89456 4440 90220 4468
rect 90266 4428 90272 4480
rect 90324 4468 90330 4480
rect 90637 4471 90695 4477
rect 90637 4468 90649 4471
rect 90324 4440 90649 4468
rect 90324 4428 90330 4440
rect 90637 4437 90649 4440
rect 90683 4437 90695 4471
rect 90637 4431 90695 4437
rect 90910 4428 90916 4480
rect 90968 4468 90974 4480
rect 92216 4468 92244 4576
rect 93029 4573 93041 4576
rect 93075 4573 93087 4607
rect 93029 4567 93087 4573
rect 92290 4496 92296 4548
rect 92348 4536 92354 4548
rect 92845 4539 92903 4545
rect 92845 4536 92857 4539
rect 92348 4508 92857 4536
rect 92348 4496 92354 4508
rect 92845 4505 92857 4508
rect 92891 4505 92903 4539
rect 92845 4499 92903 4505
rect 90968 4440 92244 4468
rect 92385 4471 92443 4477
rect 90968 4428 90974 4440
rect 92385 4437 92397 4471
rect 92431 4468 92443 4471
rect 93118 4468 93124 4480
rect 92431 4440 93124 4468
rect 92431 4437 92443 4440
rect 92385 4431 92443 4437
rect 93118 4428 93124 4440
rect 93176 4428 93182 4480
rect 93670 4468 93676 4480
rect 93631 4440 93676 4468
rect 93670 4428 93676 4440
rect 93728 4428 93734 4480
rect 94222 4468 94228 4480
rect 94183 4440 94228 4468
rect 94222 4428 94228 4440
rect 94280 4428 94286 4480
rect 1104 4378 95011 4400
rect 1104 4326 24386 4378
rect 24438 4326 24450 4378
rect 24502 4326 24514 4378
rect 24566 4326 24578 4378
rect 24630 4326 24642 4378
rect 24694 4326 47823 4378
rect 47875 4326 47887 4378
rect 47939 4326 47951 4378
rect 48003 4326 48015 4378
rect 48067 4326 48079 4378
rect 48131 4326 71260 4378
rect 71312 4326 71324 4378
rect 71376 4326 71388 4378
rect 71440 4326 71452 4378
rect 71504 4326 71516 4378
rect 71568 4326 94697 4378
rect 94749 4326 94761 4378
rect 94813 4326 94825 4378
rect 94877 4326 94889 4378
rect 94941 4326 94953 4378
rect 95005 4326 95011 4378
rect 1104 4304 95011 4326
rect 15378 4224 15384 4276
rect 15436 4264 15442 4276
rect 31386 4264 31392 4276
rect 15436 4236 31392 4264
rect 15436 4224 15442 4236
rect 31386 4224 31392 4236
rect 31444 4224 31450 4276
rect 34425 4267 34483 4273
rect 34425 4264 34437 4267
rect 33428 4236 34437 4264
rect 33428 4208 33456 4236
rect 34425 4233 34437 4236
rect 34471 4233 34483 4267
rect 34425 4227 34483 4233
rect 35342 4224 35348 4276
rect 35400 4264 35406 4276
rect 42150 4264 42156 4276
rect 35400 4236 42156 4264
rect 35400 4224 35406 4236
rect 42150 4224 42156 4236
rect 42208 4224 42214 4276
rect 43257 4267 43315 4273
rect 43257 4233 43269 4267
rect 43303 4264 43315 4267
rect 43990 4264 43996 4276
rect 43303 4236 43996 4264
rect 43303 4233 43315 4236
rect 43257 4227 43315 4233
rect 10686 4196 10692 4208
rect 9968 4168 10692 4196
rect 9122 4088 9128 4140
rect 9180 4128 9186 4140
rect 9585 4131 9643 4137
rect 9585 4128 9597 4131
rect 9180 4100 9597 4128
rect 9180 4088 9186 4100
rect 9585 4097 9597 4100
rect 9631 4097 9643 4131
rect 9858 4128 9864 4140
rect 9771 4100 9864 4128
rect 9585 4091 9643 4097
rect 9858 4088 9864 4100
rect 9916 4128 9922 4140
rect 9968 4128 9996 4168
rect 10686 4156 10692 4168
rect 10744 4156 10750 4208
rect 15470 4196 15476 4208
rect 14122 4168 15476 4196
rect 15470 4156 15476 4168
rect 15528 4156 15534 4208
rect 23017 4199 23075 4205
rect 23017 4165 23029 4199
rect 23063 4196 23075 4199
rect 24210 4196 24216 4208
rect 23063 4168 24216 4196
rect 23063 4165 23075 4168
rect 23017 4159 23075 4165
rect 24210 4156 24216 4168
rect 24268 4156 24274 4208
rect 25038 4156 25044 4208
rect 25096 4196 25102 4208
rect 25961 4199 26019 4205
rect 25961 4196 25973 4199
rect 25096 4168 25973 4196
rect 25096 4156 25102 4168
rect 25961 4165 25973 4168
rect 26007 4165 26019 4199
rect 25961 4159 26019 4165
rect 26142 4156 26148 4208
rect 26200 4196 26206 4208
rect 30006 4196 30012 4208
rect 26200 4168 30012 4196
rect 26200 4156 26206 4168
rect 30006 4156 30012 4168
rect 30064 4196 30070 4208
rect 32674 4196 32680 4208
rect 30064 4168 32680 4196
rect 30064 4156 30070 4168
rect 32674 4156 32680 4168
rect 32732 4156 32738 4208
rect 33410 4196 33416 4208
rect 33371 4168 33416 4196
rect 33410 4156 33416 4168
rect 33468 4156 33474 4208
rect 33594 4196 33600 4208
rect 33555 4168 33600 4196
rect 33594 4156 33600 4168
rect 33652 4156 33658 4208
rect 41230 4156 41236 4208
rect 41288 4196 41294 4208
rect 43272 4196 43300 4227
rect 43990 4224 43996 4236
rect 44048 4224 44054 4276
rect 51445 4267 51503 4273
rect 51445 4233 51457 4267
rect 51491 4264 51503 4267
rect 51534 4264 51540 4276
rect 51491 4236 51540 4264
rect 51491 4233 51503 4236
rect 51445 4227 51503 4233
rect 51534 4224 51540 4236
rect 51592 4224 51598 4276
rect 56597 4267 56655 4273
rect 56597 4233 56609 4267
rect 56643 4264 56655 4267
rect 57698 4264 57704 4276
rect 56643 4236 57704 4264
rect 56643 4233 56655 4236
rect 56597 4227 56655 4233
rect 57698 4224 57704 4236
rect 57756 4224 57762 4276
rect 59357 4267 59415 4273
rect 59357 4264 59369 4267
rect 57946 4236 59369 4264
rect 41288 4168 43300 4196
rect 50646 4168 51074 4196
rect 41288 4156 41294 4168
rect 10594 4128 10600 4140
rect 9916 4100 9996 4128
rect 10555 4100 10600 4128
rect 9916 4088 9922 4100
rect 10594 4088 10600 4100
rect 10652 4088 10658 4140
rect 14826 4088 14832 4140
rect 14884 4128 14890 4140
rect 25501 4131 25559 4137
rect 14884 4100 14929 4128
rect 14884 4088 14890 4100
rect 25501 4097 25513 4131
rect 25547 4128 25559 4131
rect 25682 4128 25688 4140
rect 25547 4100 25688 4128
rect 25547 4097 25559 4100
rect 25501 4091 25559 4097
rect 25682 4088 25688 4100
rect 25740 4088 25746 4140
rect 30834 4088 30840 4140
rect 30892 4128 30898 4140
rect 33229 4131 33287 4137
rect 33229 4128 33241 4131
rect 30892 4100 33241 4128
rect 30892 4088 30898 4100
rect 33229 4097 33241 4100
rect 33275 4097 33287 4131
rect 34606 4128 34612 4140
rect 34567 4100 34612 4128
rect 33229 4091 33287 4097
rect 34606 4088 34612 4100
rect 34664 4088 34670 4140
rect 38838 4088 38844 4140
rect 38896 4128 38902 4140
rect 39761 4131 39819 4137
rect 39761 4128 39773 4131
rect 38896 4100 39773 4128
rect 38896 4088 38902 4100
rect 39761 4097 39773 4100
rect 39807 4128 39819 4131
rect 39942 4128 39948 4140
rect 39807 4100 39948 4128
rect 39807 4097 39819 4100
rect 39761 4091 39819 4097
rect 39942 4088 39948 4100
rect 40000 4128 40006 4140
rect 40313 4131 40371 4137
rect 40313 4128 40325 4131
rect 40000 4100 40325 4128
rect 40000 4088 40006 4100
rect 40313 4097 40325 4100
rect 40359 4128 40371 4131
rect 41417 4131 41475 4137
rect 41417 4128 41429 4131
rect 40359 4100 41429 4128
rect 40359 4097 40371 4100
rect 40313 4091 40371 4097
rect 41417 4097 41429 4100
rect 41463 4128 41475 4131
rect 41782 4128 41788 4140
rect 41463 4100 41788 4128
rect 41463 4097 41475 4100
rect 41417 4091 41475 4097
rect 41782 4088 41788 4100
rect 41840 4088 41846 4140
rect 43806 4128 43812 4140
rect 43767 4100 43812 4128
rect 43806 4088 43812 4100
rect 43864 4088 43870 4140
rect 50430 4088 50436 4140
rect 50488 4088 50494 4140
rect 51046 4128 51074 4168
rect 52178 4156 52184 4208
rect 52236 4196 52242 4208
rect 53745 4199 53803 4205
rect 53745 4196 53757 4199
rect 52236 4168 53757 4196
rect 52236 4156 52242 4168
rect 53745 4165 53757 4168
rect 53791 4165 53803 4199
rect 55490 4196 55496 4208
rect 55451 4168 55496 4196
rect 53745 4159 53803 4165
rect 55490 4156 55496 4168
rect 55548 4156 55554 4208
rect 56410 4156 56416 4208
rect 56468 4196 56474 4208
rect 57946 4196 57974 4236
rect 59357 4233 59369 4236
rect 59403 4233 59415 4267
rect 59357 4227 59415 4233
rect 59446 4224 59452 4276
rect 59504 4264 59510 4276
rect 62206 4264 62212 4276
rect 59504 4236 62212 4264
rect 59504 4224 59510 4236
rect 62206 4224 62212 4236
rect 62264 4224 62270 4276
rect 63494 4224 63500 4276
rect 63552 4264 63558 4276
rect 64325 4267 64383 4273
rect 64325 4264 64337 4267
rect 63552 4236 64337 4264
rect 63552 4224 63558 4236
rect 64325 4233 64337 4236
rect 64371 4233 64383 4267
rect 64325 4227 64383 4233
rect 62298 4196 62304 4208
rect 56468 4168 57974 4196
rect 60398 4168 62304 4196
rect 56468 4156 56474 4168
rect 62298 4156 62304 4168
rect 62356 4156 62362 4208
rect 51258 4128 51264 4140
rect 51046 4100 51264 4128
rect 51258 4088 51264 4100
rect 51316 4088 51322 4140
rect 52270 4128 52276 4140
rect 52231 4100 52276 4128
rect 52270 4088 52276 4100
rect 52328 4088 52334 4140
rect 53190 4128 53196 4140
rect 53151 4100 53196 4128
rect 53190 4088 53196 4100
rect 53248 4128 53254 4140
rect 54662 4128 54668 4140
rect 53248 4100 54668 4128
rect 53248 4088 53254 4100
rect 54662 4088 54668 4100
rect 54720 4088 54726 4140
rect 57882 4128 57888 4140
rect 56060 4100 57888 4128
rect 13078 4060 13084 4072
rect 13039 4032 13084 4060
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 14550 4060 14556 4072
rect 14511 4032 14556 4060
rect 14550 4020 14556 4032
rect 14608 4020 14614 4072
rect 25406 4020 25412 4072
rect 25464 4060 25470 4072
rect 26329 4063 26387 4069
rect 26329 4060 26341 4063
rect 25464 4032 26341 4060
rect 25464 4020 25470 4032
rect 26329 4029 26341 4032
rect 26375 4029 26387 4063
rect 37458 4060 37464 4072
rect 37419 4032 37464 4060
rect 26329 4023 26387 4029
rect 37458 4020 37464 4032
rect 37516 4020 37522 4072
rect 37734 4060 37740 4072
rect 37695 4032 37740 4060
rect 37734 4020 37740 4032
rect 37792 4020 37798 4072
rect 38470 4020 38476 4072
rect 38528 4060 38534 4072
rect 38856 4060 38884 4088
rect 38528 4032 38884 4060
rect 39209 4063 39267 4069
rect 38528 4020 38534 4032
rect 39209 4029 39221 4063
rect 39255 4060 39267 4063
rect 40678 4060 40684 4072
rect 39255 4032 40684 4060
rect 39255 4029 39267 4032
rect 39209 4023 39267 4029
rect 40678 4020 40684 4032
rect 40736 4020 40742 4072
rect 40770 4020 40776 4072
rect 40828 4060 40834 4072
rect 40828 4032 40873 4060
rect 40828 4020 40834 4032
rect 48314 4020 48320 4072
rect 48372 4060 48378 4072
rect 49142 4060 49148 4072
rect 48372 4032 49148 4060
rect 48372 4020 48378 4032
rect 49142 4020 49148 4032
rect 49200 4020 49206 4072
rect 49421 4063 49479 4069
rect 49421 4060 49433 4063
rect 49252 4032 49433 4060
rect 10318 3952 10324 4004
rect 10376 3992 10382 4004
rect 10781 3995 10839 4001
rect 10781 3992 10793 3995
rect 10376 3964 10793 3992
rect 10376 3952 10382 3964
rect 10781 3961 10793 3964
rect 10827 3992 10839 3995
rect 13538 3992 13544 4004
rect 10827 3964 13544 3992
rect 10827 3961 10839 3964
rect 10781 3955 10839 3961
rect 13538 3952 13544 3964
rect 13596 3952 13602 4004
rect 47394 3952 47400 4004
rect 47452 3992 47458 4004
rect 49252 3992 49280 4032
rect 49421 4029 49433 4032
rect 49467 4029 49479 4063
rect 50448 4060 50476 4088
rect 50893 4063 50951 4069
rect 50893 4060 50905 4063
rect 50448 4032 50905 4060
rect 49421 4023 49479 4029
rect 50893 4029 50905 4032
rect 50939 4029 50951 4063
rect 55122 4060 55128 4072
rect 55083 4032 55128 4060
rect 50893 4023 50951 4029
rect 55122 4020 55128 4032
rect 55180 4020 55186 4072
rect 55585 4063 55643 4069
rect 55585 4029 55597 4063
rect 55631 4060 55643 4063
rect 56060 4060 56088 4100
rect 57882 4088 57888 4100
rect 57940 4088 57946 4140
rect 58066 4088 58072 4140
rect 58124 4128 58130 4140
rect 58621 4131 58679 4137
rect 58621 4128 58633 4131
rect 58124 4100 58633 4128
rect 58124 4088 58130 4100
rect 58621 4097 58633 4100
rect 58667 4097 58679 4131
rect 62022 4128 62028 4140
rect 61983 4100 62028 4128
rect 58621 4091 58679 4097
rect 62022 4088 62028 4100
rect 62080 4088 62086 4140
rect 62574 4128 62580 4140
rect 62535 4100 62580 4128
rect 62574 4088 62580 4100
rect 62632 4088 62638 4140
rect 62942 4088 62948 4140
rect 63000 4128 63006 4140
rect 63773 4131 63831 4137
rect 63773 4128 63785 4131
rect 63000 4100 63785 4128
rect 63000 4088 63006 4100
rect 63773 4097 63785 4100
rect 63819 4097 63831 4131
rect 64340 4128 64368 4227
rect 71866 4224 71872 4276
rect 71924 4224 71930 4276
rect 73982 4224 73988 4276
rect 74040 4264 74046 4276
rect 74040 4236 75868 4264
rect 74040 4224 74046 4236
rect 71501 4199 71559 4205
rect 71501 4165 71513 4199
rect 71547 4196 71559 4199
rect 71590 4196 71596 4208
rect 71547 4168 71596 4196
rect 71547 4165 71559 4168
rect 71501 4159 71559 4165
rect 71590 4156 71596 4168
rect 71648 4156 71654 4208
rect 71884 4196 71912 4224
rect 71884 4168 71990 4196
rect 73430 4156 73436 4208
rect 73488 4196 73494 4208
rect 73525 4199 73583 4205
rect 73525 4196 73537 4199
rect 73488 4168 73537 4196
rect 73488 4156 73494 4168
rect 73525 4165 73537 4168
rect 73571 4196 73583 4199
rect 74166 4196 74172 4208
rect 73571 4168 74172 4196
rect 73571 4165 73583 4168
rect 73525 4159 73583 4165
rect 74166 4156 74172 4168
rect 74224 4156 74230 4208
rect 75840 4196 75868 4236
rect 75914 4224 75920 4276
rect 75972 4264 75978 4276
rect 77294 4264 77300 4276
rect 75972 4236 76017 4264
rect 76852 4236 77300 4264
rect 75972 4224 75978 4236
rect 76852 4196 76880 4236
rect 77294 4224 77300 4236
rect 77352 4224 77358 4276
rect 77478 4264 77484 4276
rect 77439 4236 77484 4264
rect 77478 4224 77484 4236
rect 77536 4224 77542 4276
rect 79962 4264 79968 4276
rect 77588 4236 79968 4264
rect 75840 4168 76880 4196
rect 76926 4156 76932 4208
rect 76984 4196 76990 4208
rect 77588 4196 77616 4236
rect 79962 4224 79968 4236
rect 80020 4224 80026 4276
rect 80238 4224 80244 4276
rect 80296 4264 80302 4276
rect 83734 4264 83740 4276
rect 80296 4236 83740 4264
rect 80296 4224 80302 4236
rect 83734 4224 83740 4236
rect 83792 4224 83798 4276
rect 84010 4264 84016 4276
rect 83971 4236 84016 4264
rect 84010 4224 84016 4236
rect 84068 4224 84074 4276
rect 84197 4267 84255 4273
rect 84197 4233 84209 4267
rect 84243 4264 84255 4267
rect 84654 4264 84660 4276
rect 84243 4236 84660 4264
rect 84243 4233 84255 4236
rect 84197 4227 84255 4233
rect 84654 4224 84660 4236
rect 84712 4224 84718 4276
rect 85114 4224 85120 4276
rect 85172 4264 85178 4276
rect 86773 4267 86831 4273
rect 86773 4264 86785 4267
rect 85172 4236 86785 4264
rect 85172 4224 85178 4236
rect 86773 4233 86785 4236
rect 86819 4264 86831 4267
rect 87138 4264 87144 4276
rect 86819 4236 87144 4264
rect 86819 4233 86831 4236
rect 86773 4227 86831 4233
rect 87138 4224 87144 4236
rect 87196 4224 87202 4276
rect 90266 4264 90272 4276
rect 90227 4236 90272 4264
rect 90266 4224 90272 4236
rect 90324 4224 90330 4276
rect 91741 4267 91799 4273
rect 91741 4233 91753 4267
rect 91787 4264 91799 4267
rect 91922 4264 91928 4276
rect 91787 4236 91928 4264
rect 91787 4233 91799 4236
rect 91741 4227 91799 4233
rect 91922 4224 91928 4236
rect 91980 4224 91986 4276
rect 76984 4168 77616 4196
rect 76984 4156 76990 4168
rect 78398 4156 78404 4208
rect 78456 4196 78462 4208
rect 78953 4199 79011 4205
rect 78953 4196 78965 4199
rect 78456 4168 78965 4196
rect 78456 4156 78462 4168
rect 78953 4165 78965 4168
rect 78999 4165 79011 4199
rect 80606 4196 80612 4208
rect 80178 4168 80612 4196
rect 78953 4159 79011 4165
rect 80606 4156 80612 4168
rect 80664 4156 80670 4208
rect 84105 4199 84163 4205
rect 84105 4165 84117 4199
rect 84151 4196 84163 4199
rect 84562 4196 84568 4208
rect 84151 4168 84568 4196
rect 84151 4165 84163 4168
rect 84105 4159 84163 4165
rect 84562 4156 84568 4168
rect 84620 4196 84626 4208
rect 88610 4196 88616 4208
rect 84620 4168 88616 4196
rect 84620 4156 84626 4168
rect 88610 4156 88616 4168
rect 88668 4196 88674 4208
rect 88668 4168 89714 4196
rect 88668 4156 88674 4168
rect 65429 4131 65487 4137
rect 65429 4128 65441 4131
rect 64340 4100 65441 4128
rect 63773 4091 63831 4097
rect 65429 4097 65441 4100
rect 65475 4097 65487 4131
rect 71222 4128 71228 4140
rect 71183 4100 71228 4128
rect 65429 4091 65487 4097
rect 71222 4088 71228 4100
rect 71280 4088 71286 4140
rect 73706 4088 73712 4140
rect 73764 4128 73770 4140
rect 73801 4131 73859 4137
rect 73801 4128 73813 4131
rect 73764 4100 73813 4128
rect 73764 4088 73770 4100
rect 73801 4097 73813 4100
rect 73847 4128 73859 4131
rect 77389 4131 77447 4137
rect 77389 4128 77401 4131
rect 73847 4100 77401 4128
rect 73847 4097 73859 4100
rect 73801 4091 73859 4097
rect 77389 4097 77401 4100
rect 77435 4128 77447 4131
rect 77435 4100 78168 4128
rect 77435 4097 77447 4100
rect 77389 4091 77447 4097
rect 55631 4032 56088 4060
rect 56137 4063 56195 4069
rect 55631 4029 55643 4032
rect 55585 4023 55643 4029
rect 56137 4029 56149 4063
rect 56183 4060 56195 4063
rect 57054 4060 57060 4072
rect 56183 4032 56548 4060
rect 57015 4032 57060 4060
rect 56183 4029 56195 4032
rect 56137 4023 56195 4029
rect 47452 3964 49280 3992
rect 47452 3952 47458 3964
rect 55950 3952 55956 4004
rect 56008 3992 56014 4004
rect 56152 3992 56180 4023
rect 56008 3964 56180 3992
rect 56413 3995 56471 4001
rect 56008 3952 56014 3964
rect 56413 3961 56425 3995
rect 56459 3961 56471 3995
rect 56520 3992 56548 4032
rect 57054 4020 57060 4032
rect 57112 4020 57118 4072
rect 57517 4063 57575 4069
rect 57517 4029 57529 4063
rect 57563 4060 57575 4063
rect 58710 4060 58716 4072
rect 57563 4032 58716 4060
rect 57563 4029 57575 4032
rect 57517 4023 57575 4029
rect 58710 4020 58716 4032
rect 58768 4020 58774 4072
rect 60829 4063 60887 4069
rect 60829 4060 60841 4063
rect 58820 4032 60841 4060
rect 57333 3995 57391 4001
rect 57333 3992 57345 3995
rect 56520 3964 57345 3992
rect 56413 3955 56471 3961
rect 57333 3961 57345 3964
rect 57379 3961 57391 3995
rect 57333 3955 57391 3961
rect 10686 3884 10692 3936
rect 10744 3924 10750 3936
rect 11793 3927 11851 3933
rect 11793 3924 11805 3927
rect 10744 3896 11805 3924
rect 10744 3884 10750 3896
rect 11793 3893 11805 3896
rect 11839 3924 11851 3927
rect 15194 3924 15200 3936
rect 11839 3896 15200 3924
rect 11839 3893 11851 3896
rect 11793 3887 11851 3893
rect 15194 3884 15200 3896
rect 15252 3884 15258 3936
rect 36909 3927 36967 3933
rect 36909 3893 36921 3927
rect 36955 3924 36967 3927
rect 37918 3924 37924 3936
rect 36955 3896 37924 3924
rect 36955 3893 36967 3896
rect 36909 3887 36967 3893
rect 37918 3884 37924 3896
rect 37976 3884 37982 3936
rect 38102 3884 38108 3936
rect 38160 3924 38166 3936
rect 40586 3924 40592 3936
rect 38160 3896 40592 3924
rect 38160 3884 38166 3896
rect 40586 3884 40592 3896
rect 40644 3884 40650 3936
rect 49142 3884 49148 3936
rect 49200 3924 49206 3936
rect 51074 3924 51080 3936
rect 49200 3896 51080 3924
rect 49200 3884 49206 3896
rect 51074 3884 51080 3896
rect 51132 3924 51138 3936
rect 56226 3924 56232 3936
rect 51132 3896 56232 3924
rect 51132 3884 51138 3896
rect 56226 3884 56232 3896
rect 56284 3884 56290 3936
rect 56428 3924 56456 3955
rect 57790 3952 57796 4004
rect 57848 3992 57854 4004
rect 58820 3992 58848 4032
rect 60829 4029 60841 4032
rect 60875 4029 60887 4063
rect 60829 4023 60887 4029
rect 61105 4063 61163 4069
rect 61105 4029 61117 4063
rect 61151 4060 61163 4063
rect 61286 4060 61292 4072
rect 61151 4032 61292 4060
rect 61151 4029 61163 4032
rect 61105 4023 61163 4029
rect 61286 4020 61292 4032
rect 61344 4060 61350 4072
rect 61344 4032 63816 4060
rect 61344 4020 61350 4032
rect 63788 4004 63816 4032
rect 64782 4020 64788 4072
rect 64840 4060 64846 4072
rect 68646 4060 68652 4072
rect 64840 4032 68652 4060
rect 64840 4020 64846 4032
rect 68646 4020 68652 4032
rect 68704 4020 68710 4072
rect 72973 4063 73031 4069
rect 72973 4029 72985 4063
rect 73019 4060 73031 4063
rect 73522 4060 73528 4072
rect 73019 4032 73528 4060
rect 73019 4029 73031 4032
rect 72973 4023 73031 4029
rect 73522 4020 73528 4032
rect 73580 4020 73586 4072
rect 74350 4060 74356 4072
rect 74311 4032 74356 4060
rect 74350 4020 74356 4032
rect 74408 4020 74414 4072
rect 74442 4020 74448 4072
rect 74500 4060 74506 4072
rect 75178 4060 75184 4072
rect 74500 4032 75184 4060
rect 74500 4020 74506 4032
rect 75178 4020 75184 4032
rect 75236 4060 75242 4072
rect 78030 4060 78036 4072
rect 75236 4032 78036 4060
rect 75236 4020 75242 4032
rect 78030 4020 78036 4032
rect 78088 4020 78094 4072
rect 57848 3964 58848 3992
rect 57848 3952 57854 3964
rect 62022 3952 62028 4004
rect 62080 3992 62086 4004
rect 62080 3964 63724 3992
rect 62080 3952 62086 3964
rect 57054 3924 57060 3936
rect 56428 3896 57060 3924
rect 57054 3884 57060 3896
rect 57112 3884 57118 3936
rect 58161 3927 58219 3933
rect 58161 3893 58173 3927
rect 58207 3924 58219 3927
rect 59354 3924 59360 3936
rect 58207 3896 59360 3924
rect 58207 3893 58219 3896
rect 58161 3887 58219 3893
rect 59354 3884 59360 3896
rect 59412 3884 59418 3936
rect 62666 3884 62672 3936
rect 62724 3924 62730 3936
rect 63221 3927 63279 3933
rect 63221 3924 63233 3927
rect 62724 3896 63233 3924
rect 62724 3884 62730 3896
rect 63221 3893 63233 3896
rect 63267 3893 63279 3927
rect 63696 3924 63724 3964
rect 63770 3952 63776 4004
rect 63828 3992 63834 4004
rect 64874 3992 64880 4004
rect 63828 3964 64880 3992
rect 63828 3952 63834 3964
rect 64874 3952 64880 3964
rect 64932 3992 64938 4004
rect 64969 3995 65027 4001
rect 64969 3992 64981 3995
rect 64932 3964 64981 3992
rect 64932 3952 64938 3964
rect 64969 3961 64981 3964
rect 65015 3961 65027 3995
rect 73706 3992 73712 4004
rect 73667 3964 73712 3992
rect 64969 3955 65027 3961
rect 73706 3952 73712 3964
rect 73764 3952 73770 4004
rect 76190 3952 76196 4004
rect 76248 3992 76254 4004
rect 76248 3964 78076 3992
rect 76248 3952 76254 3964
rect 65981 3927 66039 3933
rect 65981 3924 65993 3927
rect 63696 3896 65993 3924
rect 63221 3887 63279 3893
rect 65981 3893 65993 3896
rect 66027 3924 66039 3927
rect 67726 3924 67732 3936
rect 66027 3896 67732 3924
rect 66027 3893 66039 3896
rect 65981 3887 66039 3893
rect 67726 3884 67732 3896
rect 67784 3924 67790 3936
rect 68373 3927 68431 3933
rect 68373 3924 68385 3927
rect 67784 3896 68385 3924
rect 67784 3884 67790 3896
rect 68373 3893 68385 3896
rect 68419 3893 68431 3927
rect 73614 3924 73620 3936
rect 73575 3896 73620 3924
rect 68373 3887 68431 3893
rect 73614 3884 73620 3896
rect 73672 3884 73678 3936
rect 76374 3884 76380 3936
rect 76432 3924 76438 3936
rect 78048 3933 78076 3964
rect 76469 3927 76527 3933
rect 76469 3924 76481 3927
rect 76432 3896 76481 3924
rect 76432 3884 76438 3896
rect 76469 3893 76481 3896
rect 76515 3893 76527 3927
rect 76469 3887 76527 3893
rect 78033 3927 78091 3933
rect 78033 3893 78045 3927
rect 78079 3893 78091 3927
rect 78140 3924 78168 4100
rect 80514 4088 80520 4140
rect 80572 4128 80578 4140
rect 80885 4131 80943 4137
rect 80885 4128 80897 4131
rect 80572 4100 80897 4128
rect 80572 4088 80578 4100
rect 80885 4097 80897 4100
rect 80931 4097 80943 4131
rect 80885 4091 80943 4097
rect 81529 4131 81587 4137
rect 81529 4097 81541 4131
rect 81575 4128 81587 4131
rect 81986 4128 81992 4140
rect 81575 4100 81992 4128
rect 81575 4097 81587 4100
rect 81529 4091 81587 4097
rect 81986 4088 81992 4100
rect 82044 4088 82050 4140
rect 83277 4131 83335 4137
rect 83277 4097 83289 4131
rect 83323 4128 83335 4131
rect 83550 4128 83556 4140
rect 83323 4100 83556 4128
rect 83323 4097 83335 4100
rect 83277 4091 83335 4097
rect 83550 4088 83556 4100
rect 83608 4088 83614 4140
rect 83826 4128 83832 4140
rect 83787 4100 83832 4128
rect 83826 4088 83832 4100
rect 83884 4088 83890 4140
rect 84838 4128 84844 4140
rect 84799 4100 84844 4128
rect 84838 4088 84844 4100
rect 84896 4088 84902 4140
rect 85482 4128 85488 4140
rect 85443 4100 85488 4128
rect 85482 4088 85488 4100
rect 85540 4088 85546 4140
rect 86126 4088 86132 4140
rect 86184 4128 86190 4140
rect 86221 4131 86279 4137
rect 86221 4128 86233 4131
rect 86184 4100 86233 4128
rect 86184 4088 86190 4100
rect 86221 4097 86233 4100
rect 86267 4097 86279 4131
rect 86954 4128 86960 4140
rect 86915 4100 86960 4128
rect 86221 4091 86279 4097
rect 86954 4088 86960 4100
rect 87012 4088 87018 4140
rect 87230 4088 87236 4140
rect 87288 4128 87294 4140
rect 87693 4131 87751 4137
rect 87693 4128 87705 4131
rect 87288 4100 87705 4128
rect 87288 4088 87294 4100
rect 87693 4097 87705 4100
rect 87739 4097 87751 4131
rect 87966 4128 87972 4140
rect 87927 4100 87972 4128
rect 87693 4091 87751 4097
rect 87966 4088 87972 4100
rect 88024 4088 88030 4140
rect 89686 4128 89714 4168
rect 89806 4156 89812 4208
rect 89864 4196 89870 4208
rect 90177 4199 90235 4205
rect 90177 4196 90189 4199
rect 89864 4168 90189 4196
rect 89864 4156 89870 4168
rect 90177 4165 90189 4168
rect 90223 4165 90235 4199
rect 90177 4159 90235 4165
rect 91020 4168 92046 4196
rect 89990 4128 89996 4140
rect 89686 4100 89996 4128
rect 89990 4088 89996 4100
rect 90048 4088 90054 4140
rect 90269 4131 90327 4137
rect 90269 4097 90281 4131
rect 90315 4128 90327 4131
rect 90729 4131 90787 4137
rect 90729 4128 90741 4131
rect 90315 4100 90741 4128
rect 90315 4097 90327 4100
rect 90269 4091 90327 4097
rect 90729 4097 90741 4100
rect 90775 4097 90787 4131
rect 90729 4091 90787 4097
rect 78582 4020 78588 4072
rect 78640 4060 78646 4072
rect 78677 4063 78735 4069
rect 78677 4060 78689 4063
rect 78640 4032 78689 4060
rect 78640 4020 78646 4032
rect 78677 4029 78689 4032
rect 78723 4029 78735 4063
rect 78677 4023 78735 4029
rect 79962 4020 79968 4072
rect 80020 4060 80026 4072
rect 80425 4063 80483 4069
rect 80425 4060 80437 4063
rect 80020 4032 80437 4060
rect 80020 4020 80026 4032
rect 80425 4029 80437 4032
rect 80471 4029 80483 4063
rect 80425 4023 80483 4029
rect 80698 4020 80704 4072
rect 80756 4060 80762 4072
rect 82173 4063 82231 4069
rect 82173 4060 82185 4063
rect 80756 4032 82185 4060
rect 80756 4020 80762 4032
rect 82173 4029 82185 4032
rect 82219 4060 82231 4063
rect 82219 4032 86908 4060
rect 82219 4029 82231 4032
rect 82173 4023 82231 4029
rect 84194 3992 84200 4004
rect 80026 3964 84200 3992
rect 80026 3924 80054 3964
rect 84194 3952 84200 3964
rect 84252 3952 84258 4004
rect 84381 3995 84439 4001
rect 84381 3961 84393 3995
rect 84427 3992 84439 3995
rect 84930 3992 84936 4004
rect 84427 3964 84936 3992
rect 84427 3961 84439 3964
rect 84381 3955 84439 3961
rect 84930 3952 84936 3964
rect 84988 3952 84994 4004
rect 78140 3896 80054 3924
rect 78033 3887 78091 3893
rect 81986 3884 81992 3936
rect 82044 3924 82050 3936
rect 82633 3927 82691 3933
rect 82633 3924 82645 3927
rect 82044 3896 82645 3924
rect 82044 3884 82050 3896
rect 82633 3893 82645 3896
rect 82679 3893 82691 3927
rect 86880 3924 86908 4032
rect 89622 4020 89628 4072
rect 89680 4060 89686 4072
rect 90284 4060 90312 4091
rect 89680 4032 90312 4060
rect 89680 4020 89686 4032
rect 89070 3992 89076 4004
rect 87892 3964 89076 3992
rect 87892 3924 87920 3964
rect 89070 3952 89076 3964
rect 89128 3952 89134 4004
rect 89898 3952 89904 4004
rect 89956 3992 89962 4004
rect 91020 3992 91048 4168
rect 93118 4020 93124 4072
rect 93176 4060 93182 4072
rect 93213 4063 93271 4069
rect 93213 4060 93225 4063
rect 93176 4032 93225 4060
rect 93176 4020 93182 4032
rect 93213 4029 93225 4032
rect 93259 4029 93271 4063
rect 93489 4063 93547 4069
rect 93489 4060 93501 4063
rect 93213 4023 93271 4029
rect 93412 4032 93501 4060
rect 89956 3964 91048 3992
rect 89956 3952 89962 3964
rect 88978 3924 88984 3936
rect 86880 3896 87920 3924
rect 88939 3896 88984 3924
rect 82633 3887 82691 3893
rect 88978 3884 88984 3896
rect 89036 3884 89042 3936
rect 91002 3884 91008 3936
rect 91060 3924 91066 3936
rect 93412 3924 93440 4032
rect 93489 4029 93501 4032
rect 93535 4060 93547 4063
rect 94133 4063 94191 4069
rect 94133 4060 94145 4063
rect 93535 4032 94145 4060
rect 93535 4029 93547 4032
rect 93489 4023 93547 4029
rect 94133 4029 94145 4032
rect 94179 4060 94191 4063
rect 94222 4060 94228 4072
rect 94179 4032 94228 4060
rect 94179 4029 94191 4032
rect 94133 4023 94191 4029
rect 94222 4020 94228 4032
rect 94280 4020 94286 4072
rect 91060 3896 93440 3924
rect 91060 3884 91066 3896
rect 1104 3834 94852 3856
rect 1104 3782 12668 3834
rect 12720 3782 12732 3834
rect 12784 3782 12796 3834
rect 12848 3782 12860 3834
rect 12912 3782 12924 3834
rect 12976 3782 36105 3834
rect 36157 3782 36169 3834
rect 36221 3782 36233 3834
rect 36285 3782 36297 3834
rect 36349 3782 36361 3834
rect 36413 3782 59542 3834
rect 59594 3782 59606 3834
rect 59658 3782 59670 3834
rect 59722 3782 59734 3834
rect 59786 3782 59798 3834
rect 59850 3782 82979 3834
rect 83031 3782 83043 3834
rect 83095 3782 83107 3834
rect 83159 3782 83171 3834
rect 83223 3782 83235 3834
rect 83287 3782 94852 3834
rect 1104 3760 94852 3782
rect 4062 3680 4068 3732
rect 4120 3720 4126 3732
rect 10962 3720 10968 3732
rect 4120 3692 10968 3720
rect 4120 3680 4126 3692
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 13538 3680 13544 3732
rect 13596 3720 13602 3732
rect 14277 3723 14335 3729
rect 14277 3720 14289 3723
rect 13596 3692 14289 3720
rect 13596 3680 13602 3692
rect 14277 3689 14289 3692
rect 14323 3689 14335 3723
rect 14277 3683 14335 3689
rect 32306 3680 32312 3732
rect 32364 3720 32370 3732
rect 32364 3692 40540 3720
rect 32364 3680 32370 3692
rect 32950 3612 32956 3664
rect 33008 3652 33014 3664
rect 38102 3652 38108 3664
rect 33008 3624 38108 3652
rect 33008 3612 33014 3624
rect 38102 3612 38108 3624
rect 38160 3612 38166 3664
rect 39942 3612 39948 3664
rect 40000 3652 40006 3664
rect 40037 3655 40095 3661
rect 40037 3652 40049 3655
rect 40000 3624 40049 3652
rect 40000 3612 40006 3624
rect 40037 3621 40049 3624
rect 40083 3621 40095 3655
rect 40037 3615 40095 3621
rect 37458 3544 37464 3596
rect 37516 3584 37522 3596
rect 39393 3587 39451 3593
rect 39393 3584 39405 3587
rect 37516 3556 39405 3584
rect 37516 3544 37522 3556
rect 39393 3553 39405 3556
rect 39439 3584 39451 3587
rect 40402 3584 40408 3596
rect 39439 3556 40408 3584
rect 39439 3553 39451 3556
rect 39393 3547 39451 3553
rect 40402 3544 40408 3556
rect 40460 3544 40466 3596
rect 40512 3584 40540 3692
rect 40586 3680 40592 3732
rect 40644 3720 40650 3732
rect 55490 3720 55496 3732
rect 40644 3692 55496 3720
rect 40644 3680 40650 3692
rect 55490 3680 55496 3692
rect 55548 3680 55554 3732
rect 58526 3720 58532 3732
rect 57900 3692 58532 3720
rect 40770 3612 40776 3664
rect 40828 3652 40834 3664
rect 49786 3652 49792 3664
rect 40828 3624 49792 3652
rect 40828 3612 40834 3624
rect 49786 3612 49792 3624
rect 49844 3612 49850 3664
rect 51074 3612 51080 3664
rect 51132 3652 51138 3664
rect 54202 3652 54208 3664
rect 51132 3624 51177 3652
rect 54163 3624 54208 3652
rect 51132 3612 51138 3624
rect 54202 3612 54208 3624
rect 54260 3612 54266 3664
rect 54662 3652 54668 3664
rect 54623 3624 54668 3652
rect 54662 3612 54668 3624
rect 54720 3612 54726 3664
rect 51905 3587 51963 3593
rect 40512 3556 51856 3584
rect 10594 3476 10600 3528
rect 10652 3516 10658 3528
rect 14461 3519 14519 3525
rect 14461 3516 14473 3519
rect 10652 3488 14473 3516
rect 10652 3476 10658 3488
rect 14461 3485 14473 3488
rect 14507 3485 14519 3519
rect 15194 3516 15200 3528
rect 15155 3488 15200 3516
rect 14461 3479 14519 3485
rect 15194 3476 15200 3488
rect 15252 3476 15258 3528
rect 15470 3516 15476 3528
rect 15431 3488 15476 3516
rect 15470 3476 15476 3488
rect 15528 3476 15534 3528
rect 15212 3448 15240 3476
rect 15933 3451 15991 3457
rect 15933 3448 15945 3451
rect 15212 3420 15945 3448
rect 15933 3417 15945 3420
rect 15979 3417 15991 3451
rect 38838 3448 38844 3460
rect 38686 3420 38844 3448
rect 15933 3411 15991 3417
rect 38838 3408 38844 3420
rect 38896 3408 38902 3460
rect 39117 3451 39175 3457
rect 39117 3417 39129 3451
rect 39163 3448 39175 3451
rect 41322 3448 41328 3460
rect 39163 3420 41328 3448
rect 39163 3417 39175 3420
rect 39117 3411 39175 3417
rect 41322 3408 41328 3420
rect 41380 3408 41386 3460
rect 24210 3340 24216 3392
rect 24268 3380 24274 3392
rect 37645 3383 37703 3389
rect 37645 3380 37657 3383
rect 24268 3352 37657 3380
rect 24268 3340 24274 3352
rect 37645 3349 37657 3352
rect 37691 3380 37703 3383
rect 39022 3380 39028 3392
rect 37691 3352 39028 3380
rect 37691 3349 37703 3352
rect 37645 3343 37703 3349
rect 39022 3340 39028 3352
rect 39080 3340 39086 3392
rect 51828 3380 51856 3556
rect 51905 3553 51917 3587
rect 51951 3584 51963 3587
rect 55950 3584 55956 3596
rect 51951 3556 55956 3584
rect 51951 3553 51963 3556
rect 51905 3547 51963 3553
rect 55950 3544 55956 3556
rect 56008 3544 56014 3596
rect 53653 3519 53711 3525
rect 53653 3485 53665 3519
rect 53699 3516 53711 3519
rect 53834 3516 53840 3528
rect 53699 3488 53840 3516
rect 53699 3485 53711 3488
rect 53653 3479 53711 3485
rect 53834 3476 53840 3488
rect 53892 3516 53898 3528
rect 55677 3519 55735 3525
rect 55677 3516 55689 3519
rect 53892 3488 55689 3516
rect 53892 3476 53898 3488
rect 55677 3485 55689 3488
rect 55723 3485 55735 3519
rect 55677 3479 55735 3485
rect 52362 3408 52368 3460
rect 52420 3408 52426 3460
rect 53374 3448 53380 3460
rect 53335 3420 53380 3448
rect 53374 3408 53380 3420
rect 53432 3408 53438 3460
rect 55122 3448 55128 3460
rect 53484 3420 55128 3448
rect 53484 3380 53512 3420
rect 55122 3408 55128 3420
rect 55180 3408 55186 3460
rect 51828 3352 53512 3380
rect 55692 3380 55720 3479
rect 57330 3476 57336 3528
rect 57388 3516 57394 3528
rect 57900 3525 57928 3692
rect 58526 3680 58532 3692
rect 58584 3680 58590 3732
rect 59262 3720 59268 3732
rect 59175 3692 59268 3720
rect 59262 3680 59268 3692
rect 59320 3720 59326 3732
rect 61194 3720 61200 3732
rect 59320 3692 61200 3720
rect 59320 3680 59326 3692
rect 61194 3680 61200 3692
rect 61252 3720 61258 3732
rect 61473 3723 61531 3729
rect 61473 3720 61485 3723
rect 61252 3692 61485 3720
rect 61252 3680 61258 3692
rect 61473 3689 61485 3692
rect 61519 3689 61531 3723
rect 64598 3720 64604 3732
rect 61473 3683 61531 3689
rect 62776 3692 64604 3720
rect 60737 3655 60795 3661
rect 60737 3621 60749 3655
rect 60783 3652 60795 3655
rect 62776 3652 62804 3692
rect 64598 3680 64604 3692
rect 64656 3680 64662 3732
rect 67174 3680 67180 3732
rect 67232 3720 67238 3732
rect 68557 3723 68615 3729
rect 68557 3720 68569 3723
rect 67232 3692 68569 3720
rect 67232 3680 67238 3692
rect 60783 3624 62804 3652
rect 64509 3655 64567 3661
rect 60783 3621 60795 3624
rect 60737 3615 60795 3621
rect 64509 3621 64521 3655
rect 64555 3652 64567 3655
rect 64690 3652 64696 3664
rect 64555 3624 64696 3652
rect 64555 3621 64567 3624
rect 64509 3615 64567 3621
rect 64690 3612 64696 3624
rect 64748 3612 64754 3664
rect 64049 3587 64107 3593
rect 64049 3584 64061 3587
rect 58452 3556 64061 3584
rect 57885 3519 57943 3525
rect 57885 3516 57897 3519
rect 57388 3488 57897 3516
rect 57388 3476 57394 3488
rect 57885 3485 57897 3488
rect 57931 3485 57943 3519
rect 57885 3479 57943 3485
rect 55858 3408 55864 3460
rect 55916 3448 55922 3460
rect 58452 3457 58480 3556
rect 64049 3553 64061 3556
rect 64095 3584 64107 3587
rect 64322 3584 64328 3596
rect 64095 3556 64328 3584
rect 64095 3553 64107 3556
rect 64049 3547 64107 3553
rect 64322 3544 64328 3556
rect 64380 3544 64386 3596
rect 62025 3519 62083 3525
rect 62025 3485 62037 3519
rect 62071 3516 62083 3519
rect 62206 3516 62212 3528
rect 62071 3488 62212 3516
rect 62071 3485 62083 3488
rect 62025 3479 62083 3485
rect 62206 3476 62212 3488
rect 62264 3476 62270 3528
rect 64598 3476 64604 3528
rect 64656 3516 64662 3528
rect 67928 3525 67956 3692
rect 68557 3689 68569 3692
rect 68603 3689 68615 3723
rect 68557 3683 68615 3689
rect 68646 3680 68652 3732
rect 68704 3720 68710 3732
rect 68704 3692 85988 3720
rect 68704 3680 68710 3692
rect 72050 3652 72056 3664
rect 72011 3624 72056 3652
rect 72050 3612 72056 3624
rect 72108 3612 72114 3664
rect 72145 3655 72203 3661
rect 72145 3621 72157 3655
rect 72191 3652 72203 3655
rect 73614 3652 73620 3664
rect 72191 3624 73620 3652
rect 72191 3621 72203 3624
rect 72145 3615 72203 3621
rect 73614 3612 73620 3624
rect 73672 3612 73678 3664
rect 75914 3612 75920 3664
rect 75972 3652 75978 3664
rect 76101 3655 76159 3661
rect 76101 3652 76113 3655
rect 75972 3624 76113 3652
rect 75972 3612 75978 3624
rect 76101 3621 76113 3624
rect 76147 3652 76159 3655
rect 76282 3652 76288 3664
rect 76147 3624 76288 3652
rect 76147 3621 76159 3624
rect 76101 3615 76159 3621
rect 76282 3612 76288 3624
rect 76340 3652 76346 3664
rect 76837 3655 76895 3661
rect 76837 3652 76849 3655
rect 76340 3624 76849 3652
rect 76340 3612 76346 3624
rect 76837 3621 76849 3624
rect 76883 3621 76895 3655
rect 80698 3652 80704 3664
rect 80659 3624 80704 3652
rect 76837 3615 76895 3621
rect 80698 3612 80704 3624
rect 80756 3612 80762 3664
rect 83461 3655 83519 3661
rect 83461 3621 83473 3655
rect 83507 3652 83519 3655
rect 84838 3652 84844 3664
rect 83507 3624 84844 3652
rect 83507 3621 83519 3624
rect 83461 3615 83519 3621
rect 84838 3612 84844 3624
rect 84896 3612 84902 3664
rect 71501 3587 71559 3593
rect 71501 3553 71513 3587
rect 71547 3584 71559 3587
rect 71961 3587 72019 3593
rect 71961 3584 71973 3587
rect 71547 3556 71973 3584
rect 71547 3553 71559 3556
rect 71501 3547 71559 3553
rect 71961 3553 71973 3556
rect 72007 3584 72019 3587
rect 74442 3584 74448 3596
rect 72007 3556 74448 3584
rect 72007 3553 72019 3556
rect 71961 3547 72019 3553
rect 74442 3544 74448 3556
rect 74500 3544 74506 3596
rect 78766 3544 78772 3596
rect 78824 3584 78830 3596
rect 80057 3587 80115 3593
rect 80057 3584 80069 3587
rect 78824 3556 80069 3584
rect 78824 3544 78830 3556
rect 80057 3553 80069 3556
rect 80103 3553 80115 3587
rect 83642 3584 83648 3596
rect 80057 3547 80115 3553
rect 82556 3556 83648 3584
rect 65153 3519 65211 3525
rect 65153 3516 65165 3519
rect 64656 3488 65165 3516
rect 64656 3476 64662 3488
rect 65153 3485 65165 3488
rect 65199 3516 65211 3519
rect 67913 3519 67971 3525
rect 65199 3488 66024 3516
rect 65199 3485 65211 3488
rect 65153 3479 65211 3485
rect 58437 3451 58495 3457
rect 58437 3448 58449 3451
rect 55916 3420 56442 3448
rect 57256 3420 58449 3448
rect 55916 3408 55922 3420
rect 57256 3380 57284 3420
rect 58437 3417 58449 3420
rect 58483 3417 58495 3451
rect 58437 3411 58495 3417
rect 62298 3408 62304 3460
rect 62356 3448 62362 3460
rect 63773 3451 63831 3457
rect 62356 3420 62606 3448
rect 62356 3408 62362 3420
rect 63773 3417 63785 3451
rect 63819 3448 63831 3451
rect 65797 3451 65855 3457
rect 65797 3448 65809 3451
rect 63819 3420 65809 3448
rect 63819 3417 63831 3420
rect 63773 3411 63831 3417
rect 65797 3417 65809 3420
rect 65843 3448 65855 3451
rect 65886 3448 65892 3460
rect 65843 3420 65892 3448
rect 65843 3417 65855 3420
rect 65797 3411 65855 3417
rect 65886 3408 65892 3420
rect 65944 3408 65950 3460
rect 65996 3448 66024 3488
rect 67913 3485 67925 3519
rect 67959 3485 67971 3519
rect 67913 3479 67971 3485
rect 72237 3519 72295 3525
rect 72237 3485 72249 3519
rect 72283 3516 72295 3519
rect 73798 3516 73804 3528
rect 72283 3488 73804 3516
rect 72283 3485 72295 3488
rect 72237 3479 72295 3485
rect 73798 3476 73804 3488
rect 73856 3476 73862 3528
rect 76374 3476 76380 3528
rect 76432 3516 76438 3528
rect 79597 3519 79655 3525
rect 76432 3488 78076 3516
rect 76432 3476 76438 3488
rect 73341 3451 73399 3457
rect 73341 3448 73353 3451
rect 65996 3420 73353 3448
rect 73341 3417 73353 3420
rect 73387 3417 73399 3451
rect 73341 3411 73399 3417
rect 57422 3380 57428 3392
rect 55692 3352 57284 3380
rect 57383 3352 57428 3380
rect 57422 3340 57428 3352
rect 57480 3340 57486 3392
rect 68097 3383 68155 3389
rect 68097 3349 68109 3383
rect 68143 3380 68155 3383
rect 68370 3380 68376 3392
rect 68143 3352 68376 3380
rect 68143 3349 68155 3352
rect 68097 3343 68155 3349
rect 68370 3340 68376 3352
rect 68428 3340 68434 3392
rect 71222 3340 71228 3392
rect 71280 3380 71286 3392
rect 72878 3380 72884 3392
rect 71280 3352 72884 3380
rect 71280 3340 71286 3352
rect 72878 3340 72884 3352
rect 72936 3340 72942 3392
rect 73356 3380 73384 3411
rect 73706 3408 73712 3460
rect 73764 3448 73770 3460
rect 73764 3420 77892 3448
rect 73764 3408 73770 3420
rect 77864 3392 77892 3420
rect 73982 3380 73988 3392
rect 73356 3352 73988 3380
rect 73982 3340 73988 3352
rect 74040 3340 74046 3392
rect 77846 3380 77852 3392
rect 77807 3352 77852 3380
rect 77846 3340 77852 3352
rect 77904 3340 77910 3392
rect 78048 3380 78076 3488
rect 79597 3485 79609 3519
rect 79643 3485 79655 3519
rect 81710 3516 81716 3528
rect 81671 3488 81716 3516
rect 79597 3479 79655 3485
rect 79042 3448 79048 3460
rect 78890 3420 79048 3448
rect 79042 3408 79048 3420
rect 79100 3408 79106 3460
rect 79226 3408 79232 3460
rect 79284 3448 79290 3460
rect 79321 3451 79379 3457
rect 79321 3448 79333 3451
rect 79284 3420 79333 3448
rect 79284 3408 79290 3420
rect 79321 3417 79333 3420
rect 79367 3417 79379 3451
rect 79321 3411 79379 3417
rect 79612 3380 79640 3479
rect 81710 3476 81716 3488
rect 81768 3476 81774 3528
rect 81986 3516 81992 3528
rect 81947 3488 81992 3516
rect 81986 3476 81992 3488
rect 82044 3516 82050 3528
rect 82556 3516 82584 3556
rect 83642 3544 83648 3556
rect 83700 3584 83706 3596
rect 83921 3587 83979 3593
rect 83921 3584 83933 3587
rect 83700 3556 83933 3584
rect 83700 3544 83706 3556
rect 83921 3553 83933 3556
rect 83967 3584 83979 3587
rect 85301 3587 85359 3593
rect 85301 3584 85313 3587
rect 83967 3556 85313 3584
rect 83967 3553 83979 3556
rect 83921 3547 83979 3553
rect 85301 3553 85313 3556
rect 85347 3584 85359 3587
rect 85666 3584 85672 3596
rect 85347 3556 85672 3584
rect 85347 3553 85359 3556
rect 85301 3547 85359 3553
rect 85666 3544 85672 3556
rect 85724 3544 85730 3596
rect 82722 3516 82728 3528
rect 82044 3488 82584 3516
rect 82683 3488 82728 3516
rect 82044 3476 82050 3488
rect 82722 3476 82728 3488
rect 82780 3476 82786 3528
rect 84841 3519 84899 3525
rect 84841 3485 84853 3519
rect 84887 3516 84899 3519
rect 84930 3516 84936 3528
rect 84887 3488 84936 3516
rect 84887 3485 84899 3488
rect 84841 3479 84899 3485
rect 84930 3476 84936 3488
rect 84988 3476 84994 3528
rect 79870 3408 79876 3460
rect 79928 3448 79934 3460
rect 82909 3451 82967 3457
rect 82909 3448 82921 3451
rect 79928 3420 82921 3448
rect 79928 3408 79934 3420
rect 82909 3417 82921 3420
rect 82955 3417 82967 3451
rect 85960 3448 85988 3692
rect 86034 3680 86040 3732
rect 86092 3720 86098 3732
rect 86405 3723 86463 3729
rect 86405 3720 86417 3723
rect 86092 3692 86417 3720
rect 86092 3680 86098 3692
rect 86405 3689 86417 3692
rect 86451 3689 86463 3723
rect 86405 3683 86463 3689
rect 87417 3723 87475 3729
rect 87417 3689 87429 3723
rect 87463 3720 87475 3723
rect 88518 3720 88524 3732
rect 87463 3692 88524 3720
rect 87463 3689 87475 3692
rect 87417 3683 87475 3689
rect 88518 3680 88524 3692
rect 88576 3680 88582 3732
rect 89990 3680 89996 3732
rect 90048 3720 90054 3732
rect 90821 3723 90879 3729
rect 90821 3720 90833 3723
rect 90048 3692 90833 3720
rect 90048 3680 90054 3692
rect 90821 3689 90833 3692
rect 90867 3720 90879 3723
rect 90910 3720 90916 3732
rect 90867 3692 90916 3720
rect 90867 3689 90879 3692
rect 90821 3683 90879 3689
rect 90910 3680 90916 3692
rect 90968 3680 90974 3732
rect 93210 3720 93216 3732
rect 93171 3692 93216 3720
rect 93210 3680 93216 3692
rect 93268 3680 93274 3732
rect 87230 3612 87236 3664
rect 87288 3652 87294 3664
rect 87877 3655 87935 3661
rect 87877 3652 87889 3655
rect 87288 3624 87889 3652
rect 87288 3612 87294 3624
rect 87877 3621 87889 3624
rect 87923 3621 87935 3655
rect 87877 3615 87935 3621
rect 88429 3655 88487 3661
rect 88429 3621 88441 3655
rect 88475 3652 88487 3655
rect 88978 3652 88984 3664
rect 88475 3624 88984 3652
rect 88475 3621 88487 3624
rect 88429 3615 88487 3621
rect 88978 3612 88984 3624
rect 89036 3612 89042 3664
rect 92661 3655 92719 3661
rect 92661 3621 92673 3655
rect 92707 3652 92719 3655
rect 93670 3652 93676 3664
rect 92707 3624 93676 3652
rect 92707 3621 92719 3624
rect 92661 3615 92719 3621
rect 93670 3612 93676 3624
rect 93728 3612 93734 3664
rect 88886 3584 88892 3596
rect 86972 3556 88892 3584
rect 86972 3525 87000 3556
rect 88886 3544 88892 3556
rect 88944 3544 88950 3596
rect 89346 3584 89352 3596
rect 89307 3556 89352 3584
rect 89346 3544 89352 3556
rect 89404 3544 89410 3596
rect 86957 3519 87015 3525
rect 86957 3485 86969 3519
rect 87003 3485 87015 3519
rect 86957 3479 87015 3485
rect 87046 3476 87052 3528
rect 87104 3516 87110 3528
rect 87233 3519 87291 3525
rect 87104 3488 87149 3516
rect 87104 3476 87110 3488
rect 87233 3485 87245 3519
rect 87279 3485 87291 3519
rect 89070 3516 89076 3528
rect 89031 3488 89076 3516
rect 87233 3479 87291 3485
rect 86862 3448 86868 3460
rect 85960 3420 86868 3448
rect 82909 3411 82967 3417
rect 86862 3408 86868 3420
rect 86920 3448 86926 3460
rect 87248 3448 87276 3479
rect 89070 3476 89076 3488
rect 89128 3476 89134 3528
rect 91922 3516 91928 3528
rect 91883 3488 91928 3516
rect 91922 3476 91928 3488
rect 91980 3476 91986 3528
rect 94041 3519 94099 3525
rect 94041 3516 94053 3519
rect 92124 3488 94053 3516
rect 86920 3420 87276 3448
rect 86920 3408 86926 3420
rect 89898 3408 89904 3460
rect 89956 3408 89962 3460
rect 80698 3380 80704 3392
rect 78048 3352 80704 3380
rect 80698 3340 80704 3352
rect 80756 3340 80762 3392
rect 92124 3389 92152 3488
rect 94041 3485 94053 3488
rect 94087 3485 94099 3519
rect 94041 3479 94099 3485
rect 92109 3383 92167 3389
rect 92109 3349 92121 3383
rect 92155 3349 92167 3383
rect 92109 3343 92167 3349
rect 93762 3340 93768 3392
rect 93820 3380 93826 3392
rect 94225 3383 94283 3389
rect 94225 3380 94237 3383
rect 93820 3352 94237 3380
rect 93820 3340 93826 3352
rect 94225 3349 94237 3352
rect 94271 3349 94283 3383
rect 94225 3343 94283 3349
rect 1104 3290 95011 3312
rect 1104 3238 24386 3290
rect 24438 3238 24450 3290
rect 24502 3238 24514 3290
rect 24566 3238 24578 3290
rect 24630 3238 24642 3290
rect 24694 3238 47823 3290
rect 47875 3238 47887 3290
rect 47939 3238 47951 3290
rect 48003 3238 48015 3290
rect 48067 3238 48079 3290
rect 48131 3238 71260 3290
rect 71312 3238 71324 3290
rect 71376 3238 71388 3290
rect 71440 3238 71452 3290
rect 71504 3238 71516 3290
rect 71568 3238 94697 3290
rect 94749 3238 94761 3290
rect 94813 3238 94825 3290
rect 94877 3238 94889 3290
rect 94941 3238 94953 3290
rect 95005 3238 95011 3290
rect 1104 3216 95011 3238
rect 37553 3179 37611 3185
rect 37553 3145 37565 3179
rect 37599 3176 37611 3179
rect 37734 3176 37740 3188
rect 37599 3148 37740 3176
rect 37599 3145 37611 3148
rect 37553 3139 37611 3145
rect 37734 3136 37740 3148
rect 37792 3136 37798 3188
rect 38838 3136 38844 3188
rect 38896 3136 38902 3188
rect 53834 3176 53840 3188
rect 53795 3148 53840 3176
rect 53834 3136 53840 3148
rect 53892 3136 53898 3188
rect 54389 3179 54447 3185
rect 54389 3145 54401 3179
rect 54435 3176 54447 3179
rect 54941 3179 54999 3185
rect 54941 3176 54953 3179
rect 54435 3148 54953 3176
rect 54435 3145 54447 3148
rect 54389 3139 54447 3145
rect 54941 3145 54953 3148
rect 54987 3176 54999 3179
rect 55030 3176 55036 3188
rect 54987 3148 55036 3176
rect 54987 3145 54999 3148
rect 54941 3139 54999 3145
rect 38856 3108 38884 3136
rect 39022 3108 39028 3120
rect 38594 3080 38884 3108
rect 38983 3080 39028 3108
rect 39022 3068 39028 3080
rect 39080 3108 39086 3120
rect 39761 3111 39819 3117
rect 39761 3108 39773 3111
rect 39080 3080 39773 3108
rect 39080 3068 39086 3080
rect 39761 3077 39773 3080
rect 39807 3077 39819 3111
rect 39761 3071 39819 3077
rect 53009 3111 53067 3117
rect 53009 3077 53021 3111
rect 53055 3108 53067 3111
rect 53926 3108 53932 3120
rect 53055 3080 53932 3108
rect 53055 3077 53067 3080
rect 53009 3071 53067 3077
rect 53926 3068 53932 3080
rect 53984 3068 53990 3120
rect 39301 3043 39359 3049
rect 39301 3009 39313 3043
rect 39347 3040 39359 3043
rect 40402 3040 40408 3052
rect 39347 3012 40408 3040
rect 39347 3009 39359 3012
rect 39301 3003 39359 3009
rect 40402 3000 40408 3012
rect 40460 3000 40466 3052
rect 51258 3040 51264 3052
rect 51171 3012 51264 3040
rect 51258 3000 51264 3012
rect 51316 3040 51322 3052
rect 51813 3043 51871 3049
rect 51813 3040 51825 3043
rect 51316 3012 51825 3040
rect 51316 3000 51322 3012
rect 51813 3009 51825 3012
rect 51859 3040 51871 3043
rect 52362 3040 52368 3052
rect 51859 3012 52368 3040
rect 51859 3009 51871 3012
rect 51813 3003 51871 3009
rect 52362 3000 52368 3012
rect 52420 3040 52426 3052
rect 54404 3040 54432 3139
rect 55030 3136 55036 3148
rect 55088 3176 55094 3188
rect 55493 3179 55551 3185
rect 55493 3176 55505 3179
rect 55088 3148 55505 3176
rect 55088 3136 55094 3148
rect 55493 3145 55505 3148
rect 55539 3176 55551 3179
rect 55858 3176 55864 3188
rect 55539 3148 55864 3176
rect 55539 3145 55551 3148
rect 55493 3139 55551 3145
rect 55858 3136 55864 3148
rect 55916 3136 55922 3188
rect 56226 3176 56232 3188
rect 56187 3148 56232 3176
rect 56226 3136 56232 3148
rect 56284 3136 56290 3188
rect 56778 3136 56784 3188
rect 56836 3176 56842 3188
rect 57149 3179 57207 3185
rect 57149 3176 57161 3179
rect 56836 3148 57161 3176
rect 56836 3136 56842 3148
rect 57149 3145 57161 3148
rect 57195 3176 57207 3179
rect 57330 3176 57336 3188
rect 57195 3148 57336 3176
rect 57195 3145 57207 3148
rect 57149 3139 57207 3145
rect 57330 3136 57336 3148
rect 57388 3136 57394 3188
rect 57422 3136 57428 3188
rect 57480 3176 57486 3188
rect 57480 3148 64736 3176
rect 57480 3136 57486 3148
rect 61286 3108 61292 3120
rect 61247 3080 61292 3108
rect 61286 3068 61292 3080
rect 61344 3068 61350 3120
rect 62298 3068 62304 3120
rect 62356 3108 62362 3120
rect 64708 3117 64736 3148
rect 64782 3136 64788 3188
rect 64840 3176 64846 3188
rect 78582 3176 78588 3188
rect 64840 3148 78588 3176
rect 64840 3136 64846 3148
rect 78582 3136 78588 3148
rect 78640 3136 78646 3188
rect 79226 3176 79232 3188
rect 79187 3148 79232 3176
rect 79226 3136 79232 3148
rect 79284 3136 79290 3188
rect 80609 3179 80667 3185
rect 80609 3176 80621 3179
rect 80026 3148 80621 3176
rect 64693 3111 64751 3117
rect 62356 3080 63526 3108
rect 62356 3068 62362 3080
rect 64693 3077 64705 3111
rect 64739 3077 64751 3111
rect 64693 3071 64751 3077
rect 72878 3068 72884 3120
rect 72936 3108 72942 3120
rect 74626 3108 74632 3120
rect 72936 3080 74632 3108
rect 72936 3068 72942 3080
rect 74626 3068 74632 3080
rect 74684 3068 74690 3120
rect 76282 3108 76288 3120
rect 76243 3080 76288 3108
rect 76282 3068 76288 3080
rect 76340 3068 76346 3120
rect 77481 3111 77539 3117
rect 77481 3077 77493 3111
rect 77527 3108 77539 3111
rect 78030 3108 78036 3120
rect 77527 3080 78036 3108
rect 77527 3077 77539 3080
rect 77481 3071 77539 3077
rect 78030 3068 78036 3080
rect 78088 3068 78094 3120
rect 78600 3108 78628 3136
rect 80026 3108 80054 3148
rect 80609 3145 80621 3148
rect 80655 3176 80667 3179
rect 81434 3176 81440 3188
rect 80655 3148 81440 3176
rect 80655 3145 80667 3148
rect 80609 3139 80667 3145
rect 81434 3136 81440 3148
rect 81492 3136 81498 3188
rect 81526 3136 81532 3188
rect 81584 3176 81590 3188
rect 81986 3176 81992 3188
rect 81584 3148 81992 3176
rect 81584 3136 81590 3148
rect 81986 3136 81992 3148
rect 82044 3136 82050 3188
rect 84930 3136 84936 3188
rect 84988 3176 84994 3188
rect 85209 3179 85267 3185
rect 85209 3176 85221 3179
rect 84988 3148 85221 3176
rect 84988 3136 84994 3148
rect 85209 3145 85221 3148
rect 85255 3176 85267 3179
rect 85945 3179 86003 3185
rect 85945 3176 85957 3179
rect 85255 3148 85957 3176
rect 85255 3145 85267 3148
rect 85209 3139 85267 3145
rect 85945 3145 85957 3148
rect 85991 3145 86003 3179
rect 85945 3139 86003 3145
rect 78600 3080 80054 3108
rect 85960 3108 85988 3139
rect 86862 3136 86868 3188
rect 86920 3176 86926 3188
rect 90453 3179 90511 3185
rect 90453 3176 90465 3179
rect 86920 3148 90465 3176
rect 86920 3136 86926 3148
rect 90453 3145 90465 3148
rect 90499 3176 90511 3179
rect 90818 3176 90824 3188
rect 90499 3148 90824 3176
rect 90499 3145 90511 3148
rect 90453 3139 90511 3145
rect 90818 3136 90824 3148
rect 90876 3136 90882 3188
rect 91002 3176 91008 3188
rect 90963 3148 91008 3176
rect 91002 3136 91008 3148
rect 91060 3136 91066 3188
rect 92017 3179 92075 3185
rect 92017 3145 92029 3179
rect 92063 3176 92075 3179
rect 92382 3176 92388 3188
rect 92063 3148 92388 3176
rect 92063 3145 92075 3148
rect 92017 3139 92075 3145
rect 92382 3136 92388 3148
rect 92440 3136 92446 3188
rect 89622 3108 89628 3120
rect 85960 3080 89628 3108
rect 89622 3068 89628 3080
rect 89680 3108 89686 3120
rect 89809 3111 89867 3117
rect 89809 3108 89821 3111
rect 89680 3080 89821 3108
rect 89680 3068 89686 3080
rect 89809 3077 89821 3080
rect 89855 3077 89867 3111
rect 89809 3071 89867 3077
rect 52420 3012 54432 3040
rect 52420 3000 52426 3012
rect 55122 3000 55128 3052
rect 55180 3040 55186 3052
rect 55180 3012 63356 3040
rect 55180 3000 55186 3012
rect 54386 2932 54392 2984
rect 54444 2972 54450 2984
rect 55490 2972 55496 2984
rect 54444 2944 55496 2972
rect 54444 2932 54450 2944
rect 55490 2932 55496 2944
rect 55548 2932 55554 2984
rect 57054 2864 57060 2916
rect 57112 2904 57118 2916
rect 63221 2907 63279 2913
rect 63221 2904 63233 2907
rect 57112 2876 63233 2904
rect 57112 2864 57118 2876
rect 63221 2873 63233 2876
rect 63267 2873 63279 2907
rect 63221 2867 63279 2873
rect 63328 2836 63356 3012
rect 77846 3000 77852 3052
rect 77904 3040 77910 3052
rect 78861 3043 78919 3049
rect 78861 3040 78873 3043
rect 77904 3012 78873 3040
rect 77904 3000 77910 3012
rect 78861 3009 78873 3012
rect 78907 3009 78919 3043
rect 79870 3040 79876 3052
rect 79831 3012 79876 3040
rect 78861 3003 78919 3009
rect 79870 3000 79876 3012
rect 79928 3000 79934 3052
rect 85666 3000 85672 3052
rect 85724 3040 85730 3052
rect 86589 3043 86647 3049
rect 86589 3040 86601 3043
rect 85724 3012 86601 3040
rect 85724 3000 85730 3012
rect 86589 3009 86601 3012
rect 86635 3040 86647 3043
rect 87141 3043 87199 3049
rect 87141 3040 87153 3043
rect 86635 3012 87153 3040
rect 86635 3009 86647 3012
rect 86589 3003 86647 3009
rect 87141 3009 87153 3012
rect 87187 3009 87199 3043
rect 87141 3003 87199 3009
rect 64966 2932 64972 2984
rect 65024 2972 65030 2984
rect 65429 2975 65487 2981
rect 65429 2972 65441 2975
rect 65024 2944 65441 2972
rect 65024 2932 65030 2944
rect 65429 2941 65441 2944
rect 65475 2941 65487 2975
rect 65429 2935 65487 2941
rect 78674 2932 78680 2984
rect 78732 2972 78738 2984
rect 78769 2975 78827 2981
rect 78769 2972 78781 2975
rect 78732 2944 78781 2972
rect 78732 2932 78738 2944
rect 78769 2941 78781 2944
rect 78815 2941 78827 2975
rect 78769 2935 78827 2941
rect 81710 2932 81716 2984
rect 81768 2972 81774 2984
rect 82633 2975 82691 2981
rect 82633 2972 82645 2975
rect 81768 2944 82645 2972
rect 81768 2932 81774 2944
rect 82633 2941 82645 2944
rect 82679 2972 82691 2975
rect 83185 2975 83243 2981
rect 83185 2972 83197 2975
rect 82679 2944 83197 2972
rect 82679 2941 82691 2944
rect 82633 2935 82691 2941
rect 83185 2941 83197 2944
rect 83231 2972 83243 2975
rect 83366 2972 83372 2984
rect 83231 2944 83372 2972
rect 83231 2941 83243 2944
rect 83185 2935 83243 2941
rect 83366 2932 83372 2944
rect 83424 2972 83430 2984
rect 84749 2975 84807 2981
rect 84749 2972 84761 2975
rect 83424 2944 84761 2972
rect 83424 2932 83430 2944
rect 84749 2941 84761 2944
rect 84795 2972 84807 2975
rect 86126 2972 86132 2984
rect 84795 2944 86132 2972
rect 84795 2941 84807 2944
rect 84749 2935 84807 2941
rect 86126 2932 86132 2944
rect 86184 2932 86190 2984
rect 89070 2932 89076 2984
rect 89128 2972 89134 2984
rect 91002 2972 91008 2984
rect 89128 2944 91008 2972
rect 89128 2932 89134 2944
rect 91002 2932 91008 2944
rect 91060 2932 91066 2984
rect 91922 2932 91928 2984
rect 91980 2932 91986 2984
rect 91940 2904 91968 2932
rect 92477 2907 92535 2913
rect 92477 2904 92489 2907
rect 67606 2876 92489 2904
rect 67606 2836 67634 2876
rect 92477 2873 92489 2876
rect 92523 2873 92535 2907
rect 92477 2867 92535 2873
rect 63328 2808 67634 2836
rect 78674 2796 78680 2848
rect 78732 2836 78738 2848
rect 79689 2839 79747 2845
rect 79689 2836 79701 2839
rect 78732 2808 79701 2836
rect 78732 2796 78738 2808
rect 79689 2805 79701 2808
rect 79735 2805 79747 2839
rect 79689 2799 79747 2805
rect 1104 2746 94852 2768
rect 1104 2694 12668 2746
rect 12720 2694 12732 2746
rect 12784 2694 12796 2746
rect 12848 2694 12860 2746
rect 12912 2694 12924 2746
rect 12976 2694 36105 2746
rect 36157 2694 36169 2746
rect 36221 2694 36233 2746
rect 36285 2694 36297 2746
rect 36349 2694 36361 2746
rect 36413 2694 59542 2746
rect 59594 2694 59606 2746
rect 59658 2694 59670 2746
rect 59722 2694 59734 2746
rect 59786 2694 59798 2746
rect 59850 2694 82979 2746
rect 83031 2694 83043 2746
rect 83095 2694 83107 2746
rect 83159 2694 83171 2746
rect 83223 2694 83235 2746
rect 83287 2694 94852 2746
rect 1104 2672 94852 2694
rect 36357 2635 36415 2641
rect 36357 2601 36369 2635
rect 36403 2632 36415 2635
rect 37366 2632 37372 2644
rect 36403 2604 37372 2632
rect 36403 2601 36415 2604
rect 36357 2595 36415 2601
rect 37366 2592 37372 2604
rect 37424 2592 37430 2644
rect 38838 2592 38844 2644
rect 38896 2632 38902 2644
rect 39393 2635 39451 2641
rect 39393 2632 39405 2635
rect 38896 2604 39405 2632
rect 38896 2592 38902 2604
rect 39393 2601 39405 2604
rect 39439 2601 39451 2635
rect 39393 2595 39451 2601
rect 41322 2592 41328 2644
rect 41380 2632 41386 2644
rect 44085 2635 44143 2641
rect 44085 2632 44097 2635
rect 41380 2604 44097 2632
rect 41380 2592 41386 2604
rect 44085 2601 44097 2604
rect 44131 2601 44143 2635
rect 54386 2632 54392 2644
rect 54347 2604 54392 2632
rect 44085 2595 44143 2601
rect 54386 2592 54392 2604
rect 54444 2592 54450 2644
rect 64322 2632 64328 2644
rect 64283 2604 64328 2632
rect 64322 2592 64328 2604
rect 64380 2632 64386 2644
rect 64966 2632 64972 2644
rect 64380 2604 64972 2632
rect 64380 2592 64386 2604
rect 64966 2592 64972 2604
rect 65024 2592 65030 2644
rect 75270 2592 75276 2644
rect 75328 2632 75334 2644
rect 78582 2632 78588 2644
rect 75328 2604 78588 2632
rect 75328 2592 75334 2604
rect 78582 2592 78588 2604
rect 78640 2592 78646 2644
rect 78766 2632 78772 2644
rect 78727 2604 78772 2632
rect 78766 2592 78772 2604
rect 78824 2592 78830 2644
rect 86862 2632 86868 2644
rect 86823 2604 86868 2632
rect 86862 2592 86868 2604
rect 86920 2592 86926 2644
rect 90910 2632 90916 2644
rect 90871 2604 90916 2632
rect 90910 2592 90916 2604
rect 90968 2592 90974 2644
rect 53377 2567 53435 2573
rect 53377 2533 53389 2567
rect 53423 2533 53435 2567
rect 53377 2527 53435 2533
rect 4154 2388 4160 2440
rect 4212 2428 4218 2440
rect 4525 2431 4583 2437
rect 4525 2428 4537 2431
rect 4212 2400 4537 2428
rect 4212 2388 4218 2400
rect 4525 2397 4537 2400
rect 4571 2397 4583 2431
rect 4525 2391 4583 2397
rect 12713 2431 12771 2437
rect 12713 2397 12725 2431
rect 12759 2428 12771 2431
rect 13354 2428 13360 2440
rect 12759 2400 13216 2428
rect 13315 2400 13360 2428
rect 12759 2397 12771 2400
rect 12713 2391 12771 2397
rect 4430 2252 4436 2304
rect 4488 2292 4494 2304
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 4488 2264 4721 2292
rect 4488 2252 4494 2264
rect 4709 2261 4721 2264
rect 4755 2261 4767 2295
rect 4709 2255 4767 2261
rect 12342 2252 12348 2304
rect 12400 2292 12406 2304
rect 13188 2301 13216 2400
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 15470 2388 15476 2440
rect 15528 2428 15534 2440
rect 20073 2431 20131 2437
rect 20073 2428 20085 2431
rect 15528 2400 20085 2428
rect 15528 2388 15534 2400
rect 20073 2397 20085 2400
rect 20119 2397 20131 2431
rect 20993 2431 21051 2437
rect 20993 2428 21005 2431
rect 20073 2391 20131 2397
rect 20272 2400 21005 2428
rect 20272 2301 20300 2400
rect 20993 2397 21005 2400
rect 21039 2397 21051 2431
rect 28442 2428 28448 2440
rect 28403 2400 28448 2428
rect 20993 2391 21051 2397
rect 28442 2388 28448 2400
rect 28500 2388 28506 2440
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 36173 2431 36231 2437
rect 36173 2428 36185 2431
rect 36136 2400 36185 2428
rect 36136 2388 36142 2400
rect 36173 2397 36185 2400
rect 36219 2428 36231 2431
rect 36817 2431 36875 2437
rect 36817 2428 36829 2431
rect 36219 2400 36829 2428
rect 36219 2397 36231 2400
rect 36173 2391 36231 2397
rect 36817 2397 36829 2400
rect 36863 2397 36875 2431
rect 44269 2431 44327 2437
rect 44269 2428 44281 2431
rect 36817 2391 36875 2397
rect 44008 2400 44281 2428
rect 44008 2304 44036 2400
rect 44269 2397 44281 2400
rect 44315 2397 44327 2431
rect 44269 2391 44327 2397
rect 52273 2431 52331 2437
rect 52273 2397 52285 2431
rect 52319 2428 52331 2431
rect 53392 2428 53420 2527
rect 64984 2496 65012 2592
rect 65886 2524 65892 2576
rect 65944 2564 65950 2576
rect 65944 2536 84194 2564
rect 65944 2524 65950 2536
rect 83829 2499 83887 2505
rect 83829 2496 83841 2499
rect 64984 2468 83841 2496
rect 83829 2465 83841 2468
rect 83875 2465 83887 2499
rect 84166 2496 84194 2536
rect 91833 2499 91891 2505
rect 91833 2496 91845 2499
rect 84166 2468 91845 2496
rect 83829 2459 83887 2465
rect 91833 2465 91845 2468
rect 91879 2465 91891 2499
rect 91833 2459 91891 2465
rect 52319 2400 53420 2428
rect 53561 2431 53619 2437
rect 52319 2397 52331 2400
rect 52273 2391 52331 2397
rect 53561 2397 53573 2431
rect 53607 2428 53619 2431
rect 56318 2428 56324 2440
rect 53607 2400 56324 2428
rect 53607 2397 53619 2400
rect 53561 2391 53619 2397
rect 56318 2388 56324 2400
rect 56376 2388 56382 2440
rect 60921 2431 60979 2437
rect 60921 2397 60933 2431
rect 60967 2428 60979 2431
rect 68370 2428 68376 2440
rect 60967 2400 61516 2428
rect 68331 2400 68376 2428
rect 60967 2397 60979 2400
rect 60921 2391 60979 2397
rect 61488 2369 61516 2400
rect 68370 2388 68376 2400
rect 68428 2388 68434 2440
rect 74810 2388 74816 2440
rect 74868 2428 74874 2440
rect 75181 2431 75239 2437
rect 75181 2428 75193 2431
rect 74868 2400 75193 2428
rect 74868 2388 74874 2400
rect 75181 2397 75193 2400
rect 75227 2397 75239 2431
rect 76101 2431 76159 2437
rect 76101 2428 76113 2431
rect 75181 2391 75239 2397
rect 75564 2400 76113 2428
rect 61473 2363 61531 2369
rect 61473 2329 61485 2363
rect 61519 2360 61531 2363
rect 75270 2360 75276 2372
rect 61519 2332 75276 2360
rect 61519 2329 61531 2332
rect 61473 2323 61531 2329
rect 75270 2320 75276 2332
rect 75328 2320 75334 2372
rect 12529 2295 12587 2301
rect 12529 2292 12541 2295
rect 12400 2264 12541 2292
rect 12400 2252 12406 2264
rect 12529 2261 12541 2264
rect 12575 2261 12587 2295
rect 12529 2255 12587 2261
rect 13173 2295 13231 2301
rect 13173 2261 13185 2295
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 20257 2295 20315 2301
rect 20257 2261 20269 2295
rect 20303 2261 20315 2295
rect 20257 2255 20315 2261
rect 20346 2252 20352 2304
rect 20404 2292 20410 2304
rect 20809 2295 20867 2301
rect 20809 2292 20821 2295
rect 20404 2264 20821 2292
rect 20404 2252 20410 2264
rect 20809 2261 20821 2264
rect 20855 2261 20867 2295
rect 20809 2255 20867 2261
rect 28166 2252 28172 2304
rect 28224 2292 28230 2304
rect 28261 2295 28319 2301
rect 28261 2292 28273 2295
rect 28224 2264 28273 2292
rect 28224 2252 28230 2264
rect 28261 2261 28273 2264
rect 28307 2261 28319 2295
rect 28261 2255 28319 2261
rect 43625 2295 43683 2301
rect 43625 2261 43637 2295
rect 43671 2292 43683 2295
rect 43990 2292 43996 2304
rect 43671 2264 43996 2292
rect 43671 2261 43683 2264
rect 43625 2255 43683 2261
rect 43990 2252 43996 2264
rect 44048 2252 44054 2304
rect 51902 2252 51908 2304
rect 51960 2292 51966 2304
rect 52089 2295 52147 2301
rect 52089 2292 52101 2295
rect 51960 2264 52101 2292
rect 51960 2252 51966 2264
rect 52089 2261 52101 2264
rect 52135 2261 52147 2295
rect 52089 2255 52147 2261
rect 59814 2252 59820 2304
rect 59872 2292 59878 2304
rect 60737 2295 60795 2301
rect 60737 2292 60749 2295
rect 59872 2264 60749 2292
rect 59872 2252 59878 2264
rect 60737 2261 60749 2264
rect 60783 2261 60795 2295
rect 60737 2255 60795 2261
rect 67726 2252 67732 2304
rect 67784 2292 67790 2304
rect 68557 2295 68615 2301
rect 68557 2292 68569 2295
rect 67784 2264 68569 2292
rect 67784 2252 67790 2264
rect 68557 2261 68569 2264
rect 68603 2261 68615 2295
rect 68557 2255 68615 2261
rect 75365 2295 75423 2301
rect 75365 2261 75377 2295
rect 75411 2292 75423 2295
rect 75564 2292 75592 2400
rect 76101 2397 76113 2400
rect 76147 2397 76159 2431
rect 76101 2391 76159 2397
rect 91462 2388 91468 2440
rect 91520 2428 91526 2440
rect 91557 2431 91615 2437
rect 91557 2428 91569 2431
rect 91520 2400 91569 2428
rect 91520 2388 91526 2400
rect 91557 2397 91569 2400
rect 91603 2428 91615 2431
rect 92845 2431 92903 2437
rect 92845 2428 92857 2431
rect 91603 2400 92857 2428
rect 91603 2397 91615 2400
rect 91557 2391 91615 2397
rect 92845 2397 92857 2400
rect 92891 2397 92903 2431
rect 92845 2391 92903 2397
rect 84013 2363 84071 2369
rect 84013 2360 84025 2363
rect 83568 2332 84025 2360
rect 83568 2304 83596 2332
rect 84013 2329 84025 2332
rect 84059 2329 84071 2363
rect 84013 2323 84071 2329
rect 75411 2264 75592 2292
rect 75411 2261 75423 2264
rect 75365 2255 75423 2261
rect 75638 2252 75644 2304
rect 75696 2292 75702 2304
rect 76285 2295 76343 2301
rect 76285 2292 76297 2295
rect 75696 2264 76297 2292
rect 75696 2252 75702 2264
rect 76285 2261 76297 2264
rect 76331 2261 76343 2295
rect 76285 2255 76343 2261
rect 83277 2295 83335 2301
rect 83277 2261 83289 2295
rect 83323 2292 83335 2295
rect 83550 2292 83556 2304
rect 83323 2264 83556 2292
rect 83323 2261 83335 2264
rect 83277 2255 83335 2261
rect 83550 2252 83556 2264
rect 83608 2252 83614 2304
rect 1104 2202 95011 2224
rect 1104 2150 24386 2202
rect 24438 2150 24450 2202
rect 24502 2150 24514 2202
rect 24566 2150 24578 2202
rect 24630 2150 24642 2202
rect 24694 2150 47823 2202
rect 47875 2150 47887 2202
rect 47939 2150 47951 2202
rect 48003 2150 48015 2202
rect 48067 2150 48079 2202
rect 48131 2150 71260 2202
rect 71312 2150 71324 2202
rect 71376 2150 71388 2202
rect 71440 2150 71452 2202
rect 71504 2150 71516 2202
rect 71568 2150 94697 2202
rect 94749 2150 94761 2202
rect 94813 2150 94825 2202
rect 94877 2150 94889 2202
rect 94941 2150 94953 2202
rect 95005 2150 95011 2202
rect 1104 2128 95011 2150
<< via1 >>
rect 20904 17484 20956 17536
rect 69664 17484 69716 17536
rect 24386 17382 24438 17434
rect 24450 17382 24502 17434
rect 24514 17382 24566 17434
rect 24578 17382 24630 17434
rect 24642 17382 24694 17434
rect 47823 17382 47875 17434
rect 47887 17382 47939 17434
rect 47951 17382 48003 17434
rect 48015 17382 48067 17434
rect 48079 17382 48131 17434
rect 71260 17382 71312 17434
rect 71324 17382 71376 17434
rect 71388 17382 71440 17434
rect 71452 17382 71504 17434
rect 71516 17382 71568 17434
rect 94697 17382 94749 17434
rect 94761 17382 94813 17434
rect 94825 17382 94877 17434
rect 94889 17382 94941 17434
rect 94953 17382 95005 17434
rect 4436 17280 4488 17332
rect 1584 17144 1636 17196
rect 12440 17280 12492 17332
rect 20260 17280 20312 17332
rect 28172 17280 28224 17332
rect 34336 17255 34388 17264
rect 6552 17144 6604 17196
rect 5080 16940 5132 16992
rect 34336 17221 34345 17255
rect 34345 17221 34379 17255
rect 34379 17221 34388 17255
rect 43996 17280 44048 17332
rect 50344 17280 50396 17332
rect 51908 17280 51960 17332
rect 59820 17280 59872 17332
rect 67732 17280 67784 17332
rect 75644 17280 75696 17332
rect 34336 17212 34388 17221
rect 11888 17144 11940 17196
rect 20536 17187 20588 17196
rect 20536 17153 20545 17187
rect 20545 17153 20579 17187
rect 20579 17153 20588 17187
rect 20536 17144 20588 17153
rect 28448 17187 28500 17196
rect 28448 17153 28457 17187
rect 28457 17153 28491 17187
rect 28491 17153 28500 17187
rect 28448 17144 28500 17153
rect 43996 17144 44048 17196
rect 34888 17119 34940 17128
rect 34888 17085 34897 17119
rect 34897 17085 34931 17119
rect 34931 17085 34940 17119
rect 34888 17076 34940 17085
rect 36912 17119 36964 17128
rect 36912 17085 36921 17119
rect 36921 17085 36955 17119
rect 36955 17085 36964 17119
rect 36912 17076 36964 17085
rect 49516 17212 49568 17264
rect 57060 17212 57112 17264
rect 52276 17187 52328 17196
rect 52276 17153 52285 17187
rect 52285 17153 52319 17187
rect 52319 17153 52328 17187
rect 52276 17144 52328 17153
rect 65892 17212 65944 17264
rect 84016 17212 84068 17264
rect 46204 17076 46256 17128
rect 59360 17076 59412 17128
rect 55128 17008 55180 17060
rect 57980 17008 58032 17060
rect 68376 17187 68428 17196
rect 68376 17153 68385 17187
rect 68385 17153 68419 17187
rect 68419 17153 68428 17187
rect 68376 17144 68428 17153
rect 76104 17187 76156 17196
rect 76104 17153 76113 17187
rect 76113 17153 76147 17187
rect 76147 17153 76156 17187
rect 76104 17144 76156 17153
rect 91468 17144 91520 17196
rect 61844 17076 61896 17128
rect 63592 17076 63644 17128
rect 65800 17119 65852 17128
rect 65800 17085 65809 17119
rect 65809 17085 65843 17119
rect 65843 17085 65852 17119
rect 65800 17076 65852 17085
rect 83372 17076 83424 17128
rect 62856 17008 62908 17060
rect 67548 17008 67600 17060
rect 83740 17008 83792 17060
rect 32220 16940 32272 16992
rect 38660 16940 38712 16992
rect 40592 16940 40644 16992
rect 46020 16940 46072 16992
rect 46480 16983 46532 16992
rect 46480 16949 46489 16983
rect 46489 16949 46523 16983
rect 46523 16949 46532 16983
rect 46480 16940 46532 16949
rect 47032 16983 47084 16992
rect 47032 16949 47041 16983
rect 47041 16949 47075 16983
rect 47075 16949 47084 16983
rect 47032 16940 47084 16949
rect 56692 16940 56744 16992
rect 60740 16940 60792 16992
rect 61108 16940 61160 16992
rect 12668 16838 12720 16890
rect 12732 16838 12784 16890
rect 12796 16838 12848 16890
rect 12860 16838 12912 16890
rect 12924 16838 12976 16890
rect 36105 16838 36157 16890
rect 36169 16838 36221 16890
rect 36233 16838 36285 16890
rect 36297 16838 36349 16890
rect 36361 16838 36413 16890
rect 59542 16838 59594 16890
rect 59606 16838 59658 16890
rect 59670 16838 59722 16890
rect 59734 16838 59786 16890
rect 59798 16838 59850 16890
rect 82979 16838 83031 16890
rect 83043 16838 83095 16890
rect 83107 16838 83159 16890
rect 83171 16838 83223 16890
rect 83235 16838 83287 16890
rect 36912 16736 36964 16788
rect 38660 16736 38712 16788
rect 46204 16736 46256 16788
rect 50344 16779 50396 16788
rect 50344 16745 50353 16779
rect 50353 16745 50387 16779
rect 50387 16745 50396 16779
rect 50344 16736 50396 16745
rect 50528 16736 50580 16788
rect 55128 16736 55180 16788
rect 57060 16736 57112 16788
rect 1584 16711 1636 16720
rect 1584 16677 1593 16711
rect 1593 16677 1627 16711
rect 1627 16677 1636 16711
rect 1584 16668 1636 16677
rect 24308 16668 24360 16720
rect 47032 16668 47084 16720
rect 54944 16711 54996 16720
rect 20352 16643 20404 16652
rect 20352 16609 20361 16643
rect 20361 16609 20395 16643
rect 20395 16609 20404 16643
rect 20352 16600 20404 16609
rect 31852 16600 31904 16652
rect 40132 16600 40184 16652
rect 42340 16643 42392 16652
rect 42340 16609 42349 16643
rect 42349 16609 42383 16643
rect 42383 16609 42392 16643
rect 42340 16600 42392 16609
rect 42432 16600 42484 16652
rect 45836 16600 45888 16652
rect 46388 16600 46440 16652
rect 46572 16600 46624 16652
rect 54944 16677 54953 16711
rect 54953 16677 54987 16711
rect 54987 16677 54996 16711
rect 54944 16668 54996 16677
rect 62028 16736 62080 16788
rect 65892 16736 65944 16788
rect 61108 16668 61160 16720
rect 68192 16668 68244 16720
rect 20628 16532 20680 16584
rect 35992 16532 36044 16584
rect 29368 16464 29420 16516
rect 53564 16600 53616 16652
rect 55956 16600 56008 16652
rect 56784 16643 56836 16652
rect 56784 16609 56793 16643
rect 56793 16609 56827 16643
rect 56827 16609 56836 16643
rect 56784 16600 56836 16609
rect 57336 16643 57388 16652
rect 57336 16609 57345 16643
rect 57345 16609 57379 16643
rect 57379 16609 57388 16643
rect 57336 16600 57388 16609
rect 59452 16600 59504 16652
rect 59912 16575 59964 16584
rect 40776 16464 40828 16516
rect 47124 16464 47176 16516
rect 19616 16439 19668 16448
rect 19616 16405 19625 16439
rect 19625 16405 19659 16439
rect 19659 16405 19668 16439
rect 19616 16396 19668 16405
rect 32220 16439 32272 16448
rect 32220 16405 32229 16439
rect 32229 16405 32263 16439
rect 32263 16405 32272 16439
rect 32220 16396 32272 16405
rect 32864 16439 32916 16448
rect 32864 16405 32873 16439
rect 32873 16405 32907 16439
rect 32907 16405 32916 16439
rect 32864 16396 32916 16405
rect 39580 16396 39632 16448
rect 43720 16396 43772 16448
rect 44824 16396 44876 16448
rect 47400 16464 47452 16516
rect 51816 16464 51868 16516
rect 48872 16396 48924 16448
rect 51172 16396 51224 16448
rect 54852 16464 54904 16516
rect 59912 16541 59921 16575
rect 59921 16541 59955 16575
rect 59955 16541 59964 16575
rect 59912 16532 59964 16541
rect 65524 16600 65576 16652
rect 83372 16668 83424 16720
rect 83740 16736 83792 16788
rect 94228 16779 94280 16788
rect 94228 16745 94237 16779
rect 94237 16745 94271 16779
rect 94271 16745 94280 16779
rect 94228 16736 94280 16745
rect 87880 16668 87932 16720
rect 77300 16600 77352 16652
rect 60832 16532 60884 16584
rect 62856 16575 62908 16584
rect 62856 16541 62865 16575
rect 62865 16541 62899 16575
rect 62899 16541 62908 16575
rect 62856 16532 62908 16541
rect 67548 16575 67600 16584
rect 67548 16541 67557 16575
rect 67557 16541 67591 16575
rect 67591 16541 67600 16575
rect 67548 16532 67600 16541
rect 83556 16532 83608 16584
rect 92572 16575 92624 16584
rect 92572 16541 92581 16575
rect 92581 16541 92615 16575
rect 92615 16541 92624 16575
rect 92572 16532 92624 16541
rect 61844 16464 61896 16516
rect 52368 16396 52420 16448
rect 55220 16396 55272 16448
rect 58164 16439 58216 16448
rect 58164 16405 58173 16439
rect 58173 16405 58207 16439
rect 58207 16405 58216 16439
rect 58164 16396 58216 16405
rect 59176 16439 59228 16448
rect 59176 16405 59185 16439
rect 59185 16405 59219 16439
rect 59219 16405 59228 16439
rect 59176 16396 59228 16405
rect 60004 16439 60056 16448
rect 60004 16405 60013 16439
rect 60013 16405 60047 16439
rect 60047 16405 60056 16439
rect 60004 16396 60056 16405
rect 60096 16396 60148 16448
rect 61936 16396 61988 16448
rect 62028 16396 62080 16448
rect 63592 16464 63644 16516
rect 65800 16464 65852 16516
rect 64604 16439 64656 16448
rect 64604 16405 64613 16439
rect 64613 16405 64647 16439
rect 64647 16405 64656 16439
rect 64604 16396 64656 16405
rect 64972 16396 65024 16448
rect 68744 16464 68796 16516
rect 71964 16439 72016 16448
rect 71964 16405 71973 16439
rect 71973 16405 72007 16439
rect 72007 16405 72016 16439
rect 71964 16396 72016 16405
rect 24386 16294 24438 16346
rect 24450 16294 24502 16346
rect 24514 16294 24566 16346
rect 24578 16294 24630 16346
rect 24642 16294 24694 16346
rect 47823 16294 47875 16346
rect 47887 16294 47939 16346
rect 47951 16294 48003 16346
rect 48015 16294 48067 16346
rect 48079 16294 48131 16346
rect 71260 16294 71312 16346
rect 71324 16294 71376 16346
rect 71388 16294 71440 16346
rect 71452 16294 71504 16346
rect 71516 16294 71568 16346
rect 94697 16294 94749 16346
rect 94761 16294 94813 16346
rect 94825 16294 94877 16346
rect 94889 16294 94941 16346
rect 94953 16294 95005 16346
rect 19616 16124 19668 16176
rect 20628 16056 20680 16108
rect 15384 15988 15436 16040
rect 20352 15988 20404 16040
rect 32864 16192 32916 16244
rect 39580 16192 39632 16244
rect 31392 16124 31444 16176
rect 29552 16056 29604 16108
rect 30104 16056 30156 16108
rect 39764 16124 39816 16176
rect 40776 16124 40828 16176
rect 41604 16192 41656 16244
rect 44824 16192 44876 16244
rect 46388 16192 46440 16244
rect 52092 16192 52144 16244
rect 52276 16192 52328 16244
rect 46480 16124 46532 16176
rect 40868 16099 40920 16108
rect 40868 16065 40877 16099
rect 40877 16065 40911 16099
rect 40911 16065 40920 16099
rect 40868 16056 40920 16065
rect 40316 15988 40368 16040
rect 40776 16031 40828 16040
rect 40776 15997 40785 16031
rect 40785 15997 40819 16031
rect 40819 15997 40828 16031
rect 40776 15988 40828 15997
rect 40960 15988 41012 16040
rect 22100 15920 22152 15972
rect 20720 15895 20772 15904
rect 20720 15861 20729 15895
rect 20729 15861 20763 15895
rect 20763 15861 20772 15895
rect 20720 15852 20772 15861
rect 27712 15852 27764 15904
rect 29552 15895 29604 15904
rect 29552 15861 29561 15895
rect 29561 15861 29595 15895
rect 29595 15861 29604 15895
rect 29552 15852 29604 15861
rect 29736 15920 29788 15972
rect 32864 15920 32916 15972
rect 34796 15963 34848 15972
rect 34796 15929 34805 15963
rect 34805 15929 34839 15963
rect 34839 15929 34848 15963
rect 34796 15920 34848 15929
rect 41880 15920 41932 15972
rect 32772 15852 32824 15904
rect 34060 15852 34112 15904
rect 34520 15852 34572 15904
rect 35808 15852 35860 15904
rect 38844 15852 38896 15904
rect 42800 16056 42852 16108
rect 44272 16056 44324 16108
rect 46020 16099 46072 16108
rect 46020 16065 46029 16099
rect 46029 16065 46063 16099
rect 46063 16065 46072 16099
rect 46020 16056 46072 16065
rect 44364 15988 44416 16040
rect 51448 16124 51500 16176
rect 53564 16167 53616 16176
rect 47032 16056 47084 16108
rect 49056 16056 49108 16108
rect 50344 16099 50396 16108
rect 50344 16065 50353 16099
rect 50353 16065 50387 16099
rect 50387 16065 50396 16099
rect 50344 16056 50396 16065
rect 50436 16056 50488 16108
rect 53564 16133 53573 16167
rect 53573 16133 53607 16167
rect 53607 16133 53616 16167
rect 53564 16124 53616 16133
rect 55864 16124 55916 16176
rect 59176 16124 59228 16176
rect 59360 16124 59412 16176
rect 60004 16124 60056 16176
rect 61936 16192 61988 16244
rect 71964 16192 72016 16244
rect 72148 16192 72200 16244
rect 77852 16192 77904 16244
rect 92572 16192 92624 16244
rect 64972 16124 65024 16176
rect 65524 16167 65576 16176
rect 65524 16133 65533 16167
rect 65533 16133 65567 16167
rect 65567 16133 65576 16167
rect 65524 16124 65576 16133
rect 66076 16124 66128 16176
rect 52368 16099 52420 16108
rect 52368 16065 52377 16099
rect 52377 16065 52411 16099
rect 52411 16065 52420 16099
rect 52368 16056 52420 16065
rect 53656 16056 53708 16108
rect 54208 16099 54260 16108
rect 54208 16065 54217 16099
rect 54217 16065 54251 16099
rect 54251 16065 54260 16099
rect 56416 16099 56468 16108
rect 54208 16056 54260 16065
rect 48688 15988 48740 16040
rect 50528 16031 50580 16040
rect 50528 15997 50537 16031
rect 50537 15997 50571 16031
rect 50571 15997 50580 16031
rect 50528 15988 50580 15997
rect 56416 16065 56425 16099
rect 56425 16065 56459 16099
rect 56459 16065 56468 16099
rect 56416 16056 56468 16065
rect 56692 16056 56744 16108
rect 60096 16056 60148 16108
rect 63592 16056 63644 16108
rect 66168 16056 66220 16108
rect 46020 15920 46072 15972
rect 46204 15920 46256 15972
rect 42892 15852 42944 15904
rect 43812 15852 43864 15904
rect 44272 15895 44324 15904
rect 44272 15861 44281 15895
rect 44281 15861 44315 15895
rect 44315 15861 44324 15895
rect 44272 15852 44324 15861
rect 45468 15895 45520 15904
rect 45468 15861 45477 15895
rect 45477 15861 45511 15895
rect 45511 15861 45520 15895
rect 45468 15852 45520 15861
rect 47032 15852 47084 15904
rect 47124 15852 47176 15904
rect 48780 15895 48832 15904
rect 48780 15861 48789 15895
rect 48789 15861 48823 15895
rect 48823 15861 48832 15895
rect 48780 15852 48832 15861
rect 48872 15852 48924 15904
rect 55312 15920 55364 15972
rect 56324 15988 56376 16040
rect 60740 15988 60792 16040
rect 61844 15988 61896 16040
rect 66352 15988 66404 16040
rect 64604 15920 64656 15972
rect 66536 15988 66588 16040
rect 72056 16124 72108 16176
rect 71136 16099 71188 16108
rect 71136 16065 71145 16099
rect 71145 16065 71179 16099
rect 71179 16065 71188 16099
rect 71136 16056 71188 16065
rect 78864 16099 78916 16108
rect 78864 16065 78873 16099
rect 78873 16065 78907 16099
rect 78907 16065 78916 16099
rect 78864 16056 78916 16065
rect 77208 15988 77260 16040
rect 53012 15895 53064 15904
rect 53012 15861 53021 15895
rect 53021 15861 53055 15895
rect 53055 15861 53064 15895
rect 53012 15852 53064 15861
rect 55956 15852 56008 15904
rect 56600 15852 56652 15904
rect 57888 15852 57940 15904
rect 58624 15895 58676 15904
rect 58624 15861 58633 15895
rect 58633 15861 58667 15895
rect 58667 15861 58676 15895
rect 58624 15852 58676 15861
rect 58716 15852 58768 15904
rect 62212 15895 62264 15904
rect 62212 15861 62221 15895
rect 62221 15861 62255 15895
rect 62255 15861 62264 15895
rect 62212 15852 62264 15861
rect 62948 15852 63000 15904
rect 65892 15852 65944 15904
rect 66076 15852 66128 15904
rect 76748 15920 76800 15972
rect 77116 15920 77168 15972
rect 80704 15920 80756 15972
rect 67916 15852 67968 15904
rect 68008 15852 68060 15904
rect 69020 15895 69072 15904
rect 69020 15861 69029 15895
rect 69029 15861 69063 15895
rect 69063 15861 69072 15895
rect 69020 15852 69072 15861
rect 69756 15852 69808 15904
rect 71044 15895 71096 15904
rect 71044 15861 71053 15895
rect 71053 15861 71087 15895
rect 71087 15861 71096 15895
rect 71044 15852 71096 15861
rect 74264 15852 74316 15904
rect 76564 15852 76616 15904
rect 77484 15852 77536 15904
rect 78772 15895 78824 15904
rect 78772 15861 78781 15895
rect 78781 15861 78815 15895
rect 78815 15861 78824 15895
rect 78772 15852 78824 15861
rect 80612 15852 80664 15904
rect 83464 15852 83516 15904
rect 83924 15895 83976 15904
rect 83924 15861 83933 15895
rect 83933 15861 83967 15895
rect 83967 15861 83976 15895
rect 83924 15852 83976 15861
rect 12668 15750 12720 15802
rect 12732 15750 12784 15802
rect 12796 15750 12848 15802
rect 12860 15750 12912 15802
rect 12924 15750 12976 15802
rect 36105 15750 36157 15802
rect 36169 15750 36221 15802
rect 36233 15750 36285 15802
rect 36297 15750 36349 15802
rect 36361 15750 36413 15802
rect 59542 15750 59594 15802
rect 59606 15750 59658 15802
rect 59670 15750 59722 15802
rect 59734 15750 59786 15802
rect 59798 15750 59850 15802
rect 82979 15750 83031 15802
rect 83043 15750 83095 15802
rect 83107 15750 83159 15802
rect 83171 15750 83223 15802
rect 83235 15750 83287 15802
rect 28080 15648 28132 15700
rect 30104 15691 30156 15700
rect 30104 15657 30113 15691
rect 30113 15657 30147 15691
rect 30147 15657 30156 15691
rect 30104 15648 30156 15657
rect 31392 15648 31444 15700
rect 27804 15580 27856 15632
rect 34980 15648 35032 15700
rect 39764 15648 39816 15700
rect 44364 15648 44416 15700
rect 45468 15648 45520 15700
rect 60832 15648 60884 15700
rect 65984 15648 66036 15700
rect 73252 15648 73304 15700
rect 19616 15512 19668 15564
rect 44272 15580 44324 15632
rect 47952 15580 48004 15632
rect 50436 15580 50488 15632
rect 60280 15580 60332 15632
rect 19340 15444 19392 15496
rect 20628 15444 20680 15496
rect 22652 15487 22704 15496
rect 22652 15453 22661 15487
rect 22661 15453 22695 15487
rect 22695 15453 22704 15487
rect 22652 15444 22704 15453
rect 27620 15444 27672 15496
rect 30472 15444 30524 15496
rect 32220 15444 32272 15496
rect 32864 15444 32916 15496
rect 34796 15444 34848 15496
rect 38752 15512 38804 15564
rect 39304 15512 39356 15564
rect 46204 15512 46256 15564
rect 46480 15512 46532 15564
rect 37096 15444 37148 15496
rect 40316 15487 40368 15496
rect 40316 15453 40325 15487
rect 40325 15453 40359 15487
rect 40359 15453 40368 15487
rect 40316 15444 40368 15453
rect 40776 15487 40828 15496
rect 40776 15453 40785 15487
rect 40785 15453 40819 15487
rect 40819 15453 40828 15487
rect 40776 15444 40828 15453
rect 40868 15444 40920 15496
rect 43720 15487 43772 15496
rect 43720 15453 43729 15487
rect 43729 15453 43763 15487
rect 43763 15453 43772 15487
rect 43720 15444 43772 15453
rect 45744 15487 45796 15496
rect 45744 15453 45753 15487
rect 45753 15453 45787 15487
rect 45787 15453 45796 15487
rect 45744 15444 45796 15453
rect 46664 15487 46716 15496
rect 46664 15453 46673 15487
rect 46673 15453 46707 15487
rect 46707 15453 46716 15487
rect 46664 15444 46716 15453
rect 61108 15555 61160 15564
rect 48688 15444 48740 15496
rect 49148 15444 49200 15496
rect 49516 15487 49568 15496
rect 49516 15453 49525 15487
rect 49525 15453 49559 15487
rect 49559 15453 49568 15487
rect 49516 15444 49568 15453
rect 51172 15487 51224 15496
rect 51172 15453 51181 15487
rect 51181 15453 51215 15487
rect 51215 15453 51224 15487
rect 51172 15444 51224 15453
rect 53656 15444 53708 15496
rect 56416 15444 56468 15496
rect 57060 15487 57112 15496
rect 57060 15453 57069 15487
rect 57069 15453 57103 15487
rect 57103 15453 57112 15487
rect 57060 15444 57112 15453
rect 59912 15444 59964 15496
rect 61108 15521 61117 15555
rect 61117 15521 61151 15555
rect 61151 15521 61160 15555
rect 61108 15512 61160 15521
rect 64696 15555 64748 15564
rect 64696 15521 64705 15555
rect 64705 15521 64739 15555
rect 64739 15521 64748 15555
rect 64696 15512 64748 15521
rect 67364 15580 67416 15632
rect 70492 15580 70544 15632
rect 72424 15580 72476 15632
rect 61016 15444 61068 15496
rect 65892 15444 65944 15496
rect 65984 15487 66036 15496
rect 65984 15453 65993 15487
rect 65993 15453 66027 15487
rect 66027 15453 66036 15487
rect 67640 15512 67692 15564
rect 70308 15512 70360 15564
rect 71136 15512 71188 15564
rect 65984 15444 66036 15453
rect 67916 15487 67968 15496
rect 20076 15351 20128 15360
rect 20076 15317 20085 15351
rect 20085 15317 20119 15351
rect 20119 15317 20128 15351
rect 20076 15308 20128 15317
rect 20812 15308 20864 15360
rect 22744 15351 22796 15360
rect 22744 15317 22753 15351
rect 22753 15317 22787 15351
rect 22787 15317 22796 15351
rect 22744 15308 22796 15317
rect 23664 15351 23716 15360
rect 23664 15317 23673 15351
rect 23673 15317 23707 15351
rect 23707 15317 23716 15351
rect 23664 15308 23716 15317
rect 24768 15308 24820 15360
rect 32404 15376 32456 15428
rect 32588 15376 32640 15428
rect 32772 15376 32824 15428
rect 41604 15376 41656 15428
rect 41880 15376 41932 15428
rect 28540 15308 28592 15360
rect 28908 15308 28960 15360
rect 32680 15308 32732 15360
rect 33140 15308 33192 15360
rect 34520 15308 34572 15360
rect 34980 15308 35032 15360
rect 35532 15351 35584 15360
rect 35532 15317 35541 15351
rect 35541 15317 35575 15351
rect 35575 15317 35584 15351
rect 35532 15308 35584 15317
rect 36268 15351 36320 15360
rect 36268 15317 36277 15351
rect 36277 15317 36311 15351
rect 36311 15317 36320 15351
rect 36268 15308 36320 15317
rect 37740 15308 37792 15360
rect 38108 15308 38160 15360
rect 40868 15308 40920 15360
rect 41144 15351 41196 15360
rect 41144 15317 41153 15351
rect 41153 15317 41187 15351
rect 41187 15317 41196 15351
rect 41144 15308 41196 15317
rect 41696 15308 41748 15360
rect 42340 15351 42392 15360
rect 42340 15317 42349 15351
rect 42349 15317 42383 15351
rect 42383 15317 42392 15351
rect 42340 15308 42392 15317
rect 43076 15376 43128 15428
rect 46940 15419 46992 15428
rect 45652 15351 45704 15360
rect 45652 15317 45661 15351
rect 45661 15317 45695 15351
rect 45695 15317 45704 15351
rect 45652 15308 45704 15317
rect 46940 15385 46949 15419
rect 46949 15385 46983 15419
rect 46983 15385 46992 15419
rect 46940 15376 46992 15385
rect 51448 15419 51500 15428
rect 48504 15308 48556 15360
rect 49700 15308 49752 15360
rect 50528 15308 50580 15360
rect 51448 15385 51457 15419
rect 51457 15385 51491 15419
rect 51491 15385 51500 15419
rect 51448 15376 51500 15385
rect 53012 15376 53064 15428
rect 56692 15376 56744 15428
rect 57980 15376 58032 15428
rect 53748 15351 53800 15360
rect 53748 15317 53757 15351
rect 53757 15317 53791 15351
rect 53791 15317 53800 15351
rect 53748 15308 53800 15317
rect 54484 15308 54536 15360
rect 54852 15351 54904 15360
rect 54852 15317 54861 15351
rect 54861 15317 54895 15351
rect 54895 15317 54904 15351
rect 54852 15308 54904 15317
rect 56048 15351 56100 15360
rect 56048 15317 56057 15351
rect 56057 15317 56091 15351
rect 56091 15317 56100 15351
rect 56048 15308 56100 15317
rect 61936 15376 61988 15428
rect 60096 15308 60148 15360
rect 63592 15308 63644 15360
rect 64972 15376 65024 15428
rect 67916 15453 67925 15487
rect 67925 15453 67959 15487
rect 67959 15453 67968 15487
rect 67916 15444 67968 15453
rect 70860 15444 70912 15496
rect 72056 15512 72108 15564
rect 72608 15580 72660 15632
rect 74632 15580 74684 15632
rect 72148 15487 72200 15496
rect 72148 15453 72157 15487
rect 72157 15453 72191 15487
rect 72191 15453 72200 15487
rect 80244 15512 80296 15564
rect 74172 15487 74224 15496
rect 72148 15444 72200 15453
rect 67824 15376 67876 15428
rect 74172 15453 74181 15487
rect 74181 15453 74215 15487
rect 74215 15453 74224 15487
rect 74172 15444 74224 15453
rect 81256 15444 81308 15496
rect 82820 15444 82872 15496
rect 66536 15308 66588 15360
rect 66720 15351 66772 15360
rect 66720 15317 66729 15351
rect 66729 15317 66763 15351
rect 66763 15317 66772 15351
rect 66720 15308 66772 15317
rect 68744 15308 68796 15360
rect 69848 15308 69900 15360
rect 70860 15308 70912 15360
rect 71596 15351 71648 15360
rect 71596 15317 71605 15351
rect 71605 15317 71639 15351
rect 71639 15317 71648 15351
rect 71596 15308 71648 15317
rect 76472 15351 76524 15360
rect 76472 15317 76481 15351
rect 76481 15317 76515 15351
rect 76515 15317 76524 15351
rect 76472 15308 76524 15317
rect 77392 15351 77444 15360
rect 77392 15317 77401 15351
rect 77401 15317 77435 15351
rect 77435 15317 77444 15351
rect 77392 15308 77444 15317
rect 78772 15376 78824 15428
rect 83004 15376 83056 15428
rect 80152 15351 80204 15360
rect 80152 15317 80161 15351
rect 80161 15317 80195 15351
rect 80195 15317 80204 15351
rect 80152 15308 80204 15317
rect 81624 15308 81676 15360
rect 83740 15351 83792 15360
rect 83740 15317 83749 15351
rect 83749 15317 83783 15351
rect 83783 15317 83792 15351
rect 83740 15308 83792 15317
rect 84108 15308 84160 15360
rect 86776 15308 86828 15360
rect 88248 15308 88300 15360
rect 88984 15308 89036 15360
rect 24386 15206 24438 15258
rect 24450 15206 24502 15258
rect 24514 15206 24566 15258
rect 24578 15206 24630 15258
rect 24642 15206 24694 15258
rect 47823 15206 47875 15258
rect 47887 15206 47939 15258
rect 47951 15206 48003 15258
rect 48015 15206 48067 15258
rect 48079 15206 48131 15258
rect 71260 15206 71312 15258
rect 71324 15206 71376 15258
rect 71388 15206 71440 15258
rect 71452 15206 71504 15258
rect 71516 15206 71568 15258
rect 94697 15206 94749 15258
rect 94761 15206 94813 15258
rect 94825 15206 94877 15258
rect 94889 15206 94941 15258
rect 94953 15206 95005 15258
rect 16304 15104 16356 15156
rect 22560 15104 22612 15156
rect 19616 15036 19668 15088
rect 20720 15036 20772 15088
rect 28080 15104 28132 15156
rect 24768 15036 24820 15088
rect 24860 15036 24912 15088
rect 27804 15036 27856 15088
rect 28908 15036 28960 15088
rect 33324 15104 33376 15156
rect 38752 15104 38804 15156
rect 15752 14900 15804 14952
rect 24584 14968 24636 15020
rect 23664 14900 23716 14952
rect 25872 14943 25924 14952
rect 25872 14909 25881 14943
rect 25881 14909 25915 14943
rect 25915 14909 25924 14943
rect 25872 14900 25924 14909
rect 30104 14968 30156 15020
rect 29644 14900 29696 14952
rect 29920 14943 29972 14952
rect 29920 14909 29929 14943
rect 29929 14909 29963 14943
rect 29963 14909 29972 14943
rect 29920 14900 29972 14909
rect 30748 14900 30800 14952
rect 35992 15036 36044 15088
rect 31392 15011 31444 15020
rect 31392 14977 31401 15011
rect 31401 14977 31435 15011
rect 31435 14977 31444 15011
rect 31392 14968 31444 14977
rect 31484 14968 31536 15020
rect 32956 14968 33008 15020
rect 34796 14968 34848 15020
rect 34980 15011 35032 15020
rect 34980 14977 34989 15011
rect 34989 14977 35023 15011
rect 35023 14977 35032 15011
rect 34980 14968 35032 14977
rect 36268 15036 36320 15088
rect 37280 14968 37332 15020
rect 32772 14900 32824 14952
rect 33232 14900 33284 14952
rect 34704 14900 34756 14952
rect 35072 14900 35124 14952
rect 38660 14968 38712 15020
rect 39304 15011 39356 15020
rect 39304 14977 39313 15011
rect 39313 14977 39347 15011
rect 39347 14977 39356 15011
rect 40316 15011 40368 15020
rect 39304 14968 39356 14977
rect 40316 14977 40325 15011
rect 40325 14977 40359 15011
rect 40359 14977 40368 15011
rect 40316 14968 40368 14977
rect 40408 14968 40460 15020
rect 43444 15011 43496 15020
rect 12532 14832 12584 14884
rect 12716 14875 12768 14884
rect 12716 14841 12725 14875
rect 12725 14841 12759 14875
rect 12759 14841 12768 14875
rect 12716 14832 12768 14841
rect 15016 14764 15068 14816
rect 16120 14764 16172 14816
rect 24400 14832 24452 14884
rect 27712 14832 27764 14884
rect 22376 14764 22428 14816
rect 24492 14764 24544 14816
rect 26792 14764 26844 14816
rect 26884 14764 26936 14816
rect 32036 14832 32088 14884
rect 41328 14900 41380 14952
rect 43444 14977 43453 15011
rect 43453 14977 43487 15011
rect 43487 14977 43496 15011
rect 43444 14968 43496 14977
rect 46020 15036 46072 15088
rect 48688 15036 48740 15088
rect 48780 15036 48832 15088
rect 49700 15036 49752 15088
rect 50712 15036 50764 15088
rect 53104 15036 53156 15088
rect 47124 14968 47176 15020
rect 47216 14968 47268 15020
rect 49148 15011 49200 15020
rect 49148 14977 49157 15011
rect 49157 14977 49191 15011
rect 49191 14977 49200 15011
rect 49148 14968 49200 14977
rect 53748 15036 53800 15088
rect 54944 15036 54996 15088
rect 55496 15036 55548 15088
rect 59084 15079 59136 15088
rect 59084 15045 59093 15079
rect 59093 15045 59127 15079
rect 59127 15045 59136 15079
rect 59084 15036 59136 15045
rect 42708 14900 42760 14952
rect 46020 14900 46072 14952
rect 46296 14900 46348 14952
rect 48320 14943 48372 14952
rect 48320 14909 48329 14943
rect 48329 14909 48363 14943
rect 48363 14909 48372 14943
rect 48320 14900 48372 14909
rect 56600 14968 56652 15020
rect 33048 14764 33100 14816
rect 35992 14807 36044 14816
rect 35992 14773 36001 14807
rect 36001 14773 36035 14807
rect 36035 14773 36044 14807
rect 35992 14764 36044 14773
rect 36084 14764 36136 14816
rect 41236 14832 41288 14884
rect 52092 14900 52144 14952
rect 55220 14943 55272 14952
rect 55220 14909 55229 14943
rect 55229 14909 55263 14943
rect 55263 14909 55272 14943
rect 55220 14900 55272 14909
rect 40224 14807 40276 14816
rect 40224 14773 40233 14807
rect 40233 14773 40267 14807
rect 40267 14773 40276 14807
rect 40224 14764 40276 14773
rect 41604 14807 41656 14816
rect 41604 14773 41613 14807
rect 41613 14773 41647 14807
rect 41647 14773 41656 14807
rect 41604 14764 41656 14773
rect 42708 14764 42760 14816
rect 44732 14807 44784 14816
rect 44732 14773 44741 14807
rect 44741 14773 44775 14807
rect 44775 14773 44784 14807
rect 44732 14764 44784 14773
rect 50896 14807 50948 14816
rect 50896 14773 50905 14807
rect 50905 14773 50939 14807
rect 50939 14773 50948 14807
rect 50896 14764 50948 14773
rect 51724 14764 51776 14816
rect 52000 14807 52052 14816
rect 52000 14773 52009 14807
rect 52009 14773 52043 14807
rect 52043 14773 52052 14807
rect 52000 14764 52052 14773
rect 55588 14900 55640 14952
rect 56692 14900 56744 14952
rect 56968 14943 57020 14952
rect 56968 14909 56977 14943
rect 56977 14909 57011 14943
rect 57011 14909 57020 14943
rect 56968 14900 57020 14909
rect 59912 15104 59964 15156
rect 61568 15104 61620 15156
rect 62304 15147 62356 15156
rect 62304 15113 62313 15147
rect 62313 15113 62347 15147
rect 62347 15113 62356 15147
rect 62304 15104 62356 15113
rect 66168 15104 66220 15156
rect 68376 15104 68428 15156
rect 60096 15036 60148 15088
rect 60832 15079 60884 15088
rect 60832 15045 60841 15079
rect 60841 15045 60875 15079
rect 60875 15045 60884 15079
rect 60832 15036 60884 15045
rect 61476 15036 61528 15088
rect 61292 14968 61344 15020
rect 61568 15011 61620 15020
rect 61568 14977 61577 15011
rect 61577 14977 61611 15011
rect 61611 14977 61620 15011
rect 61936 15036 61988 15088
rect 61568 14968 61620 14977
rect 63132 14968 63184 15020
rect 65432 15036 65484 15088
rect 66720 15036 66772 15088
rect 67180 15011 67232 15020
rect 67180 14977 67189 15011
rect 67189 14977 67223 15011
rect 67223 14977 67232 15011
rect 67180 14968 67232 14977
rect 70952 15104 71004 15156
rect 74172 15104 74224 15156
rect 74540 15104 74592 15156
rect 80612 15104 80664 15156
rect 82176 15147 82228 15156
rect 82176 15113 82185 15147
rect 82185 15113 82219 15147
rect 82219 15113 82228 15147
rect 82176 15104 82228 15113
rect 71044 15036 71096 15088
rect 76472 15036 76524 15088
rect 77300 15079 77352 15088
rect 77300 15045 77309 15079
rect 77309 15045 77343 15079
rect 77343 15045 77352 15079
rect 77852 15079 77904 15088
rect 77300 15036 77352 15045
rect 77852 15045 77861 15079
rect 77861 15045 77895 15079
rect 77895 15045 77904 15079
rect 77852 15036 77904 15045
rect 78680 15036 78732 15088
rect 80152 15036 80204 15088
rect 69020 14968 69072 15020
rect 64880 14943 64932 14952
rect 55496 14764 55548 14816
rect 58808 14764 58860 14816
rect 59452 14764 59504 14816
rect 62304 14832 62356 14884
rect 61660 14807 61712 14816
rect 61660 14773 61669 14807
rect 61669 14773 61703 14807
rect 61703 14773 61712 14807
rect 61660 14764 61712 14773
rect 64236 14764 64288 14816
rect 64880 14909 64889 14943
rect 64889 14909 64923 14943
rect 64923 14909 64932 14943
rect 64880 14900 64932 14909
rect 65892 14900 65944 14952
rect 66444 14900 66496 14952
rect 71504 14968 71556 15020
rect 72056 14968 72108 15020
rect 74264 14968 74316 15020
rect 75828 15011 75880 15020
rect 75828 14977 75837 15011
rect 75837 14977 75871 15011
rect 75871 14977 75880 15011
rect 75828 14968 75880 14977
rect 78864 15011 78916 15020
rect 78864 14977 78873 15011
rect 78873 14977 78907 15011
rect 78907 14977 78916 15011
rect 78864 14968 78916 14977
rect 79600 14968 79652 15020
rect 80612 15011 80664 15020
rect 80612 14977 80621 15011
rect 80621 14977 80655 15011
rect 80655 14977 80664 15011
rect 80612 14968 80664 14977
rect 82544 15011 82596 15020
rect 82544 14977 82553 15011
rect 82553 14977 82587 15011
rect 82587 14977 82596 15011
rect 82544 14968 82596 14977
rect 84936 15104 84988 15156
rect 83924 15036 83976 15088
rect 86500 14968 86552 15020
rect 69756 14943 69808 14952
rect 69756 14909 69765 14943
rect 69765 14909 69799 14943
rect 69799 14909 69808 14943
rect 69756 14900 69808 14909
rect 71044 14900 71096 14952
rect 73252 14900 73304 14952
rect 80704 14943 80756 14952
rect 67732 14764 67784 14816
rect 68468 14807 68520 14816
rect 68468 14773 68477 14807
rect 68477 14773 68511 14807
rect 68511 14773 68520 14807
rect 68468 14764 68520 14773
rect 72148 14832 72200 14884
rect 75276 14875 75328 14884
rect 75276 14841 75285 14875
rect 75285 14841 75319 14875
rect 75319 14841 75328 14875
rect 75276 14832 75328 14841
rect 80704 14909 80713 14943
rect 80713 14909 80747 14943
rect 80747 14909 80756 14943
rect 80704 14900 80756 14909
rect 82820 14900 82872 14952
rect 83004 14900 83056 14952
rect 85028 14900 85080 14952
rect 86776 14900 86828 14952
rect 92664 14832 92716 14884
rect 74540 14764 74592 14816
rect 74632 14764 74684 14816
rect 75920 14764 75972 14816
rect 78220 14764 78272 14816
rect 79324 14807 79376 14816
rect 79324 14773 79333 14807
rect 79333 14773 79367 14807
rect 79367 14773 79376 14807
rect 79324 14764 79376 14773
rect 80336 14807 80388 14816
rect 80336 14773 80345 14807
rect 80345 14773 80379 14807
rect 80379 14773 80388 14807
rect 80336 14764 80388 14773
rect 81716 14764 81768 14816
rect 85212 14807 85264 14816
rect 85212 14773 85221 14807
rect 85221 14773 85255 14807
rect 85255 14773 85264 14807
rect 85212 14764 85264 14773
rect 86776 14764 86828 14816
rect 86960 14764 87012 14816
rect 89076 14807 89128 14816
rect 89076 14773 89085 14807
rect 89085 14773 89119 14807
rect 89119 14773 89128 14807
rect 89076 14764 89128 14773
rect 90456 14764 90508 14816
rect 12668 14662 12720 14714
rect 12732 14662 12784 14714
rect 12796 14662 12848 14714
rect 12860 14662 12912 14714
rect 12924 14662 12976 14714
rect 36105 14662 36157 14714
rect 36169 14662 36221 14714
rect 36233 14662 36285 14714
rect 36297 14662 36349 14714
rect 36361 14662 36413 14714
rect 59542 14662 59594 14714
rect 59606 14662 59658 14714
rect 59670 14662 59722 14714
rect 59734 14662 59786 14714
rect 59798 14662 59850 14714
rect 82979 14662 83031 14714
rect 83043 14662 83095 14714
rect 83107 14662 83159 14714
rect 83171 14662 83223 14714
rect 83235 14662 83287 14714
rect 8024 14492 8076 14544
rect 7288 14399 7340 14408
rect 7288 14365 7297 14399
rect 7297 14365 7331 14399
rect 7331 14365 7340 14399
rect 7288 14356 7340 14365
rect 8024 14399 8076 14408
rect 8024 14365 8033 14399
rect 8033 14365 8067 14399
rect 8067 14365 8076 14399
rect 8024 14356 8076 14365
rect 9128 14288 9180 14340
rect 15384 14492 15436 14544
rect 11336 14467 11388 14476
rect 11336 14433 11345 14467
rect 11345 14433 11379 14467
rect 11379 14433 11388 14467
rect 11336 14424 11388 14433
rect 14556 14424 14608 14476
rect 15200 14424 15252 14476
rect 24400 14560 24452 14612
rect 24584 14603 24636 14612
rect 24584 14569 24593 14603
rect 24593 14569 24627 14603
rect 24627 14569 24636 14603
rect 24584 14560 24636 14569
rect 25044 14560 25096 14612
rect 28724 14560 28776 14612
rect 23756 14492 23808 14544
rect 27160 14492 27212 14544
rect 35992 14560 36044 14612
rect 26884 14424 26936 14476
rect 28816 14424 28868 14476
rect 30656 14424 30708 14476
rect 11428 14399 11480 14408
rect 11428 14365 11437 14399
rect 11437 14365 11471 14399
rect 11471 14365 11480 14399
rect 11428 14356 11480 14365
rect 12532 14399 12584 14408
rect 12532 14365 12541 14399
rect 12541 14365 12575 14399
rect 12575 14365 12584 14399
rect 12532 14356 12584 14365
rect 15108 14356 15160 14408
rect 20812 14356 20864 14408
rect 24492 14356 24544 14408
rect 24768 14399 24820 14408
rect 24768 14365 24777 14399
rect 24777 14365 24811 14399
rect 24811 14365 24820 14399
rect 24768 14356 24820 14365
rect 12440 14288 12492 14340
rect 13084 14331 13136 14340
rect 13084 14297 13093 14331
rect 13093 14297 13127 14331
rect 13127 14297 13136 14331
rect 13084 14288 13136 14297
rect 22744 14288 22796 14340
rect 24860 14288 24912 14340
rect 14004 14220 14056 14272
rect 15568 14263 15620 14272
rect 15568 14229 15577 14263
rect 15577 14229 15611 14263
rect 15611 14229 15620 14263
rect 15568 14220 15620 14229
rect 16212 14263 16264 14272
rect 16212 14229 16221 14263
rect 16221 14229 16255 14263
rect 16255 14229 16264 14263
rect 16212 14220 16264 14229
rect 20628 14220 20680 14272
rect 25596 14356 25648 14408
rect 27160 14399 27212 14408
rect 25596 14263 25648 14272
rect 25596 14229 25605 14263
rect 25605 14229 25639 14263
rect 25639 14229 25648 14263
rect 25596 14220 25648 14229
rect 26240 14220 26292 14272
rect 27160 14365 27169 14399
rect 27169 14365 27203 14399
rect 27203 14365 27212 14399
rect 27160 14356 27212 14365
rect 28540 14356 28592 14408
rect 30472 14399 30524 14408
rect 27344 14288 27396 14340
rect 30472 14365 30481 14399
rect 30481 14365 30515 14399
rect 30515 14365 30524 14399
rect 30472 14356 30524 14365
rect 27620 14220 27672 14272
rect 31852 14467 31904 14476
rect 31852 14433 31861 14467
rect 31861 14433 31895 14467
rect 31895 14433 31904 14467
rect 32036 14467 32088 14476
rect 31852 14424 31904 14433
rect 32036 14433 32045 14467
rect 32045 14433 32079 14467
rect 32079 14433 32088 14467
rect 32036 14424 32088 14433
rect 32772 14424 32824 14476
rect 42708 14560 42760 14612
rect 46664 14560 46716 14612
rect 47124 14560 47176 14612
rect 50712 14560 50764 14612
rect 50896 14560 50948 14612
rect 51448 14560 51500 14612
rect 51540 14560 51592 14612
rect 54208 14560 54260 14612
rect 41880 14492 41932 14544
rect 40592 14467 40644 14476
rect 34888 14356 34940 14408
rect 40592 14433 40601 14467
rect 40601 14433 40635 14467
rect 40635 14433 40644 14467
rect 40592 14424 40644 14433
rect 40684 14424 40736 14476
rect 41328 14424 41380 14476
rect 49332 14492 49384 14544
rect 53104 14492 53156 14544
rect 64880 14560 64932 14612
rect 59268 14492 59320 14544
rect 59360 14492 59412 14544
rect 60464 14492 60516 14544
rect 63040 14492 63092 14544
rect 32956 14288 33008 14340
rect 33968 14288 34020 14340
rect 37096 14399 37148 14408
rect 37096 14365 37105 14399
rect 37105 14365 37139 14399
rect 37139 14365 37148 14399
rect 37372 14399 37424 14408
rect 37096 14356 37148 14365
rect 37372 14365 37381 14399
rect 37381 14365 37415 14399
rect 37415 14365 37424 14399
rect 37372 14356 37424 14365
rect 38844 14399 38896 14408
rect 30012 14220 30064 14272
rect 30196 14220 30248 14272
rect 31392 14263 31444 14272
rect 31392 14229 31401 14263
rect 31401 14229 31435 14263
rect 31435 14229 31444 14263
rect 31392 14220 31444 14229
rect 34244 14263 34296 14272
rect 34244 14229 34253 14263
rect 34253 14229 34287 14263
rect 34287 14229 34296 14263
rect 34244 14220 34296 14229
rect 35072 14263 35124 14272
rect 35072 14229 35081 14263
rect 35081 14229 35115 14263
rect 35115 14229 35124 14263
rect 35072 14220 35124 14229
rect 35440 14220 35492 14272
rect 38844 14365 38853 14399
rect 38853 14365 38887 14399
rect 38887 14365 38896 14399
rect 38844 14356 38896 14365
rect 38568 14288 38620 14340
rect 40132 14356 40184 14408
rect 55772 14424 55824 14476
rect 43812 14399 43864 14408
rect 43812 14365 43821 14399
rect 43821 14365 43855 14399
rect 43855 14365 43864 14399
rect 43812 14356 43864 14365
rect 45468 14399 45520 14408
rect 45468 14365 45477 14399
rect 45477 14365 45511 14399
rect 45511 14365 45520 14399
rect 45468 14356 45520 14365
rect 45744 14356 45796 14408
rect 49240 14399 49292 14408
rect 49240 14365 49249 14399
rect 49249 14365 49283 14399
rect 49283 14365 49292 14399
rect 49240 14356 49292 14365
rect 50620 14356 50672 14408
rect 51540 14399 51592 14408
rect 51540 14365 51549 14399
rect 51549 14365 51583 14399
rect 51583 14365 51592 14399
rect 51540 14356 51592 14365
rect 53748 14356 53800 14408
rect 54944 14356 54996 14408
rect 55588 14356 55640 14408
rect 39120 14331 39172 14340
rect 39120 14297 39129 14331
rect 39129 14297 39163 14331
rect 39163 14297 39172 14331
rect 39120 14288 39172 14297
rect 41604 14288 41656 14340
rect 46848 14331 46900 14340
rect 41880 14220 41932 14272
rect 42708 14263 42760 14272
rect 42708 14229 42717 14263
rect 42717 14229 42751 14263
rect 42751 14229 42760 14263
rect 42708 14220 42760 14229
rect 44916 14220 44968 14272
rect 45192 14220 45244 14272
rect 46848 14297 46857 14331
rect 46857 14297 46891 14331
rect 46891 14297 46900 14331
rect 46848 14288 46900 14297
rect 47032 14288 47084 14340
rect 51816 14331 51868 14340
rect 47308 14220 47360 14272
rect 48320 14220 48372 14272
rect 49700 14263 49752 14272
rect 49700 14229 49709 14263
rect 49709 14229 49743 14263
rect 49743 14229 49752 14263
rect 49700 14220 49752 14229
rect 50068 14220 50120 14272
rect 50252 14220 50304 14272
rect 51816 14297 51825 14331
rect 51825 14297 51859 14331
rect 51859 14297 51868 14331
rect 51816 14288 51868 14297
rect 54852 14288 54904 14340
rect 56324 14424 56376 14476
rect 55956 14399 56008 14408
rect 55956 14365 55965 14399
rect 55965 14365 55999 14399
rect 55999 14365 56008 14399
rect 55956 14356 56008 14365
rect 58992 14356 59044 14408
rect 59912 14399 59964 14408
rect 59912 14365 59921 14399
rect 59921 14365 59955 14399
rect 59955 14365 59964 14399
rect 59912 14356 59964 14365
rect 60556 14424 60608 14476
rect 56232 14288 56284 14340
rect 57244 14331 57296 14340
rect 57244 14297 57253 14331
rect 57253 14297 57287 14331
rect 57287 14297 57296 14331
rect 57244 14288 57296 14297
rect 58256 14288 58308 14340
rect 60556 14288 60608 14340
rect 54484 14220 54536 14272
rect 57336 14220 57388 14272
rect 60004 14263 60056 14272
rect 60004 14229 60013 14263
rect 60013 14229 60047 14263
rect 60047 14229 60056 14263
rect 60004 14220 60056 14229
rect 62948 14356 63000 14408
rect 67640 14424 67692 14476
rect 68560 14424 68612 14476
rect 71044 14467 71096 14476
rect 71044 14433 71053 14467
rect 71053 14433 71087 14467
rect 71087 14433 71096 14467
rect 71044 14424 71096 14433
rect 71504 14535 71556 14544
rect 71504 14501 71513 14535
rect 71513 14501 71547 14535
rect 71547 14501 71556 14535
rect 75828 14560 75880 14612
rect 77116 14560 77168 14612
rect 77668 14560 77720 14612
rect 78496 14560 78548 14612
rect 92664 14603 92716 14612
rect 92664 14569 92673 14603
rect 92673 14569 92707 14603
rect 92707 14569 92716 14603
rect 92664 14560 92716 14569
rect 71504 14492 71556 14501
rect 77392 14492 77444 14544
rect 88524 14492 88576 14544
rect 65432 14356 65484 14408
rect 65984 14356 66036 14408
rect 66076 14399 66128 14408
rect 66076 14365 66085 14399
rect 66085 14365 66119 14399
rect 66119 14365 66128 14399
rect 66076 14356 66128 14365
rect 66536 14356 66588 14408
rect 67272 14356 67324 14408
rect 67732 14399 67784 14408
rect 67732 14365 67741 14399
rect 67741 14365 67775 14399
rect 67775 14365 67784 14399
rect 67732 14356 67784 14365
rect 68192 14399 68244 14408
rect 68192 14365 68201 14399
rect 68201 14365 68235 14399
rect 68235 14365 68244 14399
rect 68192 14356 68244 14365
rect 70952 14356 71004 14408
rect 73528 14356 73580 14408
rect 74816 14356 74868 14408
rect 78588 14424 78640 14476
rect 80336 14424 80388 14476
rect 80612 14424 80664 14476
rect 84108 14424 84160 14476
rect 79600 14399 79652 14408
rect 79600 14365 79609 14399
rect 79609 14365 79643 14399
rect 79643 14365 79652 14399
rect 79600 14356 79652 14365
rect 81808 14356 81860 14408
rect 83464 14399 83516 14408
rect 83464 14365 83473 14399
rect 83473 14365 83507 14399
rect 83507 14365 83516 14399
rect 83464 14356 83516 14365
rect 84936 14399 84988 14408
rect 84936 14365 84945 14399
rect 84945 14365 84979 14399
rect 84979 14365 84988 14399
rect 84936 14356 84988 14365
rect 86776 14399 86828 14408
rect 86776 14365 86785 14399
rect 86785 14365 86819 14399
rect 86819 14365 86828 14399
rect 86776 14356 86828 14365
rect 86960 14356 87012 14408
rect 88248 14356 88300 14408
rect 89352 14399 89404 14408
rect 89352 14365 89361 14399
rect 89361 14365 89395 14399
rect 89395 14365 89404 14399
rect 89352 14356 89404 14365
rect 61660 14288 61712 14340
rect 68468 14331 68520 14340
rect 68468 14297 68477 14331
rect 68477 14297 68511 14331
rect 68511 14297 68520 14331
rect 68468 14288 68520 14297
rect 71044 14288 71096 14340
rect 71872 14288 71924 14340
rect 63224 14220 63276 14272
rect 63684 14263 63736 14272
rect 63684 14229 63693 14263
rect 63693 14229 63727 14263
rect 63727 14229 63736 14263
rect 63684 14220 63736 14229
rect 64236 14263 64288 14272
rect 64236 14229 64245 14263
rect 64245 14229 64279 14263
rect 64279 14229 64288 14263
rect 64236 14220 64288 14229
rect 65156 14263 65208 14272
rect 65156 14229 65165 14263
rect 65165 14229 65199 14263
rect 65199 14229 65208 14263
rect 65156 14220 65208 14229
rect 65892 14263 65944 14272
rect 65892 14229 65901 14263
rect 65901 14229 65935 14263
rect 65935 14229 65944 14263
rect 65892 14220 65944 14229
rect 65984 14220 66036 14272
rect 69296 14220 69348 14272
rect 69940 14263 69992 14272
rect 69940 14229 69949 14263
rect 69949 14229 69983 14263
rect 69983 14229 69992 14263
rect 69940 14220 69992 14229
rect 72056 14263 72108 14272
rect 72056 14229 72065 14263
rect 72065 14229 72099 14263
rect 72099 14229 72108 14263
rect 72056 14220 72108 14229
rect 72332 14220 72384 14272
rect 76932 14288 76984 14340
rect 78220 14288 78272 14340
rect 78404 14288 78456 14340
rect 79232 14288 79284 14340
rect 82544 14288 82596 14340
rect 85672 14288 85724 14340
rect 89260 14331 89312 14340
rect 73988 14263 74040 14272
rect 73988 14229 73997 14263
rect 73997 14229 74031 14263
rect 74031 14229 74040 14263
rect 73988 14220 74040 14229
rect 75092 14220 75144 14272
rect 75184 14220 75236 14272
rect 75920 14220 75972 14272
rect 76196 14263 76248 14272
rect 76196 14229 76205 14263
rect 76205 14229 76239 14263
rect 76239 14229 76248 14263
rect 76196 14220 76248 14229
rect 78864 14220 78916 14272
rect 79508 14263 79560 14272
rect 79508 14229 79517 14263
rect 79517 14229 79551 14263
rect 79551 14229 79560 14263
rect 79508 14220 79560 14229
rect 80060 14220 80112 14272
rect 80612 14220 80664 14272
rect 81348 14220 81400 14272
rect 85028 14263 85080 14272
rect 85028 14229 85037 14263
rect 85037 14229 85071 14263
rect 85071 14229 85080 14263
rect 85028 14220 85080 14229
rect 85856 14220 85908 14272
rect 86408 14263 86460 14272
rect 86408 14229 86417 14263
rect 86417 14229 86451 14263
rect 86451 14229 86460 14263
rect 86408 14220 86460 14229
rect 88156 14263 88208 14272
rect 88156 14229 88165 14263
rect 88165 14229 88199 14263
rect 88199 14229 88208 14263
rect 88156 14220 88208 14229
rect 89260 14297 89269 14331
rect 89269 14297 89303 14331
rect 89303 14297 89312 14331
rect 89260 14288 89312 14297
rect 89536 14220 89588 14272
rect 91100 14220 91152 14272
rect 92480 14220 92532 14272
rect 24386 14118 24438 14170
rect 24450 14118 24502 14170
rect 24514 14118 24566 14170
rect 24578 14118 24630 14170
rect 24642 14118 24694 14170
rect 47823 14118 47875 14170
rect 47887 14118 47939 14170
rect 47951 14118 48003 14170
rect 48015 14118 48067 14170
rect 48079 14118 48131 14170
rect 71260 14118 71312 14170
rect 71324 14118 71376 14170
rect 71388 14118 71440 14170
rect 71452 14118 71504 14170
rect 71516 14118 71568 14170
rect 94697 14118 94749 14170
rect 94761 14118 94813 14170
rect 94825 14118 94877 14170
rect 94889 14118 94941 14170
rect 94953 14118 95005 14170
rect 9128 14016 9180 14068
rect 20444 14016 20496 14068
rect 8024 13948 8076 14000
rect 9312 13991 9364 14000
rect 2964 13923 3016 13932
rect 2964 13889 2973 13923
rect 2973 13889 3007 13923
rect 3007 13889 3016 13923
rect 2964 13880 3016 13889
rect 4160 13880 4212 13932
rect 7288 13880 7340 13932
rect 9312 13957 9321 13991
rect 9321 13957 9355 13991
rect 9355 13957 9364 13991
rect 9312 13948 9364 13957
rect 8208 13855 8260 13864
rect 8208 13821 8217 13855
rect 8217 13821 8251 13855
rect 8251 13821 8260 13855
rect 8208 13812 8260 13821
rect 12440 13880 12492 13932
rect 13912 13923 13964 13932
rect 13912 13889 13921 13923
rect 13921 13889 13955 13923
rect 13955 13889 13964 13923
rect 13912 13880 13964 13889
rect 16212 13948 16264 14000
rect 16948 13991 17000 14000
rect 16948 13957 16957 13991
rect 16957 13957 16991 13991
rect 16991 13957 17000 13991
rect 16948 13948 17000 13957
rect 20076 13948 20128 14000
rect 22652 14016 22704 14068
rect 15108 13880 15160 13932
rect 11980 13855 12032 13864
rect 11980 13821 11989 13855
rect 11989 13821 12023 13855
rect 12023 13821 12032 13855
rect 11980 13812 12032 13821
rect 14004 13855 14056 13864
rect 14004 13821 14013 13855
rect 14013 13821 14047 13855
rect 14047 13821 14056 13855
rect 14004 13812 14056 13821
rect 14464 13812 14516 13864
rect 15016 13855 15068 13864
rect 15016 13821 15025 13855
rect 15025 13821 15059 13855
rect 15059 13821 15068 13855
rect 15016 13812 15068 13821
rect 15844 13855 15896 13864
rect 15844 13821 15853 13855
rect 15853 13821 15887 13855
rect 15887 13821 15896 13855
rect 15844 13812 15896 13821
rect 4804 13719 4856 13728
rect 4804 13685 4813 13719
rect 4813 13685 4847 13719
rect 4847 13685 4856 13719
rect 4804 13676 4856 13685
rect 6828 13676 6880 13728
rect 10140 13676 10192 13728
rect 11336 13676 11388 13728
rect 15200 13744 15252 13796
rect 21272 13923 21324 13932
rect 21272 13889 21281 13923
rect 21281 13889 21315 13923
rect 21315 13889 21324 13923
rect 21272 13880 21324 13889
rect 23664 13948 23716 14000
rect 25688 14016 25740 14068
rect 26148 14016 26200 14068
rect 30288 14016 30340 14068
rect 37372 14016 37424 14068
rect 41420 14016 41472 14068
rect 47216 14059 47268 14068
rect 24308 13948 24360 14000
rect 25596 13948 25648 14000
rect 25044 13880 25096 13932
rect 30196 13948 30248 14000
rect 32404 13948 32456 14000
rect 27896 13880 27948 13932
rect 30104 13923 30156 13932
rect 30104 13889 30113 13923
rect 30113 13889 30147 13923
rect 30147 13889 30156 13923
rect 30104 13880 30156 13889
rect 31484 13880 31536 13932
rect 31760 13923 31812 13932
rect 31760 13889 31769 13923
rect 31769 13889 31803 13923
rect 31803 13889 31812 13923
rect 31760 13880 31812 13889
rect 32588 13880 32640 13932
rect 34244 13948 34296 14000
rect 35440 13991 35492 14000
rect 35440 13957 35449 13991
rect 35449 13957 35483 13991
rect 35483 13957 35492 13991
rect 35440 13948 35492 13957
rect 35624 13948 35676 14000
rect 36728 13948 36780 14000
rect 37464 13880 37516 13932
rect 22192 13812 22244 13864
rect 22560 13812 22612 13864
rect 25964 13812 26016 13864
rect 20076 13744 20128 13796
rect 25320 13744 25372 13796
rect 28264 13812 28316 13864
rect 29828 13812 29880 13864
rect 15752 13676 15804 13728
rect 17408 13719 17460 13728
rect 17408 13685 17417 13719
rect 17417 13685 17451 13719
rect 17451 13685 17460 13719
rect 17408 13676 17460 13685
rect 17500 13676 17552 13728
rect 19616 13676 19668 13728
rect 19708 13676 19760 13728
rect 28540 13676 28592 13728
rect 29644 13676 29696 13728
rect 30196 13744 30248 13796
rect 30104 13676 30156 13728
rect 30748 13812 30800 13864
rect 30932 13812 30984 13864
rect 33968 13855 34020 13864
rect 33968 13821 33977 13855
rect 33977 13821 34011 13855
rect 34011 13821 34020 13855
rect 33968 13812 34020 13821
rect 34060 13812 34112 13864
rect 35072 13812 35124 13864
rect 37280 13812 37332 13864
rect 38568 13948 38620 14000
rect 38476 13923 38528 13932
rect 38476 13889 38485 13923
rect 38485 13889 38519 13923
rect 38519 13889 38528 13923
rect 38476 13880 38528 13889
rect 39120 13948 39172 14000
rect 40224 13948 40276 14000
rect 40500 13948 40552 14000
rect 40960 13923 41012 13932
rect 40960 13889 40969 13923
rect 40969 13889 41003 13923
rect 41003 13889 41012 13923
rect 40960 13880 41012 13889
rect 41788 13880 41840 13932
rect 42432 13880 42484 13932
rect 44088 13948 44140 14000
rect 42800 13880 42852 13932
rect 47216 14025 47225 14059
rect 47225 14025 47259 14059
rect 47259 14025 47268 14059
rect 47216 14016 47268 14025
rect 47308 14016 47360 14068
rect 45652 13948 45704 14000
rect 46480 13948 46532 14000
rect 48320 13948 48372 14000
rect 48780 13948 48832 14000
rect 49516 13948 49568 14000
rect 50068 13948 50120 14000
rect 49332 13880 49384 13932
rect 52368 13880 52420 13932
rect 53564 13880 53616 13932
rect 53748 13923 53800 13932
rect 53748 13889 53757 13923
rect 53757 13889 53791 13923
rect 53791 13889 53800 13923
rect 53748 13880 53800 13889
rect 38200 13812 38252 13864
rect 44824 13855 44876 13864
rect 30472 13744 30524 13796
rect 38660 13744 38712 13796
rect 30656 13676 30708 13728
rect 31024 13676 31076 13728
rect 33140 13676 33192 13728
rect 33324 13676 33376 13728
rect 33416 13676 33468 13728
rect 35992 13676 36044 13728
rect 36452 13676 36504 13728
rect 38844 13676 38896 13728
rect 44824 13821 44833 13855
rect 44833 13821 44867 13855
rect 44867 13821 44876 13855
rect 44824 13812 44876 13821
rect 45744 13855 45796 13864
rect 45744 13821 45753 13855
rect 45753 13821 45787 13855
rect 45787 13821 45796 13855
rect 45744 13812 45796 13821
rect 46112 13812 46164 13864
rect 50344 13812 50396 13864
rect 51448 13812 51500 13864
rect 54944 13880 54996 13932
rect 55312 13880 55364 13932
rect 54208 13855 54260 13864
rect 54208 13821 54217 13855
rect 54217 13821 54251 13855
rect 54251 13821 54260 13855
rect 54208 13812 54260 13821
rect 42248 13676 42300 13728
rect 49792 13744 49844 13796
rect 52276 13744 52328 13796
rect 53840 13744 53892 13796
rect 48780 13676 48832 13728
rect 49700 13676 49752 13728
rect 50436 13676 50488 13728
rect 51632 13719 51684 13728
rect 51632 13685 51641 13719
rect 51641 13685 51675 13719
rect 51675 13685 51684 13719
rect 51632 13676 51684 13685
rect 52184 13719 52236 13728
rect 52184 13685 52193 13719
rect 52193 13685 52227 13719
rect 52227 13685 52236 13719
rect 52184 13676 52236 13685
rect 53656 13719 53708 13728
rect 53656 13685 53665 13719
rect 53665 13685 53699 13719
rect 53699 13685 53708 13719
rect 53656 13676 53708 13685
rect 55772 14016 55824 14068
rect 58256 14059 58308 14068
rect 56048 13948 56100 14000
rect 56692 13948 56744 14000
rect 57980 13948 58032 14000
rect 57336 13880 57388 13932
rect 58256 14025 58265 14059
rect 58265 14025 58299 14059
rect 58299 14025 58308 14059
rect 58256 14016 58308 14025
rect 58348 14016 58400 14068
rect 59268 13991 59320 14000
rect 59268 13957 59277 13991
rect 59277 13957 59311 13991
rect 59311 13957 59320 13991
rect 59268 13948 59320 13957
rect 60004 13948 60056 14000
rect 61108 13948 61160 14000
rect 61660 14016 61712 14068
rect 62212 14016 62264 14068
rect 67456 14059 67508 14068
rect 63868 13948 63920 14000
rect 65156 13948 65208 14000
rect 67456 14025 67465 14059
rect 67465 14025 67499 14059
rect 67499 14025 67508 14059
rect 67456 14016 67508 14025
rect 74816 14059 74868 14068
rect 67732 13948 67784 14000
rect 59452 13880 59504 13932
rect 61476 13880 61528 13932
rect 56692 13812 56744 13864
rect 57152 13812 57204 13864
rect 60464 13812 60516 13864
rect 60004 13744 60056 13796
rect 61568 13812 61620 13864
rect 64604 13880 64656 13932
rect 66536 13880 66588 13932
rect 64236 13812 64288 13864
rect 66628 13812 66680 13864
rect 74816 14025 74825 14059
rect 74825 14025 74859 14059
rect 74859 14025 74868 14059
rect 74816 14016 74868 14025
rect 78404 14016 78456 14068
rect 78588 14016 78640 14068
rect 81348 14016 81400 14068
rect 83464 14016 83516 14068
rect 71596 13948 71648 14000
rect 73712 13948 73764 14000
rect 72608 13923 72660 13932
rect 72608 13889 72617 13923
rect 72617 13889 72651 13923
rect 72651 13889 72660 13923
rect 73528 13923 73580 13932
rect 72608 13880 72660 13889
rect 73528 13889 73537 13923
rect 73537 13889 73571 13923
rect 73571 13889 73580 13923
rect 73528 13880 73580 13889
rect 73804 13880 73856 13932
rect 74356 13880 74408 13932
rect 75184 13880 75236 13932
rect 76932 13923 76984 13932
rect 56968 13676 57020 13728
rect 68652 13744 68704 13796
rect 70676 13744 70728 13796
rect 70768 13744 70820 13796
rect 72976 13812 73028 13864
rect 73896 13812 73948 13864
rect 76932 13889 76941 13923
rect 76941 13889 76975 13923
rect 76975 13889 76984 13923
rect 76932 13880 76984 13889
rect 73712 13744 73764 13796
rect 74264 13787 74316 13796
rect 74264 13753 74273 13787
rect 74273 13753 74307 13787
rect 74307 13753 74316 13787
rect 74264 13744 74316 13753
rect 78220 13880 78272 13932
rect 78128 13855 78180 13864
rect 78128 13821 78137 13855
rect 78137 13821 78171 13855
rect 78171 13821 78180 13855
rect 78128 13812 78180 13821
rect 79048 13948 79100 14000
rect 78680 13923 78732 13932
rect 78680 13889 78689 13923
rect 78689 13889 78723 13923
rect 78723 13889 78732 13923
rect 78680 13880 78732 13889
rect 80060 13880 80112 13932
rect 81348 13880 81400 13932
rect 84108 13880 84160 13932
rect 86960 14016 87012 14068
rect 88248 14059 88300 14068
rect 88248 14025 88257 14059
rect 88257 14025 88291 14059
rect 88291 14025 88300 14059
rect 88248 14016 88300 14025
rect 94044 14016 94096 14068
rect 89260 13991 89312 14000
rect 89260 13957 89269 13991
rect 89269 13957 89303 13991
rect 89303 13957 89312 13991
rect 89260 13948 89312 13957
rect 89812 13948 89864 14000
rect 90732 13880 90784 13932
rect 92664 13880 92716 13932
rect 83556 13812 83608 13864
rect 84660 13812 84712 13864
rect 84936 13855 84988 13864
rect 84936 13821 84945 13855
rect 84945 13821 84979 13855
rect 84979 13821 84988 13855
rect 84936 13812 84988 13821
rect 63500 13719 63552 13728
rect 63500 13685 63509 13719
rect 63509 13685 63543 13719
rect 63543 13685 63552 13719
rect 63500 13676 63552 13685
rect 64696 13719 64748 13728
rect 64696 13685 64705 13719
rect 64705 13685 64739 13719
rect 64739 13685 64748 13719
rect 64696 13676 64748 13685
rect 66536 13676 66588 13728
rect 68008 13676 68060 13728
rect 70860 13676 70912 13728
rect 73068 13676 73120 13728
rect 76840 13719 76892 13728
rect 76840 13685 76849 13719
rect 76849 13685 76883 13719
rect 76883 13685 76892 13719
rect 76840 13676 76892 13685
rect 77208 13676 77260 13728
rect 79692 13676 79744 13728
rect 80796 13744 80848 13796
rect 85028 13744 85080 13796
rect 87972 13812 88024 13864
rect 88984 13855 89036 13864
rect 88984 13821 88993 13855
rect 88993 13821 89027 13855
rect 89027 13821 89036 13855
rect 88984 13812 89036 13821
rect 80520 13676 80572 13728
rect 81072 13676 81124 13728
rect 85856 13676 85908 13728
rect 90548 13676 90600 13728
rect 92664 13676 92716 13728
rect 94136 13719 94188 13728
rect 94136 13685 94145 13719
rect 94145 13685 94179 13719
rect 94179 13685 94188 13719
rect 94136 13676 94188 13685
rect 12668 13574 12720 13626
rect 12732 13574 12784 13626
rect 12796 13574 12848 13626
rect 12860 13574 12912 13626
rect 12924 13574 12976 13626
rect 36105 13574 36157 13626
rect 36169 13574 36221 13626
rect 36233 13574 36285 13626
rect 36297 13574 36349 13626
rect 36361 13574 36413 13626
rect 59542 13574 59594 13626
rect 59606 13574 59658 13626
rect 59670 13574 59722 13626
rect 59734 13574 59786 13626
rect 59798 13574 59850 13626
rect 82979 13574 83031 13626
rect 83043 13574 83095 13626
rect 83107 13574 83159 13626
rect 83171 13574 83223 13626
rect 83235 13574 83287 13626
rect 5080 13515 5132 13524
rect 5080 13481 5089 13515
rect 5089 13481 5123 13515
rect 5123 13481 5132 13515
rect 5080 13472 5132 13481
rect 6828 13472 6880 13524
rect 7288 13404 7340 13456
rect 8116 13472 8168 13524
rect 19432 13472 19484 13524
rect 11244 13404 11296 13456
rect 13360 13404 13412 13456
rect 14004 13404 14056 13456
rect 21088 13472 21140 13524
rect 21916 13472 21968 13524
rect 22008 13472 22060 13524
rect 22100 13472 22152 13524
rect 2964 13379 3016 13388
rect 2964 13345 2973 13379
rect 2973 13345 3007 13379
rect 3007 13345 3016 13379
rect 2964 13336 3016 13345
rect 4068 13379 4120 13388
rect 4068 13345 4077 13379
rect 4077 13345 4111 13379
rect 4111 13345 4120 13379
rect 4068 13336 4120 13345
rect 7380 13336 7432 13388
rect 8484 13336 8536 13388
rect 9772 13379 9824 13388
rect 4160 13311 4212 13320
rect 4160 13277 4169 13311
rect 4169 13277 4203 13311
rect 4203 13277 4212 13311
rect 4160 13268 4212 13277
rect 5816 13311 5868 13320
rect 5816 13277 5825 13311
rect 5825 13277 5859 13311
rect 5859 13277 5868 13311
rect 5816 13268 5868 13277
rect 6828 13268 6880 13320
rect 9312 13268 9364 13320
rect 9772 13345 9781 13379
rect 9781 13345 9815 13379
rect 9815 13345 9824 13379
rect 9772 13336 9824 13345
rect 11428 13336 11480 13388
rect 14556 13379 14608 13388
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 10508 13311 10560 13320
rect 10508 13277 10517 13311
rect 10517 13277 10551 13311
rect 10551 13277 10560 13311
rect 10508 13268 10560 13277
rect 4436 13200 4488 13252
rect 14004 13268 14056 13320
rect 10692 13200 10744 13252
rect 11428 13200 11480 13252
rect 3424 13175 3476 13184
rect 3424 13141 3433 13175
rect 3433 13141 3467 13175
rect 3467 13141 3476 13175
rect 3424 13132 3476 13141
rect 4528 13175 4580 13184
rect 4528 13141 4537 13175
rect 4537 13141 4571 13175
rect 4571 13141 4580 13175
rect 4528 13132 4580 13141
rect 7012 13132 7064 13184
rect 7656 13132 7708 13184
rect 8484 13132 8536 13184
rect 13268 13132 13320 13184
rect 14556 13345 14565 13379
rect 14565 13345 14599 13379
rect 14599 13345 14608 13379
rect 14556 13336 14608 13345
rect 15016 13336 15068 13388
rect 16120 13336 16172 13388
rect 20720 13404 20772 13456
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 16764 13268 16816 13320
rect 17408 13268 17460 13320
rect 21272 13336 21324 13388
rect 22100 13336 22152 13388
rect 19248 13268 19300 13320
rect 19432 13311 19484 13320
rect 19432 13277 19441 13311
rect 19441 13277 19475 13311
rect 19475 13277 19484 13311
rect 19432 13268 19484 13277
rect 22192 13311 22244 13320
rect 22192 13277 22201 13311
rect 22201 13277 22235 13311
rect 22235 13277 22244 13311
rect 22192 13268 22244 13277
rect 15568 13200 15620 13252
rect 17500 13200 17552 13252
rect 19340 13200 19392 13252
rect 19708 13243 19760 13252
rect 19708 13209 19717 13243
rect 19717 13209 19751 13243
rect 19751 13209 19760 13243
rect 19708 13200 19760 13209
rect 16856 13175 16908 13184
rect 16856 13141 16865 13175
rect 16865 13141 16899 13175
rect 16899 13141 16908 13175
rect 16856 13132 16908 13141
rect 17960 13132 18012 13184
rect 21456 13200 21508 13252
rect 23204 13200 23256 13252
rect 25320 13472 25372 13524
rect 27436 13472 27488 13524
rect 27620 13472 27672 13524
rect 28448 13515 28500 13524
rect 28448 13481 28457 13515
rect 28457 13481 28491 13515
rect 28491 13481 28500 13515
rect 28448 13472 28500 13481
rect 28540 13472 28592 13524
rect 29460 13472 29512 13524
rect 30196 13472 30248 13524
rect 31024 13472 31076 13524
rect 31484 13515 31536 13524
rect 31484 13481 31493 13515
rect 31493 13481 31527 13515
rect 31527 13481 31536 13515
rect 31484 13472 31536 13481
rect 31760 13472 31812 13524
rect 32772 13472 32824 13524
rect 32864 13472 32916 13524
rect 33416 13472 33468 13524
rect 35900 13472 35952 13524
rect 37280 13515 37332 13524
rect 37280 13481 37289 13515
rect 37289 13481 37323 13515
rect 37323 13481 37332 13515
rect 37280 13472 37332 13481
rect 38476 13472 38528 13524
rect 42432 13472 42484 13524
rect 46848 13472 46900 13524
rect 26792 13404 26844 13456
rect 29552 13404 29604 13456
rect 30564 13336 30616 13388
rect 25964 13268 26016 13320
rect 27712 13268 27764 13320
rect 29736 13311 29788 13320
rect 29736 13277 29745 13311
rect 29745 13277 29779 13311
rect 29779 13277 29788 13311
rect 29736 13268 29788 13277
rect 26332 13200 26384 13252
rect 30012 13243 30064 13252
rect 21088 13132 21140 13184
rect 27436 13132 27488 13184
rect 29092 13132 29144 13184
rect 29644 13132 29696 13184
rect 30012 13209 30021 13243
rect 30021 13209 30055 13243
rect 30055 13209 30064 13243
rect 30012 13200 30064 13209
rect 30472 13200 30524 13252
rect 36452 13404 36504 13456
rect 36636 13404 36688 13456
rect 42524 13404 42576 13456
rect 32680 13379 32732 13388
rect 32680 13345 32689 13379
rect 32689 13345 32723 13379
rect 32723 13345 32732 13379
rect 32680 13336 32732 13345
rect 32772 13336 32824 13388
rect 32496 13311 32548 13320
rect 32496 13277 32505 13311
rect 32505 13277 32539 13311
rect 32539 13277 32548 13311
rect 32496 13268 32548 13277
rect 35440 13311 35492 13320
rect 35440 13277 35449 13311
rect 35449 13277 35483 13311
rect 35483 13277 35492 13311
rect 35440 13268 35492 13277
rect 31484 13200 31536 13252
rect 33968 13200 34020 13252
rect 35716 13200 35768 13252
rect 35992 13336 36044 13388
rect 45192 13379 45244 13388
rect 45192 13345 45201 13379
rect 45201 13345 45235 13379
rect 45235 13345 45244 13379
rect 45192 13336 45244 13345
rect 49332 13472 49384 13524
rect 52368 13472 52420 13524
rect 49608 13404 49660 13456
rect 51724 13404 51776 13456
rect 51540 13336 51592 13388
rect 36452 13268 36504 13320
rect 38292 13268 38344 13320
rect 38476 13268 38528 13320
rect 40316 13268 40368 13320
rect 42432 13311 42484 13320
rect 42432 13277 42441 13311
rect 42441 13277 42475 13311
rect 42475 13277 42484 13311
rect 42432 13268 42484 13277
rect 48780 13268 48832 13320
rect 49240 13268 49292 13320
rect 50344 13268 50396 13320
rect 39396 13200 39448 13252
rect 42892 13243 42944 13252
rect 32220 13132 32272 13184
rect 32864 13132 32916 13184
rect 35624 13132 35676 13184
rect 39948 13132 40000 13184
rect 40132 13175 40184 13184
rect 40132 13141 40141 13175
rect 40141 13141 40175 13175
rect 40175 13141 40184 13175
rect 40132 13132 40184 13141
rect 42892 13209 42901 13243
rect 42901 13209 42935 13243
rect 42935 13209 42944 13243
rect 42892 13200 42944 13209
rect 43168 13200 43220 13252
rect 46480 13200 46532 13252
rect 47676 13243 47728 13252
rect 47676 13209 47685 13243
rect 47685 13209 47719 13243
rect 47719 13209 47728 13243
rect 47676 13200 47728 13209
rect 49056 13200 49108 13252
rect 52092 13243 52144 13252
rect 52092 13209 52101 13243
rect 52101 13209 52135 13243
rect 52135 13209 52144 13243
rect 52092 13200 52144 13209
rect 53656 13200 53708 13252
rect 44732 13132 44784 13184
rect 46756 13132 46808 13184
rect 48964 13132 49016 13184
rect 51264 13132 51316 13184
rect 52184 13132 52236 13184
rect 56600 13472 56652 13524
rect 57244 13472 57296 13524
rect 57888 13472 57940 13524
rect 60464 13472 60516 13524
rect 61016 13472 61068 13524
rect 62120 13404 62172 13456
rect 64236 13404 64288 13456
rect 69020 13472 69072 13524
rect 70860 13472 70912 13524
rect 71044 13515 71096 13524
rect 71044 13481 71053 13515
rect 71053 13481 71087 13515
rect 71087 13481 71096 13515
rect 71044 13472 71096 13481
rect 71872 13472 71924 13524
rect 72516 13472 72568 13524
rect 76104 13515 76156 13524
rect 73068 13404 73120 13456
rect 76104 13481 76113 13515
rect 76113 13481 76147 13515
rect 76147 13481 76156 13515
rect 76104 13472 76156 13481
rect 78956 13472 79008 13524
rect 79048 13472 79100 13524
rect 79692 13472 79744 13524
rect 84200 13472 84252 13524
rect 85212 13515 85264 13524
rect 85212 13481 85221 13515
rect 85221 13481 85255 13515
rect 85255 13481 85264 13515
rect 85212 13472 85264 13481
rect 78312 13404 78364 13456
rect 79968 13404 80020 13456
rect 81164 13404 81216 13456
rect 88984 13472 89036 13524
rect 89352 13472 89404 13524
rect 89812 13515 89864 13524
rect 89812 13481 89821 13515
rect 89821 13481 89855 13515
rect 89855 13481 89864 13515
rect 89812 13472 89864 13481
rect 56232 13336 56284 13388
rect 58440 13336 58492 13388
rect 58992 13379 59044 13388
rect 58992 13345 59001 13379
rect 59001 13345 59035 13379
rect 59035 13345 59044 13379
rect 58992 13336 59044 13345
rect 57244 13243 57296 13252
rect 55864 13132 55916 13184
rect 56968 13132 57020 13184
rect 57244 13209 57253 13243
rect 57253 13209 57287 13243
rect 57287 13209 57296 13243
rect 57244 13200 57296 13209
rect 59176 13200 59228 13252
rect 59452 13268 59504 13320
rect 60648 13311 60700 13320
rect 60648 13277 60657 13311
rect 60657 13277 60691 13311
rect 60691 13277 60700 13311
rect 60648 13268 60700 13277
rect 61660 13268 61712 13320
rect 62488 13336 62540 13388
rect 62948 13336 63000 13388
rect 64604 13268 64656 13320
rect 65984 13311 66036 13320
rect 65984 13277 65993 13311
rect 65993 13277 66027 13311
rect 66027 13277 66036 13311
rect 65984 13268 66036 13277
rect 66168 13268 66220 13320
rect 61752 13200 61804 13252
rect 63500 13200 63552 13252
rect 59084 13132 59136 13184
rect 60740 13175 60792 13184
rect 60740 13141 60749 13175
rect 60749 13141 60783 13175
rect 60783 13141 60792 13175
rect 60740 13132 60792 13141
rect 63316 13132 63368 13184
rect 63408 13132 63460 13184
rect 66628 13200 66680 13252
rect 64696 13132 64748 13184
rect 65892 13175 65944 13184
rect 65892 13141 65901 13175
rect 65901 13141 65935 13175
rect 65935 13141 65944 13175
rect 65892 13132 65944 13141
rect 67088 13175 67140 13184
rect 67088 13141 67097 13175
rect 67097 13141 67131 13175
rect 67131 13141 67140 13175
rect 67088 13132 67140 13141
rect 69848 13311 69900 13320
rect 69848 13277 69857 13311
rect 69857 13277 69891 13311
rect 69891 13277 69900 13311
rect 69848 13268 69900 13277
rect 70308 13268 70360 13320
rect 72976 13268 73028 13320
rect 73988 13336 74040 13388
rect 79600 13336 79652 13388
rect 76564 13268 76616 13320
rect 77024 13311 77076 13320
rect 77024 13277 77033 13311
rect 77033 13277 77067 13311
rect 77067 13277 77076 13311
rect 77024 13268 77076 13277
rect 78956 13268 79008 13320
rect 79416 13268 79468 13320
rect 71780 13200 71832 13252
rect 71688 13132 71740 13184
rect 76840 13200 76892 13252
rect 76932 13200 76984 13252
rect 80336 13336 80388 13388
rect 86224 13336 86276 13388
rect 84476 13268 84528 13320
rect 92572 13336 92624 13388
rect 86408 13268 86460 13320
rect 86684 13311 86736 13320
rect 86684 13277 86693 13311
rect 86693 13277 86727 13311
rect 86727 13277 86736 13311
rect 86684 13268 86736 13277
rect 89076 13268 89128 13320
rect 90548 13311 90600 13320
rect 90548 13277 90557 13311
rect 90557 13277 90591 13311
rect 90591 13277 90600 13311
rect 90548 13268 90600 13277
rect 73252 13132 73304 13184
rect 79876 13132 79928 13184
rect 79968 13132 80020 13184
rect 83188 13243 83240 13252
rect 83188 13209 83197 13243
rect 83197 13209 83231 13243
rect 83231 13209 83240 13243
rect 83188 13200 83240 13209
rect 84568 13200 84620 13252
rect 87788 13200 87840 13252
rect 89444 13200 89496 13252
rect 93308 13243 93360 13252
rect 80612 13175 80664 13184
rect 80612 13141 80621 13175
rect 80621 13141 80655 13175
rect 80655 13141 80664 13175
rect 80612 13132 80664 13141
rect 81164 13132 81216 13184
rect 86500 13132 86552 13184
rect 91836 13175 91888 13184
rect 91836 13141 91845 13175
rect 91845 13141 91879 13175
rect 91879 13141 91888 13175
rect 91836 13132 91888 13141
rect 93308 13209 93317 13243
rect 93317 13209 93351 13243
rect 93351 13209 93360 13243
rect 93308 13200 93360 13209
rect 92572 13132 92624 13184
rect 24386 13030 24438 13082
rect 24450 13030 24502 13082
rect 24514 13030 24566 13082
rect 24578 13030 24630 13082
rect 24642 13030 24694 13082
rect 47823 13030 47875 13082
rect 47887 13030 47939 13082
rect 47951 13030 48003 13082
rect 48015 13030 48067 13082
rect 48079 13030 48131 13082
rect 71260 13030 71312 13082
rect 71324 13030 71376 13082
rect 71388 13030 71440 13082
rect 71452 13030 71504 13082
rect 71516 13030 71568 13082
rect 94697 13030 94749 13082
rect 94761 13030 94813 13082
rect 94825 13030 94877 13082
rect 94889 13030 94941 13082
rect 94953 13030 95005 13082
rect 4436 12971 4488 12980
rect 4436 12937 4445 12971
rect 4445 12937 4479 12971
rect 4479 12937 4488 12971
rect 4436 12928 4488 12937
rect 6552 12971 6604 12980
rect 6552 12937 6561 12971
rect 6561 12937 6595 12971
rect 6595 12937 6604 12971
rect 6552 12928 6604 12937
rect 4160 12860 4212 12912
rect 9588 12928 9640 12980
rect 11888 12971 11940 12980
rect 5080 12792 5132 12844
rect 5172 12724 5224 12776
rect 7656 12860 7708 12912
rect 8944 12860 8996 12912
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 13268 12928 13320 12980
rect 21456 12928 21508 12980
rect 6828 12792 6880 12844
rect 8668 12792 8720 12844
rect 9588 12835 9640 12844
rect 9588 12801 9597 12835
rect 9597 12801 9631 12835
rect 9631 12801 9640 12835
rect 9588 12792 9640 12801
rect 14280 12860 14332 12912
rect 15016 12860 15068 12912
rect 16856 12860 16908 12912
rect 13912 12835 13964 12844
rect 13912 12801 13921 12835
rect 13921 12801 13955 12835
rect 13955 12801 13964 12835
rect 13912 12792 13964 12801
rect 15844 12792 15896 12844
rect 7012 12767 7064 12776
rect 7012 12733 7021 12767
rect 7021 12733 7055 12767
rect 7055 12733 7064 12767
rect 7012 12724 7064 12733
rect 7932 12724 7984 12776
rect 8116 12767 8168 12776
rect 8116 12733 8125 12767
rect 8125 12733 8159 12767
rect 8159 12733 8168 12767
rect 8116 12724 8168 12733
rect 8484 12724 8536 12776
rect 10508 12724 10560 12776
rect 3424 12656 3476 12708
rect 15108 12724 15160 12776
rect 20444 12792 20496 12844
rect 22376 12860 22428 12912
rect 21272 12792 21324 12844
rect 23204 12860 23256 12912
rect 25136 12860 25188 12912
rect 26148 12928 26200 12980
rect 30472 12971 30524 12980
rect 25320 12860 25372 12912
rect 30472 12937 30481 12971
rect 30481 12937 30515 12971
rect 30515 12937 30524 12971
rect 30472 12928 30524 12937
rect 30564 12928 30616 12980
rect 45468 12971 45520 12980
rect 26240 12835 26292 12844
rect 26240 12801 26249 12835
rect 26249 12801 26283 12835
rect 26283 12801 26292 12835
rect 26240 12792 26292 12801
rect 27344 12792 27396 12844
rect 22192 12724 22244 12776
rect 5632 12588 5684 12640
rect 5816 12588 5868 12640
rect 11152 12588 11204 12640
rect 12532 12588 12584 12640
rect 13820 12631 13872 12640
rect 13820 12597 13829 12631
rect 13829 12597 13863 12631
rect 13863 12597 13872 12631
rect 13820 12588 13872 12597
rect 14004 12588 14056 12640
rect 19156 12656 19208 12708
rect 26332 12767 26384 12776
rect 26332 12733 26341 12767
rect 26341 12733 26375 12767
rect 26375 12733 26384 12767
rect 26332 12724 26384 12733
rect 27160 12724 27212 12776
rect 16304 12588 16356 12640
rect 16856 12588 16908 12640
rect 17500 12588 17552 12640
rect 18604 12631 18656 12640
rect 18604 12597 18613 12631
rect 18613 12597 18647 12631
rect 18647 12597 18656 12631
rect 18604 12588 18656 12597
rect 19616 12631 19668 12640
rect 19616 12597 19625 12631
rect 19625 12597 19659 12631
rect 19659 12597 19668 12631
rect 19616 12588 19668 12597
rect 22284 12588 22336 12640
rect 27252 12588 27304 12640
rect 27620 12588 27672 12640
rect 29552 12792 29604 12844
rect 30104 12792 30156 12844
rect 29276 12724 29328 12776
rect 29828 12767 29880 12776
rect 29828 12733 29837 12767
rect 29837 12733 29871 12767
rect 29871 12733 29880 12767
rect 29828 12724 29880 12733
rect 32404 12860 32456 12912
rect 32864 12903 32916 12912
rect 32864 12869 32873 12903
rect 32873 12869 32907 12903
rect 32907 12869 32916 12903
rect 32864 12860 32916 12869
rect 33324 12860 33376 12912
rect 38660 12903 38712 12912
rect 38660 12869 38669 12903
rect 38669 12869 38703 12903
rect 38703 12869 38712 12903
rect 38660 12860 38712 12869
rect 40132 12860 40184 12912
rect 30472 12792 30524 12844
rect 31300 12792 31352 12844
rect 31392 12792 31444 12844
rect 32588 12835 32640 12844
rect 31484 12724 31536 12776
rect 31668 12767 31720 12776
rect 31668 12733 31677 12767
rect 31677 12733 31711 12767
rect 31711 12733 31720 12767
rect 31668 12724 31720 12733
rect 32588 12801 32597 12835
rect 32597 12801 32631 12835
rect 32631 12801 32640 12835
rect 32588 12792 32640 12801
rect 34980 12835 35032 12844
rect 34980 12801 34989 12835
rect 34989 12801 35023 12835
rect 35023 12801 35032 12835
rect 34980 12792 35032 12801
rect 35532 12792 35584 12844
rect 37740 12835 37792 12844
rect 35624 12724 35676 12776
rect 31392 12656 31444 12708
rect 30840 12588 30892 12640
rect 31300 12631 31352 12640
rect 31300 12597 31309 12631
rect 31309 12597 31343 12631
rect 31343 12597 31352 12631
rect 31300 12588 31352 12597
rect 33600 12588 33652 12640
rect 33968 12588 34020 12640
rect 37740 12801 37749 12835
rect 37749 12801 37783 12835
rect 37783 12801 37792 12835
rect 37740 12792 37792 12801
rect 39948 12792 40000 12844
rect 41696 12835 41748 12844
rect 41696 12801 41705 12835
rect 41705 12801 41739 12835
rect 41739 12801 41748 12835
rect 41696 12792 41748 12801
rect 43076 12792 43128 12844
rect 43996 12792 44048 12844
rect 44732 12860 44784 12912
rect 45468 12937 45477 12971
rect 45477 12937 45511 12971
rect 45511 12937 45520 12971
rect 45468 12928 45520 12937
rect 45928 12928 45980 12980
rect 46480 12928 46532 12980
rect 46940 12928 46992 12980
rect 50344 12928 50396 12980
rect 52000 12928 52052 12980
rect 53748 12928 53800 12980
rect 55036 12928 55088 12980
rect 55956 12928 56008 12980
rect 56600 12860 56652 12912
rect 57152 12928 57204 12980
rect 60372 12928 60424 12980
rect 60648 12928 60700 12980
rect 61292 12928 61344 12980
rect 61568 12971 61620 12980
rect 61568 12937 61577 12971
rect 61577 12937 61611 12971
rect 61611 12937 61620 12971
rect 61568 12928 61620 12937
rect 62120 12928 62172 12980
rect 66536 12971 66588 12980
rect 59360 12860 59412 12912
rect 60740 12860 60792 12912
rect 65892 12860 65944 12912
rect 44272 12792 44324 12844
rect 44824 12792 44876 12844
rect 46756 12835 46808 12844
rect 46756 12801 46765 12835
rect 46765 12801 46799 12835
rect 46799 12801 46808 12835
rect 46756 12792 46808 12801
rect 48136 12835 48188 12844
rect 37004 12724 37056 12776
rect 37280 12724 37332 12776
rect 39304 12724 39356 12776
rect 39396 12724 39448 12776
rect 41604 12724 41656 12776
rect 42340 12724 42392 12776
rect 42892 12767 42944 12776
rect 42892 12733 42901 12767
rect 42901 12733 42935 12767
rect 42935 12733 42944 12767
rect 42892 12724 42944 12733
rect 47032 12767 47084 12776
rect 40040 12656 40092 12708
rect 47032 12733 47041 12767
rect 47041 12733 47075 12767
rect 47075 12733 47084 12767
rect 47032 12724 47084 12733
rect 48136 12801 48145 12835
rect 48145 12801 48179 12835
rect 48179 12801 48188 12835
rect 48136 12792 48188 12801
rect 48964 12835 49016 12844
rect 48964 12801 48973 12835
rect 48973 12801 49007 12835
rect 49007 12801 49016 12835
rect 48964 12792 49016 12801
rect 49332 12835 49384 12844
rect 49332 12801 49341 12835
rect 49341 12801 49375 12835
rect 49375 12801 49384 12835
rect 49332 12792 49384 12801
rect 51724 12792 51776 12844
rect 52000 12792 52052 12844
rect 55036 12792 55088 12844
rect 58716 12792 58768 12844
rect 59084 12835 59136 12844
rect 59084 12801 59093 12835
rect 59093 12801 59127 12835
rect 59127 12801 59136 12835
rect 59084 12792 59136 12801
rect 61016 12792 61068 12844
rect 62028 12792 62080 12844
rect 63224 12835 63276 12844
rect 63224 12801 63233 12835
rect 63233 12801 63267 12835
rect 63267 12801 63276 12835
rect 63224 12792 63276 12801
rect 66168 12792 66220 12844
rect 66536 12937 66545 12971
rect 66545 12937 66579 12971
rect 66579 12937 66588 12971
rect 66536 12928 66588 12937
rect 66628 12928 66680 12980
rect 76932 12971 76984 12980
rect 66720 12860 66772 12912
rect 66904 12792 66956 12844
rect 67824 12792 67876 12844
rect 67916 12792 67968 12844
rect 68468 12792 68520 12844
rect 69020 12860 69072 12912
rect 70768 12903 70820 12912
rect 49700 12724 49752 12776
rect 49976 12724 50028 12776
rect 51172 12724 51224 12776
rect 51632 12724 51684 12776
rect 52184 12724 52236 12776
rect 54852 12724 54904 12776
rect 56232 12767 56284 12776
rect 56232 12733 56241 12767
rect 56241 12733 56275 12767
rect 56275 12733 56284 12767
rect 56232 12724 56284 12733
rect 43168 12699 43220 12708
rect 43168 12665 43177 12699
rect 43177 12665 43211 12699
rect 43211 12665 43220 12699
rect 43168 12656 43220 12665
rect 43260 12656 43312 12708
rect 55404 12656 55456 12708
rect 36912 12631 36964 12640
rect 36912 12597 36921 12631
rect 36921 12597 36955 12631
rect 36955 12597 36964 12631
rect 36912 12588 36964 12597
rect 39212 12588 39264 12640
rect 41696 12588 41748 12640
rect 41788 12588 41840 12640
rect 43904 12588 43956 12640
rect 43996 12588 44048 12640
rect 47032 12588 47084 12640
rect 50344 12588 50396 12640
rect 56876 12724 56928 12776
rect 61660 12724 61712 12776
rect 67088 12724 67140 12776
rect 68284 12724 68336 12776
rect 56416 12656 56468 12708
rect 57704 12656 57756 12708
rect 58256 12588 58308 12640
rect 58440 12656 58492 12708
rect 59084 12656 59136 12708
rect 60464 12656 60516 12708
rect 60648 12588 60700 12640
rect 61016 12588 61068 12640
rect 61936 12588 61988 12640
rect 62212 12588 62264 12640
rect 68376 12656 68428 12708
rect 68652 12699 68704 12708
rect 68652 12665 68661 12699
rect 68661 12665 68695 12699
rect 68695 12665 68704 12699
rect 68652 12656 68704 12665
rect 68836 12792 68888 12844
rect 70768 12869 70777 12903
rect 70777 12869 70811 12903
rect 70811 12869 70820 12903
rect 70768 12860 70820 12869
rect 72056 12860 72108 12912
rect 72424 12860 72476 12912
rect 70492 12835 70544 12844
rect 70492 12801 70501 12835
rect 70501 12801 70535 12835
rect 70535 12801 70544 12835
rect 70492 12792 70544 12801
rect 73528 12792 73580 12844
rect 75276 12792 75328 12844
rect 75736 12903 75788 12912
rect 75736 12869 75745 12903
rect 75745 12869 75779 12903
rect 75779 12869 75788 12903
rect 75736 12860 75788 12869
rect 76932 12937 76941 12971
rect 76941 12937 76975 12971
rect 76975 12937 76984 12971
rect 76932 12928 76984 12937
rect 77024 12928 77076 12980
rect 77208 12860 77260 12912
rect 79508 12860 79560 12912
rect 79876 12928 79928 12980
rect 83188 12928 83240 12980
rect 84568 12928 84620 12980
rect 87788 12971 87840 12980
rect 87788 12937 87797 12971
rect 87797 12937 87831 12971
rect 87831 12937 87840 12971
rect 87788 12928 87840 12937
rect 93308 12971 93360 12980
rect 93308 12937 93317 12971
rect 93317 12937 93351 12971
rect 93351 12937 93360 12971
rect 93308 12928 93360 12937
rect 77116 12792 77168 12844
rect 78680 12792 78732 12844
rect 80520 12792 80572 12844
rect 82268 12835 82320 12844
rect 82268 12801 82277 12835
rect 82277 12801 82311 12835
rect 82311 12801 82320 12835
rect 82268 12792 82320 12801
rect 85028 12860 85080 12912
rect 84108 12835 84160 12844
rect 69296 12767 69348 12776
rect 69296 12733 69305 12767
rect 69305 12733 69339 12767
rect 69339 12733 69348 12767
rect 69296 12724 69348 12733
rect 71964 12724 72016 12776
rect 72516 12767 72568 12776
rect 72516 12733 72525 12767
rect 72525 12733 72559 12767
rect 72559 12733 72568 12767
rect 72516 12724 72568 12733
rect 78220 12724 78272 12776
rect 70124 12588 70176 12640
rect 70952 12588 71004 12640
rect 71228 12588 71280 12640
rect 73896 12656 73948 12708
rect 75828 12656 75880 12708
rect 73528 12588 73580 12640
rect 73988 12588 74040 12640
rect 75000 12631 75052 12640
rect 75000 12597 75009 12631
rect 75009 12597 75043 12631
rect 75043 12597 75052 12631
rect 75000 12588 75052 12597
rect 75184 12588 75236 12640
rect 78312 12588 78364 12640
rect 78588 12588 78640 12640
rect 83832 12656 83884 12708
rect 84108 12801 84117 12835
rect 84117 12801 84151 12835
rect 84151 12801 84160 12835
rect 84108 12792 84160 12801
rect 84476 12656 84528 12708
rect 85212 12792 85264 12844
rect 86224 12835 86276 12844
rect 86224 12801 86233 12835
rect 86233 12801 86267 12835
rect 86267 12801 86276 12835
rect 86224 12792 86276 12801
rect 86868 12835 86920 12844
rect 86868 12801 86877 12835
rect 86877 12801 86911 12835
rect 86911 12801 86920 12835
rect 86868 12792 86920 12801
rect 89352 12860 89404 12912
rect 87788 12792 87840 12844
rect 89444 12835 89496 12844
rect 89444 12801 89453 12835
rect 89453 12801 89487 12835
rect 89487 12801 89496 12835
rect 89444 12792 89496 12801
rect 89536 12835 89588 12844
rect 89536 12801 89545 12835
rect 89545 12801 89579 12835
rect 89579 12801 89588 12835
rect 89536 12792 89588 12801
rect 90548 12792 90600 12844
rect 92480 12860 92532 12912
rect 92572 12835 92624 12844
rect 92572 12801 92581 12835
rect 92581 12801 92615 12835
rect 92615 12801 92624 12835
rect 92572 12792 92624 12801
rect 86776 12767 86828 12776
rect 86776 12733 86785 12767
rect 86785 12733 86819 12767
rect 86819 12733 86828 12767
rect 86776 12724 86828 12733
rect 89076 12724 89128 12776
rect 92112 12724 92164 12776
rect 93308 12792 93360 12844
rect 89628 12656 89680 12708
rect 80152 12588 80204 12640
rect 81532 12631 81584 12640
rect 81532 12597 81541 12631
rect 81541 12597 81575 12631
rect 81575 12597 81584 12631
rect 81532 12588 81584 12597
rect 85120 12588 85172 12640
rect 85580 12588 85632 12640
rect 90180 12631 90232 12640
rect 90180 12597 90189 12631
rect 90189 12597 90223 12631
rect 90223 12597 90232 12631
rect 90180 12588 90232 12597
rect 92940 12588 92992 12640
rect 12668 12486 12720 12538
rect 12732 12486 12784 12538
rect 12796 12486 12848 12538
rect 12860 12486 12912 12538
rect 12924 12486 12976 12538
rect 36105 12486 36157 12538
rect 36169 12486 36221 12538
rect 36233 12486 36285 12538
rect 36297 12486 36349 12538
rect 36361 12486 36413 12538
rect 59542 12486 59594 12538
rect 59606 12486 59658 12538
rect 59670 12486 59722 12538
rect 59734 12486 59786 12538
rect 59798 12486 59850 12538
rect 82979 12486 83031 12538
rect 83043 12486 83095 12538
rect 83107 12486 83159 12538
rect 83171 12486 83223 12538
rect 83235 12486 83287 12538
rect 4528 12384 4580 12436
rect 13912 12384 13964 12436
rect 15108 12384 15160 12436
rect 15752 12384 15804 12436
rect 4068 12248 4120 12300
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 13820 12248 13872 12300
rect 16120 12316 16172 12368
rect 15752 12248 15804 12300
rect 16948 12248 17000 12300
rect 19248 12316 19300 12368
rect 18604 12248 18656 12300
rect 19340 12248 19392 12300
rect 20444 12384 20496 12436
rect 22100 12384 22152 12436
rect 22192 12384 22244 12436
rect 22744 12384 22796 12436
rect 26424 12384 26476 12436
rect 29920 12427 29972 12436
rect 24032 12359 24084 12368
rect 24032 12325 24041 12359
rect 24041 12325 24075 12359
rect 24075 12325 24084 12359
rect 24032 12316 24084 12325
rect 26240 12316 26292 12368
rect 27160 12316 27212 12368
rect 22284 12291 22336 12300
rect 22284 12257 22293 12291
rect 22293 12257 22327 12291
rect 22327 12257 22336 12291
rect 22284 12248 22336 12257
rect 2964 12180 3016 12232
rect 5172 12180 5224 12232
rect 9680 12180 9732 12232
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 21640 12223 21692 12232
rect 16120 12180 16172 12189
rect 21640 12189 21649 12223
rect 21649 12189 21683 12223
rect 21683 12189 21692 12223
rect 21640 12180 21692 12189
rect 4528 12112 4580 12164
rect 5540 12112 5592 12164
rect 12992 12112 13044 12164
rect 13452 12155 13504 12164
rect 13452 12121 13461 12155
rect 13461 12121 13495 12155
rect 13495 12121 13504 12155
rect 13452 12112 13504 12121
rect 14004 12112 14056 12164
rect 15568 12112 15620 12164
rect 16856 12112 16908 12164
rect 18236 12155 18288 12164
rect 3056 12044 3108 12096
rect 6000 12087 6052 12096
rect 6000 12053 6009 12087
rect 6009 12053 6043 12087
rect 6043 12053 6052 12087
rect 6000 12044 6052 12053
rect 6828 12087 6880 12096
rect 6828 12053 6837 12087
rect 6837 12053 6871 12087
rect 6871 12053 6880 12087
rect 6828 12044 6880 12053
rect 7288 12087 7340 12096
rect 7288 12053 7297 12087
rect 7297 12053 7331 12087
rect 7331 12053 7340 12087
rect 7288 12044 7340 12053
rect 7932 12044 7984 12096
rect 11980 12087 12032 12096
rect 11980 12053 11989 12087
rect 11989 12053 12023 12087
rect 12023 12053 12032 12087
rect 11980 12044 12032 12053
rect 14372 12087 14424 12096
rect 14372 12053 14381 12087
rect 14381 12053 14415 12087
rect 14415 12053 14424 12087
rect 14372 12044 14424 12053
rect 15476 12044 15528 12096
rect 18236 12121 18245 12155
rect 18245 12121 18279 12155
rect 18279 12121 18288 12155
rect 18236 12112 18288 12121
rect 29920 12393 29929 12427
rect 29929 12393 29963 12427
rect 29963 12393 29972 12427
rect 29920 12384 29972 12393
rect 30748 12384 30800 12436
rect 34980 12427 35032 12436
rect 34980 12393 34989 12427
rect 34989 12393 35023 12427
rect 35023 12393 35032 12427
rect 34980 12384 35032 12393
rect 36452 12384 36504 12436
rect 37832 12384 37884 12436
rect 30656 12316 30708 12368
rect 26424 12180 26476 12232
rect 18420 12044 18472 12096
rect 26884 12112 26936 12164
rect 22744 12044 22796 12096
rect 23204 12044 23256 12096
rect 25412 12087 25464 12096
rect 25412 12053 25421 12087
rect 25421 12053 25455 12087
rect 25455 12053 25464 12087
rect 25412 12044 25464 12053
rect 25872 12087 25924 12096
rect 25872 12053 25881 12087
rect 25881 12053 25915 12087
rect 25915 12053 25924 12087
rect 25872 12044 25924 12053
rect 30288 12291 30340 12300
rect 27068 12223 27120 12232
rect 27068 12189 27077 12223
rect 27077 12189 27111 12223
rect 27111 12189 27120 12223
rect 27068 12180 27120 12189
rect 27252 12180 27304 12232
rect 30288 12257 30297 12291
rect 30297 12257 30331 12291
rect 30331 12257 30340 12291
rect 30288 12248 30340 12257
rect 31116 12291 31168 12300
rect 31116 12257 31125 12291
rect 31125 12257 31159 12291
rect 31159 12257 31168 12291
rect 31392 12316 31444 12368
rect 40500 12384 40552 12436
rect 42616 12384 42668 12436
rect 43444 12384 43496 12436
rect 31116 12248 31168 12257
rect 32404 12248 32456 12300
rect 28356 12180 28408 12232
rect 30196 12223 30248 12232
rect 30196 12189 30205 12223
rect 30205 12189 30239 12223
rect 30239 12189 30248 12223
rect 30196 12180 30248 12189
rect 31300 12180 31352 12232
rect 31760 12180 31812 12232
rect 32128 12223 32180 12232
rect 32128 12189 32137 12223
rect 32137 12189 32171 12223
rect 32171 12189 32180 12223
rect 32128 12180 32180 12189
rect 32220 12180 32272 12232
rect 33784 12223 33836 12232
rect 33784 12189 33793 12223
rect 33793 12189 33827 12223
rect 33827 12189 33836 12223
rect 33784 12180 33836 12189
rect 27160 12112 27212 12164
rect 32404 12112 32456 12164
rect 27896 12044 27948 12096
rect 33048 12112 33100 12164
rect 34244 12180 34296 12232
rect 36636 12248 36688 12300
rect 37004 12291 37056 12300
rect 37004 12257 37013 12291
rect 37013 12257 37047 12291
rect 37047 12257 37056 12291
rect 37004 12248 37056 12257
rect 39212 12291 39264 12300
rect 39212 12257 39221 12291
rect 39221 12257 39255 12291
rect 39255 12257 39264 12291
rect 39212 12248 39264 12257
rect 39488 12291 39540 12300
rect 39488 12257 39497 12291
rect 39497 12257 39531 12291
rect 39531 12257 39540 12291
rect 45284 12316 45336 12368
rect 39488 12248 39540 12257
rect 42708 12248 42760 12300
rect 47584 12384 47636 12436
rect 49608 12427 49660 12436
rect 49608 12393 49617 12427
rect 49617 12393 49651 12427
rect 49651 12393 49660 12427
rect 49608 12384 49660 12393
rect 49700 12384 49752 12436
rect 59360 12427 59412 12436
rect 45560 12316 45612 12368
rect 37280 12223 37332 12232
rect 37280 12189 37289 12223
rect 37289 12189 37323 12223
rect 37323 12189 37332 12223
rect 42524 12223 42576 12232
rect 37280 12180 37332 12189
rect 42524 12189 42533 12223
rect 42533 12189 42567 12223
rect 42567 12189 42576 12223
rect 42524 12180 42576 12189
rect 42616 12180 42668 12232
rect 46296 12248 46348 12300
rect 46756 12248 46808 12300
rect 48136 12248 48188 12300
rect 43812 12223 43864 12232
rect 43812 12189 43821 12223
rect 43821 12189 43855 12223
rect 43855 12189 43864 12223
rect 43812 12180 43864 12189
rect 43996 12223 44048 12232
rect 43996 12189 44005 12223
rect 44005 12189 44039 12223
rect 44039 12189 44048 12223
rect 43996 12180 44048 12189
rect 32864 12044 32916 12096
rect 34980 12044 35032 12096
rect 35440 12044 35492 12096
rect 36544 12112 36596 12164
rect 38200 12112 38252 12164
rect 38936 12112 38988 12164
rect 41788 12155 41840 12164
rect 41788 12121 41797 12155
rect 41797 12121 41831 12155
rect 41831 12121 41840 12155
rect 41788 12112 41840 12121
rect 44548 12155 44600 12164
rect 44548 12121 44557 12155
rect 44557 12121 44591 12155
rect 44591 12121 44600 12155
rect 44548 12112 44600 12121
rect 46020 12223 46072 12232
rect 46020 12189 46029 12223
rect 46029 12189 46063 12223
rect 46063 12189 46072 12223
rect 46020 12180 46072 12189
rect 48504 12223 48556 12232
rect 48504 12189 48513 12223
rect 48513 12189 48547 12223
rect 48547 12189 48556 12223
rect 48504 12180 48556 12189
rect 51540 12316 51592 12368
rect 51724 12316 51776 12368
rect 56140 12316 56192 12368
rect 56416 12316 56468 12368
rect 49516 12223 49568 12232
rect 49516 12189 49525 12223
rect 49525 12189 49559 12223
rect 49559 12189 49568 12223
rect 49516 12180 49568 12189
rect 36728 12044 36780 12096
rect 37004 12044 37056 12096
rect 43720 12044 43772 12096
rect 47124 12112 47176 12164
rect 48780 12155 48832 12164
rect 48780 12121 48789 12155
rect 48789 12121 48823 12155
rect 48823 12121 48832 12155
rect 48780 12112 48832 12121
rect 49240 12112 49292 12164
rect 45468 12087 45520 12096
rect 45468 12053 45477 12087
rect 45477 12053 45511 12087
rect 45511 12053 45520 12087
rect 45468 12044 45520 12053
rect 45652 12044 45704 12096
rect 50344 12180 50396 12232
rect 52184 12248 52236 12300
rect 55956 12248 56008 12300
rect 51264 12180 51316 12232
rect 51632 12180 51684 12232
rect 52828 12180 52880 12232
rect 52920 12180 52972 12232
rect 53288 12180 53340 12232
rect 57060 12180 57112 12232
rect 58072 12316 58124 12368
rect 59360 12393 59369 12427
rect 59369 12393 59403 12427
rect 59403 12393 59412 12427
rect 59360 12384 59412 12393
rect 60832 12384 60884 12436
rect 61752 12316 61804 12368
rect 62580 12316 62632 12368
rect 62120 12248 62172 12300
rect 67088 12384 67140 12436
rect 67640 12384 67692 12436
rect 69940 12384 69992 12436
rect 69204 12316 69256 12368
rect 71228 12316 71280 12368
rect 50160 12112 50212 12164
rect 50896 12112 50948 12164
rect 50068 12044 50120 12096
rect 50344 12044 50396 12096
rect 54208 12112 54260 12164
rect 54300 12112 54352 12164
rect 52000 12044 52052 12096
rect 52368 12044 52420 12096
rect 54484 12044 54536 12096
rect 55220 12044 55272 12096
rect 55772 12112 55824 12164
rect 57704 12180 57756 12232
rect 57520 12112 57572 12164
rect 57980 12223 58032 12232
rect 57980 12189 57989 12223
rect 57989 12189 58023 12223
rect 58023 12189 58032 12223
rect 57980 12180 58032 12189
rect 58348 12180 58400 12232
rect 58716 12180 58768 12232
rect 58900 12223 58952 12232
rect 58900 12189 58909 12223
rect 58909 12189 58943 12223
rect 58943 12189 58952 12223
rect 58900 12180 58952 12189
rect 60004 12180 60056 12232
rect 60648 12223 60700 12232
rect 60648 12189 60657 12223
rect 60657 12189 60691 12223
rect 60691 12189 60700 12223
rect 60648 12180 60700 12189
rect 61660 12180 61712 12232
rect 64696 12248 64748 12300
rect 65984 12223 66036 12232
rect 58532 12112 58584 12164
rect 65984 12189 65993 12223
rect 65993 12189 66027 12223
rect 66027 12189 66036 12223
rect 66628 12223 66680 12232
rect 65984 12180 66036 12189
rect 66628 12189 66637 12223
rect 66637 12189 66671 12223
rect 66671 12189 66680 12223
rect 66628 12180 66680 12189
rect 67548 12248 67600 12300
rect 71044 12248 71096 12300
rect 72240 12248 72292 12300
rect 73528 12291 73580 12300
rect 73528 12257 73537 12291
rect 73537 12257 73571 12291
rect 73571 12257 73580 12291
rect 73528 12248 73580 12257
rect 74816 12248 74868 12300
rect 75000 12384 75052 12436
rect 78588 12384 78640 12436
rect 78680 12384 78732 12436
rect 79968 12384 80020 12436
rect 80244 12427 80296 12436
rect 80244 12393 80253 12427
rect 80253 12393 80287 12427
rect 80287 12393 80296 12427
rect 80244 12384 80296 12393
rect 80796 12384 80848 12436
rect 84108 12427 84160 12436
rect 84108 12393 84117 12427
rect 84117 12393 84151 12427
rect 84151 12393 84160 12427
rect 84108 12384 84160 12393
rect 71504 12180 71556 12232
rect 75368 12248 75420 12300
rect 75644 12248 75696 12300
rect 77116 12291 77168 12300
rect 77116 12257 77125 12291
rect 77125 12257 77159 12291
rect 77159 12257 77168 12291
rect 77116 12248 77168 12257
rect 56600 12044 56652 12096
rect 59452 12044 59504 12096
rect 60648 12044 60700 12096
rect 61752 12044 61804 12096
rect 61936 12044 61988 12096
rect 63684 12044 63736 12096
rect 64788 12044 64840 12096
rect 65892 12087 65944 12096
rect 65892 12053 65901 12087
rect 65901 12053 65935 12087
rect 65935 12053 65944 12087
rect 65892 12044 65944 12053
rect 66536 12112 66588 12164
rect 68744 12112 68796 12164
rect 70768 12112 70820 12164
rect 67640 12044 67692 12096
rect 67732 12044 67784 12096
rect 70308 12087 70360 12096
rect 70308 12053 70317 12087
rect 70317 12053 70351 12087
rect 70351 12053 70360 12087
rect 70308 12044 70360 12053
rect 71136 12044 71188 12096
rect 71320 12087 71372 12096
rect 71320 12053 71329 12087
rect 71329 12053 71363 12087
rect 71363 12053 71372 12087
rect 71320 12044 71372 12053
rect 72516 12112 72568 12164
rect 72700 12112 72752 12164
rect 76380 12223 76432 12232
rect 76380 12189 76389 12223
rect 76389 12189 76423 12223
rect 76423 12189 76432 12223
rect 76380 12180 76432 12189
rect 76656 12180 76708 12232
rect 77024 12223 77076 12232
rect 77024 12189 77033 12223
rect 77033 12189 77067 12223
rect 77067 12189 77076 12223
rect 77024 12180 77076 12189
rect 77944 12316 77996 12368
rect 77576 12248 77628 12300
rect 78496 12291 78548 12300
rect 73896 12112 73948 12164
rect 74540 12112 74592 12164
rect 75552 12112 75604 12164
rect 75092 12044 75144 12096
rect 75644 12044 75696 12096
rect 75920 12112 75972 12164
rect 77484 12180 77536 12232
rect 78496 12257 78505 12291
rect 78505 12257 78539 12291
rect 78539 12257 78548 12291
rect 78496 12248 78548 12257
rect 78956 12316 79008 12368
rect 79600 12359 79652 12368
rect 79600 12325 79609 12359
rect 79609 12325 79643 12359
rect 79643 12325 79652 12359
rect 79600 12316 79652 12325
rect 79876 12316 79928 12368
rect 81072 12316 81124 12368
rect 81256 12359 81308 12368
rect 81256 12325 81265 12359
rect 81265 12325 81299 12359
rect 81299 12325 81308 12359
rect 81256 12316 81308 12325
rect 79232 12248 79284 12300
rect 79784 12248 79836 12300
rect 80336 12248 80388 12300
rect 78404 12180 78456 12232
rect 79876 12180 79928 12232
rect 84016 12316 84068 12368
rect 84568 12316 84620 12368
rect 81716 12291 81768 12300
rect 81716 12257 81725 12291
rect 81725 12257 81759 12291
rect 81759 12257 81768 12291
rect 81716 12248 81768 12257
rect 76196 12044 76248 12096
rect 79048 12155 79100 12164
rect 79048 12121 79057 12155
rect 79057 12121 79091 12155
rect 79091 12121 79100 12155
rect 79048 12112 79100 12121
rect 79784 12112 79836 12164
rect 77852 12044 77904 12096
rect 77944 12044 77996 12096
rect 78680 12044 78732 12096
rect 79600 12044 79652 12096
rect 81808 12180 81860 12232
rect 81164 12112 81216 12164
rect 85212 12248 85264 12300
rect 85580 12291 85632 12300
rect 85580 12257 85589 12291
rect 85589 12257 85623 12291
rect 85623 12257 85632 12291
rect 85580 12248 85632 12257
rect 85856 12291 85908 12300
rect 85856 12257 85865 12291
rect 85865 12257 85899 12291
rect 85899 12257 85908 12291
rect 85856 12248 85908 12257
rect 87788 12384 87840 12436
rect 93308 12427 93360 12436
rect 93308 12393 93317 12427
rect 93317 12393 93351 12427
rect 93351 12393 93360 12427
rect 93308 12384 93360 12393
rect 94228 12427 94280 12436
rect 94228 12393 94237 12427
rect 94237 12393 94271 12427
rect 94271 12393 94280 12427
rect 94228 12384 94280 12393
rect 86224 12316 86276 12368
rect 84108 12180 84160 12232
rect 84200 12180 84252 12232
rect 86224 12180 86276 12232
rect 92480 12248 92532 12300
rect 89536 12180 89588 12232
rect 94044 12223 94096 12232
rect 94044 12189 94053 12223
rect 94053 12189 94087 12223
rect 94087 12189 94096 12223
rect 94044 12180 94096 12189
rect 83648 12112 83700 12164
rect 85120 12112 85172 12164
rect 85580 12112 85632 12164
rect 91100 12112 91152 12164
rect 82360 12087 82412 12096
rect 82360 12053 82369 12087
rect 82369 12053 82403 12087
rect 82403 12053 82412 12087
rect 82360 12044 82412 12053
rect 84200 12044 84252 12096
rect 86960 12044 87012 12096
rect 89168 12087 89220 12096
rect 89168 12053 89177 12087
rect 89177 12053 89211 12087
rect 89211 12053 89220 12087
rect 89168 12044 89220 12053
rect 24386 11942 24438 11994
rect 24450 11942 24502 11994
rect 24514 11942 24566 11994
rect 24578 11942 24630 11994
rect 24642 11942 24694 11994
rect 47823 11942 47875 11994
rect 47887 11942 47939 11994
rect 47951 11942 48003 11994
rect 48015 11942 48067 11994
rect 48079 11942 48131 11994
rect 71260 11942 71312 11994
rect 71324 11942 71376 11994
rect 71388 11942 71440 11994
rect 71452 11942 71504 11994
rect 71516 11942 71568 11994
rect 94697 11942 94749 11994
rect 94761 11942 94813 11994
rect 94825 11942 94877 11994
rect 94889 11942 94941 11994
rect 94953 11942 95005 11994
rect 3976 11840 4028 11892
rect 4528 11883 4580 11892
rect 3056 11815 3108 11824
rect 3056 11781 3065 11815
rect 3065 11781 3099 11815
rect 3099 11781 3108 11815
rect 3056 11772 3108 11781
rect 4528 11849 4537 11883
rect 4537 11849 4571 11883
rect 4571 11849 4580 11883
rect 4528 11840 4580 11849
rect 9680 11883 9732 11892
rect 9680 11849 9689 11883
rect 9689 11849 9723 11883
rect 9723 11849 9732 11883
rect 9680 11840 9732 11849
rect 14004 11883 14056 11892
rect 14004 11849 14013 11883
rect 14013 11849 14047 11883
rect 14047 11849 14056 11883
rect 14004 11840 14056 11849
rect 6000 11772 6052 11824
rect 8208 11815 8260 11824
rect 8208 11781 8217 11815
rect 8217 11781 8251 11815
rect 8251 11781 8260 11815
rect 8208 11772 8260 11781
rect 8852 11772 8904 11824
rect 15384 11772 15436 11824
rect 18052 11772 18104 11824
rect 18420 11772 18472 11824
rect 6828 11704 6880 11756
rect 10140 11747 10192 11756
rect 2320 11636 2372 11688
rect 6920 11636 6972 11688
rect 7104 11611 7156 11620
rect 7104 11577 7113 11611
rect 7113 11577 7147 11611
rect 7147 11577 7156 11611
rect 7104 11568 7156 11577
rect 10140 11713 10149 11747
rect 10149 11713 10183 11747
rect 10183 11713 10192 11747
rect 10140 11704 10192 11713
rect 13360 11704 13412 11756
rect 13912 11747 13964 11756
rect 13912 11713 13921 11747
rect 13921 11713 13955 11747
rect 13955 11713 13964 11747
rect 13912 11704 13964 11713
rect 17132 11747 17184 11756
rect 17132 11713 17141 11747
rect 17141 11713 17175 11747
rect 17175 11713 17184 11747
rect 17132 11704 17184 11713
rect 17500 11704 17552 11756
rect 19248 11704 19300 11756
rect 7932 11679 7984 11688
rect 7932 11645 7941 11679
rect 7941 11645 7975 11679
rect 7975 11645 7984 11679
rect 7932 11636 7984 11645
rect 13176 11679 13228 11688
rect 13176 11645 13185 11679
rect 13185 11645 13219 11679
rect 13219 11645 13228 11679
rect 13176 11636 13228 11645
rect 13544 11636 13596 11688
rect 14832 11679 14884 11688
rect 14464 11568 14516 11620
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 5080 11543 5132 11552
rect 5080 11509 5089 11543
rect 5089 11509 5123 11543
rect 5123 11509 5132 11543
rect 5080 11500 5132 11509
rect 5540 11543 5592 11552
rect 5540 11509 5549 11543
rect 5549 11509 5583 11543
rect 5583 11509 5592 11543
rect 5540 11500 5592 11509
rect 11888 11500 11940 11552
rect 12992 11500 13044 11552
rect 14832 11645 14841 11679
rect 14841 11645 14875 11679
rect 14875 11645 14884 11679
rect 14832 11636 14884 11645
rect 15200 11636 15252 11688
rect 16120 11636 16172 11688
rect 18052 11636 18104 11688
rect 22560 11772 22612 11824
rect 22836 11772 22888 11824
rect 26240 11772 26292 11824
rect 26976 11840 27028 11892
rect 32496 11840 32548 11892
rect 36360 11840 36412 11892
rect 36544 11883 36596 11892
rect 36544 11849 36553 11883
rect 36553 11849 36587 11883
rect 36587 11849 36596 11883
rect 36544 11840 36596 11849
rect 36728 11840 36780 11892
rect 41972 11840 42024 11892
rect 42616 11883 42668 11892
rect 42616 11849 42625 11883
rect 42625 11849 42659 11883
rect 42659 11849 42668 11883
rect 42616 11840 42668 11849
rect 43720 11840 43772 11892
rect 21916 11704 21968 11756
rect 21640 11636 21692 11688
rect 25044 11679 25096 11688
rect 25044 11645 25053 11679
rect 25053 11645 25087 11679
rect 25087 11645 25096 11679
rect 25044 11636 25096 11645
rect 26056 11636 26108 11688
rect 26608 11679 26660 11688
rect 26608 11645 26617 11679
rect 26617 11645 26651 11679
rect 26651 11645 26660 11679
rect 26608 11636 26660 11645
rect 28816 11772 28868 11824
rect 30656 11815 30708 11824
rect 30656 11781 30665 11815
rect 30665 11781 30699 11815
rect 30699 11781 30708 11815
rect 30656 11772 30708 11781
rect 31116 11772 31168 11824
rect 33784 11772 33836 11824
rect 37188 11772 37240 11824
rect 37464 11772 37516 11824
rect 27160 11704 27212 11756
rect 29000 11704 29052 11756
rect 29460 11747 29512 11756
rect 29460 11713 29469 11747
rect 29469 11713 29503 11747
rect 29503 11713 29512 11747
rect 29460 11704 29512 11713
rect 19984 11500 20036 11552
rect 20168 11500 20220 11552
rect 27436 11679 27488 11688
rect 27436 11645 27445 11679
rect 27445 11645 27479 11679
rect 27479 11645 27488 11679
rect 27436 11636 27488 11645
rect 27804 11636 27856 11688
rect 28816 11636 28868 11688
rect 28908 11636 28960 11688
rect 29184 11636 29236 11688
rect 29368 11679 29420 11688
rect 29368 11645 29377 11679
rect 29377 11645 29411 11679
rect 29411 11645 29420 11679
rect 31576 11704 31628 11756
rect 33968 11747 34020 11756
rect 29368 11636 29420 11645
rect 27896 11568 27948 11620
rect 33508 11636 33560 11688
rect 33968 11713 33977 11747
rect 33977 11713 34011 11747
rect 34011 11713 34020 11747
rect 33968 11704 34020 11713
rect 34980 11704 35032 11756
rect 36452 11704 36504 11756
rect 36636 11747 36688 11756
rect 36636 11713 36645 11747
rect 36645 11713 36679 11747
rect 36679 11713 36688 11747
rect 36636 11704 36688 11713
rect 38844 11772 38896 11824
rect 39028 11815 39080 11824
rect 39028 11781 39037 11815
rect 39037 11781 39071 11815
rect 39071 11781 39080 11815
rect 39028 11772 39080 11781
rect 40592 11815 40644 11824
rect 40592 11781 40601 11815
rect 40601 11781 40635 11815
rect 40635 11781 40644 11815
rect 40592 11772 40644 11781
rect 44364 11840 44416 11892
rect 44088 11772 44140 11824
rect 52828 11840 52880 11892
rect 53748 11840 53800 11892
rect 31484 11568 31536 11620
rect 35440 11636 35492 11688
rect 36360 11636 36412 11688
rect 40224 11704 40276 11756
rect 41420 11704 41472 11756
rect 45652 11772 45704 11824
rect 46572 11815 46624 11824
rect 46572 11781 46581 11815
rect 46581 11781 46615 11815
rect 46615 11781 46624 11815
rect 46572 11772 46624 11781
rect 28632 11500 28684 11552
rect 31576 11500 31628 11552
rect 37740 11568 37792 11620
rect 38384 11636 38436 11688
rect 39580 11636 39632 11688
rect 39764 11679 39816 11688
rect 39764 11645 39773 11679
rect 39773 11645 39807 11679
rect 39807 11645 39816 11679
rect 39764 11636 39816 11645
rect 41604 11679 41656 11688
rect 41604 11645 41613 11679
rect 41613 11645 41647 11679
rect 41647 11645 41656 11679
rect 41604 11636 41656 11645
rect 42892 11636 42944 11688
rect 44088 11636 44140 11688
rect 44364 11679 44416 11688
rect 44364 11645 44373 11679
rect 44373 11645 44407 11679
rect 44407 11645 44416 11679
rect 44364 11636 44416 11645
rect 46848 11704 46900 11756
rect 50252 11772 50304 11824
rect 38200 11568 38252 11620
rect 38292 11568 38344 11620
rect 46020 11636 46072 11688
rect 46296 11636 46348 11688
rect 47584 11636 47636 11688
rect 50160 11704 50212 11756
rect 52276 11772 52328 11824
rect 49332 11679 49384 11688
rect 49332 11645 49341 11679
rect 49341 11645 49375 11679
rect 49375 11645 49384 11679
rect 49332 11636 49384 11645
rect 51908 11704 51960 11756
rect 52184 11747 52236 11756
rect 52184 11713 52193 11747
rect 52193 11713 52227 11747
rect 52227 11713 52236 11747
rect 52184 11704 52236 11713
rect 52368 11747 52420 11756
rect 52368 11713 52377 11747
rect 52377 11713 52411 11747
rect 52411 11713 52420 11747
rect 52368 11704 52420 11713
rect 52920 11747 52972 11756
rect 52920 11713 52929 11747
rect 52929 11713 52963 11747
rect 52963 11713 52972 11747
rect 52920 11704 52972 11713
rect 53012 11704 53064 11756
rect 50528 11636 50580 11688
rect 45192 11568 45244 11620
rect 45560 11568 45612 11620
rect 33416 11500 33468 11552
rect 35716 11500 35768 11552
rect 37464 11500 37516 11552
rect 41972 11500 42024 11552
rect 49608 11568 49660 11620
rect 51264 11636 51316 11688
rect 52276 11636 52328 11688
rect 54300 11772 54352 11824
rect 54852 11704 54904 11756
rect 55036 11747 55088 11756
rect 55036 11713 55045 11747
rect 55045 11713 55079 11747
rect 55079 11713 55088 11747
rect 55036 11704 55088 11713
rect 58808 11840 58860 11892
rect 57520 11815 57572 11824
rect 57520 11781 57529 11815
rect 57529 11781 57563 11815
rect 57563 11781 57572 11815
rect 57520 11772 57572 11781
rect 62304 11840 62356 11892
rect 63316 11840 63368 11892
rect 63684 11840 63736 11892
rect 62120 11772 62172 11824
rect 56692 11747 56744 11756
rect 56692 11713 56701 11747
rect 56701 11713 56735 11747
rect 56735 11713 56744 11747
rect 56692 11704 56744 11713
rect 57796 11704 57848 11756
rect 58256 11747 58308 11756
rect 58256 11713 58265 11747
rect 58265 11713 58299 11747
rect 58299 11713 58308 11747
rect 58256 11704 58308 11713
rect 56324 11636 56376 11688
rect 58532 11747 58584 11756
rect 58532 11713 58541 11747
rect 58541 11713 58575 11747
rect 58575 11713 58584 11747
rect 58532 11704 58584 11713
rect 58716 11704 58768 11756
rect 58900 11704 58952 11756
rect 63224 11772 63276 11824
rect 65892 11772 65944 11824
rect 63132 11704 63184 11756
rect 63592 11636 63644 11688
rect 64788 11636 64840 11688
rect 65064 11679 65116 11688
rect 65064 11645 65073 11679
rect 65073 11645 65107 11679
rect 65107 11645 65116 11679
rect 69848 11840 69900 11892
rect 71780 11840 71832 11892
rect 72608 11840 72660 11892
rect 73620 11883 73672 11892
rect 73620 11849 73629 11883
rect 73629 11849 73663 11883
rect 73663 11849 73672 11883
rect 73620 11840 73672 11849
rect 75368 11840 75420 11892
rect 77116 11840 77168 11892
rect 78680 11840 78732 11892
rect 79324 11840 79376 11892
rect 80612 11840 80664 11892
rect 66076 11772 66128 11824
rect 67732 11772 67784 11824
rect 68376 11815 68428 11824
rect 68376 11781 68385 11815
rect 68385 11781 68419 11815
rect 68419 11781 68428 11815
rect 68376 11772 68428 11781
rect 69940 11772 69992 11824
rect 67364 11747 67416 11756
rect 67364 11713 67373 11747
rect 67373 11713 67407 11747
rect 67407 11713 67416 11747
rect 67364 11704 67416 11713
rect 67824 11704 67876 11756
rect 68008 11704 68060 11756
rect 71136 11747 71188 11756
rect 65064 11636 65116 11645
rect 66168 11636 66220 11688
rect 52920 11568 52972 11620
rect 56508 11568 56560 11620
rect 60096 11568 60148 11620
rect 45744 11500 45796 11552
rect 46848 11500 46900 11552
rect 50436 11500 50488 11552
rect 51172 11500 51224 11552
rect 51264 11500 51316 11552
rect 52276 11500 52328 11552
rect 53012 11500 53064 11552
rect 53656 11500 53708 11552
rect 56140 11500 56192 11552
rect 57888 11500 57940 11552
rect 57980 11500 58032 11552
rect 58624 11500 58676 11552
rect 58900 11543 58952 11552
rect 58900 11509 58909 11543
rect 58909 11509 58943 11543
rect 58943 11509 58952 11543
rect 58900 11500 58952 11509
rect 58992 11500 59044 11552
rect 59360 11543 59412 11552
rect 59360 11509 59369 11543
rect 59369 11509 59403 11543
rect 59403 11509 59412 11543
rect 59360 11500 59412 11509
rect 60004 11500 60056 11552
rect 64972 11568 65024 11620
rect 65892 11568 65944 11620
rect 67272 11636 67324 11688
rect 71136 11713 71145 11747
rect 71145 11713 71179 11747
rect 71179 11713 71188 11747
rect 71136 11704 71188 11713
rect 70676 11636 70728 11688
rect 73988 11772 74040 11824
rect 74172 11815 74224 11824
rect 74172 11781 74181 11815
rect 74181 11781 74215 11815
rect 74215 11781 74224 11815
rect 74172 11772 74224 11781
rect 75736 11772 75788 11824
rect 79600 11815 79652 11824
rect 72056 11704 72108 11756
rect 72240 11704 72292 11756
rect 72608 11704 72660 11756
rect 72792 11704 72844 11756
rect 73528 11747 73580 11756
rect 73528 11713 73537 11747
rect 73537 11713 73571 11747
rect 73571 11713 73580 11747
rect 73528 11704 73580 11713
rect 75368 11747 75420 11756
rect 75368 11713 75377 11747
rect 75377 11713 75411 11747
rect 75411 11713 75420 11747
rect 75368 11704 75420 11713
rect 75552 11747 75604 11756
rect 75552 11713 75561 11747
rect 75561 11713 75595 11747
rect 75595 11713 75604 11747
rect 75552 11704 75604 11713
rect 75920 11704 75972 11756
rect 74080 11636 74132 11688
rect 74724 11679 74776 11688
rect 74724 11645 74733 11679
rect 74733 11645 74767 11679
rect 74767 11645 74776 11679
rect 74724 11636 74776 11645
rect 75828 11636 75880 11688
rect 66904 11568 66956 11620
rect 67088 11568 67140 11620
rect 76748 11747 76800 11756
rect 76748 11713 76757 11747
rect 76757 11713 76791 11747
rect 76791 11713 76800 11747
rect 76748 11704 76800 11713
rect 77116 11704 77168 11756
rect 79600 11781 79609 11815
rect 79609 11781 79643 11815
rect 79643 11781 79652 11815
rect 79600 11772 79652 11781
rect 80152 11815 80204 11824
rect 80152 11781 80161 11815
rect 80161 11781 80195 11815
rect 80195 11781 80204 11815
rect 80152 11772 80204 11781
rect 81256 11772 81308 11824
rect 84200 11840 84252 11892
rect 84292 11840 84344 11892
rect 85672 11840 85724 11892
rect 86132 11840 86184 11892
rect 82360 11772 82412 11824
rect 77484 11704 77536 11756
rect 77944 11704 77996 11756
rect 79048 11747 79100 11756
rect 76196 11636 76248 11688
rect 79048 11713 79057 11747
rect 79057 11713 79091 11747
rect 79091 11713 79100 11747
rect 79048 11704 79100 11713
rect 79508 11704 79560 11756
rect 80244 11636 80296 11688
rect 60372 11500 60424 11552
rect 62580 11500 62632 11552
rect 63592 11500 63644 11552
rect 67272 11500 67324 11552
rect 69480 11500 69532 11552
rect 69664 11543 69716 11552
rect 69664 11509 69673 11543
rect 69673 11509 69707 11543
rect 69707 11509 69716 11543
rect 69664 11500 69716 11509
rect 71596 11500 71648 11552
rect 72700 11500 72752 11552
rect 72884 11543 72936 11552
rect 72884 11509 72893 11543
rect 72893 11509 72927 11543
rect 72927 11509 72936 11543
rect 72884 11500 72936 11509
rect 73988 11500 74040 11552
rect 76932 11568 76984 11620
rect 78864 11568 78916 11620
rect 76196 11543 76248 11552
rect 76196 11509 76205 11543
rect 76205 11509 76239 11543
rect 76239 11509 76248 11543
rect 76196 11500 76248 11509
rect 77208 11500 77260 11552
rect 80704 11747 80756 11756
rect 80704 11713 80713 11747
rect 80713 11713 80747 11747
rect 80747 11713 80756 11747
rect 80704 11704 80756 11713
rect 83740 11704 83792 11756
rect 85948 11772 86000 11824
rect 84384 11704 84436 11756
rect 89168 11840 89220 11892
rect 90548 11772 90600 11824
rect 89168 11747 89220 11756
rect 89168 11713 89177 11747
rect 89177 11713 89211 11747
rect 89211 11713 89220 11747
rect 89168 11704 89220 11713
rect 92112 11747 92164 11756
rect 92112 11713 92121 11747
rect 92121 11713 92155 11747
rect 92155 11713 92164 11747
rect 92112 11704 92164 11713
rect 92296 11747 92348 11756
rect 92296 11713 92305 11747
rect 92305 11713 92339 11747
rect 92339 11713 92348 11747
rect 92296 11704 92348 11713
rect 93308 11704 93360 11756
rect 83004 11636 83056 11688
rect 83556 11636 83608 11688
rect 83832 11679 83884 11688
rect 83832 11645 83841 11679
rect 83841 11645 83875 11679
rect 83875 11645 83884 11679
rect 83832 11636 83884 11645
rect 84292 11679 84344 11688
rect 84292 11645 84301 11679
rect 84301 11645 84335 11679
rect 84335 11645 84344 11679
rect 84292 11636 84344 11645
rect 86960 11636 87012 11688
rect 87696 11679 87748 11688
rect 87696 11645 87705 11679
rect 87705 11645 87739 11679
rect 87739 11645 87748 11679
rect 87696 11636 87748 11645
rect 87972 11679 88024 11688
rect 87972 11645 87981 11679
rect 87981 11645 88015 11679
rect 88015 11645 88024 11679
rect 87972 11636 88024 11645
rect 88984 11636 89036 11688
rect 92480 11636 92532 11688
rect 93400 11636 93452 11688
rect 84660 11568 84712 11620
rect 84752 11568 84804 11620
rect 83004 11500 83056 11552
rect 86040 11500 86092 11552
rect 86224 11543 86276 11552
rect 86224 11509 86233 11543
rect 86233 11509 86267 11543
rect 86267 11509 86276 11543
rect 86224 11500 86276 11509
rect 89720 11568 89772 11620
rect 91100 11500 91152 11552
rect 12668 11398 12720 11450
rect 12732 11398 12784 11450
rect 12796 11398 12848 11450
rect 12860 11398 12912 11450
rect 12924 11398 12976 11450
rect 36105 11398 36157 11450
rect 36169 11398 36221 11450
rect 36233 11398 36285 11450
rect 36297 11398 36349 11450
rect 36361 11398 36413 11450
rect 59542 11398 59594 11450
rect 59606 11398 59658 11450
rect 59670 11398 59722 11450
rect 59734 11398 59786 11450
rect 59798 11398 59850 11450
rect 82979 11398 83031 11450
rect 83043 11398 83095 11450
rect 83107 11398 83159 11450
rect 83171 11398 83223 11450
rect 83235 11398 83287 11450
rect 1768 11339 1820 11348
rect 1768 11305 1777 11339
rect 1777 11305 1811 11339
rect 1811 11305 1820 11339
rect 1768 11296 1820 11305
rect 2504 11296 2556 11348
rect 5080 11296 5132 11348
rect 2504 11135 2556 11144
rect 2504 11101 2513 11135
rect 2513 11101 2547 11135
rect 2547 11101 2556 11135
rect 2504 11092 2556 11101
rect 3884 11092 3936 11144
rect 2320 11024 2372 11076
rect 3424 10999 3476 11008
rect 3424 10965 3433 10999
rect 3433 10965 3467 10999
rect 3467 10965 3476 10999
rect 3424 10956 3476 10965
rect 5448 11228 5500 11280
rect 6920 11296 6972 11348
rect 7380 11296 7432 11348
rect 9496 11296 9548 11348
rect 11888 11296 11940 11348
rect 6920 11160 6972 11212
rect 8484 11203 8536 11212
rect 8484 11169 8493 11203
rect 8493 11169 8527 11203
rect 8527 11169 8536 11203
rect 8484 11160 8536 11169
rect 4988 11092 5040 11144
rect 9772 11160 9824 11212
rect 12532 11228 12584 11280
rect 13452 11296 13504 11348
rect 14832 11296 14884 11348
rect 20168 11296 20220 11348
rect 20536 11296 20588 11348
rect 27620 11296 27672 11348
rect 28356 11296 28408 11348
rect 30012 11339 30064 11348
rect 30012 11305 30021 11339
rect 30021 11305 30055 11339
rect 30055 11305 30064 11339
rect 30012 11296 30064 11305
rect 31484 11339 31536 11348
rect 31484 11305 31493 11339
rect 31493 11305 31527 11339
rect 31527 11305 31536 11339
rect 31484 11296 31536 11305
rect 34520 11296 34572 11348
rect 37096 11296 37148 11348
rect 37188 11296 37240 11348
rect 39120 11296 39172 11348
rect 41696 11296 41748 11348
rect 41972 11339 42024 11348
rect 41972 11305 41981 11339
rect 41981 11305 42015 11339
rect 42015 11305 42024 11339
rect 41972 11296 42024 11305
rect 42892 11296 42944 11348
rect 43904 11296 43956 11348
rect 45468 11296 45520 11348
rect 51816 11296 51868 11348
rect 52000 11296 52052 11348
rect 14096 11228 14148 11280
rect 14372 11228 14424 11280
rect 19340 11228 19392 11280
rect 19432 11228 19484 11280
rect 12256 11160 12308 11212
rect 13360 11160 13412 11212
rect 15936 11160 15988 11212
rect 6000 11024 6052 11076
rect 4620 10956 4672 11008
rect 7288 11024 7340 11076
rect 8484 11024 8536 11076
rect 11796 11092 11848 11144
rect 8024 10999 8076 11008
rect 8024 10965 8033 10999
rect 8033 10965 8067 10999
rect 8067 10965 8076 10999
rect 8024 10956 8076 10965
rect 12532 11024 12584 11076
rect 15200 11092 15252 11144
rect 15476 11092 15528 11144
rect 15568 11092 15620 11144
rect 17132 11135 17184 11144
rect 17132 11101 17141 11135
rect 17141 11101 17175 11135
rect 17175 11101 17184 11135
rect 17132 11092 17184 11101
rect 16488 11024 16540 11076
rect 18328 11092 18380 11144
rect 18420 11092 18472 11144
rect 20812 11160 20864 11212
rect 25872 11228 25924 11280
rect 28816 11228 28868 11280
rect 30472 11228 30524 11280
rect 31300 11228 31352 11280
rect 32496 11228 32548 11280
rect 19340 11092 19392 11144
rect 17868 11024 17920 11076
rect 19616 11135 19668 11144
rect 19616 11101 19625 11135
rect 19625 11101 19659 11135
rect 19659 11101 19668 11135
rect 19616 11092 19668 11101
rect 19984 11092 20036 11144
rect 22744 11092 22796 11144
rect 22928 11024 22980 11076
rect 27436 11160 27488 11212
rect 29368 11160 29420 11212
rect 25872 11092 25924 11144
rect 27528 11092 27580 11144
rect 29460 11092 29512 11144
rect 36544 11160 36596 11212
rect 36820 11160 36872 11212
rect 37556 11160 37608 11212
rect 38016 11203 38068 11212
rect 38016 11169 38025 11203
rect 38025 11169 38059 11203
rect 38059 11169 38068 11203
rect 38016 11160 38068 11169
rect 38292 11203 38344 11212
rect 38292 11169 38301 11203
rect 38301 11169 38335 11203
rect 38335 11169 38344 11203
rect 38292 11160 38344 11169
rect 38660 11160 38712 11212
rect 44456 11228 44508 11280
rect 52368 11228 52420 11280
rect 53472 11228 53524 11280
rect 53656 11228 53708 11280
rect 32496 11135 32548 11144
rect 32496 11101 32505 11135
rect 32505 11101 32539 11135
rect 32539 11101 32548 11135
rect 32496 11092 32548 11101
rect 35256 11092 35308 11144
rect 38844 11092 38896 11144
rect 39764 11092 39816 11144
rect 40500 11135 40552 11144
rect 40500 11101 40509 11135
rect 40509 11101 40543 11135
rect 40543 11101 40552 11135
rect 40500 11092 40552 11101
rect 41788 11092 41840 11144
rect 42156 11092 42208 11144
rect 43812 11135 43864 11144
rect 43812 11101 43821 11135
rect 43821 11101 43855 11135
rect 43855 11101 43864 11135
rect 43812 11092 43864 11101
rect 43996 11203 44048 11212
rect 43996 11169 44005 11203
rect 44005 11169 44039 11203
rect 44039 11169 44048 11203
rect 44640 11203 44692 11212
rect 43996 11160 44048 11169
rect 44640 11169 44649 11203
rect 44649 11169 44683 11203
rect 44683 11169 44692 11203
rect 44640 11160 44692 11169
rect 48964 11203 49016 11212
rect 48964 11169 48973 11203
rect 48973 11169 49007 11203
rect 49007 11169 49016 11203
rect 48964 11160 49016 11169
rect 45744 11092 45796 11144
rect 46756 11135 46808 11144
rect 46756 11101 46765 11135
rect 46765 11101 46799 11135
rect 46799 11101 46808 11135
rect 46756 11092 46808 11101
rect 13636 10956 13688 11008
rect 15016 10956 15068 11008
rect 19064 10956 19116 11008
rect 19294 10956 19346 11008
rect 19432 10956 19484 11008
rect 19800 10956 19852 11008
rect 20996 10956 21048 11008
rect 23940 10956 23992 11008
rect 24768 10956 24820 11008
rect 26240 10956 26292 11008
rect 26700 11024 26752 11076
rect 29092 11024 29144 11076
rect 30288 11024 30340 11076
rect 30380 11024 30432 11076
rect 33048 11024 33100 11076
rect 34336 11024 34388 11076
rect 34796 11024 34848 11076
rect 35624 11024 35676 11076
rect 38200 11024 38252 11076
rect 41972 11024 42024 11076
rect 29000 10956 29052 11008
rect 30012 10956 30064 11008
rect 31760 10956 31812 11008
rect 31852 10956 31904 11008
rect 37372 10956 37424 11008
rect 37464 10956 37516 11008
rect 38292 10956 38344 11008
rect 38384 10956 38436 11008
rect 39764 10956 39816 11008
rect 42800 11024 42852 11076
rect 48780 11092 48832 11144
rect 50436 11160 50488 11212
rect 51908 11160 51960 11212
rect 49608 11135 49660 11144
rect 49608 11101 49617 11135
rect 49617 11101 49651 11135
rect 49651 11101 49660 11135
rect 49608 11092 49660 11101
rect 49700 11135 49752 11144
rect 49700 11101 49709 11135
rect 49709 11101 49743 11135
rect 49743 11101 49752 11135
rect 49700 11092 49752 11101
rect 50068 11092 50120 11144
rect 50620 11135 50672 11144
rect 50620 11101 50629 11135
rect 50629 11101 50663 11135
rect 50663 11101 50672 11135
rect 50620 11092 50672 11101
rect 50712 11092 50764 11144
rect 51264 11135 51316 11144
rect 51264 11101 51273 11135
rect 51273 11101 51307 11135
rect 51307 11101 51316 11135
rect 51264 11092 51316 11101
rect 51724 11092 51776 11144
rect 53564 11160 53616 11212
rect 54392 11160 54444 11212
rect 57336 11296 57388 11348
rect 57612 11296 57664 11348
rect 59636 11296 59688 11348
rect 62488 11296 62540 11348
rect 63592 11339 63644 11348
rect 63592 11305 63601 11339
rect 63601 11305 63635 11339
rect 63635 11305 63644 11339
rect 63592 11296 63644 11305
rect 64420 11296 64472 11348
rect 64972 11296 65024 11348
rect 54668 11271 54720 11280
rect 54668 11237 54677 11271
rect 54677 11237 54711 11271
rect 54711 11237 54720 11271
rect 54668 11228 54720 11237
rect 54760 11228 54812 11280
rect 55956 11228 56008 11280
rect 57428 11228 57480 11280
rect 59176 11228 59228 11280
rect 58164 11160 58216 11212
rect 58440 11160 58492 11212
rect 58624 11203 58676 11212
rect 58624 11169 58633 11203
rect 58633 11169 58667 11203
rect 58667 11169 58676 11203
rect 58624 11160 58676 11169
rect 59084 11160 59136 11212
rect 50528 11024 50580 11076
rect 50896 11024 50948 11076
rect 51356 11067 51408 11076
rect 42708 10956 42760 11008
rect 49240 10956 49292 11008
rect 49700 10956 49752 11008
rect 50804 10999 50856 11008
rect 50804 10965 50813 10999
rect 50813 10965 50847 10999
rect 50847 10965 50856 10999
rect 50804 10956 50856 10965
rect 51356 11033 51365 11067
rect 51365 11033 51399 11067
rect 51399 11033 51408 11067
rect 51356 11024 51408 11033
rect 52736 11024 52788 11076
rect 53012 11024 53064 11076
rect 54392 11024 54444 11076
rect 54668 11092 54720 11144
rect 55128 11092 55180 11144
rect 56048 11135 56100 11144
rect 56048 11101 56057 11135
rect 56057 11101 56091 11135
rect 56091 11101 56100 11135
rect 56048 11092 56100 11101
rect 56140 11135 56192 11144
rect 56140 11101 56149 11135
rect 56149 11101 56183 11135
rect 56183 11101 56192 11135
rect 56140 11092 56192 11101
rect 56324 11135 56376 11144
rect 56324 11101 56333 11135
rect 56333 11101 56367 11135
rect 56367 11101 56376 11135
rect 57336 11135 57388 11144
rect 56324 11092 56376 11101
rect 57336 11101 57345 11135
rect 57345 11101 57379 11135
rect 57379 11101 57388 11135
rect 57336 11092 57388 11101
rect 57704 11092 57756 11144
rect 61660 11228 61712 11280
rect 61752 11228 61804 11280
rect 60740 11203 60792 11212
rect 60740 11169 60749 11203
rect 60749 11169 60783 11203
rect 60783 11169 60792 11203
rect 60740 11160 60792 11169
rect 60924 11203 60976 11212
rect 60924 11169 60933 11203
rect 60933 11169 60967 11203
rect 60967 11169 60976 11203
rect 61844 11203 61896 11212
rect 60924 11160 60976 11169
rect 61844 11169 61853 11203
rect 61853 11169 61887 11203
rect 61887 11169 61896 11203
rect 61844 11160 61896 11169
rect 63224 11228 63276 11280
rect 66536 11296 66588 11348
rect 67272 11296 67324 11348
rect 67456 11296 67508 11348
rect 66444 11228 66496 11280
rect 62488 11160 62540 11212
rect 66628 11160 66680 11212
rect 69756 11203 69808 11212
rect 59636 11135 59688 11144
rect 59636 11101 59645 11135
rect 59645 11101 59679 11135
rect 59679 11101 59688 11135
rect 59636 11092 59688 11101
rect 56508 11024 56560 11076
rect 57980 11024 58032 11076
rect 58256 11067 58308 11076
rect 58256 11033 58265 11067
rect 58265 11033 58299 11067
rect 58299 11033 58308 11067
rect 58256 11024 58308 11033
rect 58440 11024 58492 11076
rect 58992 11067 59044 11076
rect 58992 11033 59001 11067
rect 59001 11033 59035 11067
rect 59035 11033 59044 11067
rect 58992 11024 59044 11033
rect 59084 11024 59136 11076
rect 51816 10956 51868 11008
rect 53564 10956 53616 11008
rect 54208 10956 54260 11008
rect 54944 10956 54996 11008
rect 59452 10956 59504 11008
rect 60556 10956 60608 11008
rect 61476 11092 61528 11144
rect 64604 11092 64656 11144
rect 65432 11092 65484 11144
rect 65984 11135 66036 11144
rect 65984 11101 65993 11135
rect 65993 11101 66027 11135
rect 66027 11101 66036 11135
rect 65984 11092 66036 11101
rect 62120 11024 62172 11076
rect 62396 11024 62448 11076
rect 67088 11067 67140 11076
rect 67088 11033 67097 11067
rect 67097 11033 67131 11067
rect 67131 11033 67140 11067
rect 67088 11024 67140 11033
rect 69756 11169 69765 11203
rect 69765 11169 69799 11203
rect 69799 11169 69808 11203
rect 69756 11160 69808 11169
rect 72700 11296 72752 11348
rect 74080 11339 74132 11348
rect 73804 11228 73856 11280
rect 74080 11305 74089 11339
rect 74089 11305 74123 11339
rect 74123 11305 74132 11339
rect 74080 11296 74132 11305
rect 74448 11296 74500 11348
rect 75276 11296 75328 11348
rect 76656 11296 76708 11348
rect 76932 11339 76984 11348
rect 76932 11305 76941 11339
rect 76941 11305 76975 11339
rect 76975 11305 76984 11339
rect 76932 11296 76984 11305
rect 77116 11296 77168 11348
rect 77484 11296 77536 11348
rect 78128 11296 78180 11348
rect 78588 11296 78640 11348
rect 78864 11339 78916 11348
rect 78864 11305 78873 11339
rect 78873 11305 78907 11339
rect 78907 11305 78916 11339
rect 78864 11296 78916 11305
rect 79968 11296 80020 11348
rect 85028 11296 85080 11348
rect 85212 11339 85264 11348
rect 85212 11305 85221 11339
rect 85221 11305 85255 11339
rect 85255 11305 85264 11339
rect 85212 11296 85264 11305
rect 87696 11296 87748 11348
rect 90548 11339 90600 11348
rect 90548 11305 90557 11339
rect 90557 11305 90591 11339
rect 90591 11305 90600 11339
rect 90548 11296 90600 11305
rect 74172 11228 74224 11280
rect 74356 11271 74408 11280
rect 74356 11237 74365 11271
rect 74365 11237 74399 11271
rect 74399 11237 74408 11271
rect 74356 11228 74408 11237
rect 68560 11135 68612 11144
rect 68560 11101 68569 11135
rect 68569 11101 68603 11135
rect 68603 11101 68612 11135
rect 68560 11092 68612 11101
rect 69204 11092 69256 11144
rect 69480 11092 69532 11144
rect 70676 11092 70728 11144
rect 71136 11135 71188 11144
rect 71136 11101 71145 11135
rect 71145 11101 71179 11135
rect 71179 11101 71188 11135
rect 71136 11092 71188 11101
rect 72792 11160 72844 11212
rect 75368 11160 75420 11212
rect 75736 11160 75788 11212
rect 76840 11160 76892 11212
rect 77760 11228 77812 11280
rect 78496 11228 78548 11280
rect 80704 11228 80756 11280
rect 77852 11203 77904 11212
rect 77852 11169 77861 11203
rect 77861 11169 77895 11203
rect 77895 11169 77904 11203
rect 77852 11160 77904 11169
rect 72332 11135 72384 11144
rect 72332 11101 72341 11135
rect 72341 11101 72375 11135
rect 72375 11101 72384 11135
rect 72332 11092 72384 11101
rect 73068 11092 73120 11144
rect 73620 11092 73672 11144
rect 73988 11092 74040 11144
rect 74356 11092 74408 11144
rect 75276 11135 75328 11144
rect 71872 11067 71924 11076
rect 71872 11033 71881 11067
rect 71881 11033 71915 11067
rect 71915 11033 71924 11067
rect 71872 11024 71924 11033
rect 75276 11101 75285 11135
rect 75285 11101 75319 11135
rect 75319 11101 75328 11135
rect 75276 11092 75328 11101
rect 76104 11092 76156 11144
rect 77208 11092 77260 11144
rect 77760 11135 77812 11144
rect 75184 11024 75236 11076
rect 75644 11024 75696 11076
rect 61476 10956 61528 11008
rect 67456 10956 67508 11008
rect 71044 10956 71096 11008
rect 71136 10999 71188 11008
rect 71136 10965 71145 10999
rect 71145 10965 71179 10999
rect 71179 10965 71188 10999
rect 77484 11024 77536 11076
rect 77760 11101 77769 11135
rect 77769 11101 77803 11135
rect 77803 11101 77812 11135
rect 80152 11160 80204 11212
rect 81164 11160 81216 11212
rect 81440 11160 81492 11212
rect 77760 11092 77812 11101
rect 78588 11092 78640 11144
rect 78680 11135 78732 11144
rect 78680 11101 78689 11135
rect 78689 11101 78723 11135
rect 78723 11101 78732 11135
rect 79600 11135 79652 11144
rect 78680 11092 78732 11101
rect 79600 11101 79609 11135
rect 79609 11101 79643 11135
rect 79643 11101 79652 11135
rect 79600 11092 79652 11101
rect 78864 11024 78916 11076
rect 79692 11024 79744 11076
rect 82544 11135 82596 11144
rect 82544 11101 82553 11135
rect 82553 11101 82587 11135
rect 82587 11101 82596 11135
rect 82544 11092 82596 11101
rect 84292 11228 84344 11280
rect 85764 11271 85816 11280
rect 85764 11237 85773 11271
rect 85773 11237 85807 11271
rect 85807 11237 85816 11271
rect 85764 11228 85816 11237
rect 85948 11228 86000 11280
rect 91836 11296 91888 11348
rect 92296 11296 92348 11348
rect 93308 11339 93360 11348
rect 93308 11305 93317 11339
rect 93317 11305 93351 11339
rect 93351 11305 93360 11339
rect 93308 11296 93360 11305
rect 83740 11160 83792 11212
rect 84016 11160 84068 11212
rect 84108 11160 84160 11212
rect 86224 11160 86276 11212
rect 86868 11160 86920 11212
rect 71136 10956 71188 10965
rect 77116 10956 77168 11008
rect 80428 10999 80480 11008
rect 80428 10965 80437 10999
rect 80437 10965 80471 10999
rect 80471 10965 80480 10999
rect 80428 10956 80480 10965
rect 82176 11024 82228 11076
rect 84016 11067 84068 11076
rect 84016 11033 84025 11067
rect 84025 11033 84059 11067
rect 84059 11033 84068 11067
rect 84016 11024 84068 11033
rect 86040 11092 86092 11144
rect 86592 11024 86644 11076
rect 90456 11135 90508 11144
rect 90456 11101 90465 11135
rect 90465 11101 90499 11135
rect 90499 11101 90508 11135
rect 90456 11092 90508 11101
rect 93768 11135 93820 11144
rect 88156 11024 88208 11076
rect 89628 11024 89680 11076
rect 93768 11101 93777 11135
rect 93777 11101 93811 11135
rect 93811 11101 93820 11135
rect 93768 11092 93820 11101
rect 94228 11024 94280 11076
rect 84108 10956 84160 11008
rect 84292 10956 84344 11008
rect 86868 10956 86920 11008
rect 89904 10999 89956 11008
rect 89904 10965 89913 10999
rect 89913 10965 89947 10999
rect 89947 10965 89956 10999
rect 89904 10956 89956 10965
rect 92480 10956 92532 11008
rect 93768 10956 93820 11008
rect 24386 10854 24438 10906
rect 24450 10854 24502 10906
rect 24514 10854 24566 10906
rect 24578 10854 24630 10906
rect 24642 10854 24694 10906
rect 47823 10854 47875 10906
rect 47887 10854 47939 10906
rect 47951 10854 48003 10906
rect 48015 10854 48067 10906
rect 48079 10854 48131 10906
rect 71260 10854 71312 10906
rect 71324 10854 71376 10906
rect 71388 10854 71440 10906
rect 71452 10854 71504 10906
rect 71516 10854 71568 10906
rect 94697 10854 94749 10906
rect 94761 10854 94813 10906
rect 94825 10854 94877 10906
rect 94889 10854 94941 10906
rect 94953 10854 95005 10906
rect 1768 10795 1820 10804
rect 1768 10761 1777 10795
rect 1777 10761 1811 10795
rect 1811 10761 1820 10795
rect 1768 10752 1820 10761
rect 4988 10752 5040 10804
rect 3976 10684 4028 10736
rect 4528 10659 4580 10668
rect 4528 10625 4537 10659
rect 4537 10625 4571 10659
rect 4571 10625 4580 10659
rect 4528 10616 4580 10625
rect 8024 10752 8076 10804
rect 10140 10752 10192 10804
rect 11152 10795 11204 10804
rect 11152 10761 11161 10795
rect 11161 10761 11195 10795
rect 11195 10761 11204 10795
rect 11152 10752 11204 10761
rect 12256 10795 12308 10804
rect 12256 10761 12265 10795
rect 12265 10761 12299 10795
rect 12299 10761 12308 10795
rect 12256 10752 12308 10761
rect 7104 10684 7156 10736
rect 12992 10727 13044 10736
rect 6736 10659 6788 10668
rect 2320 10591 2372 10600
rect 2320 10557 2329 10591
rect 2329 10557 2363 10591
rect 2363 10557 2372 10591
rect 2320 10548 2372 10557
rect 6736 10625 6745 10659
rect 6745 10625 6779 10659
rect 6779 10625 6788 10659
rect 7472 10659 7524 10668
rect 6736 10616 6788 10625
rect 4804 10591 4856 10600
rect 4804 10557 4813 10591
rect 4813 10557 4847 10591
rect 4847 10557 4856 10591
rect 4804 10548 4856 10557
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 8852 10616 8904 10668
rect 12992 10693 13001 10727
rect 13001 10693 13035 10727
rect 13035 10693 13044 10727
rect 12992 10684 13044 10693
rect 14832 10684 14884 10736
rect 15200 10795 15252 10804
rect 15200 10761 15230 10795
rect 15230 10761 15252 10795
rect 15384 10795 15436 10804
rect 15200 10752 15252 10761
rect 15384 10761 15393 10795
rect 15393 10761 15427 10795
rect 15427 10761 15436 10795
rect 15384 10752 15436 10761
rect 18236 10752 18288 10804
rect 18788 10752 18840 10804
rect 24308 10752 24360 10804
rect 24492 10752 24544 10804
rect 15476 10684 15528 10736
rect 16764 10684 16816 10736
rect 20996 10684 21048 10736
rect 21272 10727 21324 10736
rect 21272 10693 21281 10727
rect 21281 10693 21315 10727
rect 21315 10693 21324 10727
rect 21272 10684 21324 10693
rect 22744 10684 22796 10736
rect 11060 10616 11112 10668
rect 12072 10616 12124 10668
rect 14096 10616 14148 10668
rect 12164 10548 12216 10600
rect 5448 10480 5500 10532
rect 7104 10480 7156 10532
rect 10968 10480 11020 10532
rect 11152 10480 11204 10532
rect 11888 10480 11940 10532
rect 6644 10455 6696 10464
rect 6644 10421 6653 10455
rect 6653 10421 6687 10455
rect 6687 10421 6696 10455
rect 6644 10412 6696 10421
rect 7472 10412 7524 10464
rect 8116 10412 8168 10464
rect 12532 10548 12584 10600
rect 16488 10616 16540 10668
rect 18052 10659 18104 10668
rect 18052 10625 18061 10659
rect 18061 10625 18095 10659
rect 18095 10625 18104 10659
rect 18052 10616 18104 10625
rect 15936 10548 15988 10600
rect 16120 10548 16172 10600
rect 17960 10548 18012 10600
rect 18328 10616 18380 10668
rect 19064 10659 19116 10668
rect 18604 10548 18656 10600
rect 19064 10625 19073 10659
rect 19073 10625 19107 10659
rect 19107 10625 19116 10659
rect 19064 10616 19116 10625
rect 19708 10659 19760 10668
rect 19708 10625 19717 10659
rect 19717 10625 19751 10659
rect 19751 10625 19760 10659
rect 19708 10616 19760 10625
rect 19892 10548 19944 10600
rect 19984 10548 20036 10600
rect 24952 10684 25004 10736
rect 25136 10684 25188 10736
rect 27528 10684 27580 10736
rect 28908 10752 28960 10804
rect 31208 10795 31260 10804
rect 29000 10684 29052 10736
rect 31208 10761 31217 10795
rect 31217 10761 31251 10795
rect 31251 10761 31260 10795
rect 37464 10795 37516 10804
rect 31208 10752 31260 10761
rect 31300 10684 31352 10736
rect 27436 10616 27488 10668
rect 27712 10659 27764 10668
rect 27712 10625 27721 10659
rect 27721 10625 27755 10659
rect 27755 10625 27764 10659
rect 27712 10616 27764 10625
rect 29644 10616 29696 10668
rect 30288 10616 30340 10668
rect 24860 10591 24912 10600
rect 16764 10480 16816 10532
rect 12992 10412 13044 10464
rect 13636 10412 13688 10464
rect 18144 10412 18196 10464
rect 19248 10412 19300 10464
rect 24492 10480 24544 10532
rect 23756 10455 23808 10464
rect 23756 10421 23765 10455
rect 23765 10421 23799 10455
rect 23799 10421 23808 10455
rect 23756 10412 23808 10421
rect 24860 10557 24869 10591
rect 24869 10557 24903 10591
rect 24903 10557 24912 10591
rect 24860 10548 24912 10557
rect 24952 10548 25004 10600
rect 31852 10616 31904 10668
rect 31944 10616 31996 10668
rect 32772 10616 32824 10668
rect 31484 10548 31536 10600
rect 32680 10591 32732 10600
rect 32680 10557 32689 10591
rect 32689 10557 32723 10591
rect 32723 10557 32732 10591
rect 32680 10548 32732 10557
rect 33508 10684 33560 10736
rect 35624 10684 35676 10736
rect 33692 10659 33744 10668
rect 33692 10625 33701 10659
rect 33701 10625 33735 10659
rect 33735 10625 33744 10659
rect 33692 10616 33744 10625
rect 37464 10761 37473 10795
rect 37473 10761 37507 10795
rect 37507 10761 37516 10795
rect 37464 10752 37516 10761
rect 37556 10752 37608 10804
rect 40132 10684 40184 10736
rect 41144 10684 41196 10736
rect 36636 10659 36688 10668
rect 36636 10625 36645 10659
rect 36645 10625 36679 10659
rect 36679 10625 36688 10659
rect 36636 10616 36688 10625
rect 37372 10616 37424 10668
rect 38200 10616 38252 10668
rect 38292 10616 38344 10668
rect 38752 10616 38804 10668
rect 38844 10659 38896 10668
rect 38844 10625 38867 10659
rect 38867 10625 38896 10659
rect 38844 10616 38896 10625
rect 34520 10548 34572 10600
rect 35716 10548 35768 10600
rect 29736 10480 29788 10532
rect 31852 10480 31904 10532
rect 32956 10523 33008 10532
rect 32956 10489 32965 10523
rect 32965 10489 32999 10523
rect 32999 10489 33008 10523
rect 32956 10480 33008 10489
rect 33692 10480 33744 10532
rect 36820 10480 36872 10532
rect 37096 10480 37148 10532
rect 40040 10616 40092 10668
rect 41604 10684 41656 10736
rect 42524 10752 42576 10804
rect 44272 10752 44324 10804
rect 48320 10795 48372 10804
rect 44916 10727 44968 10736
rect 39672 10591 39724 10600
rect 39672 10557 39681 10591
rect 39681 10557 39715 10591
rect 39715 10557 39724 10591
rect 39672 10548 39724 10557
rect 39764 10548 39816 10600
rect 42432 10616 42484 10668
rect 42800 10659 42852 10668
rect 42800 10625 42809 10659
rect 42809 10625 42843 10659
rect 42843 10625 42852 10659
rect 42800 10616 42852 10625
rect 44916 10693 44925 10727
rect 44925 10693 44959 10727
rect 44959 10693 44968 10727
rect 44916 10684 44968 10693
rect 48320 10761 48329 10795
rect 48329 10761 48363 10795
rect 48363 10761 48372 10795
rect 48320 10752 48372 10761
rect 48412 10684 48464 10736
rect 50068 10752 50120 10804
rect 50160 10752 50212 10804
rect 62488 10752 62540 10804
rect 62764 10752 62816 10804
rect 44456 10616 44508 10668
rect 48504 10659 48556 10668
rect 48504 10625 48513 10659
rect 48513 10625 48547 10659
rect 48547 10625 48556 10659
rect 48504 10616 48556 10625
rect 50804 10684 50856 10736
rect 54024 10684 54076 10736
rect 54208 10727 54260 10736
rect 54208 10693 54217 10727
rect 54217 10693 54251 10727
rect 54251 10693 54260 10727
rect 54208 10684 54260 10693
rect 54392 10684 54444 10736
rect 41880 10548 41932 10600
rect 42708 10548 42760 10600
rect 42892 10591 42944 10600
rect 42892 10557 42901 10591
rect 42901 10557 42935 10591
rect 42935 10557 42944 10591
rect 42892 10548 42944 10557
rect 43260 10548 43312 10600
rect 43904 10591 43956 10600
rect 43904 10557 43913 10591
rect 43913 10557 43947 10591
rect 43947 10557 43956 10591
rect 43904 10548 43956 10557
rect 45192 10591 45244 10600
rect 45192 10557 45201 10591
rect 45201 10557 45235 10591
rect 45235 10557 45244 10591
rect 45192 10548 45244 10557
rect 48780 10523 48832 10532
rect 48780 10489 48789 10523
rect 48789 10489 48823 10523
rect 48823 10489 48832 10523
rect 49700 10548 49752 10600
rect 50344 10616 50396 10668
rect 50436 10591 50488 10600
rect 50436 10557 50445 10591
rect 50445 10557 50479 10591
rect 50479 10557 50488 10591
rect 50436 10548 50488 10557
rect 50712 10591 50764 10600
rect 50712 10557 50721 10591
rect 50721 10557 50755 10591
rect 50755 10557 50764 10591
rect 50712 10548 50764 10557
rect 53104 10548 53156 10600
rect 53288 10659 53340 10668
rect 53288 10625 53297 10659
rect 53297 10625 53331 10659
rect 53331 10625 53340 10659
rect 53472 10659 53524 10668
rect 53288 10616 53340 10625
rect 53472 10625 53481 10659
rect 53481 10625 53515 10659
rect 53515 10625 53524 10659
rect 53472 10616 53524 10625
rect 53564 10616 53616 10668
rect 53748 10616 53800 10668
rect 48780 10480 48832 10489
rect 25872 10412 25924 10464
rect 26700 10412 26752 10464
rect 27528 10412 27580 10464
rect 28080 10412 28132 10464
rect 31208 10412 31260 10464
rect 33048 10412 33100 10464
rect 35716 10412 35768 10464
rect 37280 10412 37332 10464
rect 37372 10412 37424 10464
rect 41880 10412 41932 10464
rect 41972 10412 42024 10464
rect 45192 10412 45244 10464
rect 48320 10412 48372 10464
rect 49884 10412 49936 10464
rect 50068 10412 50120 10464
rect 53380 10523 53432 10532
rect 53380 10489 53389 10523
rect 53389 10489 53423 10523
rect 53423 10489 53432 10523
rect 53380 10480 53432 10489
rect 54208 10480 54260 10532
rect 54484 10616 54536 10668
rect 54944 10659 54996 10668
rect 54944 10625 54953 10659
rect 54953 10625 54987 10659
rect 54987 10625 54996 10659
rect 54944 10616 54996 10625
rect 55772 10659 55824 10668
rect 55772 10625 55781 10659
rect 55781 10625 55815 10659
rect 55815 10625 55824 10659
rect 55772 10616 55824 10625
rect 56600 10684 56652 10736
rect 57796 10684 57848 10736
rect 58808 10684 58860 10736
rect 59636 10684 59688 10736
rect 61660 10684 61712 10736
rect 56508 10659 56560 10668
rect 56508 10625 56517 10659
rect 56517 10625 56551 10659
rect 56551 10625 56560 10659
rect 56508 10616 56560 10625
rect 57336 10659 57388 10668
rect 57336 10625 57345 10659
rect 57345 10625 57379 10659
rect 57379 10625 57388 10659
rect 57336 10616 57388 10625
rect 54576 10548 54628 10600
rect 55496 10548 55548 10600
rect 57428 10591 57480 10600
rect 52184 10455 52236 10464
rect 52184 10421 52193 10455
rect 52193 10421 52227 10455
rect 52227 10421 52236 10455
rect 52184 10412 52236 10421
rect 52276 10412 52328 10464
rect 55312 10455 55364 10464
rect 55312 10421 55321 10455
rect 55321 10421 55355 10455
rect 55355 10421 55364 10455
rect 55312 10412 55364 10421
rect 56324 10480 56376 10532
rect 57428 10557 57437 10591
rect 57437 10557 57471 10591
rect 57471 10557 57480 10591
rect 57428 10548 57480 10557
rect 61568 10591 61620 10600
rect 61568 10557 61577 10591
rect 61577 10557 61611 10591
rect 61611 10557 61620 10591
rect 61568 10548 61620 10557
rect 62120 10591 62172 10600
rect 62120 10557 62129 10591
rect 62129 10557 62163 10591
rect 62163 10557 62172 10591
rect 62120 10548 62172 10557
rect 61936 10480 61988 10532
rect 62672 10684 62724 10736
rect 63224 10659 63276 10668
rect 63224 10625 63233 10659
rect 63233 10625 63267 10659
rect 63267 10625 63276 10659
rect 63224 10616 63276 10625
rect 65432 10727 65484 10736
rect 65432 10693 65441 10727
rect 65441 10693 65475 10727
rect 65475 10693 65484 10727
rect 65432 10684 65484 10693
rect 69664 10752 69716 10804
rect 68744 10684 68796 10736
rect 70308 10684 70360 10736
rect 71044 10752 71096 10804
rect 79508 10752 79560 10804
rect 70676 10684 70728 10736
rect 72240 10684 72292 10736
rect 73528 10684 73580 10736
rect 76012 10684 76064 10736
rect 80428 10752 80480 10804
rect 82268 10752 82320 10804
rect 92112 10752 92164 10804
rect 94228 10795 94280 10804
rect 94228 10761 94237 10795
rect 94237 10761 94271 10795
rect 94271 10761 94280 10795
rect 94228 10752 94280 10761
rect 81348 10684 81400 10736
rect 67732 10616 67784 10668
rect 68284 10616 68336 10668
rect 62396 10548 62448 10600
rect 63132 10480 63184 10532
rect 67364 10548 67416 10600
rect 68376 10591 68428 10600
rect 68376 10557 68385 10591
rect 68385 10557 68419 10591
rect 68419 10557 68428 10591
rect 68376 10548 68428 10557
rect 68652 10591 68704 10600
rect 68652 10557 68661 10591
rect 68661 10557 68695 10591
rect 68695 10557 68704 10591
rect 68652 10548 68704 10557
rect 68744 10548 68796 10600
rect 71780 10616 71832 10668
rect 74080 10616 74132 10668
rect 76748 10616 76800 10668
rect 77116 10616 77168 10668
rect 78496 10616 78548 10668
rect 78864 10616 78916 10668
rect 70400 10548 70452 10600
rect 74448 10548 74500 10600
rect 66076 10480 66128 10532
rect 59084 10412 59136 10464
rect 63316 10412 63368 10464
rect 63868 10412 63920 10464
rect 69664 10480 69716 10532
rect 73528 10480 73580 10532
rect 67640 10412 67692 10464
rect 67824 10412 67876 10464
rect 70492 10412 70544 10464
rect 72976 10412 73028 10464
rect 74172 10455 74224 10464
rect 74172 10421 74181 10455
rect 74181 10421 74215 10455
rect 74215 10421 74224 10455
rect 74172 10412 74224 10421
rect 77944 10480 77996 10532
rect 78772 10480 78824 10532
rect 76932 10455 76984 10464
rect 76932 10421 76941 10455
rect 76941 10421 76975 10455
rect 76975 10421 76984 10455
rect 76932 10412 76984 10421
rect 77576 10412 77628 10464
rect 79600 10548 79652 10600
rect 82268 10659 82320 10668
rect 82268 10625 82277 10659
rect 82277 10625 82311 10659
rect 82311 10625 82320 10659
rect 82268 10616 82320 10625
rect 83372 10616 83424 10668
rect 83556 10616 83608 10668
rect 84016 10548 84068 10600
rect 84200 10659 84252 10668
rect 84200 10625 84209 10659
rect 84209 10625 84243 10659
rect 84243 10625 84252 10659
rect 84660 10659 84712 10668
rect 84200 10616 84252 10625
rect 84660 10625 84669 10659
rect 84669 10625 84703 10659
rect 84703 10625 84712 10659
rect 84660 10616 84712 10625
rect 89904 10684 89956 10736
rect 90640 10684 90692 10736
rect 88984 10616 89036 10668
rect 89168 10659 89220 10668
rect 89168 10625 89177 10659
rect 89177 10625 89211 10659
rect 89211 10625 89220 10659
rect 89168 10616 89220 10625
rect 93308 10616 93360 10668
rect 94136 10659 94188 10668
rect 94136 10625 94145 10659
rect 94145 10625 94179 10659
rect 94179 10625 94188 10659
rect 94136 10616 94188 10625
rect 84292 10548 84344 10600
rect 84568 10548 84620 10600
rect 86500 10548 86552 10600
rect 90732 10548 90784 10600
rect 92480 10591 92532 10600
rect 92480 10557 92489 10591
rect 92489 10557 92523 10591
rect 92523 10557 92532 10591
rect 92480 10548 92532 10557
rect 93216 10591 93268 10600
rect 93216 10557 93225 10591
rect 93225 10557 93259 10591
rect 93259 10557 93268 10591
rect 93216 10548 93268 10557
rect 82360 10412 82412 10464
rect 84844 10480 84896 10532
rect 84752 10455 84804 10464
rect 84752 10421 84761 10455
rect 84761 10421 84795 10455
rect 84795 10421 84804 10455
rect 84752 10412 84804 10421
rect 85304 10455 85356 10464
rect 85304 10421 85313 10455
rect 85313 10421 85347 10455
rect 85347 10421 85356 10455
rect 85304 10412 85356 10421
rect 12668 10310 12720 10362
rect 12732 10310 12784 10362
rect 12796 10310 12848 10362
rect 12860 10310 12912 10362
rect 12924 10310 12976 10362
rect 36105 10310 36157 10362
rect 36169 10310 36221 10362
rect 36233 10310 36285 10362
rect 36297 10310 36349 10362
rect 36361 10310 36413 10362
rect 59542 10310 59594 10362
rect 59606 10310 59658 10362
rect 59670 10310 59722 10362
rect 59734 10310 59786 10362
rect 59798 10310 59850 10362
rect 82979 10310 83031 10362
rect 83043 10310 83095 10362
rect 83107 10310 83159 10362
rect 83171 10310 83223 10362
rect 83235 10310 83287 10362
rect 4528 10208 4580 10260
rect 3424 10183 3476 10192
rect 3424 10149 3433 10183
rect 3433 10149 3467 10183
rect 3467 10149 3476 10183
rect 3424 10140 3476 10149
rect 4068 10183 4120 10192
rect 4068 10149 4077 10183
rect 4077 10149 4111 10183
rect 4111 10149 4120 10183
rect 4068 10140 4120 10149
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 2228 10047 2280 10056
rect 2228 10013 2237 10047
rect 2237 10013 2271 10047
rect 2271 10013 2280 10047
rect 2228 10004 2280 10013
rect 2504 10047 2556 10056
rect 2504 10013 2513 10047
rect 2513 10013 2547 10047
rect 2547 10013 2556 10047
rect 2504 10004 2556 10013
rect 3884 10004 3936 10056
rect 4528 10072 4580 10124
rect 5080 10208 5132 10260
rect 11796 10251 11848 10260
rect 6644 10072 6696 10124
rect 11796 10217 11805 10251
rect 11805 10217 11839 10251
rect 11839 10217 11848 10251
rect 11796 10208 11848 10217
rect 12532 10072 12584 10124
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 13544 10072 13596 10081
rect 15108 10115 15160 10124
rect 15108 10081 15117 10115
rect 15117 10081 15151 10115
rect 15151 10081 15160 10115
rect 15108 10072 15160 10081
rect 4620 10047 4672 10056
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 4620 10004 4672 10013
rect 6000 10004 6052 10056
rect 6736 9936 6788 9988
rect 7656 10004 7708 10056
rect 8024 10047 8076 10056
rect 8024 10013 8033 10047
rect 8033 10013 8067 10047
rect 8067 10013 8076 10047
rect 8024 10004 8076 10013
rect 8116 10004 8168 10056
rect 8300 10047 8352 10056
rect 8300 10013 8309 10047
rect 8309 10013 8343 10047
rect 8343 10013 8352 10047
rect 8300 10004 8352 10013
rect 11060 10004 11112 10056
rect 11980 10004 12032 10056
rect 13820 10004 13872 10056
rect 18696 10208 18748 10260
rect 20720 10208 20772 10260
rect 22560 10251 22612 10260
rect 22560 10217 22569 10251
rect 22569 10217 22603 10251
rect 22603 10217 22612 10251
rect 22560 10208 22612 10217
rect 23756 10208 23808 10260
rect 30380 10208 30432 10260
rect 33692 10208 33744 10260
rect 34336 10208 34388 10260
rect 35164 10208 35216 10260
rect 36544 10251 36596 10260
rect 36544 10217 36553 10251
rect 36553 10217 36587 10251
rect 36587 10217 36596 10251
rect 36544 10208 36596 10217
rect 18052 10140 18104 10192
rect 19064 10140 19116 10192
rect 26792 10140 26844 10192
rect 29092 10183 29144 10192
rect 17960 10072 18012 10124
rect 19156 10072 19208 10124
rect 19984 10115 20036 10124
rect 19984 10081 19993 10115
rect 19993 10081 20027 10115
rect 20027 10081 20036 10115
rect 19984 10072 20036 10081
rect 22008 10115 22060 10124
rect 19708 10004 19760 10056
rect 22008 10081 22017 10115
rect 22017 10081 22051 10115
rect 22051 10081 22060 10115
rect 22008 10072 22060 10081
rect 25780 10072 25832 10124
rect 29092 10149 29101 10183
rect 29101 10149 29135 10183
rect 29135 10149 29144 10183
rect 29092 10140 29144 10149
rect 29644 10072 29696 10124
rect 33140 10140 33192 10192
rect 35072 10140 35124 10192
rect 36452 10140 36504 10192
rect 32496 10072 32548 10124
rect 35716 10072 35768 10124
rect 41880 10208 41932 10260
rect 42064 10208 42116 10260
rect 43904 10208 43956 10260
rect 44456 10251 44508 10260
rect 44456 10217 44465 10251
rect 44465 10217 44499 10251
rect 44499 10217 44508 10251
rect 44456 10208 44508 10217
rect 47032 10251 47084 10260
rect 47032 10217 47041 10251
rect 47041 10217 47075 10251
rect 47075 10217 47084 10251
rect 47032 10208 47084 10217
rect 47584 10208 47636 10260
rect 49700 10208 49752 10260
rect 50712 10208 50764 10260
rect 50804 10208 50856 10260
rect 53288 10208 53340 10260
rect 53472 10251 53524 10260
rect 53472 10217 53481 10251
rect 53481 10217 53515 10251
rect 53515 10217 53524 10251
rect 53472 10208 53524 10217
rect 53656 10208 53708 10260
rect 54024 10208 54076 10260
rect 54576 10208 54628 10260
rect 40224 10140 40276 10192
rect 41788 10140 41840 10192
rect 42432 10140 42484 10192
rect 44916 10140 44968 10192
rect 22560 10004 22612 10056
rect 22652 10004 22704 10056
rect 27436 10047 27488 10056
rect 8852 9936 8904 9988
rect 3976 9868 4028 9920
rect 6920 9868 6972 9920
rect 7840 9868 7892 9920
rect 8944 9868 8996 9920
rect 9404 9868 9456 9920
rect 9772 9911 9824 9920
rect 9772 9877 9781 9911
rect 9781 9877 9815 9911
rect 9815 9877 9824 9911
rect 9772 9868 9824 9877
rect 10508 9911 10560 9920
rect 10508 9877 10517 9911
rect 10517 9877 10551 9911
rect 10551 9877 10560 9911
rect 10508 9868 10560 9877
rect 10968 9868 11020 9920
rect 13912 9936 13964 9988
rect 18052 9936 18104 9988
rect 22468 9936 22520 9988
rect 22836 9936 22888 9988
rect 24676 9979 24728 9988
rect 24676 9945 24685 9979
rect 24685 9945 24719 9979
rect 24719 9945 24728 9979
rect 24676 9936 24728 9945
rect 27436 10013 27445 10047
rect 27445 10013 27479 10047
rect 27479 10013 27488 10047
rect 27436 10004 27488 10013
rect 29828 10004 29880 10056
rect 29920 10004 29972 10056
rect 33140 10004 33192 10056
rect 36544 10004 36596 10056
rect 36728 10047 36780 10056
rect 36728 10013 36751 10047
rect 36751 10013 36780 10047
rect 38568 10047 38620 10056
rect 36728 10004 36780 10013
rect 38568 10013 38577 10047
rect 38577 10013 38611 10047
rect 38611 10013 38620 10047
rect 38568 10004 38620 10013
rect 13544 9868 13596 9920
rect 15384 9868 15436 9920
rect 16396 9868 16448 9920
rect 18328 9868 18380 9920
rect 18604 9911 18656 9920
rect 18604 9877 18613 9911
rect 18613 9877 18647 9911
rect 18647 9877 18656 9911
rect 18604 9868 18656 9877
rect 19064 9868 19116 9920
rect 23388 9868 23440 9920
rect 24584 9868 24636 9920
rect 27988 9979 28040 9988
rect 27988 9945 27997 9979
rect 27997 9945 28031 9979
rect 28031 9945 28040 9979
rect 27988 9936 28040 9945
rect 32772 9936 32824 9988
rect 33416 9936 33468 9988
rect 25320 9868 25372 9920
rect 26056 9868 26108 9920
rect 29000 9868 29052 9920
rect 33140 9868 33192 9920
rect 34612 9868 34664 9920
rect 35164 9936 35216 9988
rect 39948 10004 40000 10056
rect 35992 9911 36044 9920
rect 35992 9877 36001 9911
rect 36001 9877 36035 9911
rect 36035 9877 36044 9911
rect 35992 9868 36044 9877
rect 39764 9936 39816 9988
rect 40316 10047 40368 10056
rect 40316 10013 40325 10047
rect 40325 10013 40359 10047
rect 40359 10013 40368 10047
rect 41144 10047 41196 10056
rect 40316 10004 40368 10013
rect 41144 10013 41153 10047
rect 41153 10013 41187 10047
rect 41187 10013 41196 10047
rect 41144 10004 41196 10013
rect 40592 9936 40644 9988
rect 41236 9936 41288 9988
rect 39856 9868 39908 9920
rect 40224 9868 40276 9920
rect 40316 9868 40368 9920
rect 41972 10004 42024 10056
rect 43352 10072 43404 10124
rect 44548 10072 44600 10124
rect 44732 10072 44784 10124
rect 42616 10047 42668 10056
rect 42616 10013 42625 10047
rect 42625 10013 42659 10047
rect 42659 10013 42668 10047
rect 42616 10004 42668 10013
rect 43536 10047 43588 10056
rect 43536 10013 43545 10047
rect 43545 10013 43579 10047
rect 43579 10013 43588 10047
rect 43812 10047 43864 10056
rect 43536 10004 43588 10013
rect 43812 10013 43821 10047
rect 43821 10013 43855 10047
rect 43855 10013 43864 10047
rect 43812 10004 43864 10013
rect 44364 10004 44416 10056
rect 41788 9979 41840 9988
rect 41788 9945 41797 9979
rect 41797 9945 41831 9979
rect 41831 9945 41840 9979
rect 41788 9936 41840 9945
rect 44824 10004 44876 10056
rect 46112 10004 46164 10056
rect 46296 10047 46348 10056
rect 46296 10013 46305 10047
rect 46305 10013 46339 10047
rect 46339 10013 46348 10047
rect 46296 10004 46348 10013
rect 48780 10140 48832 10192
rect 49884 10140 49936 10192
rect 54760 10140 54812 10192
rect 54852 10140 54904 10192
rect 56600 10140 56652 10192
rect 57336 10208 57388 10260
rect 60740 10208 60792 10260
rect 62672 10251 62724 10260
rect 62672 10217 62681 10251
rect 62681 10217 62715 10251
rect 62715 10217 62724 10251
rect 62672 10208 62724 10217
rect 63316 10251 63368 10260
rect 63316 10217 63325 10251
rect 63325 10217 63359 10251
rect 63359 10217 63368 10251
rect 63316 10208 63368 10217
rect 67456 10251 67508 10260
rect 67456 10217 67465 10251
rect 67465 10217 67499 10251
rect 67499 10217 67508 10251
rect 67456 10208 67508 10217
rect 68652 10208 68704 10260
rect 60372 10140 60424 10192
rect 60464 10140 60516 10192
rect 65432 10140 65484 10192
rect 49608 10072 49660 10124
rect 52276 10072 52328 10124
rect 53288 10072 53340 10124
rect 53656 10072 53708 10124
rect 56968 10115 57020 10124
rect 56968 10081 56977 10115
rect 56977 10081 57011 10115
rect 57011 10081 57020 10115
rect 56968 10072 57020 10081
rect 59360 10115 59412 10124
rect 59360 10081 59369 10115
rect 59369 10081 59403 10115
rect 59403 10081 59412 10115
rect 59360 10072 59412 10081
rect 48780 10047 48832 10056
rect 44916 9936 44968 9988
rect 48780 10013 48789 10047
rect 48789 10013 48823 10047
rect 48823 10013 48832 10047
rect 48780 10004 48832 10013
rect 49240 10004 49292 10056
rect 49516 10004 49568 10056
rect 49792 10047 49844 10056
rect 49792 10013 49801 10047
rect 49801 10013 49835 10047
rect 49835 10013 49844 10047
rect 49792 10004 49844 10013
rect 50252 10004 50304 10056
rect 53380 10004 53432 10056
rect 46572 9936 46624 9988
rect 49424 9936 49476 9988
rect 50804 9936 50856 9988
rect 51264 9936 51316 9988
rect 52552 9979 52604 9988
rect 52552 9945 52561 9979
rect 52561 9945 52595 9979
rect 52595 9945 52604 9979
rect 52552 9936 52604 9945
rect 53012 9936 53064 9988
rect 53748 10004 53800 10056
rect 41972 9911 42024 9920
rect 41972 9877 41997 9911
rect 41997 9877 42024 9911
rect 41972 9868 42024 9877
rect 42616 9868 42668 9920
rect 42708 9868 42760 9920
rect 43904 9868 43956 9920
rect 49332 9868 49384 9920
rect 55680 10004 55732 10056
rect 55864 10047 55916 10056
rect 55864 10013 55873 10047
rect 55873 10013 55907 10047
rect 55907 10013 55916 10047
rect 55864 10004 55916 10013
rect 56784 10047 56836 10056
rect 56784 10013 56793 10047
rect 56793 10013 56827 10047
rect 56827 10013 56836 10047
rect 56784 10004 56836 10013
rect 62396 10072 62448 10124
rect 62488 10072 62540 10124
rect 63408 10072 63460 10124
rect 67824 10140 67876 10192
rect 71688 10208 71740 10260
rect 72240 10208 72292 10260
rect 74172 10208 74224 10260
rect 75920 10208 75972 10260
rect 61108 10047 61160 10056
rect 58624 9979 58676 9988
rect 58624 9945 58633 9979
rect 58633 9945 58667 9979
rect 58667 9945 58676 9979
rect 58624 9936 58676 9945
rect 58900 9936 58952 9988
rect 61108 10013 61117 10047
rect 61117 10013 61151 10047
rect 61151 10013 61160 10047
rect 61108 10004 61160 10013
rect 54484 9868 54536 9920
rect 54852 9868 54904 9920
rect 55496 9911 55548 9920
rect 55496 9877 55505 9911
rect 55505 9877 55539 9911
rect 55539 9877 55548 9911
rect 55496 9868 55548 9877
rect 57796 9868 57848 9920
rect 60372 9868 60424 9920
rect 60464 9868 60516 9920
rect 62764 10004 62816 10056
rect 63684 10004 63736 10056
rect 64696 9979 64748 9988
rect 61936 9868 61988 9920
rect 63500 9868 63552 9920
rect 64696 9945 64705 9979
rect 64705 9945 64739 9979
rect 64739 9945 64748 9979
rect 64696 9936 64748 9945
rect 66628 9936 66680 9988
rect 65432 9868 65484 9920
rect 67364 10004 67416 10056
rect 68376 10004 68428 10056
rect 69664 10072 69716 10124
rect 70124 10072 70176 10124
rect 71688 10072 71740 10124
rect 77116 10208 77168 10260
rect 81348 10251 81400 10260
rect 81348 10217 81357 10251
rect 81357 10217 81391 10251
rect 81391 10217 81400 10251
rect 81348 10208 81400 10217
rect 78680 10140 78732 10192
rect 85304 10208 85356 10260
rect 85396 10208 85448 10260
rect 90640 10208 90692 10260
rect 87880 10140 87932 10192
rect 79784 10115 79836 10124
rect 79784 10081 79793 10115
rect 79793 10081 79827 10115
rect 79827 10081 79836 10115
rect 79784 10072 79836 10081
rect 80796 10072 80848 10124
rect 81716 10072 81768 10124
rect 83372 10072 83424 10124
rect 84752 10072 84804 10124
rect 85488 10072 85540 10124
rect 70676 10004 70728 10056
rect 70952 10047 71004 10056
rect 70952 10013 70961 10047
rect 70961 10013 70995 10047
rect 70995 10013 71004 10047
rect 70952 10004 71004 10013
rect 72976 10004 73028 10056
rect 73160 10047 73212 10056
rect 73160 10013 73169 10047
rect 73169 10013 73203 10047
rect 73203 10013 73212 10047
rect 73160 10004 73212 10013
rect 75920 10004 75972 10056
rect 76104 10047 76156 10056
rect 76104 10013 76113 10047
rect 76113 10013 76147 10047
rect 76147 10013 76156 10047
rect 76104 10004 76156 10013
rect 77668 10004 77720 10056
rect 79140 10047 79192 10056
rect 79140 10013 79149 10047
rect 79149 10013 79183 10047
rect 79183 10013 79192 10047
rect 79140 10004 79192 10013
rect 79968 10047 80020 10056
rect 79968 10013 79997 10047
rect 79997 10013 80020 10047
rect 79968 10004 80020 10013
rect 68468 9936 68520 9988
rect 68836 9868 68888 9920
rect 70860 9936 70912 9988
rect 73436 9979 73488 9988
rect 73436 9945 73445 9979
rect 73445 9945 73479 9979
rect 73479 9945 73488 9979
rect 73436 9936 73488 9945
rect 75276 9936 75328 9988
rect 71596 9868 71648 9920
rect 74816 9868 74868 9920
rect 77392 9936 77444 9988
rect 77760 9936 77812 9988
rect 82360 10004 82412 10056
rect 84200 10047 84252 10056
rect 84200 10013 84209 10047
rect 84209 10013 84243 10047
rect 84243 10013 84252 10047
rect 84844 10047 84896 10056
rect 84200 10004 84252 10013
rect 84844 10013 84853 10047
rect 84853 10013 84887 10047
rect 84887 10013 84896 10047
rect 84844 10004 84896 10013
rect 85764 10047 85816 10056
rect 85764 10013 85773 10047
rect 85773 10013 85807 10047
rect 85807 10013 85816 10047
rect 85764 10004 85816 10013
rect 86408 10047 86460 10056
rect 86408 10013 86417 10047
rect 86417 10013 86451 10047
rect 86451 10013 86460 10047
rect 86408 10004 86460 10013
rect 87788 10004 87840 10056
rect 88524 10004 88576 10056
rect 93860 10072 93912 10124
rect 89812 10047 89864 10056
rect 89812 10013 89821 10047
rect 89821 10013 89855 10047
rect 89855 10013 89864 10047
rect 89812 10004 89864 10013
rect 90456 10004 90508 10056
rect 94136 10004 94188 10056
rect 83832 9936 83884 9988
rect 90732 9936 90784 9988
rect 91100 9936 91152 9988
rect 94228 9936 94280 9988
rect 77668 9868 77720 9920
rect 78128 9868 78180 9920
rect 79048 9868 79100 9920
rect 79416 9868 79468 9920
rect 80244 9911 80296 9920
rect 80244 9877 80253 9911
rect 80253 9877 80287 9911
rect 80287 9877 80296 9911
rect 80244 9868 80296 9877
rect 84752 9911 84804 9920
rect 84752 9877 84761 9911
rect 84761 9877 84795 9911
rect 84795 9877 84804 9911
rect 84752 9868 84804 9877
rect 87696 9868 87748 9920
rect 93768 9868 93820 9920
rect 24386 9766 24438 9818
rect 24450 9766 24502 9818
rect 24514 9766 24566 9818
rect 24578 9766 24630 9818
rect 24642 9766 24694 9818
rect 47823 9766 47875 9818
rect 47887 9766 47939 9818
rect 47951 9766 48003 9818
rect 48015 9766 48067 9818
rect 48079 9766 48131 9818
rect 71260 9766 71312 9818
rect 71324 9766 71376 9818
rect 71388 9766 71440 9818
rect 71452 9766 71504 9818
rect 71516 9766 71568 9818
rect 94697 9766 94749 9818
rect 94761 9766 94813 9818
rect 94825 9766 94877 9818
rect 94889 9766 94941 9818
rect 94953 9766 95005 9818
rect 4804 9664 4856 9716
rect 14924 9664 14976 9716
rect 17868 9707 17920 9716
rect 17868 9673 17877 9707
rect 17877 9673 17911 9707
rect 17911 9673 17920 9707
rect 17868 9664 17920 9673
rect 18420 9664 18472 9716
rect 2320 9596 2372 9648
rect 2136 9571 2188 9580
rect 2136 9537 2145 9571
rect 2145 9537 2179 9571
rect 2179 9537 2188 9571
rect 2136 9528 2188 9537
rect 4620 9596 4672 9648
rect 3884 9528 3936 9580
rect 4344 9571 4396 9580
rect 4344 9537 4353 9571
rect 4353 9537 4387 9571
rect 4387 9537 4396 9571
rect 4344 9528 4396 9537
rect 5448 9528 5500 9580
rect 5816 9571 5868 9580
rect 5816 9537 5825 9571
rect 5825 9537 5859 9571
rect 5859 9537 5868 9571
rect 5816 9528 5868 9537
rect 7472 9596 7524 9648
rect 7104 9528 7156 9580
rect 8024 9596 8076 9648
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 11244 9596 11296 9648
rect 7656 9528 7708 9537
rect 4620 9460 4672 9512
rect 9220 9528 9272 9580
rect 8300 9503 8352 9512
rect 3240 9324 3292 9376
rect 3424 9324 3476 9376
rect 6920 9324 6972 9376
rect 7012 9324 7064 9376
rect 8300 9469 8309 9503
rect 8309 9469 8343 9503
rect 8343 9469 8352 9503
rect 8300 9460 8352 9469
rect 7840 9435 7892 9444
rect 7840 9401 7849 9435
rect 7849 9401 7883 9435
rect 7883 9401 7892 9435
rect 7840 9392 7892 9401
rect 10048 9528 10100 9580
rect 11704 9571 11756 9580
rect 9404 9460 9456 9512
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 12992 9596 13044 9648
rect 13636 9596 13688 9648
rect 16120 9596 16172 9648
rect 17040 9596 17092 9648
rect 10508 9460 10560 9512
rect 12072 9460 12124 9512
rect 13452 9528 13504 9580
rect 14188 9571 14240 9580
rect 14188 9537 14197 9571
rect 14197 9537 14231 9571
rect 14231 9537 14240 9571
rect 14188 9528 14240 9537
rect 16028 9571 16080 9580
rect 16028 9537 16037 9571
rect 16037 9537 16071 9571
rect 16071 9537 16080 9571
rect 16028 9528 16080 9537
rect 16212 9571 16264 9580
rect 16212 9537 16221 9571
rect 16221 9537 16255 9571
rect 16255 9537 16264 9571
rect 16212 9528 16264 9537
rect 16304 9571 16356 9580
rect 16304 9537 16313 9571
rect 16313 9537 16347 9571
rect 16347 9537 16356 9571
rect 16304 9528 16356 9537
rect 11980 9392 12032 9444
rect 11888 9367 11940 9376
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 11888 9324 11940 9333
rect 14648 9460 14700 9512
rect 16120 9460 16172 9512
rect 17960 9528 18012 9580
rect 19248 9596 19300 9648
rect 20720 9664 20772 9716
rect 22652 9664 22704 9716
rect 20996 9596 21048 9648
rect 21180 9596 21232 9648
rect 20076 9571 20128 9580
rect 20076 9537 20085 9571
rect 20085 9537 20119 9571
rect 20119 9537 20128 9571
rect 20076 9528 20128 9537
rect 16948 9460 17000 9512
rect 19064 9503 19116 9512
rect 19064 9469 19073 9503
rect 19073 9469 19107 9503
rect 19107 9469 19116 9503
rect 19340 9503 19392 9512
rect 19064 9460 19116 9469
rect 19340 9469 19349 9503
rect 19349 9469 19383 9503
rect 19383 9469 19392 9503
rect 19340 9460 19392 9469
rect 20812 9503 20864 9512
rect 14556 9435 14608 9444
rect 14556 9401 14565 9435
rect 14565 9401 14599 9435
rect 14599 9401 14608 9435
rect 14556 9392 14608 9401
rect 18328 9392 18380 9444
rect 20812 9469 20821 9503
rect 20821 9469 20855 9503
rect 20855 9469 20864 9503
rect 20812 9460 20864 9469
rect 20996 9460 21048 9512
rect 21824 9460 21876 9512
rect 22100 9503 22152 9512
rect 22100 9469 22109 9503
rect 22109 9469 22143 9503
rect 22143 9469 22152 9503
rect 23388 9596 23440 9648
rect 25872 9664 25924 9716
rect 24860 9596 24912 9648
rect 26240 9664 26292 9716
rect 33140 9664 33192 9716
rect 27068 9528 27120 9580
rect 27712 9596 27764 9648
rect 30196 9639 30248 9648
rect 30196 9605 30205 9639
rect 30205 9605 30239 9639
rect 30239 9605 30248 9639
rect 30196 9596 30248 9605
rect 35716 9664 35768 9716
rect 33508 9596 33560 9648
rect 33692 9596 33744 9648
rect 35348 9639 35400 9648
rect 35348 9605 35357 9639
rect 35357 9605 35391 9639
rect 35391 9605 35400 9639
rect 35348 9596 35400 9605
rect 22100 9460 22152 9469
rect 25320 9460 25372 9512
rect 26056 9460 26108 9512
rect 22928 9392 22980 9444
rect 21916 9324 21968 9376
rect 22652 9367 22704 9376
rect 22652 9333 22661 9367
rect 22661 9333 22695 9367
rect 22695 9333 22704 9367
rect 22652 9324 22704 9333
rect 23388 9324 23440 9376
rect 27528 9460 27580 9512
rect 29920 9503 29972 9512
rect 26608 9392 26660 9444
rect 29920 9469 29929 9503
rect 29929 9469 29963 9503
rect 29963 9469 29972 9503
rect 29920 9460 29972 9469
rect 30656 9460 30708 9512
rect 32496 9528 32548 9580
rect 29000 9324 29052 9376
rect 34520 9460 34572 9512
rect 36452 9664 36504 9716
rect 38384 9664 38436 9716
rect 37004 9596 37056 9648
rect 39028 9596 39080 9648
rect 40224 9664 40276 9716
rect 41788 9664 41840 9716
rect 44272 9664 44324 9716
rect 46296 9664 46348 9716
rect 40592 9596 40644 9648
rect 41880 9596 41932 9648
rect 36544 9528 36596 9580
rect 36820 9571 36872 9580
rect 36820 9537 36829 9571
rect 36829 9537 36863 9571
rect 36863 9537 36872 9571
rect 36820 9528 36872 9537
rect 36452 9460 36504 9512
rect 37464 9528 37516 9580
rect 37740 9571 37792 9580
rect 37740 9537 37749 9571
rect 37749 9537 37783 9571
rect 37783 9537 37792 9571
rect 37740 9528 37792 9537
rect 38752 9528 38804 9580
rect 37372 9460 37424 9512
rect 38568 9460 38620 9512
rect 38936 9503 38988 9512
rect 38936 9469 38945 9503
rect 38945 9469 38979 9503
rect 38979 9469 38988 9503
rect 38936 9460 38988 9469
rect 41512 9528 41564 9580
rect 42156 9528 42208 9580
rect 42800 9528 42852 9580
rect 43536 9528 43588 9580
rect 43812 9571 43864 9580
rect 43812 9537 43821 9571
rect 43821 9537 43855 9571
rect 43855 9537 43864 9571
rect 43812 9528 43864 9537
rect 43904 9571 43956 9580
rect 43904 9537 43913 9571
rect 43913 9537 43947 9571
rect 43947 9537 43956 9571
rect 44640 9596 44692 9648
rect 47124 9639 47176 9648
rect 43904 9528 43956 9537
rect 39396 9460 39448 9512
rect 31484 9392 31536 9444
rect 34704 9435 34756 9444
rect 34704 9401 34713 9435
rect 34713 9401 34747 9435
rect 34747 9401 34756 9435
rect 34704 9392 34756 9401
rect 35532 9392 35584 9444
rect 35624 9392 35676 9444
rect 36084 9392 36136 9444
rect 36544 9392 36596 9444
rect 37924 9392 37976 9444
rect 41052 9460 41104 9512
rect 41236 9503 41288 9512
rect 41236 9469 41245 9503
rect 41245 9469 41279 9503
rect 41279 9469 41288 9503
rect 41236 9460 41288 9469
rect 42064 9460 42116 9512
rect 44364 9528 44416 9580
rect 47124 9605 47133 9639
rect 47133 9605 47167 9639
rect 47167 9605 47176 9639
rect 48780 9664 48832 9716
rect 48320 9639 48372 9648
rect 47124 9596 47176 9605
rect 48320 9605 48329 9639
rect 48329 9605 48363 9639
rect 48363 9605 48372 9639
rect 48320 9596 48372 9605
rect 48504 9639 48556 9648
rect 48504 9605 48513 9639
rect 48513 9605 48547 9639
rect 48547 9605 48556 9639
rect 48504 9596 48556 9605
rect 50344 9664 50396 9716
rect 49608 9596 49660 9648
rect 49976 9639 50028 9648
rect 49976 9605 49985 9639
rect 49985 9605 50019 9639
rect 50019 9605 50028 9639
rect 49976 9596 50028 9605
rect 51356 9596 51408 9648
rect 53104 9639 53156 9648
rect 53104 9605 53113 9639
rect 53113 9605 53147 9639
rect 53147 9605 53156 9639
rect 53104 9596 53156 9605
rect 62396 9664 62448 9716
rect 53840 9639 53892 9648
rect 53840 9605 53849 9639
rect 53849 9605 53883 9639
rect 53883 9605 53892 9639
rect 53840 9596 53892 9605
rect 46204 9460 46256 9512
rect 46296 9460 46348 9512
rect 46572 9503 46624 9512
rect 46572 9469 46581 9503
rect 46581 9469 46615 9503
rect 46615 9469 46624 9503
rect 46572 9460 46624 9469
rect 48228 9460 48280 9512
rect 48688 9460 48740 9512
rect 49332 9571 49384 9580
rect 49332 9537 49341 9571
rect 49341 9537 49375 9571
rect 49375 9537 49384 9571
rect 49332 9528 49384 9537
rect 51448 9528 51500 9580
rect 52184 9571 52236 9580
rect 52184 9537 52193 9571
rect 52193 9537 52227 9571
rect 52227 9537 52236 9571
rect 52184 9528 52236 9537
rect 52276 9528 52328 9580
rect 52460 9528 52512 9580
rect 53288 9571 53340 9580
rect 53288 9537 53297 9571
rect 53297 9537 53331 9571
rect 53331 9537 53340 9571
rect 53288 9528 53340 9537
rect 61108 9596 61160 9648
rect 58072 9571 58124 9580
rect 58072 9537 58081 9571
rect 58081 9537 58115 9571
rect 58115 9537 58124 9571
rect 58072 9528 58124 9537
rect 58808 9528 58860 9580
rect 58992 9528 59044 9580
rect 62396 9571 62448 9580
rect 62396 9537 62405 9571
rect 62405 9537 62439 9571
rect 62439 9537 62448 9571
rect 63316 9639 63368 9648
rect 63316 9605 63325 9639
rect 63325 9605 63359 9639
rect 63359 9605 63368 9639
rect 63316 9596 63368 9605
rect 65432 9664 65484 9716
rect 70400 9664 70452 9716
rect 62396 9528 62448 9537
rect 63040 9528 63092 9580
rect 63224 9571 63276 9580
rect 63224 9537 63233 9571
rect 63233 9537 63267 9571
rect 63267 9537 63276 9571
rect 63224 9528 63276 9537
rect 64328 9596 64380 9648
rect 64696 9596 64748 9648
rect 67640 9596 67692 9648
rect 67916 9596 67968 9648
rect 70492 9596 70544 9648
rect 73160 9664 73212 9716
rect 73620 9664 73672 9716
rect 75920 9664 75972 9716
rect 76840 9664 76892 9716
rect 76932 9664 76984 9716
rect 84476 9664 84528 9716
rect 84660 9664 84712 9716
rect 84844 9664 84896 9716
rect 73436 9596 73488 9648
rect 74172 9596 74224 9648
rect 66444 9528 66496 9580
rect 67824 9571 67876 9580
rect 67824 9537 67833 9571
rect 67833 9537 67867 9571
rect 67867 9537 67876 9571
rect 67824 9528 67876 9537
rect 70400 9528 70452 9580
rect 72700 9571 72752 9580
rect 72700 9537 72709 9571
rect 72709 9537 72743 9571
rect 72743 9537 72752 9571
rect 72700 9528 72752 9537
rect 73620 9528 73672 9580
rect 74816 9571 74868 9580
rect 74816 9537 74825 9571
rect 74825 9537 74859 9571
rect 74859 9537 74868 9571
rect 74816 9528 74868 9537
rect 40040 9392 40092 9444
rect 40224 9392 40276 9444
rect 45008 9435 45060 9444
rect 45008 9401 45017 9435
rect 45017 9401 45051 9435
rect 45051 9401 45060 9435
rect 45008 9392 45060 9401
rect 47492 9392 47544 9444
rect 49700 9460 49752 9512
rect 51356 9460 51408 9512
rect 55772 9503 55824 9512
rect 55772 9469 55781 9503
rect 55781 9469 55815 9503
rect 55815 9469 55824 9503
rect 55772 9460 55824 9469
rect 56048 9503 56100 9512
rect 56048 9469 56057 9503
rect 56057 9469 56091 9503
rect 56091 9469 56100 9503
rect 56048 9460 56100 9469
rect 56508 9460 56560 9512
rect 58624 9460 58676 9512
rect 60648 9503 60700 9512
rect 60648 9469 60657 9503
rect 60657 9469 60691 9503
rect 60691 9469 60700 9503
rect 60648 9460 60700 9469
rect 61292 9503 61344 9512
rect 31668 9367 31720 9376
rect 31668 9333 31677 9367
rect 31677 9333 31711 9367
rect 31711 9333 31720 9367
rect 31668 9324 31720 9333
rect 33048 9324 33100 9376
rect 33324 9324 33376 9376
rect 35164 9324 35216 9376
rect 36268 9367 36320 9376
rect 36268 9333 36277 9367
rect 36277 9333 36311 9367
rect 36311 9333 36320 9367
rect 36268 9324 36320 9333
rect 38200 9324 38252 9376
rect 38384 9324 38436 9376
rect 38936 9324 38988 9376
rect 41788 9324 41840 9376
rect 45560 9324 45612 9376
rect 48872 9324 48924 9376
rect 49056 9367 49108 9376
rect 49056 9333 49065 9367
rect 49065 9333 49099 9367
rect 49099 9333 49108 9367
rect 49056 9324 49108 9333
rect 49424 9392 49476 9444
rect 61016 9392 61068 9444
rect 61292 9469 61301 9503
rect 61301 9469 61335 9503
rect 61335 9469 61344 9503
rect 61292 9460 61344 9469
rect 62120 9460 62172 9512
rect 64144 9460 64196 9512
rect 64420 9460 64472 9512
rect 68836 9503 68888 9512
rect 63132 9392 63184 9444
rect 68836 9469 68845 9503
rect 68845 9469 68879 9503
rect 68879 9469 68888 9503
rect 68836 9460 68888 9469
rect 65800 9392 65852 9444
rect 71412 9460 71464 9512
rect 75276 9596 75328 9648
rect 76012 9639 76064 9648
rect 76012 9605 76021 9639
rect 76021 9605 76055 9639
rect 76055 9605 76064 9639
rect 76012 9596 76064 9605
rect 75460 9571 75512 9580
rect 75460 9537 75469 9571
rect 75469 9537 75503 9571
rect 75503 9537 75512 9571
rect 75460 9528 75512 9537
rect 78956 9596 79008 9648
rect 79232 9596 79284 9648
rect 78128 9571 78180 9580
rect 78128 9537 78137 9571
rect 78137 9537 78171 9571
rect 78171 9537 78180 9571
rect 78128 9528 78180 9537
rect 79140 9528 79192 9580
rect 76932 9503 76984 9512
rect 55864 9324 55916 9376
rect 57152 9367 57204 9376
rect 57152 9333 57161 9367
rect 57161 9333 57195 9367
rect 57195 9333 57204 9367
rect 57152 9324 57204 9333
rect 58808 9367 58860 9376
rect 58808 9333 58817 9367
rect 58817 9333 58851 9367
rect 58851 9333 58860 9367
rect 58808 9324 58860 9333
rect 58992 9324 59044 9376
rect 61752 9324 61804 9376
rect 61936 9324 61988 9376
rect 62580 9367 62632 9376
rect 62580 9333 62589 9367
rect 62589 9333 62623 9367
rect 62623 9333 62632 9367
rect 62580 9324 62632 9333
rect 63776 9324 63828 9376
rect 66720 9367 66772 9376
rect 66720 9333 66729 9367
rect 66729 9333 66763 9367
rect 66763 9333 66772 9367
rect 66720 9324 66772 9333
rect 67364 9367 67416 9376
rect 67364 9333 67373 9367
rect 67373 9333 67407 9367
rect 67407 9333 67416 9367
rect 67364 9324 67416 9333
rect 70400 9324 70452 9376
rect 71044 9367 71096 9376
rect 71044 9333 71053 9367
rect 71053 9333 71087 9367
rect 71087 9333 71096 9367
rect 71044 9324 71096 9333
rect 71136 9324 71188 9376
rect 72148 9324 72200 9376
rect 74080 9367 74132 9376
rect 74080 9333 74089 9367
rect 74089 9333 74123 9367
rect 74123 9333 74132 9367
rect 74080 9324 74132 9333
rect 75920 9392 75972 9444
rect 76932 9469 76941 9503
rect 76941 9469 76975 9503
rect 76975 9469 76984 9503
rect 76932 9460 76984 9469
rect 77760 9460 77812 9512
rect 77944 9460 77996 9512
rect 79232 9392 79284 9444
rect 78128 9324 78180 9376
rect 78864 9324 78916 9376
rect 79600 9324 79652 9376
rect 85580 9596 85632 9648
rect 85948 9596 86000 9648
rect 87788 9639 87840 9648
rect 87788 9605 87797 9639
rect 87797 9605 87831 9639
rect 87831 9605 87840 9639
rect 87788 9596 87840 9605
rect 82820 9528 82872 9580
rect 83372 9528 83424 9580
rect 84476 9571 84528 9580
rect 84476 9537 84485 9571
rect 84485 9537 84519 9571
rect 84519 9537 84528 9571
rect 84476 9528 84528 9537
rect 88248 9528 88300 9580
rect 91192 9596 91244 9648
rect 93768 9596 93820 9648
rect 94228 9639 94280 9648
rect 94228 9605 94237 9639
rect 94237 9605 94271 9639
rect 94271 9605 94280 9639
rect 94228 9596 94280 9605
rect 80704 9460 80756 9512
rect 80612 9392 80664 9444
rect 82728 9460 82780 9512
rect 83832 9503 83884 9512
rect 83832 9469 83841 9503
rect 83841 9469 83875 9503
rect 83875 9469 83884 9503
rect 83832 9460 83884 9469
rect 81440 9392 81492 9444
rect 85396 9392 85448 9444
rect 87236 9503 87288 9512
rect 87236 9469 87245 9503
rect 87245 9469 87279 9503
rect 87279 9469 87288 9503
rect 87236 9460 87288 9469
rect 87696 9460 87748 9512
rect 92848 9528 92900 9580
rect 94044 9528 94096 9580
rect 89720 9460 89772 9512
rect 90640 9503 90692 9512
rect 90640 9469 90649 9503
rect 90649 9469 90683 9503
rect 90683 9469 90692 9503
rect 90640 9460 90692 9469
rect 93952 9460 94004 9512
rect 84108 9324 84160 9376
rect 85764 9324 85816 9376
rect 86500 9324 86552 9376
rect 86592 9324 86644 9376
rect 88064 9324 88116 9376
rect 88248 9324 88300 9376
rect 91100 9324 91152 9376
rect 91284 9324 91336 9376
rect 92388 9367 92440 9376
rect 92388 9333 92397 9367
rect 92397 9333 92431 9367
rect 92431 9333 92440 9367
rect 92388 9324 92440 9333
rect 92480 9324 92532 9376
rect 12668 9222 12720 9274
rect 12732 9222 12784 9274
rect 12796 9222 12848 9274
rect 12860 9222 12912 9274
rect 12924 9222 12976 9274
rect 36105 9222 36157 9274
rect 36169 9222 36221 9274
rect 36233 9222 36285 9274
rect 36297 9222 36349 9274
rect 36361 9222 36413 9274
rect 59542 9222 59594 9274
rect 59606 9222 59658 9274
rect 59670 9222 59722 9274
rect 59734 9222 59786 9274
rect 59798 9222 59850 9274
rect 82979 9222 83031 9274
rect 83043 9222 83095 9274
rect 83107 9222 83159 9274
rect 83171 9222 83223 9274
rect 83235 9222 83287 9274
rect 2504 9120 2556 9172
rect 3424 9163 3476 9172
rect 3424 9129 3433 9163
rect 3433 9129 3467 9163
rect 3467 9129 3476 9163
rect 3424 9120 3476 9129
rect 5816 9120 5868 9172
rect 7012 9120 7064 9172
rect 14648 9163 14700 9172
rect 4068 9052 4120 9104
rect 2228 9027 2280 9036
rect 2228 8993 2237 9027
rect 2237 8993 2271 9027
rect 2271 8993 2280 9027
rect 2228 8984 2280 8993
rect 4252 9027 4304 9036
rect 4252 8993 4261 9027
rect 4261 8993 4295 9027
rect 4295 8993 4304 9027
rect 4252 8984 4304 8993
rect 8024 9052 8076 9104
rect 9220 9052 9272 9104
rect 9128 8984 9180 9036
rect 9404 9027 9456 9036
rect 9404 8993 9413 9027
rect 9413 8993 9447 9027
rect 9447 8993 9456 9027
rect 9404 8984 9456 8993
rect 9772 8984 9824 9036
rect 11244 8984 11296 9036
rect 13452 9052 13504 9104
rect 14648 9129 14657 9163
rect 14657 9129 14691 9163
rect 14691 9129 14700 9163
rect 14648 9120 14700 9129
rect 16028 9120 16080 9172
rect 16212 9163 16264 9172
rect 16212 9129 16221 9163
rect 16221 9129 16255 9163
rect 16255 9129 16264 9163
rect 16212 9120 16264 9129
rect 16948 9163 17000 9172
rect 16948 9129 16957 9163
rect 16957 9129 16991 9163
rect 16991 9129 17000 9163
rect 16948 9120 17000 9129
rect 17224 9120 17276 9172
rect 17776 9120 17828 9172
rect 14832 9052 14884 9104
rect 14924 9052 14976 9104
rect 16764 9052 16816 9104
rect 18420 9120 18472 9172
rect 18512 9120 18564 9172
rect 19708 9163 19760 9172
rect 19708 9129 19717 9163
rect 19717 9129 19751 9163
rect 19751 9129 19760 9163
rect 19708 9120 19760 9129
rect 19892 9163 19944 9172
rect 19892 9129 19901 9163
rect 19901 9129 19935 9163
rect 19935 9129 19944 9163
rect 19892 9120 19944 9129
rect 21180 9120 21232 9172
rect 21824 9163 21876 9172
rect 21824 9129 21833 9163
rect 21833 9129 21867 9163
rect 21867 9129 21876 9163
rect 21824 9120 21876 9129
rect 22100 9120 22152 9172
rect 27436 9120 27488 9172
rect 27528 9120 27580 9172
rect 29000 9120 29052 9172
rect 29368 9120 29420 9172
rect 31668 9120 31720 9172
rect 41236 9120 41288 9172
rect 41328 9120 41380 9172
rect 42892 9120 42944 9172
rect 43812 9120 43864 9172
rect 45100 9120 45152 9172
rect 46204 9163 46256 9172
rect 46204 9129 46213 9163
rect 46213 9129 46247 9163
rect 46247 9129 46256 9163
rect 46204 9120 46256 9129
rect 46296 9120 46348 9172
rect 49424 9120 49476 9172
rect 50620 9120 50672 9172
rect 18052 9052 18104 9104
rect 12532 8984 12584 9036
rect 2504 8959 2556 8968
rect 2504 8925 2513 8959
rect 2513 8925 2547 8959
rect 2547 8925 2556 8959
rect 2504 8916 2556 8925
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 4068 8916 4120 8968
rect 4436 8959 4488 8968
rect 4436 8925 4445 8959
rect 4445 8925 4479 8959
rect 4479 8925 4488 8959
rect 4436 8916 4488 8925
rect 4712 8916 4764 8968
rect 8300 8916 8352 8968
rect 10508 8916 10560 8968
rect 10876 8916 10928 8968
rect 6276 8891 6328 8900
rect 6276 8857 6285 8891
rect 6285 8857 6319 8891
rect 6319 8857 6328 8891
rect 6276 8848 6328 8857
rect 2136 8780 2188 8832
rect 5540 8780 5592 8832
rect 7104 8780 7156 8832
rect 7656 8780 7708 8832
rect 8576 8780 8628 8832
rect 13544 8984 13596 9036
rect 15108 8984 15160 9036
rect 16534 8984 16586 9036
rect 16672 8984 16724 9036
rect 16948 8984 17000 9036
rect 13820 8916 13872 8968
rect 16120 8959 16172 8968
rect 13544 8848 13596 8900
rect 16120 8925 16129 8959
rect 16129 8925 16163 8959
rect 16163 8925 16172 8959
rect 16120 8916 16172 8925
rect 16764 8959 16816 8968
rect 16764 8925 16773 8959
rect 16773 8925 16807 8959
rect 16807 8925 16816 8959
rect 16764 8916 16816 8925
rect 16856 8959 16908 8968
rect 16856 8925 16865 8959
rect 16865 8925 16899 8959
rect 16899 8925 16908 8959
rect 16856 8916 16908 8925
rect 17316 8916 17368 8968
rect 17592 8984 17644 9036
rect 18052 8916 18104 8968
rect 16672 8848 16724 8900
rect 18328 8891 18380 8900
rect 15292 8780 15344 8832
rect 15844 8780 15896 8832
rect 18328 8857 18337 8891
rect 18337 8857 18371 8891
rect 18371 8857 18380 8891
rect 18328 8848 18380 8857
rect 18420 8823 18472 8832
rect 18420 8789 18429 8823
rect 18429 8789 18463 8823
rect 18463 8789 18472 8823
rect 18420 8780 18472 8789
rect 19156 8984 19208 9036
rect 20536 9027 20588 9036
rect 20536 8993 20545 9027
rect 20545 8993 20579 9027
rect 20579 8993 20588 9027
rect 20536 8984 20588 8993
rect 25320 9095 25372 9104
rect 25320 9061 25329 9095
rect 25329 9061 25363 9095
rect 25363 9061 25372 9095
rect 25320 9052 25372 9061
rect 27068 9052 27120 9104
rect 19616 8916 19668 8968
rect 19708 8959 19760 8968
rect 19708 8925 19717 8959
rect 19717 8925 19751 8959
rect 19751 8925 19760 8959
rect 20628 8959 20680 8968
rect 19708 8916 19760 8925
rect 20628 8925 20637 8959
rect 20637 8925 20671 8959
rect 20671 8925 20680 8959
rect 20628 8916 20680 8925
rect 20720 8916 20772 8968
rect 22100 8984 22152 9036
rect 22192 8984 22244 9036
rect 25044 8984 25096 9036
rect 25780 9027 25832 9036
rect 25780 8993 25789 9027
rect 25789 8993 25823 9027
rect 25823 8993 25832 9027
rect 25780 8984 25832 8993
rect 28540 9027 28592 9036
rect 22376 8959 22428 8968
rect 18696 8891 18748 8900
rect 18696 8857 18705 8891
rect 18705 8857 18739 8891
rect 18739 8857 18748 8891
rect 18696 8848 18748 8857
rect 19524 8848 19576 8900
rect 19800 8848 19852 8900
rect 22376 8925 22385 8959
rect 22385 8925 22419 8959
rect 22419 8925 22428 8959
rect 22376 8916 22428 8925
rect 22560 8959 22612 8968
rect 22560 8925 22569 8959
rect 22569 8925 22603 8959
rect 22603 8925 22612 8959
rect 22560 8916 22612 8925
rect 21916 8891 21968 8900
rect 21916 8857 21925 8891
rect 21925 8857 21959 8891
rect 21959 8857 21968 8891
rect 21916 8848 21968 8857
rect 26516 8848 26568 8900
rect 28540 8993 28549 9027
rect 28549 8993 28583 9027
rect 28583 8993 28592 9027
rect 28540 8984 28592 8993
rect 28448 8959 28500 8968
rect 28448 8925 28457 8959
rect 28457 8925 28491 8959
rect 28491 8925 28500 8959
rect 28448 8916 28500 8925
rect 29736 9052 29788 9104
rect 31484 9052 31536 9104
rect 33232 9052 33284 9104
rect 29920 8984 29972 9036
rect 32496 8984 32548 9036
rect 38844 9052 38896 9104
rect 19708 8780 19760 8832
rect 20260 8780 20312 8832
rect 22652 8780 22704 8832
rect 27068 8780 27120 8832
rect 31484 8848 31536 8900
rect 32864 8916 32916 8968
rect 33508 8916 33560 8968
rect 33692 8916 33744 8968
rect 33968 8916 34020 8968
rect 34336 8959 34388 8968
rect 34336 8925 34345 8959
rect 34345 8925 34379 8959
rect 34379 8925 34388 8959
rect 34336 8916 34388 8925
rect 31760 8848 31812 8900
rect 28724 8780 28776 8832
rect 29644 8780 29696 8832
rect 30012 8780 30064 8832
rect 31668 8780 31720 8832
rect 34520 8848 34572 8900
rect 35164 8891 35216 8900
rect 35164 8857 35173 8891
rect 35173 8857 35207 8891
rect 35207 8857 35216 8891
rect 35164 8848 35216 8857
rect 35624 8848 35676 8900
rect 36820 8848 36872 8900
rect 37556 8959 37608 8968
rect 37556 8925 37565 8959
rect 37565 8925 37599 8959
rect 37599 8925 37608 8959
rect 37556 8916 37608 8925
rect 38108 8916 38160 8968
rect 38384 8959 38436 8968
rect 38384 8925 38393 8959
rect 38393 8925 38427 8959
rect 38427 8925 38436 8959
rect 38384 8916 38436 8925
rect 41512 9052 41564 9104
rect 41604 9052 41656 9104
rect 43536 9052 43588 9104
rect 55220 9120 55272 9172
rect 56140 9120 56192 9172
rect 57888 9120 57940 9172
rect 58164 9120 58216 9172
rect 58992 9120 59044 9172
rect 62396 9120 62448 9172
rect 67272 9120 67324 9172
rect 70216 9120 70268 9172
rect 70308 9120 70360 9172
rect 71044 9120 71096 9172
rect 71596 9120 71648 9172
rect 39304 9027 39356 9036
rect 39304 8993 39313 9027
rect 39313 8993 39347 9027
rect 39347 8993 39356 9027
rect 39304 8984 39356 8993
rect 39764 8984 39816 9036
rect 39028 8916 39080 8968
rect 40500 8959 40552 8968
rect 40500 8925 40509 8959
rect 40509 8925 40543 8959
rect 40543 8925 40552 8959
rect 40500 8916 40552 8925
rect 40684 8959 40736 8968
rect 40684 8925 40693 8959
rect 40693 8925 40727 8959
rect 40727 8925 40736 8959
rect 40684 8916 40736 8925
rect 43444 8984 43496 9036
rect 44272 9027 44324 9036
rect 44272 8993 44281 9027
rect 44281 8993 44315 9027
rect 44315 8993 44324 9027
rect 44272 8984 44324 8993
rect 33324 8823 33376 8832
rect 33324 8789 33333 8823
rect 33333 8789 33367 8823
rect 33367 8789 33376 8823
rect 33324 8780 33376 8789
rect 33876 8823 33928 8832
rect 33876 8789 33885 8823
rect 33885 8789 33919 8823
rect 33919 8789 33928 8823
rect 33876 8780 33928 8789
rect 34152 8780 34204 8832
rect 34888 8780 34940 8832
rect 36728 8780 36780 8832
rect 37188 8823 37240 8832
rect 37188 8789 37197 8823
rect 37197 8789 37231 8823
rect 37231 8789 37240 8823
rect 37188 8780 37240 8789
rect 41604 8848 41656 8900
rect 38660 8780 38712 8832
rect 38844 8823 38896 8832
rect 38844 8789 38853 8823
rect 38853 8789 38887 8823
rect 38887 8789 38896 8823
rect 38844 8780 38896 8789
rect 40960 8780 41012 8832
rect 41420 8823 41472 8832
rect 41420 8789 41429 8823
rect 41429 8789 41463 8823
rect 41463 8789 41472 8823
rect 43812 8959 43864 8968
rect 43812 8925 43821 8959
rect 43821 8925 43855 8959
rect 43855 8925 43864 8959
rect 43812 8916 43864 8925
rect 44456 8916 44508 8968
rect 44732 8916 44784 8968
rect 45192 8916 45244 8968
rect 45468 8959 45520 8968
rect 45468 8925 45477 8959
rect 45477 8925 45511 8959
rect 45511 8925 45520 8959
rect 45652 8959 45704 8968
rect 45468 8916 45520 8925
rect 45652 8925 45661 8959
rect 45661 8925 45695 8959
rect 45695 8925 45704 8959
rect 45652 8916 45704 8925
rect 46204 8916 46256 8968
rect 46388 8959 46440 8968
rect 46388 8925 46397 8959
rect 46397 8925 46431 8959
rect 46431 8925 46440 8959
rect 46388 8916 46440 8925
rect 49056 8984 49108 9036
rect 50712 8984 50764 9036
rect 52460 9052 52512 9104
rect 58532 9052 58584 9104
rect 59636 9052 59688 9104
rect 60096 9052 60148 9104
rect 61292 9052 61344 9104
rect 61752 9052 61804 9104
rect 66720 9052 66772 9104
rect 55772 8984 55824 9036
rect 58624 8984 58676 9036
rect 47400 8959 47452 8968
rect 47400 8925 47409 8959
rect 47409 8925 47443 8959
rect 47443 8925 47452 8959
rect 47400 8916 47452 8925
rect 49792 8916 49844 8968
rect 50620 8916 50672 8968
rect 51448 8916 51500 8968
rect 52276 8916 52328 8968
rect 54944 8916 54996 8968
rect 47584 8891 47636 8900
rect 47584 8857 47593 8891
rect 47593 8857 47627 8891
rect 47627 8857 47636 8891
rect 47584 8848 47636 8857
rect 41420 8780 41472 8789
rect 44364 8780 44416 8832
rect 44916 8780 44968 8832
rect 45468 8780 45520 8832
rect 46572 8823 46624 8832
rect 46572 8789 46581 8823
rect 46581 8789 46615 8823
rect 46615 8789 46624 8823
rect 46572 8780 46624 8789
rect 46756 8780 46808 8832
rect 51356 8848 51408 8900
rect 49424 8780 49476 8832
rect 51632 8780 51684 8832
rect 57612 8891 57664 8900
rect 57612 8857 57621 8891
rect 57621 8857 57655 8891
rect 57655 8857 57664 8891
rect 57612 8848 57664 8857
rect 57888 8916 57940 8968
rect 59912 8984 59964 9036
rect 60648 9027 60700 9036
rect 60648 8993 60657 9027
rect 60657 8993 60691 9027
rect 60691 8993 60700 9027
rect 60648 8984 60700 8993
rect 58900 8959 58952 8968
rect 58900 8925 58909 8959
rect 58909 8925 58943 8959
rect 58943 8925 58952 8959
rect 58900 8916 58952 8925
rect 60924 8916 60976 8968
rect 59636 8848 59688 8900
rect 62120 8984 62172 9036
rect 62304 9027 62356 9036
rect 62304 8993 62313 9027
rect 62313 8993 62347 9027
rect 62347 8993 62356 9027
rect 62304 8984 62356 8993
rect 63500 9027 63552 9036
rect 63500 8993 63509 9027
rect 63509 8993 63543 9027
rect 63543 8993 63552 9027
rect 63500 8984 63552 8993
rect 66168 9027 66220 9036
rect 66168 8993 66177 9027
rect 66177 8993 66211 9027
rect 66211 8993 66220 9027
rect 66168 8984 66220 8993
rect 66260 8984 66312 9036
rect 68192 8984 68244 9036
rect 68468 9027 68520 9036
rect 68468 8993 68477 9027
rect 68477 8993 68511 9027
rect 68511 8993 68520 9027
rect 68468 8984 68520 8993
rect 70860 8984 70912 9036
rect 71412 8984 71464 9036
rect 72700 8984 72752 9036
rect 61292 8848 61344 8900
rect 63776 8916 63828 8968
rect 64236 8959 64288 8968
rect 64236 8925 64245 8959
rect 64245 8925 64279 8959
rect 64279 8925 64288 8959
rect 64236 8916 64288 8925
rect 64328 8916 64380 8968
rect 66536 8848 66588 8900
rect 66996 8848 67048 8900
rect 69940 8916 69992 8968
rect 68192 8848 68244 8900
rect 70768 8848 70820 8900
rect 71688 8916 71740 8968
rect 71780 8959 71832 8968
rect 71780 8925 71789 8959
rect 71789 8925 71823 8959
rect 71823 8925 71832 8959
rect 71780 8916 71832 8925
rect 74816 9120 74868 9172
rect 77392 9120 77444 9172
rect 74080 9027 74132 9036
rect 74080 8993 74089 9027
rect 74089 8993 74123 9027
rect 74123 8993 74132 9027
rect 74080 8984 74132 8993
rect 74540 8984 74592 9036
rect 76656 9052 76708 9104
rect 75276 8984 75328 9036
rect 76196 8984 76248 9036
rect 73804 8959 73856 8968
rect 73068 8848 73120 8900
rect 73804 8925 73813 8959
rect 73813 8925 73847 8959
rect 73847 8925 73856 8959
rect 73804 8916 73856 8925
rect 75184 8916 75236 8968
rect 76564 8916 76616 8968
rect 76932 8959 76984 8968
rect 76932 8925 76941 8959
rect 76941 8925 76975 8959
rect 76975 8925 76984 8959
rect 76932 8916 76984 8925
rect 74356 8848 74408 8900
rect 79140 9120 79192 9172
rect 79416 9120 79468 9172
rect 80612 9052 80664 9104
rect 85672 9120 85724 9172
rect 86592 9120 86644 9172
rect 88064 9120 88116 9172
rect 88432 9120 88484 9172
rect 93952 9163 94004 9172
rect 93952 9129 93961 9163
rect 93961 9129 93995 9163
rect 93995 9129 94004 9163
rect 93952 9120 94004 9129
rect 87236 9052 87288 9104
rect 77852 9027 77904 9036
rect 77852 8993 77861 9027
rect 77861 8993 77895 9027
rect 77895 8993 77904 9027
rect 77852 8984 77904 8993
rect 77944 8984 77996 9036
rect 79140 8916 79192 8968
rect 80520 8961 80572 8968
rect 80520 8927 80529 8961
rect 80529 8927 80563 8961
rect 80563 8927 80572 8961
rect 81256 8959 81308 8968
rect 80520 8916 80572 8927
rect 81256 8925 81265 8959
rect 81265 8925 81299 8959
rect 81299 8925 81308 8959
rect 81256 8916 81308 8925
rect 86040 8984 86092 9036
rect 88156 9027 88208 9036
rect 88156 8993 88165 9027
rect 88165 8993 88199 9027
rect 88199 8993 88208 9027
rect 88156 8984 88208 8993
rect 88432 9027 88484 9036
rect 88432 8993 88441 9027
rect 88441 8993 88475 9027
rect 88475 8993 88484 9027
rect 88432 8984 88484 8993
rect 89812 8984 89864 9036
rect 94136 9052 94188 9104
rect 93216 9027 93268 9036
rect 93216 8993 93225 9027
rect 93225 8993 93259 9027
rect 93259 8993 93268 9027
rect 93216 8984 93268 8993
rect 86500 8959 86552 8968
rect 86500 8925 86509 8959
rect 86509 8925 86543 8959
rect 86543 8925 86552 8959
rect 86500 8916 86552 8925
rect 87696 8916 87748 8968
rect 87880 8916 87932 8968
rect 89444 8916 89496 8968
rect 91284 8916 91336 8968
rect 93860 8959 93912 8968
rect 58440 8780 58492 8832
rect 59360 8780 59412 8832
rect 60556 8780 60608 8832
rect 63224 8780 63276 8832
rect 66628 8780 66680 8832
rect 67548 8780 67600 8832
rect 67640 8780 67692 8832
rect 69940 8780 69992 8832
rect 72516 8780 72568 8832
rect 78128 8848 78180 8900
rect 81532 8891 81584 8900
rect 81532 8857 81541 8891
rect 81541 8857 81575 8891
rect 81575 8857 81584 8891
rect 81532 8848 81584 8857
rect 75552 8823 75604 8832
rect 75552 8789 75561 8823
rect 75561 8789 75595 8823
rect 75595 8789 75604 8823
rect 75552 8780 75604 8789
rect 75736 8780 75788 8832
rect 84016 8848 84068 8900
rect 85672 8848 85724 8900
rect 82820 8780 82872 8832
rect 83464 8780 83516 8832
rect 90180 8848 90232 8900
rect 89168 8780 89220 8832
rect 91008 8780 91060 8832
rect 93124 8848 93176 8900
rect 93860 8925 93869 8959
rect 93869 8925 93903 8959
rect 93903 8925 93912 8959
rect 93860 8916 93912 8925
rect 24386 8678 24438 8730
rect 24450 8678 24502 8730
rect 24514 8678 24566 8730
rect 24578 8678 24630 8730
rect 24642 8678 24694 8730
rect 47823 8678 47875 8730
rect 47887 8678 47939 8730
rect 47951 8678 48003 8730
rect 48015 8678 48067 8730
rect 48079 8678 48131 8730
rect 71260 8678 71312 8730
rect 71324 8678 71376 8730
rect 71388 8678 71440 8730
rect 71452 8678 71504 8730
rect 71516 8678 71568 8730
rect 94697 8678 94749 8730
rect 94761 8678 94813 8730
rect 94825 8678 94877 8730
rect 94889 8678 94941 8730
rect 94953 8678 95005 8730
rect 2136 8619 2188 8628
rect 2136 8585 2145 8619
rect 2145 8585 2179 8619
rect 2179 8585 2188 8619
rect 2136 8576 2188 8585
rect 4712 8619 4764 8628
rect 4712 8585 4721 8619
rect 4721 8585 4755 8619
rect 4755 8585 4764 8619
rect 4712 8576 4764 8585
rect 6276 8576 6328 8628
rect 8576 8576 8628 8628
rect 4436 8508 4488 8560
rect 5080 8508 5132 8560
rect 2228 8304 2280 8356
rect 2872 8304 2924 8356
rect 3976 8372 4028 8424
rect 4252 8415 4304 8424
rect 4252 8381 4261 8415
rect 4261 8381 4295 8415
rect 4295 8381 4304 8415
rect 4252 8372 4304 8381
rect 4528 8304 4580 8356
rect 5724 8508 5776 8560
rect 6736 8440 6788 8492
rect 7012 8440 7064 8492
rect 7472 8440 7524 8492
rect 7564 8483 7616 8492
rect 7564 8449 7573 8483
rect 7573 8449 7607 8483
rect 7607 8449 7616 8483
rect 7564 8440 7616 8449
rect 8208 8440 8260 8492
rect 9128 8483 9180 8492
rect 9128 8449 9137 8483
rect 9137 8449 9171 8483
rect 9171 8449 9180 8483
rect 9128 8440 9180 8449
rect 10876 8415 10928 8424
rect 10876 8381 10885 8415
rect 10885 8381 10919 8415
rect 10919 8381 10928 8415
rect 10876 8372 10928 8381
rect 11888 8576 11940 8628
rect 12348 8440 12400 8492
rect 13728 8483 13780 8492
rect 13728 8449 13737 8483
rect 13737 8449 13771 8483
rect 13771 8449 13780 8483
rect 13728 8440 13780 8449
rect 15016 8576 15068 8628
rect 16856 8576 16908 8628
rect 17040 8619 17092 8628
rect 17040 8585 17049 8619
rect 17049 8585 17083 8619
rect 17083 8585 17092 8619
rect 17040 8576 17092 8585
rect 20536 8576 20588 8628
rect 14188 8508 14240 8560
rect 15844 8551 15896 8560
rect 15844 8517 15853 8551
rect 15853 8517 15887 8551
rect 15887 8517 15896 8551
rect 15844 8508 15896 8517
rect 16028 8508 16080 8560
rect 17132 8508 17184 8560
rect 20260 8551 20312 8560
rect 20260 8517 20269 8551
rect 20269 8517 20303 8551
rect 20303 8517 20312 8551
rect 20260 8508 20312 8517
rect 21456 8551 21508 8560
rect 5264 8279 5316 8288
rect 5264 8245 5273 8279
rect 5273 8245 5307 8279
rect 5307 8245 5316 8279
rect 5264 8236 5316 8245
rect 11336 8304 11388 8356
rect 17500 8440 17552 8492
rect 17592 8440 17644 8492
rect 17684 8483 17736 8492
rect 17684 8449 17694 8483
rect 17694 8449 17728 8483
rect 17728 8449 17736 8483
rect 17684 8440 17736 8449
rect 18696 8440 18748 8492
rect 17408 8372 17460 8424
rect 17960 8415 18012 8424
rect 17960 8381 17969 8415
rect 17969 8381 18003 8415
rect 18003 8381 18012 8415
rect 17960 8372 18012 8381
rect 18328 8372 18380 8424
rect 19616 8440 19668 8492
rect 20444 8483 20496 8492
rect 20444 8449 20453 8483
rect 20453 8449 20487 8483
rect 20487 8449 20496 8483
rect 21456 8517 21465 8551
rect 21465 8517 21499 8551
rect 21499 8517 21508 8551
rect 21456 8508 21508 8517
rect 20444 8440 20496 8449
rect 22100 8440 22152 8492
rect 22376 8508 22428 8560
rect 22560 8440 22612 8492
rect 21824 8372 21876 8424
rect 15108 8347 15160 8356
rect 15108 8313 15117 8347
rect 15117 8313 15151 8347
rect 15151 8313 15160 8347
rect 15108 8304 15160 8313
rect 17224 8304 17276 8356
rect 17592 8304 17644 8356
rect 22928 8372 22980 8424
rect 23296 8415 23348 8424
rect 23296 8381 23305 8415
rect 23305 8381 23339 8415
rect 23339 8381 23348 8415
rect 23296 8372 23348 8381
rect 24860 8508 24912 8560
rect 23756 8483 23808 8492
rect 23756 8449 23765 8483
rect 23765 8449 23799 8483
rect 23799 8449 23808 8483
rect 23756 8440 23808 8449
rect 27712 8576 27764 8628
rect 28540 8576 28592 8628
rect 33876 8576 33928 8628
rect 29828 8508 29880 8560
rect 30656 8508 30708 8560
rect 31484 8508 31536 8560
rect 34520 8508 34572 8560
rect 35716 8576 35768 8628
rect 36268 8576 36320 8628
rect 36452 8619 36504 8628
rect 36452 8585 36461 8619
rect 36461 8585 36495 8619
rect 36495 8585 36504 8619
rect 36452 8576 36504 8585
rect 37096 8576 37148 8628
rect 38384 8576 38436 8628
rect 42432 8576 42484 8628
rect 37188 8508 37240 8560
rect 37556 8508 37608 8560
rect 41328 8508 41380 8560
rect 29920 8483 29972 8492
rect 29920 8449 29929 8483
rect 29929 8449 29963 8483
rect 29963 8449 29972 8483
rect 29920 8440 29972 8449
rect 32496 8440 32548 8492
rect 33324 8440 33376 8492
rect 29736 8372 29788 8424
rect 33876 8415 33928 8424
rect 16304 8236 16356 8288
rect 19892 8236 19944 8288
rect 29460 8347 29512 8356
rect 29460 8313 29469 8347
rect 29469 8313 29503 8347
rect 29503 8313 29512 8347
rect 29460 8304 29512 8313
rect 29920 8304 29972 8356
rect 31852 8304 31904 8356
rect 32404 8304 32456 8356
rect 33416 8304 33468 8356
rect 26148 8236 26200 8288
rect 31668 8279 31720 8288
rect 31668 8245 31677 8279
rect 31677 8245 31711 8279
rect 31711 8245 31720 8279
rect 31668 8236 31720 8245
rect 32772 8236 32824 8288
rect 33876 8381 33885 8415
rect 33885 8381 33919 8415
rect 33919 8381 33928 8415
rect 33876 8372 33928 8381
rect 33968 8372 34020 8424
rect 36360 8440 36412 8492
rect 35808 8372 35860 8424
rect 37648 8483 37700 8492
rect 37648 8449 37657 8483
rect 37657 8449 37691 8483
rect 37691 8449 37700 8483
rect 37648 8440 37700 8449
rect 38660 8440 38712 8492
rect 40316 8440 40368 8492
rect 40500 8483 40552 8492
rect 40500 8449 40509 8483
rect 40509 8449 40543 8483
rect 40543 8449 40552 8483
rect 40500 8440 40552 8449
rect 40776 8483 40828 8492
rect 40776 8449 40785 8483
rect 40785 8449 40819 8483
rect 40819 8449 40828 8483
rect 40776 8440 40828 8449
rect 41052 8440 41104 8492
rect 40408 8372 40460 8424
rect 37832 8304 37884 8356
rect 39764 8347 39816 8356
rect 39764 8313 39773 8347
rect 39773 8313 39807 8347
rect 39807 8313 39816 8347
rect 39764 8304 39816 8313
rect 40684 8415 40736 8424
rect 40684 8381 40693 8415
rect 40693 8381 40727 8415
rect 40727 8381 40736 8415
rect 41604 8415 41656 8424
rect 40684 8372 40736 8381
rect 41604 8381 41613 8415
rect 41613 8381 41647 8415
rect 41647 8381 41656 8415
rect 41604 8372 41656 8381
rect 42064 8415 42116 8424
rect 42064 8381 42073 8415
rect 42073 8381 42107 8415
rect 42107 8381 42116 8415
rect 42064 8372 42116 8381
rect 42708 8372 42760 8424
rect 42892 8483 42944 8492
rect 42892 8449 42901 8483
rect 42901 8449 42935 8483
rect 42935 8449 42944 8483
rect 44180 8576 44232 8628
rect 45192 8619 45244 8628
rect 45192 8585 45201 8619
rect 45201 8585 45235 8619
rect 45235 8585 45244 8619
rect 45192 8576 45244 8585
rect 45376 8576 45428 8628
rect 47400 8576 47452 8628
rect 46572 8508 46624 8560
rect 49516 8619 49568 8628
rect 49516 8585 49525 8619
rect 49525 8585 49559 8619
rect 49559 8585 49568 8619
rect 49516 8576 49568 8585
rect 50620 8619 50672 8628
rect 50620 8585 50629 8619
rect 50629 8585 50663 8619
rect 50663 8585 50672 8619
rect 50620 8576 50672 8585
rect 42892 8440 42944 8449
rect 43168 8440 43220 8492
rect 44916 8440 44968 8492
rect 46848 8440 46900 8492
rect 43444 8372 43496 8424
rect 43536 8372 43588 8424
rect 44088 8372 44140 8424
rect 45652 8372 45704 8424
rect 47032 8372 47084 8424
rect 35808 8236 35860 8288
rect 35900 8236 35952 8288
rect 36268 8236 36320 8288
rect 37556 8236 37608 8288
rect 38752 8279 38804 8288
rect 38752 8245 38761 8279
rect 38761 8245 38795 8279
rect 38795 8245 38804 8279
rect 38752 8236 38804 8245
rect 40684 8236 40736 8288
rect 42892 8236 42944 8288
rect 45744 8279 45796 8288
rect 45744 8245 45753 8279
rect 45753 8245 45787 8279
rect 45787 8245 45796 8279
rect 45744 8236 45796 8245
rect 46572 8304 46624 8356
rect 46756 8236 46808 8288
rect 47308 8372 47360 8424
rect 49424 8440 49476 8492
rect 49608 8440 49660 8492
rect 53656 8576 53708 8628
rect 53748 8576 53800 8628
rect 57244 8576 57296 8628
rect 59268 8576 59320 8628
rect 62580 8576 62632 8628
rect 73804 8576 73856 8628
rect 75184 8619 75236 8628
rect 75184 8585 75193 8619
rect 75193 8585 75227 8619
rect 75227 8585 75236 8619
rect 75184 8576 75236 8585
rect 51632 8508 51684 8560
rect 52092 8551 52144 8560
rect 52092 8517 52101 8551
rect 52101 8517 52135 8551
rect 52135 8517 52144 8551
rect 52092 8508 52144 8517
rect 52184 8508 52236 8560
rect 53196 8483 53248 8492
rect 53196 8449 53205 8483
rect 53205 8449 53239 8483
rect 53239 8449 53248 8483
rect 53196 8440 53248 8449
rect 58624 8508 58676 8560
rect 53932 8483 53984 8492
rect 48688 8415 48740 8424
rect 48688 8381 48697 8415
rect 48697 8381 48731 8415
rect 48731 8381 48740 8415
rect 48688 8372 48740 8381
rect 49976 8415 50028 8424
rect 49976 8381 49985 8415
rect 49985 8381 50019 8415
rect 50019 8381 50028 8415
rect 49976 8372 50028 8381
rect 52368 8415 52420 8424
rect 52368 8381 52377 8415
rect 52377 8381 52411 8415
rect 52411 8381 52420 8415
rect 52368 8372 52420 8381
rect 52644 8372 52696 8424
rect 53472 8415 53524 8424
rect 53472 8381 53481 8415
rect 53481 8381 53515 8415
rect 53515 8381 53524 8415
rect 53472 8372 53524 8381
rect 53932 8449 53941 8483
rect 53941 8449 53975 8483
rect 53975 8449 53984 8483
rect 53932 8440 53984 8449
rect 58164 8440 58216 8492
rect 55220 8415 55272 8424
rect 48320 8304 48372 8356
rect 48872 8236 48924 8288
rect 51448 8236 51500 8288
rect 55220 8381 55229 8415
rect 55229 8381 55263 8415
rect 55263 8381 55272 8415
rect 55220 8372 55272 8381
rect 55496 8415 55548 8424
rect 55496 8381 55505 8415
rect 55505 8381 55539 8415
rect 55539 8381 55548 8415
rect 55496 8372 55548 8381
rect 55864 8372 55916 8424
rect 58256 8372 58308 8424
rect 60096 8508 60148 8560
rect 66812 8508 66864 8560
rect 67548 8508 67600 8560
rect 69756 8508 69808 8560
rect 59360 8483 59412 8492
rect 59360 8449 59369 8483
rect 59369 8449 59403 8483
rect 59403 8449 59412 8483
rect 59360 8440 59412 8449
rect 62212 8483 62264 8492
rect 59084 8415 59136 8424
rect 59084 8381 59093 8415
rect 59093 8381 59127 8415
rect 59127 8381 59136 8415
rect 59084 8372 59136 8381
rect 59268 8415 59320 8424
rect 59268 8381 59277 8415
rect 59277 8381 59311 8415
rect 59311 8381 59320 8415
rect 59268 8372 59320 8381
rect 59820 8415 59872 8424
rect 59820 8381 59829 8415
rect 59829 8381 59863 8415
rect 59863 8381 59872 8415
rect 59820 8372 59872 8381
rect 60096 8415 60148 8424
rect 60096 8381 60105 8415
rect 60105 8381 60139 8415
rect 60139 8381 60148 8415
rect 60096 8372 60148 8381
rect 59360 8304 59412 8356
rect 62212 8449 62221 8483
rect 62221 8449 62255 8483
rect 62255 8449 62264 8483
rect 62212 8440 62264 8449
rect 63684 8483 63736 8492
rect 63684 8449 63693 8483
rect 63693 8449 63727 8483
rect 63727 8449 63736 8483
rect 64512 8483 64564 8492
rect 63684 8440 63736 8449
rect 64512 8449 64521 8483
rect 64521 8449 64555 8483
rect 64555 8449 64564 8483
rect 64512 8440 64564 8449
rect 73620 8483 73672 8492
rect 73620 8449 73629 8483
rect 73629 8449 73663 8483
rect 73663 8449 73672 8483
rect 73620 8440 73672 8449
rect 75552 8508 75604 8560
rect 74356 8440 74408 8492
rect 75276 8483 75328 8492
rect 75276 8449 75285 8483
rect 75285 8449 75319 8483
rect 75319 8449 75328 8483
rect 75276 8440 75328 8449
rect 75736 8483 75788 8492
rect 63776 8415 63828 8424
rect 63776 8381 63785 8415
rect 63785 8381 63819 8415
rect 63819 8381 63828 8415
rect 63776 8372 63828 8381
rect 64788 8415 64840 8424
rect 64788 8381 64797 8415
rect 64797 8381 64831 8415
rect 64831 8381 64840 8415
rect 64788 8372 64840 8381
rect 67548 8415 67600 8424
rect 67548 8381 67557 8415
rect 67557 8381 67591 8415
rect 67591 8381 67600 8415
rect 67548 8372 67600 8381
rect 68192 8372 68244 8424
rect 68560 8372 68612 8424
rect 63408 8304 63460 8356
rect 70768 8372 70820 8424
rect 72516 8415 72568 8424
rect 72516 8381 72525 8415
rect 72525 8381 72559 8415
rect 72559 8381 72568 8415
rect 72516 8372 72568 8381
rect 72792 8415 72844 8424
rect 72792 8381 72801 8415
rect 72801 8381 72835 8415
rect 72835 8381 72844 8415
rect 72792 8372 72844 8381
rect 72976 8415 73028 8424
rect 72976 8381 72985 8415
rect 72985 8381 73019 8415
rect 73019 8381 73028 8415
rect 72976 8372 73028 8381
rect 73068 8372 73120 8424
rect 73160 8304 73212 8356
rect 74724 8372 74776 8424
rect 74816 8372 74868 8424
rect 75736 8449 75745 8483
rect 75745 8449 75779 8483
rect 75779 8449 75788 8483
rect 75736 8440 75788 8449
rect 80520 8576 80572 8628
rect 81532 8576 81584 8628
rect 82636 8576 82688 8628
rect 76472 8508 76524 8560
rect 76104 8415 76156 8424
rect 76104 8381 76113 8415
rect 76113 8381 76147 8415
rect 76147 8381 76156 8415
rect 76104 8372 76156 8381
rect 76380 8372 76432 8424
rect 77944 8508 77996 8560
rect 78864 8551 78916 8560
rect 78864 8517 78873 8551
rect 78873 8517 78907 8551
rect 78907 8517 78916 8551
rect 78864 8508 78916 8517
rect 80244 8440 80296 8492
rect 78680 8415 78732 8424
rect 78680 8381 78689 8415
rect 78689 8381 78723 8415
rect 78723 8381 78732 8415
rect 78680 8372 78732 8381
rect 78864 8372 78916 8424
rect 81716 8372 81768 8424
rect 56508 8236 56560 8288
rect 57244 8236 57296 8288
rect 59176 8279 59228 8288
rect 59176 8245 59185 8279
rect 59185 8245 59219 8279
rect 59219 8245 59228 8279
rect 59176 8236 59228 8245
rect 60188 8236 60240 8288
rect 63316 8236 63368 8288
rect 64144 8236 64196 8288
rect 66076 8279 66128 8288
rect 66076 8245 66085 8279
rect 66085 8245 66119 8279
rect 66119 8245 66128 8279
rect 66076 8236 66128 8245
rect 66996 8236 67048 8288
rect 67456 8236 67508 8288
rect 69112 8236 69164 8288
rect 73620 8236 73672 8288
rect 74356 8236 74408 8288
rect 81256 8347 81308 8356
rect 81256 8313 81265 8347
rect 81265 8313 81299 8347
rect 81299 8313 81308 8347
rect 82636 8440 82688 8492
rect 83556 8508 83608 8560
rect 84292 8508 84344 8560
rect 88984 8576 89036 8628
rect 83372 8440 83424 8492
rect 83648 8440 83700 8492
rect 84200 8440 84252 8492
rect 85396 8415 85448 8424
rect 85396 8381 85405 8415
rect 85405 8381 85439 8415
rect 85439 8381 85448 8415
rect 85396 8372 85448 8381
rect 85488 8372 85540 8424
rect 88340 8508 88392 8560
rect 93400 8551 93452 8560
rect 89260 8483 89312 8492
rect 81256 8304 81308 8313
rect 84660 8304 84712 8356
rect 82728 8236 82780 8288
rect 84292 8236 84344 8288
rect 86684 8236 86736 8288
rect 89260 8449 89269 8483
rect 89269 8449 89303 8483
rect 89303 8449 89312 8483
rect 89260 8440 89312 8449
rect 89720 8440 89772 8492
rect 89444 8372 89496 8424
rect 90180 8415 90232 8424
rect 90180 8381 90189 8415
rect 90189 8381 90223 8415
rect 90223 8381 90232 8415
rect 90180 8372 90232 8381
rect 93400 8517 93409 8551
rect 93409 8517 93443 8551
rect 93443 8517 93452 8551
rect 93400 8508 93452 8517
rect 91008 8372 91060 8424
rect 93584 8415 93636 8424
rect 93584 8381 93593 8415
rect 93593 8381 93627 8415
rect 93627 8381 93636 8415
rect 93584 8372 93636 8381
rect 91192 8347 91244 8356
rect 91192 8313 91201 8347
rect 91201 8313 91235 8347
rect 91235 8313 91244 8347
rect 91192 8304 91244 8313
rect 94136 8347 94188 8356
rect 94136 8313 94145 8347
rect 94145 8313 94179 8347
rect 94179 8313 94188 8347
rect 94136 8304 94188 8313
rect 89812 8236 89864 8288
rect 12668 8134 12720 8186
rect 12732 8134 12784 8186
rect 12796 8134 12848 8186
rect 12860 8134 12912 8186
rect 12924 8134 12976 8186
rect 36105 8134 36157 8186
rect 36169 8134 36221 8186
rect 36233 8134 36285 8186
rect 36297 8134 36349 8186
rect 36361 8134 36413 8186
rect 59542 8134 59594 8186
rect 59606 8134 59658 8186
rect 59670 8134 59722 8186
rect 59734 8134 59786 8186
rect 59798 8134 59850 8186
rect 82979 8134 83031 8186
rect 83043 8134 83095 8186
rect 83107 8134 83159 8186
rect 83171 8134 83223 8186
rect 83235 8134 83287 8186
rect 2872 8075 2924 8084
rect 2872 8041 2881 8075
rect 2881 8041 2915 8075
rect 2915 8041 2924 8075
rect 2872 8032 2924 8041
rect 4344 8032 4396 8084
rect 6828 8032 6880 8084
rect 5264 7939 5316 7948
rect 5264 7905 5273 7939
rect 5273 7905 5307 7939
rect 5307 7905 5316 7939
rect 5264 7896 5316 7905
rect 11704 8032 11756 8084
rect 12532 8032 12584 8084
rect 17316 8032 17368 8084
rect 17500 8032 17552 8084
rect 18880 8032 18932 8084
rect 21640 8075 21692 8084
rect 21640 8041 21649 8075
rect 21649 8041 21683 8075
rect 21683 8041 21692 8075
rect 21640 8032 21692 8041
rect 21824 8075 21876 8084
rect 21824 8041 21833 8075
rect 21833 8041 21867 8075
rect 21867 8041 21876 8075
rect 21824 8032 21876 8041
rect 21916 8032 21968 8084
rect 28632 8032 28684 8084
rect 33140 8032 33192 8084
rect 33324 8075 33376 8084
rect 33324 8041 33333 8075
rect 33333 8041 33367 8075
rect 33367 8041 33376 8075
rect 33324 8032 33376 8041
rect 7656 8007 7708 8016
rect 7656 7973 7665 8007
rect 7665 7973 7699 8007
rect 7699 7973 7708 8007
rect 7656 7964 7708 7973
rect 13544 7964 13596 8016
rect 15108 7964 15160 8016
rect 17960 7896 18012 7948
rect 20720 7896 20772 7948
rect 20904 7939 20956 7948
rect 20904 7905 20913 7939
rect 20913 7905 20947 7939
rect 20947 7905 20956 7939
rect 20904 7896 20956 7905
rect 3700 7828 3752 7880
rect 9128 7828 9180 7880
rect 9680 7828 9732 7880
rect 10140 7828 10192 7880
rect 11336 7871 11388 7880
rect 5724 7760 5776 7812
rect 4252 7692 4304 7744
rect 4436 7692 4488 7744
rect 11336 7837 11345 7871
rect 11345 7837 11379 7871
rect 11379 7837 11388 7871
rect 11336 7828 11388 7837
rect 11704 7871 11756 7880
rect 11704 7837 11713 7871
rect 11713 7837 11747 7871
rect 11747 7837 11756 7871
rect 11704 7828 11756 7837
rect 18144 7828 18196 7880
rect 18696 7871 18748 7880
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 12348 7760 12400 7812
rect 13176 7803 13228 7812
rect 13176 7769 13185 7803
rect 13185 7769 13219 7803
rect 13219 7769 13228 7803
rect 13176 7760 13228 7769
rect 13728 7760 13780 7812
rect 20260 7828 20312 7880
rect 21272 7828 21324 7880
rect 21916 7896 21968 7948
rect 27988 7964 28040 8016
rect 29000 7964 29052 8016
rect 35716 8032 35768 8084
rect 35808 8032 35860 8084
rect 24860 7896 24912 7948
rect 26240 7896 26292 7948
rect 26516 7896 26568 7948
rect 27160 7939 27212 7948
rect 27160 7905 27169 7939
rect 27169 7905 27203 7939
rect 27203 7905 27212 7939
rect 27160 7896 27212 7905
rect 27252 7896 27304 7948
rect 33048 7896 33100 7948
rect 33140 7896 33192 7948
rect 40040 7964 40092 8016
rect 40684 7964 40736 8016
rect 40132 7896 40184 7948
rect 40776 7939 40828 7948
rect 40776 7905 40785 7939
rect 40785 7905 40819 7939
rect 40819 7905 40828 7939
rect 40776 7896 40828 7905
rect 22192 7760 22244 7812
rect 8576 7692 8628 7744
rect 16948 7735 17000 7744
rect 16948 7701 16957 7735
rect 16957 7701 16991 7735
rect 16991 7701 17000 7735
rect 16948 7692 17000 7701
rect 18604 7692 18656 7744
rect 22928 7735 22980 7744
rect 22928 7701 22937 7735
rect 22937 7701 22971 7735
rect 22971 7701 22980 7735
rect 22928 7692 22980 7701
rect 23296 7692 23348 7744
rect 28448 7828 28500 7880
rect 27712 7760 27764 7812
rect 30472 7828 30524 7880
rect 33600 7828 33652 7880
rect 34888 7871 34940 7880
rect 34888 7837 34897 7871
rect 34897 7837 34931 7871
rect 34931 7837 34940 7871
rect 34888 7828 34940 7837
rect 37740 7828 37792 7880
rect 40040 7828 40092 7880
rect 43076 8032 43128 8084
rect 45652 8032 45704 8084
rect 47216 8032 47268 8084
rect 48228 8075 48280 8084
rect 48228 8041 48237 8075
rect 48237 8041 48271 8075
rect 48271 8041 48280 8075
rect 48228 8032 48280 8041
rect 49240 8075 49292 8084
rect 49240 8041 49249 8075
rect 49249 8041 49283 8075
rect 49283 8041 49292 8075
rect 49240 8032 49292 8041
rect 49700 8075 49752 8084
rect 49700 8041 49709 8075
rect 49709 8041 49743 8075
rect 49743 8041 49752 8075
rect 49700 8032 49752 8041
rect 49976 8032 50028 8084
rect 52184 8075 52236 8084
rect 52184 8041 52193 8075
rect 52193 8041 52227 8075
rect 52227 8041 52236 8075
rect 52184 8032 52236 8041
rect 53196 8032 53248 8084
rect 55496 8032 55548 8084
rect 58900 8032 58952 8084
rect 42616 7964 42668 8016
rect 41604 7871 41656 7880
rect 41604 7837 41613 7871
rect 41613 7837 41647 7871
rect 41647 7837 41656 7871
rect 41604 7828 41656 7837
rect 42524 7828 42576 7880
rect 29828 7803 29880 7812
rect 29828 7769 29837 7803
rect 29837 7769 29871 7803
rect 29871 7769 29880 7803
rect 29828 7760 29880 7769
rect 28724 7692 28776 7744
rect 28908 7735 28960 7744
rect 28908 7701 28917 7735
rect 28917 7701 28951 7735
rect 28951 7701 28960 7735
rect 33508 7760 33560 7812
rect 34520 7760 34572 7812
rect 35624 7760 35676 7812
rect 37464 7760 37516 7812
rect 28908 7692 28960 7701
rect 36544 7692 36596 7744
rect 36636 7692 36688 7744
rect 40960 7760 41012 7812
rect 39120 7692 39172 7744
rect 41328 7692 41380 7744
rect 42892 7939 42944 7948
rect 42892 7905 42901 7939
rect 42901 7905 42935 7939
rect 42935 7905 42944 7939
rect 42892 7896 42944 7905
rect 45376 7896 45428 7948
rect 47032 8007 47084 8016
rect 47032 7973 47041 8007
rect 47041 7973 47075 8007
rect 47075 7973 47084 8007
rect 47032 7964 47084 7973
rect 47400 7964 47452 8016
rect 45836 7896 45888 7948
rect 47216 7896 47268 7948
rect 42984 7871 43036 7880
rect 42984 7837 42993 7871
rect 42993 7837 43027 7871
rect 43027 7837 43036 7871
rect 42984 7828 43036 7837
rect 43812 7828 43864 7880
rect 45652 7871 45704 7880
rect 45652 7837 45661 7871
rect 45661 7837 45695 7871
rect 45695 7837 45704 7871
rect 45652 7828 45704 7837
rect 47032 7828 47084 7880
rect 49332 7896 49384 7948
rect 49700 7896 49752 7948
rect 53380 7964 53432 8016
rect 57704 7964 57756 8016
rect 61016 8032 61068 8084
rect 61108 8032 61160 8084
rect 60096 7964 60148 8016
rect 48228 7871 48280 7880
rect 48228 7837 48237 7871
rect 48237 7837 48271 7871
rect 48271 7837 48280 7871
rect 48228 7828 48280 7837
rect 48320 7871 48372 7880
rect 48320 7837 48329 7871
rect 48329 7837 48363 7871
rect 48363 7837 48372 7871
rect 48320 7828 48372 7837
rect 42892 7692 42944 7744
rect 46848 7760 46900 7812
rect 47216 7760 47268 7812
rect 52644 7896 52696 7948
rect 52736 7896 52788 7948
rect 55312 7896 55364 7948
rect 57152 7896 57204 7948
rect 57336 7896 57388 7948
rect 51172 7871 51224 7880
rect 51172 7837 51200 7871
rect 51200 7837 51224 7871
rect 51172 7828 51224 7837
rect 51448 7871 51500 7880
rect 51448 7837 51457 7871
rect 51457 7837 51491 7871
rect 51491 7837 51500 7871
rect 51448 7828 51500 7837
rect 50436 7803 50488 7812
rect 50436 7769 50445 7803
rect 50445 7769 50479 7803
rect 50479 7769 50488 7803
rect 50436 7760 50488 7769
rect 50988 7760 51040 7812
rect 51356 7803 51408 7812
rect 51356 7769 51365 7803
rect 51365 7769 51399 7803
rect 51399 7769 51408 7803
rect 51356 7760 51408 7769
rect 51816 7760 51868 7812
rect 53196 7828 53248 7880
rect 54852 7828 54904 7880
rect 53932 7760 53984 7812
rect 55680 7828 55732 7880
rect 55956 7760 56008 7812
rect 44088 7735 44140 7744
rect 44088 7701 44097 7735
rect 44097 7701 44131 7735
rect 44131 7701 44140 7735
rect 44088 7692 44140 7701
rect 44180 7692 44232 7744
rect 48872 7692 48924 7744
rect 51908 7692 51960 7744
rect 52092 7692 52144 7744
rect 52920 7735 52972 7744
rect 52920 7701 52929 7735
rect 52929 7701 52963 7735
rect 52963 7701 52972 7735
rect 52920 7692 52972 7701
rect 55864 7692 55916 7744
rect 58808 7760 58860 7812
rect 59176 7896 59228 7948
rect 60924 7939 60976 7948
rect 60924 7905 60933 7939
rect 60933 7905 60967 7939
rect 60967 7905 60976 7939
rect 60924 7896 60976 7905
rect 61016 7896 61068 7948
rect 66260 7964 66312 8016
rect 69112 8007 69164 8016
rect 69112 7973 69121 8007
rect 69121 7973 69155 8007
rect 69155 7973 69164 8007
rect 69112 7964 69164 7973
rect 71872 7964 71924 8016
rect 66076 7939 66128 7948
rect 60188 7828 60240 7880
rect 60648 7871 60700 7880
rect 60648 7837 60657 7871
rect 60657 7837 60691 7871
rect 60691 7837 60700 7871
rect 60648 7828 60700 7837
rect 62212 7828 62264 7880
rect 65156 7871 65208 7880
rect 65156 7837 65165 7871
rect 65165 7837 65199 7871
rect 65199 7837 65208 7871
rect 66076 7905 66085 7939
rect 66085 7905 66119 7939
rect 66119 7905 66128 7939
rect 66076 7896 66128 7905
rect 66352 7896 66404 7948
rect 67272 7896 67324 7948
rect 65156 7828 65208 7837
rect 69756 7871 69808 7880
rect 69756 7837 69765 7871
rect 69765 7837 69799 7871
rect 69799 7837 69808 7871
rect 69756 7828 69808 7837
rect 70584 7828 70636 7880
rect 71504 7871 71556 7880
rect 71504 7837 71513 7871
rect 71513 7837 71547 7871
rect 71547 7837 71556 7871
rect 71504 7828 71556 7837
rect 71872 7828 71924 7880
rect 73160 8032 73212 8084
rect 72976 7964 73028 8016
rect 76472 8032 76524 8084
rect 79048 8032 79100 8084
rect 74724 7939 74776 7948
rect 74724 7905 74733 7939
rect 74733 7905 74767 7939
rect 74767 7905 74776 7939
rect 74724 7896 74776 7905
rect 78864 7964 78916 8016
rect 81716 7964 81768 8016
rect 76288 7896 76340 7948
rect 78128 7896 78180 7948
rect 81440 7939 81492 7948
rect 81440 7905 81449 7939
rect 81449 7905 81483 7939
rect 81483 7905 81492 7939
rect 81440 7896 81492 7905
rect 83832 7939 83884 7948
rect 83832 7905 83841 7939
rect 83841 7905 83875 7939
rect 83875 7905 83884 7939
rect 83832 7896 83884 7905
rect 84108 7939 84160 7948
rect 84108 7905 84117 7939
rect 84117 7905 84151 7939
rect 84151 7905 84160 7939
rect 84108 7896 84160 7905
rect 84844 8032 84896 8084
rect 86684 8007 86736 8016
rect 86684 7973 86693 8007
rect 86693 7973 86727 8007
rect 86727 7973 86736 8007
rect 86684 7964 86736 7973
rect 92848 8032 92900 8084
rect 93584 8032 93636 8084
rect 89444 7939 89496 7948
rect 89444 7905 89453 7939
rect 89453 7905 89487 7939
rect 89487 7905 89496 7939
rect 89444 7896 89496 7905
rect 91192 7896 91244 7948
rect 58348 7692 58400 7744
rect 59176 7692 59228 7744
rect 61936 7760 61988 7812
rect 62672 7760 62724 7812
rect 64788 7692 64840 7744
rect 67640 7760 67692 7812
rect 67732 7692 67784 7744
rect 67916 7692 67968 7744
rect 72424 7871 72476 7880
rect 72424 7837 72433 7871
rect 72433 7837 72467 7871
rect 72467 7837 72476 7871
rect 72424 7828 72476 7837
rect 73160 7828 73212 7880
rect 74908 7871 74960 7880
rect 74908 7837 74917 7871
rect 74917 7837 74951 7871
rect 74951 7837 74960 7871
rect 74908 7828 74960 7837
rect 78680 7828 78732 7880
rect 79876 7828 79928 7880
rect 76472 7760 76524 7812
rect 78588 7760 78640 7812
rect 80060 7828 80112 7880
rect 80520 7828 80572 7880
rect 82636 7871 82688 7880
rect 82636 7837 82645 7871
rect 82645 7837 82679 7871
rect 82679 7837 82688 7871
rect 82636 7828 82688 7837
rect 82820 7828 82872 7880
rect 83648 7871 83700 7880
rect 83648 7837 83657 7871
rect 83657 7837 83691 7871
rect 83691 7837 83700 7871
rect 83648 7828 83700 7837
rect 86132 7828 86184 7880
rect 89720 7871 89772 7880
rect 89720 7837 89729 7871
rect 89729 7837 89763 7871
rect 89763 7837 89772 7871
rect 90456 7871 90508 7880
rect 89720 7828 89772 7837
rect 90456 7837 90465 7871
rect 90465 7837 90499 7871
rect 90499 7837 90508 7871
rect 90456 7828 90508 7837
rect 92480 7896 92532 7948
rect 72424 7692 72476 7744
rect 74632 7692 74684 7744
rect 77668 7692 77720 7744
rect 80428 7692 80480 7744
rect 82176 7760 82228 7812
rect 84844 7760 84896 7812
rect 88432 7760 88484 7812
rect 89260 7760 89312 7812
rect 89628 7760 89680 7812
rect 90824 7760 90876 7812
rect 93400 7828 93452 7880
rect 93032 7760 93084 7812
rect 84384 7692 84436 7744
rect 87236 7735 87288 7744
rect 87236 7701 87245 7735
rect 87245 7701 87279 7735
rect 87279 7701 87288 7735
rect 87236 7692 87288 7701
rect 90732 7692 90784 7744
rect 95148 7692 95200 7744
rect 24386 7590 24438 7642
rect 24450 7590 24502 7642
rect 24514 7590 24566 7642
rect 24578 7590 24630 7642
rect 24642 7590 24694 7642
rect 47823 7590 47875 7642
rect 47887 7590 47939 7642
rect 47951 7590 48003 7642
rect 48015 7590 48067 7642
rect 48079 7590 48131 7642
rect 71260 7590 71312 7642
rect 71324 7590 71376 7642
rect 71388 7590 71440 7642
rect 71452 7590 71504 7642
rect 71516 7590 71568 7642
rect 94697 7590 94749 7642
rect 94761 7590 94813 7642
rect 94825 7590 94877 7642
rect 94889 7590 94941 7642
rect 94953 7590 95005 7642
rect 2228 7463 2280 7472
rect 2228 7429 2237 7463
rect 2237 7429 2271 7463
rect 2271 7429 2280 7463
rect 2228 7420 2280 7429
rect 4068 7420 4120 7472
rect 4436 7463 4488 7472
rect 4436 7429 4445 7463
rect 4445 7429 4479 7463
rect 4479 7429 4488 7463
rect 4436 7420 4488 7429
rect 5724 7488 5776 7540
rect 8208 7488 8260 7540
rect 18328 7531 18380 7540
rect 9588 7463 9640 7472
rect 9588 7429 9597 7463
rect 9597 7429 9631 7463
rect 9631 7429 9640 7463
rect 9588 7420 9640 7429
rect 12992 7420 13044 7472
rect 13728 7463 13780 7472
rect 13728 7429 13737 7463
rect 13737 7429 13771 7463
rect 13771 7429 13780 7463
rect 13728 7420 13780 7429
rect 16304 7420 16356 7472
rect 17316 7420 17368 7472
rect 18328 7497 18337 7531
rect 18337 7497 18371 7531
rect 18371 7497 18380 7531
rect 18328 7488 18380 7497
rect 18696 7488 18748 7540
rect 21824 7488 21876 7540
rect 27528 7531 27580 7540
rect 27528 7497 27537 7531
rect 27537 7497 27571 7531
rect 27571 7497 27580 7531
rect 27528 7488 27580 7497
rect 28448 7531 28500 7540
rect 18880 7420 18932 7472
rect 3700 7327 3752 7336
rect 3700 7293 3709 7327
rect 3709 7293 3743 7327
rect 3743 7293 3752 7327
rect 3700 7284 3752 7293
rect 3976 7284 4028 7336
rect 6828 7352 6880 7404
rect 9496 7352 9548 7404
rect 10048 7395 10100 7404
rect 10048 7361 10057 7395
rect 10057 7361 10091 7395
rect 10091 7361 10100 7395
rect 10048 7352 10100 7361
rect 10692 7352 10744 7404
rect 8300 7191 8352 7200
rect 8300 7157 8309 7191
rect 8309 7157 8343 7191
rect 8343 7157 8352 7191
rect 8300 7148 8352 7157
rect 9680 7148 9732 7200
rect 10784 7148 10836 7200
rect 10968 7148 11020 7200
rect 18236 7395 18288 7404
rect 13728 7284 13780 7336
rect 18236 7361 18245 7395
rect 18245 7361 18279 7395
rect 18279 7361 18288 7395
rect 18236 7352 18288 7361
rect 18604 7352 18656 7404
rect 20076 7420 20128 7472
rect 20996 7420 21048 7472
rect 20260 7352 20312 7404
rect 22284 7420 22336 7472
rect 26148 7463 26200 7472
rect 21272 7352 21324 7404
rect 22468 7284 22520 7336
rect 26148 7429 26157 7463
rect 26157 7429 26191 7463
rect 26191 7429 26200 7463
rect 26148 7420 26200 7429
rect 26240 7420 26292 7472
rect 28448 7497 28457 7531
rect 28457 7497 28491 7531
rect 28491 7497 28500 7531
rect 28448 7488 28500 7497
rect 30748 7488 30800 7540
rect 36544 7488 36596 7540
rect 39856 7488 39908 7540
rect 41604 7488 41656 7540
rect 42432 7488 42484 7540
rect 42984 7531 43036 7540
rect 42984 7497 42993 7531
rect 42993 7497 43027 7531
rect 43027 7497 43036 7531
rect 42984 7488 43036 7497
rect 44364 7488 44416 7540
rect 44916 7488 44968 7540
rect 45468 7531 45520 7540
rect 45468 7497 45477 7531
rect 45477 7497 45511 7531
rect 45511 7497 45520 7531
rect 45468 7488 45520 7497
rect 46572 7531 46624 7540
rect 46572 7497 46581 7531
rect 46581 7497 46615 7531
rect 46615 7497 46624 7531
rect 46572 7488 46624 7497
rect 47308 7488 47360 7540
rect 50344 7488 50396 7540
rect 51356 7488 51408 7540
rect 52276 7488 52328 7540
rect 57704 7488 57756 7540
rect 58624 7488 58676 7540
rect 60556 7531 60608 7540
rect 23664 7352 23716 7404
rect 23112 7327 23164 7336
rect 23112 7293 23121 7327
rect 23121 7293 23155 7327
rect 23155 7293 23164 7327
rect 23112 7284 23164 7293
rect 23388 7284 23440 7336
rect 25136 7352 25188 7404
rect 27712 7395 27764 7404
rect 27712 7361 27721 7395
rect 27721 7361 27755 7395
rect 27755 7361 27764 7395
rect 27712 7352 27764 7361
rect 29644 7420 29696 7472
rect 31760 7420 31812 7472
rect 32404 7463 32456 7472
rect 32404 7429 32413 7463
rect 32413 7429 32447 7463
rect 32447 7429 32456 7463
rect 32404 7420 32456 7429
rect 33140 7463 33192 7472
rect 33140 7429 33149 7463
rect 33149 7429 33183 7463
rect 33183 7429 33192 7463
rect 33140 7420 33192 7429
rect 33600 7420 33652 7472
rect 35808 7395 35860 7404
rect 35808 7361 35817 7395
rect 35817 7361 35851 7395
rect 35851 7361 35860 7395
rect 35808 7352 35860 7361
rect 35900 7352 35952 7404
rect 41512 7420 41564 7472
rect 36728 7352 36780 7404
rect 26608 7284 26660 7336
rect 27160 7284 27212 7336
rect 28724 7284 28776 7336
rect 30196 7327 30248 7336
rect 30196 7293 30205 7327
rect 30205 7293 30239 7327
rect 30239 7293 30248 7327
rect 30196 7284 30248 7293
rect 32864 7327 32916 7336
rect 32864 7293 32873 7327
rect 32873 7293 32907 7327
rect 32907 7293 32916 7327
rect 32864 7284 32916 7293
rect 19340 7148 19392 7200
rect 28632 7216 28684 7268
rect 31668 7216 31720 7268
rect 36636 7284 36688 7336
rect 38108 7352 38160 7404
rect 38844 7352 38896 7404
rect 40132 7395 40184 7404
rect 39028 7327 39080 7336
rect 36544 7216 36596 7268
rect 39028 7293 39037 7327
rect 39037 7293 39071 7327
rect 39071 7293 39080 7327
rect 39028 7284 39080 7293
rect 39396 7216 39448 7268
rect 40132 7361 40141 7395
rect 40141 7361 40175 7395
rect 40175 7361 40184 7395
rect 40132 7352 40184 7361
rect 40592 7284 40644 7336
rect 40132 7216 40184 7268
rect 43076 7420 43128 7472
rect 44088 7420 44140 7472
rect 49700 7420 49752 7472
rect 55864 7420 55916 7472
rect 59360 7420 59412 7472
rect 60556 7497 60565 7531
rect 60565 7497 60599 7531
rect 60599 7497 60608 7531
rect 60556 7488 60608 7497
rect 60832 7531 60884 7540
rect 60832 7497 60841 7531
rect 60841 7497 60875 7531
rect 60875 7497 60884 7531
rect 60832 7488 60884 7497
rect 61568 7488 61620 7540
rect 63040 7488 63092 7540
rect 63500 7463 63552 7472
rect 63500 7429 63509 7463
rect 63509 7429 63543 7463
rect 63543 7429 63552 7463
rect 63500 7420 63552 7429
rect 67548 7488 67600 7540
rect 67640 7488 67692 7540
rect 68008 7488 68060 7540
rect 42432 7352 42484 7404
rect 40868 7327 40920 7336
rect 40868 7293 40877 7327
rect 40877 7293 40911 7327
rect 40911 7293 40920 7327
rect 40868 7284 40920 7293
rect 40960 7327 41012 7336
rect 40960 7293 40969 7327
rect 40969 7293 41003 7327
rect 41003 7293 41012 7327
rect 40960 7284 41012 7293
rect 41236 7284 41288 7336
rect 41604 7284 41656 7336
rect 46572 7352 46624 7404
rect 49148 7395 49200 7404
rect 49148 7361 49157 7395
rect 49157 7361 49191 7395
rect 49191 7361 49200 7395
rect 49148 7352 49200 7361
rect 49516 7352 49568 7404
rect 52092 7395 52144 7404
rect 43076 7284 43128 7336
rect 43444 7284 43496 7336
rect 47308 7284 47360 7336
rect 49332 7284 49384 7336
rect 52092 7361 52101 7395
rect 52101 7361 52135 7395
rect 52135 7361 52144 7395
rect 52092 7352 52144 7361
rect 53564 7395 53616 7404
rect 51632 7327 51684 7336
rect 51632 7293 51641 7327
rect 51641 7293 51675 7327
rect 51675 7293 51684 7327
rect 51632 7284 51684 7293
rect 52184 7284 52236 7336
rect 41880 7259 41932 7268
rect 41880 7225 41889 7259
rect 41889 7225 41923 7259
rect 41923 7225 41932 7259
rect 41880 7216 41932 7225
rect 42064 7216 42116 7268
rect 45560 7216 45612 7268
rect 22468 7148 22520 7200
rect 23388 7148 23440 7200
rect 23664 7191 23716 7200
rect 23664 7157 23673 7191
rect 23673 7157 23707 7191
rect 23707 7157 23716 7191
rect 23664 7148 23716 7157
rect 24216 7191 24268 7200
rect 24216 7157 24225 7191
rect 24225 7157 24259 7191
rect 24259 7157 24268 7191
rect 24216 7148 24268 7157
rect 25136 7148 25188 7200
rect 27252 7148 27304 7200
rect 28080 7148 28132 7200
rect 28908 7148 28960 7200
rect 32772 7148 32824 7200
rect 33784 7148 33836 7200
rect 33876 7148 33928 7200
rect 35808 7148 35860 7200
rect 37648 7148 37700 7200
rect 37832 7148 37884 7200
rect 38292 7148 38344 7200
rect 38844 7148 38896 7200
rect 39856 7148 39908 7200
rect 41144 7148 41196 7200
rect 41972 7191 42024 7200
rect 41972 7157 41981 7191
rect 41981 7157 42015 7191
rect 42015 7157 42024 7191
rect 41972 7148 42024 7157
rect 44916 7191 44968 7200
rect 44916 7157 44925 7191
rect 44925 7157 44959 7191
rect 44959 7157 44968 7191
rect 44916 7148 44968 7157
rect 45468 7148 45520 7200
rect 48228 7216 48280 7268
rect 45744 7148 45796 7200
rect 48688 7216 48740 7268
rect 51816 7216 51868 7268
rect 52092 7216 52144 7268
rect 53564 7361 53573 7395
rect 53573 7361 53607 7395
rect 53607 7361 53616 7395
rect 53564 7352 53616 7361
rect 57244 7395 57296 7404
rect 57244 7361 57253 7395
rect 57253 7361 57287 7395
rect 57287 7361 57296 7395
rect 57244 7352 57296 7361
rect 58072 7395 58124 7404
rect 58072 7361 58081 7395
rect 58081 7361 58115 7395
rect 58115 7361 58124 7395
rect 58072 7352 58124 7361
rect 53656 7148 53708 7200
rect 54208 7284 54260 7336
rect 54852 7327 54904 7336
rect 54852 7293 54861 7327
rect 54861 7293 54895 7327
rect 54895 7293 54904 7327
rect 54852 7284 54904 7293
rect 54944 7284 54996 7336
rect 60464 7284 60516 7336
rect 55956 7216 56008 7268
rect 59360 7216 59412 7268
rect 61936 7352 61988 7404
rect 62672 7395 62724 7404
rect 62672 7361 62681 7395
rect 62681 7361 62715 7395
rect 62715 7361 62724 7395
rect 62672 7352 62724 7361
rect 63868 7395 63920 7404
rect 63868 7361 63877 7395
rect 63877 7361 63911 7395
rect 63911 7361 63920 7395
rect 63868 7352 63920 7361
rect 64512 7352 64564 7404
rect 64696 7352 64748 7404
rect 61568 7327 61620 7336
rect 61568 7293 61577 7327
rect 61577 7293 61611 7327
rect 61611 7293 61620 7327
rect 61568 7284 61620 7293
rect 60924 7216 60976 7268
rect 61108 7259 61160 7268
rect 61108 7225 61117 7259
rect 61117 7225 61151 7259
rect 61151 7225 61160 7259
rect 61108 7216 61160 7225
rect 62120 7216 62172 7268
rect 64144 7284 64196 7336
rect 65340 7284 65392 7336
rect 65616 7395 65668 7404
rect 65616 7361 65625 7395
rect 65625 7361 65659 7395
rect 65659 7361 65668 7395
rect 65616 7352 65668 7361
rect 66352 7352 66404 7404
rect 74356 7488 74408 7540
rect 71964 7420 72016 7472
rect 72424 7420 72476 7472
rect 66720 7352 66772 7404
rect 67456 7352 67508 7404
rect 68100 7352 68152 7404
rect 69572 7395 69624 7404
rect 69572 7361 69581 7395
rect 69581 7361 69615 7395
rect 69615 7361 69624 7395
rect 69572 7352 69624 7361
rect 74816 7488 74868 7540
rect 76104 7488 76156 7540
rect 76380 7420 76432 7472
rect 76012 7395 76064 7404
rect 76012 7361 76021 7395
rect 76021 7361 76055 7395
rect 76055 7361 76064 7395
rect 76012 7352 76064 7361
rect 76288 7395 76340 7404
rect 76288 7361 76297 7395
rect 76297 7361 76331 7395
rect 76331 7361 76340 7395
rect 76288 7352 76340 7361
rect 76656 7488 76708 7540
rect 78128 7531 78180 7540
rect 78128 7497 78137 7531
rect 78137 7497 78171 7531
rect 78171 7497 78180 7531
rect 78128 7488 78180 7497
rect 78680 7488 78732 7540
rect 77668 7395 77720 7404
rect 77668 7361 77677 7395
rect 77677 7361 77711 7395
rect 77711 7361 77720 7395
rect 77668 7352 77720 7361
rect 77944 7395 77996 7404
rect 77944 7361 77953 7395
rect 77953 7361 77987 7395
rect 77987 7361 77996 7395
rect 77944 7352 77996 7361
rect 78680 7395 78732 7404
rect 78680 7361 78689 7395
rect 78689 7361 78723 7395
rect 78723 7361 78732 7395
rect 78680 7352 78732 7361
rect 78864 7395 78916 7404
rect 78864 7361 78873 7395
rect 78873 7361 78907 7395
rect 78907 7361 78916 7395
rect 78864 7352 78916 7361
rect 80336 7352 80388 7404
rect 67364 7327 67416 7336
rect 67364 7293 67373 7327
rect 67373 7293 67407 7327
rect 67407 7293 67416 7327
rect 68652 7327 68704 7336
rect 67364 7284 67416 7293
rect 68652 7293 68661 7327
rect 68661 7293 68695 7327
rect 68695 7293 68704 7327
rect 68652 7284 68704 7293
rect 68836 7284 68888 7336
rect 56416 7148 56468 7200
rect 62488 7148 62540 7200
rect 67088 7216 67140 7268
rect 65156 7148 65208 7200
rect 66628 7191 66680 7200
rect 66628 7157 66637 7191
rect 66637 7157 66671 7191
rect 66671 7157 66680 7191
rect 66628 7148 66680 7157
rect 67272 7148 67324 7200
rect 68284 7148 68336 7200
rect 68468 7191 68520 7200
rect 68468 7157 68477 7191
rect 68477 7157 68511 7191
rect 68511 7157 68520 7191
rect 68468 7148 68520 7157
rect 73528 7327 73580 7336
rect 73528 7293 73537 7327
rect 73537 7293 73571 7327
rect 73571 7293 73580 7327
rect 73528 7284 73580 7293
rect 74632 7327 74684 7336
rect 74632 7293 74641 7327
rect 74641 7293 74675 7327
rect 74675 7293 74684 7327
rect 74632 7284 74684 7293
rect 82636 7488 82688 7540
rect 83280 7488 83332 7540
rect 80704 7463 80756 7472
rect 80704 7429 80713 7463
rect 80713 7429 80747 7463
rect 80747 7429 80756 7463
rect 80704 7420 80756 7429
rect 81348 7420 81400 7472
rect 83280 7395 83332 7404
rect 83280 7361 83289 7395
rect 83289 7361 83323 7395
rect 83323 7361 83332 7395
rect 83280 7352 83332 7361
rect 84476 7395 84528 7404
rect 74540 7216 74592 7268
rect 81624 7284 81676 7336
rect 81716 7327 81768 7336
rect 81716 7293 81725 7327
rect 81725 7293 81759 7327
rect 81759 7293 81768 7327
rect 81716 7284 81768 7293
rect 71964 7148 72016 7200
rect 84200 7216 84252 7268
rect 84476 7361 84485 7395
rect 84485 7361 84519 7395
rect 84519 7361 84528 7395
rect 84476 7352 84528 7361
rect 85488 7488 85540 7540
rect 85948 7488 86000 7540
rect 86592 7531 86644 7540
rect 86592 7497 86601 7531
rect 86601 7497 86635 7531
rect 86635 7497 86644 7531
rect 86592 7488 86644 7497
rect 92848 7488 92900 7540
rect 88340 7420 88392 7472
rect 89168 7463 89220 7472
rect 89168 7429 89177 7463
rect 89177 7429 89211 7463
rect 89211 7429 89220 7463
rect 89168 7420 89220 7429
rect 90456 7420 90508 7472
rect 86040 7352 86092 7404
rect 85028 7284 85080 7336
rect 87144 7284 87196 7336
rect 84660 7216 84712 7268
rect 88432 7352 88484 7404
rect 91008 7352 91060 7404
rect 93032 7420 93084 7472
rect 88892 7284 88944 7336
rect 89076 7216 89128 7268
rect 90180 7284 90232 7336
rect 92940 7395 92992 7404
rect 92940 7361 92949 7395
rect 92949 7361 92983 7395
rect 92983 7361 92992 7395
rect 92940 7352 92992 7361
rect 89720 7216 89772 7268
rect 76472 7148 76524 7200
rect 79876 7191 79928 7200
rect 79876 7157 79885 7191
rect 79885 7157 79919 7191
rect 79919 7157 79928 7191
rect 79876 7148 79928 7157
rect 80060 7191 80112 7200
rect 80060 7157 80069 7191
rect 80069 7157 80103 7191
rect 80103 7157 80112 7191
rect 82820 7191 82872 7200
rect 80060 7148 80112 7157
rect 82820 7157 82829 7191
rect 82829 7157 82863 7191
rect 82863 7157 82872 7191
rect 82820 7148 82872 7157
rect 89812 7148 89864 7200
rect 92756 7148 92808 7200
rect 12668 7046 12720 7098
rect 12732 7046 12784 7098
rect 12796 7046 12848 7098
rect 12860 7046 12912 7098
rect 12924 7046 12976 7098
rect 36105 7046 36157 7098
rect 36169 7046 36221 7098
rect 36233 7046 36285 7098
rect 36297 7046 36349 7098
rect 36361 7046 36413 7098
rect 59542 7046 59594 7098
rect 59606 7046 59658 7098
rect 59670 7046 59722 7098
rect 59734 7046 59786 7098
rect 59798 7046 59850 7098
rect 82979 7046 83031 7098
rect 83043 7046 83095 7098
rect 83107 7046 83159 7098
rect 83171 7046 83223 7098
rect 83235 7046 83287 7098
rect 4252 6851 4304 6860
rect 4252 6817 4261 6851
rect 4261 6817 4295 6851
rect 4295 6817 4304 6851
rect 4252 6808 4304 6817
rect 5172 6808 5224 6860
rect 9680 6808 9732 6860
rect 9864 6808 9916 6860
rect 12348 6944 12400 6996
rect 10692 6876 10744 6928
rect 13728 6944 13780 6996
rect 20904 6944 20956 6996
rect 22284 6944 22336 6996
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 6920 6740 6972 6792
rect 4160 6604 4212 6656
rect 6736 6672 6788 6724
rect 7564 6740 7616 6792
rect 8116 6783 8168 6792
rect 8116 6749 8125 6783
rect 8125 6749 8159 6783
rect 8159 6749 8168 6783
rect 8116 6740 8168 6749
rect 8300 6672 8352 6724
rect 8576 6672 8628 6724
rect 5080 6647 5132 6656
rect 5080 6613 5089 6647
rect 5089 6613 5123 6647
rect 5123 6613 5132 6647
rect 5080 6604 5132 6613
rect 6644 6647 6696 6656
rect 6644 6613 6653 6647
rect 6653 6613 6687 6647
rect 6687 6613 6696 6647
rect 6644 6604 6696 6613
rect 10140 6604 10192 6656
rect 10784 6740 10836 6792
rect 16948 6876 17000 6928
rect 17960 6876 18012 6928
rect 18236 6876 18288 6928
rect 22192 6876 22244 6928
rect 25136 6944 25188 6996
rect 28080 6987 28132 6996
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 10508 6672 10560 6724
rect 15016 6740 15068 6792
rect 15292 6783 15344 6792
rect 15292 6749 15301 6783
rect 15301 6749 15335 6783
rect 15335 6749 15344 6783
rect 15292 6740 15344 6749
rect 17316 6740 17368 6792
rect 10416 6604 10468 6656
rect 13636 6604 13688 6656
rect 17960 6672 18012 6724
rect 20444 6808 20496 6860
rect 20536 6808 20588 6860
rect 23020 6783 23072 6792
rect 22100 6672 22152 6724
rect 22744 6715 22796 6724
rect 22744 6681 22753 6715
rect 22753 6681 22787 6715
rect 22787 6681 22796 6715
rect 22744 6672 22796 6681
rect 23020 6749 23029 6783
rect 23029 6749 23063 6783
rect 23063 6749 23072 6783
rect 23020 6740 23072 6749
rect 24860 6851 24912 6860
rect 24860 6817 24869 6851
rect 24869 6817 24903 6851
rect 24903 6817 24912 6851
rect 24860 6808 24912 6817
rect 23756 6740 23808 6792
rect 26332 6808 26384 6860
rect 28080 6953 28089 6987
rect 28089 6953 28123 6987
rect 28123 6953 28132 6987
rect 28080 6944 28132 6953
rect 28448 6944 28500 6996
rect 34060 6944 34112 6996
rect 35164 6987 35216 6996
rect 35164 6953 35194 6987
rect 35194 6953 35216 6987
rect 35164 6944 35216 6953
rect 35256 6944 35308 6996
rect 37004 6944 37056 6996
rect 37832 6987 37884 6996
rect 37832 6953 37841 6987
rect 37841 6953 37875 6987
rect 37875 6953 37884 6987
rect 37832 6944 37884 6953
rect 39028 6944 39080 6996
rect 40776 6944 40828 6996
rect 41512 6944 41564 6996
rect 45744 6944 45796 6996
rect 26700 6876 26752 6928
rect 31208 6876 31260 6928
rect 28448 6808 28500 6860
rect 29460 6808 29512 6860
rect 30196 6808 30248 6860
rect 32864 6876 32916 6928
rect 33140 6808 33192 6860
rect 33416 6851 33468 6860
rect 33416 6817 33425 6851
rect 33425 6817 33459 6851
rect 33459 6817 33468 6851
rect 33416 6808 33468 6817
rect 34152 6919 34204 6928
rect 34152 6885 34161 6919
rect 34161 6885 34195 6919
rect 34195 6885 34204 6919
rect 34152 6876 34204 6885
rect 36176 6876 36228 6928
rect 37372 6876 37424 6928
rect 38016 6876 38068 6928
rect 34888 6851 34940 6860
rect 34888 6817 34897 6851
rect 34897 6817 34931 6851
rect 34931 6817 34940 6851
rect 34888 6808 34940 6817
rect 35808 6808 35860 6860
rect 37280 6851 37332 6860
rect 30104 6740 30156 6792
rect 33324 6783 33376 6792
rect 33324 6749 33333 6783
rect 33333 6749 33367 6783
rect 33367 6749 33376 6783
rect 33324 6740 33376 6749
rect 33784 6740 33836 6792
rect 34704 6740 34756 6792
rect 37280 6817 37289 6851
rect 37289 6817 37323 6851
rect 37323 6817 37332 6851
rect 37280 6808 37332 6817
rect 38476 6851 38528 6860
rect 38476 6817 38485 6851
rect 38485 6817 38519 6851
rect 38519 6817 38528 6851
rect 38476 6808 38528 6817
rect 38844 6808 38896 6860
rect 40224 6876 40276 6928
rect 40868 6876 40920 6928
rect 41236 6876 41288 6928
rect 43076 6876 43128 6928
rect 40040 6851 40092 6860
rect 39028 6740 39080 6792
rect 40040 6817 40049 6851
rect 40049 6817 40083 6851
rect 40083 6817 40092 6851
rect 40040 6808 40092 6817
rect 41972 6808 42024 6860
rect 42892 6851 42944 6860
rect 42892 6817 42901 6851
rect 42901 6817 42935 6851
rect 42935 6817 42944 6851
rect 42892 6808 42944 6817
rect 25596 6715 25648 6724
rect 18236 6647 18288 6656
rect 18236 6613 18245 6647
rect 18245 6613 18279 6647
rect 18279 6613 18288 6647
rect 18236 6604 18288 6613
rect 22928 6604 22980 6656
rect 23388 6604 23440 6656
rect 24124 6604 24176 6656
rect 25596 6681 25605 6715
rect 25605 6681 25639 6715
rect 25639 6681 25648 6715
rect 25596 6672 25648 6681
rect 26240 6672 26292 6724
rect 28172 6672 28224 6724
rect 30472 6715 30524 6724
rect 28724 6647 28776 6656
rect 28724 6613 28749 6647
rect 28749 6613 28776 6647
rect 28724 6604 28776 6613
rect 29736 6604 29788 6656
rect 30472 6681 30481 6715
rect 30481 6681 30515 6715
rect 30515 6681 30524 6715
rect 30472 6672 30524 6681
rect 31668 6672 31720 6724
rect 33048 6672 33100 6724
rect 33876 6672 33928 6724
rect 34244 6715 34296 6724
rect 34244 6681 34253 6715
rect 34253 6681 34287 6715
rect 34287 6681 34296 6715
rect 34244 6672 34296 6681
rect 34520 6672 34572 6724
rect 35624 6672 35676 6724
rect 40776 6740 40828 6792
rect 41144 6783 41196 6792
rect 41144 6749 41153 6783
rect 41153 6749 41187 6783
rect 41187 6749 41196 6783
rect 41144 6740 41196 6749
rect 33416 6604 33468 6656
rect 34888 6604 34940 6656
rect 36728 6604 36780 6656
rect 38936 6604 38988 6656
rect 39304 6647 39356 6656
rect 39304 6613 39313 6647
rect 39313 6613 39347 6647
rect 39347 6613 39356 6647
rect 39304 6604 39356 6613
rect 40316 6672 40368 6724
rect 40868 6672 40920 6724
rect 43444 6808 43496 6860
rect 44640 6851 44692 6860
rect 44640 6817 44649 6851
rect 44649 6817 44683 6851
rect 44683 6817 44692 6851
rect 44640 6808 44692 6817
rect 44916 6808 44968 6860
rect 45836 6808 45888 6860
rect 49608 6944 49660 6996
rect 53288 6944 53340 6996
rect 54852 6944 54904 6996
rect 58532 6987 58584 6996
rect 58532 6953 58541 6987
rect 58541 6953 58575 6987
rect 58575 6953 58584 6987
rect 58532 6944 58584 6953
rect 61108 6944 61160 6996
rect 51908 6876 51960 6928
rect 56784 6876 56836 6928
rect 48780 6851 48832 6860
rect 43076 6740 43128 6792
rect 45284 6783 45336 6792
rect 45284 6749 45293 6783
rect 45293 6749 45327 6783
rect 45327 6749 45336 6783
rect 48780 6817 48789 6851
rect 48789 6817 48823 6851
rect 48823 6817 48832 6851
rect 48780 6808 48832 6817
rect 50068 6808 50120 6860
rect 50344 6851 50396 6860
rect 50344 6817 50353 6851
rect 50353 6817 50387 6851
rect 50387 6817 50396 6851
rect 50344 6808 50396 6817
rect 50988 6808 51040 6860
rect 53472 6808 53524 6860
rect 56416 6851 56468 6860
rect 45284 6740 45336 6749
rect 43168 6672 43220 6724
rect 43352 6672 43404 6724
rect 44640 6672 44692 6724
rect 49148 6672 49200 6724
rect 49516 6783 49568 6792
rect 49516 6749 49525 6783
rect 49525 6749 49559 6783
rect 49559 6749 49568 6783
rect 49516 6740 49568 6749
rect 53656 6740 53708 6792
rect 42432 6647 42484 6656
rect 42432 6613 42441 6647
rect 42441 6613 42475 6647
rect 42475 6613 42484 6647
rect 42432 6604 42484 6613
rect 42892 6604 42944 6656
rect 44916 6604 44968 6656
rect 45468 6647 45520 6656
rect 45468 6613 45477 6647
rect 45477 6613 45511 6647
rect 45511 6613 45520 6647
rect 45468 6604 45520 6613
rect 47308 6604 47360 6656
rect 49700 6647 49752 6656
rect 49700 6613 49709 6647
rect 49709 6613 49743 6647
rect 49743 6613 49752 6647
rect 49700 6604 49752 6613
rect 52920 6672 52972 6724
rect 51632 6604 51684 6656
rect 53564 6604 53616 6656
rect 56416 6817 56425 6851
rect 56425 6817 56459 6851
rect 56459 6817 56468 6851
rect 56416 6808 56468 6817
rect 56508 6808 56560 6860
rect 60648 6808 60700 6860
rect 60924 6808 60976 6860
rect 65156 6944 65208 6996
rect 67824 6944 67876 6996
rect 68468 6944 68520 6996
rect 68744 6944 68796 6996
rect 72976 6944 73028 6996
rect 77944 6944 77996 6996
rect 79968 6944 80020 6996
rect 80336 6944 80388 6996
rect 68284 6876 68336 6928
rect 69204 6876 69256 6928
rect 62488 6808 62540 6860
rect 62948 6851 63000 6860
rect 62948 6817 62957 6851
rect 62957 6817 62991 6851
rect 62991 6817 63000 6851
rect 62948 6808 63000 6817
rect 57244 6740 57296 6792
rect 59452 6740 59504 6792
rect 59912 6740 59964 6792
rect 60004 6740 60056 6792
rect 60280 6740 60332 6792
rect 60832 6783 60884 6792
rect 60832 6749 60841 6783
rect 60841 6749 60875 6783
rect 60875 6749 60884 6783
rect 60832 6740 60884 6749
rect 61016 6740 61068 6792
rect 61660 6740 61712 6792
rect 61936 6783 61988 6792
rect 61936 6749 61945 6783
rect 61945 6749 61979 6783
rect 61979 6749 61988 6783
rect 61936 6740 61988 6749
rect 62120 6783 62172 6792
rect 62120 6749 62129 6783
rect 62129 6749 62163 6783
rect 62163 6749 62172 6783
rect 62120 6740 62172 6749
rect 63224 6808 63276 6860
rect 65156 6808 65208 6860
rect 65432 6808 65484 6860
rect 68652 6808 68704 6860
rect 69296 6851 69348 6860
rect 69296 6817 69305 6851
rect 69305 6817 69339 6851
rect 69339 6817 69348 6851
rect 69296 6808 69348 6817
rect 74356 6808 74408 6860
rect 78036 6876 78088 6928
rect 80520 6876 80572 6928
rect 63500 6783 63552 6792
rect 63500 6749 63509 6783
rect 63509 6749 63543 6783
rect 63543 6749 63552 6783
rect 63500 6740 63552 6749
rect 64880 6740 64932 6792
rect 56968 6715 57020 6724
rect 56968 6681 56977 6715
rect 56977 6681 57011 6715
rect 57011 6681 57020 6715
rect 56968 6672 57020 6681
rect 61108 6672 61160 6724
rect 59544 6604 59596 6656
rect 60004 6647 60056 6656
rect 60004 6613 60013 6647
rect 60013 6613 60047 6647
rect 60047 6613 60056 6647
rect 60004 6604 60056 6613
rect 61660 6647 61712 6656
rect 61660 6613 61669 6647
rect 61669 6613 61703 6647
rect 61703 6613 61712 6647
rect 61660 6604 61712 6613
rect 65432 6672 65484 6724
rect 66812 6740 66864 6792
rect 68192 6783 68244 6792
rect 68192 6749 68201 6783
rect 68201 6749 68235 6783
rect 68235 6749 68244 6783
rect 68192 6740 68244 6749
rect 70308 6740 70360 6792
rect 71136 6740 71188 6792
rect 74540 6783 74592 6792
rect 74540 6749 74549 6783
rect 74549 6749 74583 6783
rect 74583 6749 74592 6783
rect 74540 6740 74592 6749
rect 66076 6672 66128 6724
rect 65248 6604 65300 6656
rect 67640 6604 67692 6656
rect 71872 6672 71924 6724
rect 72056 6672 72108 6724
rect 73160 6672 73212 6724
rect 70400 6647 70452 6656
rect 70400 6613 70409 6647
rect 70409 6613 70443 6647
rect 70443 6613 70452 6647
rect 70400 6604 70452 6613
rect 70676 6604 70728 6656
rect 70768 6604 70820 6656
rect 72424 6604 72476 6656
rect 75184 6740 75236 6792
rect 75460 6783 75512 6792
rect 75460 6749 75469 6783
rect 75469 6749 75503 6783
rect 75503 6749 75512 6783
rect 75460 6740 75512 6749
rect 78864 6808 78916 6860
rect 80428 6851 80480 6860
rect 80428 6817 80437 6851
rect 80437 6817 80471 6851
rect 80471 6817 80480 6851
rect 80428 6808 80480 6817
rect 82636 6944 82688 6996
rect 83648 6944 83700 6996
rect 84016 6944 84068 6996
rect 84476 6944 84528 6996
rect 88432 6944 88484 6996
rect 84108 6876 84160 6928
rect 85028 6876 85080 6928
rect 87144 6876 87196 6928
rect 87972 6876 88024 6928
rect 89720 6944 89772 6996
rect 90180 6944 90232 6996
rect 92848 6944 92900 6996
rect 93768 6944 93820 6996
rect 82544 6808 82596 6860
rect 87236 6808 87288 6860
rect 75644 6672 75696 6724
rect 76932 6740 76984 6792
rect 77300 6783 77352 6792
rect 77300 6749 77309 6783
rect 77309 6749 77343 6783
rect 77343 6749 77352 6783
rect 77300 6740 77352 6749
rect 77760 6740 77812 6792
rect 78956 6740 79008 6792
rect 79784 6740 79836 6792
rect 80336 6783 80388 6792
rect 80336 6749 80345 6783
rect 80345 6749 80379 6783
rect 80379 6749 80388 6783
rect 80336 6740 80388 6749
rect 81624 6783 81676 6792
rect 81624 6749 81633 6783
rect 81633 6749 81667 6783
rect 81667 6749 81676 6783
rect 81624 6740 81676 6749
rect 82176 6783 82228 6792
rect 82176 6749 82185 6783
rect 82185 6749 82219 6783
rect 82219 6749 82228 6783
rect 82176 6740 82228 6749
rect 84384 6783 84436 6792
rect 84384 6749 84393 6783
rect 84393 6749 84427 6783
rect 84427 6749 84436 6783
rect 84384 6740 84436 6749
rect 84568 6740 84620 6792
rect 86684 6740 86736 6792
rect 86960 6740 87012 6792
rect 88248 6808 88300 6860
rect 89812 6876 89864 6928
rect 90732 6876 90784 6928
rect 89444 6808 89496 6860
rect 92388 6851 92440 6860
rect 92388 6817 92397 6851
rect 92397 6817 92431 6851
rect 92431 6817 92440 6851
rect 92388 6808 92440 6817
rect 87420 6740 87472 6792
rect 89076 6740 89128 6792
rect 89628 6783 89680 6792
rect 89628 6749 89637 6783
rect 89637 6749 89671 6783
rect 89671 6749 89680 6783
rect 89628 6740 89680 6749
rect 89904 6740 89956 6792
rect 94044 6808 94096 6860
rect 93860 6740 93912 6792
rect 76748 6715 76800 6724
rect 76748 6681 76757 6715
rect 76757 6681 76791 6715
rect 76791 6681 76800 6715
rect 76748 6672 76800 6681
rect 78496 6672 78548 6724
rect 81716 6672 81768 6724
rect 74632 6604 74684 6656
rect 76472 6647 76524 6656
rect 76472 6613 76481 6647
rect 76481 6613 76515 6647
rect 76515 6613 76524 6647
rect 76472 6604 76524 6613
rect 76564 6647 76616 6656
rect 76564 6613 76573 6647
rect 76573 6613 76607 6647
rect 76607 6613 76616 6647
rect 76564 6604 76616 6613
rect 76840 6604 76892 6656
rect 79876 6604 79928 6656
rect 82544 6604 82596 6656
rect 83832 6672 83884 6724
rect 84108 6672 84160 6724
rect 88892 6672 88944 6724
rect 84016 6604 84068 6656
rect 86960 6604 87012 6656
rect 87052 6604 87104 6656
rect 93124 6672 93176 6724
rect 90732 6604 90784 6656
rect 92756 6604 92808 6656
rect 24386 6502 24438 6554
rect 24450 6502 24502 6554
rect 24514 6502 24566 6554
rect 24578 6502 24630 6554
rect 24642 6502 24694 6554
rect 47823 6502 47875 6554
rect 47887 6502 47939 6554
rect 47951 6502 48003 6554
rect 48015 6502 48067 6554
rect 48079 6502 48131 6554
rect 71260 6502 71312 6554
rect 71324 6502 71376 6554
rect 71388 6502 71440 6554
rect 71452 6502 71504 6554
rect 71516 6502 71568 6554
rect 94697 6502 94749 6554
rect 94761 6502 94813 6554
rect 94825 6502 94877 6554
rect 94889 6502 94941 6554
rect 94953 6502 95005 6554
rect 4252 6400 4304 6452
rect 5080 6400 5132 6452
rect 5172 6400 5224 6452
rect 10508 6400 10560 6452
rect 15016 6443 15068 6452
rect 15016 6409 15025 6443
rect 15025 6409 15059 6443
rect 15059 6409 15068 6443
rect 15016 6400 15068 6409
rect 17960 6443 18012 6452
rect 17960 6409 17969 6443
rect 17969 6409 18003 6443
rect 18003 6409 18012 6443
rect 17960 6400 18012 6409
rect 19432 6443 19484 6452
rect 6644 6332 6696 6384
rect 7564 6332 7616 6384
rect 8116 6264 8168 6316
rect 8392 6264 8444 6316
rect 9680 6264 9732 6316
rect 9864 6307 9916 6316
rect 9864 6273 9873 6307
rect 9873 6273 9907 6307
rect 9907 6273 9916 6307
rect 9864 6264 9916 6273
rect 10140 6307 10192 6316
rect 10140 6273 10149 6307
rect 10149 6273 10183 6307
rect 10183 6273 10192 6307
rect 10140 6264 10192 6273
rect 5724 6196 5776 6248
rect 10600 6264 10652 6316
rect 10784 6307 10836 6316
rect 10784 6273 10793 6307
rect 10793 6273 10827 6307
rect 10827 6273 10836 6307
rect 10784 6264 10836 6273
rect 14832 6264 14884 6316
rect 19432 6409 19441 6443
rect 19441 6409 19475 6443
rect 19475 6409 19484 6443
rect 19432 6400 19484 6409
rect 20536 6443 20588 6452
rect 20536 6409 20545 6443
rect 20545 6409 20579 6443
rect 20579 6409 20588 6443
rect 20536 6400 20588 6409
rect 19248 6332 19300 6384
rect 20904 6332 20956 6384
rect 10692 6196 10744 6248
rect 10784 6128 10836 6180
rect 12624 6128 12676 6180
rect 17960 6196 18012 6248
rect 19708 6264 19760 6316
rect 19248 6128 19300 6180
rect 20444 6264 20496 6316
rect 22192 6400 22244 6452
rect 22744 6400 22796 6452
rect 22652 6332 22704 6384
rect 21180 6264 21232 6316
rect 23204 6264 23256 6316
rect 28172 6400 28224 6452
rect 25228 6332 25280 6384
rect 25596 6332 25648 6384
rect 26424 6332 26476 6384
rect 32312 6400 32364 6452
rect 33324 6400 33376 6452
rect 39304 6443 39356 6452
rect 29736 6332 29788 6384
rect 33140 6375 33192 6384
rect 23020 6196 23072 6248
rect 26516 6264 26568 6316
rect 24216 6196 24268 6248
rect 24768 6196 24820 6248
rect 25136 6239 25188 6248
rect 8576 6060 8628 6112
rect 10416 6060 10468 6112
rect 18512 6103 18564 6112
rect 18512 6069 18521 6103
rect 18521 6069 18555 6103
rect 18555 6069 18564 6103
rect 18512 6060 18564 6069
rect 19616 6060 19668 6112
rect 22744 6128 22796 6180
rect 22836 6060 22888 6112
rect 23756 6103 23808 6112
rect 23756 6069 23765 6103
rect 23765 6069 23799 6103
rect 23799 6069 23808 6103
rect 23756 6060 23808 6069
rect 24308 6060 24360 6112
rect 25136 6205 25145 6239
rect 25145 6205 25179 6239
rect 25179 6205 25188 6239
rect 25136 6196 25188 6205
rect 25872 6196 25924 6248
rect 26240 6128 26292 6180
rect 30196 6264 30248 6316
rect 30748 6196 30800 6248
rect 33140 6341 33149 6375
rect 33149 6341 33183 6375
rect 33183 6341 33192 6375
rect 33140 6332 33192 6341
rect 33232 6332 33284 6384
rect 33600 6332 33652 6384
rect 34888 6375 34940 6384
rect 34888 6341 34897 6375
rect 34897 6341 34931 6375
rect 34931 6341 34940 6375
rect 34888 6332 34940 6341
rect 32496 6264 32548 6316
rect 32864 6307 32916 6316
rect 32864 6273 32873 6307
rect 32873 6273 32907 6307
rect 32907 6273 32916 6307
rect 32864 6264 32916 6273
rect 34704 6264 34756 6316
rect 35624 6196 35676 6248
rect 35900 6264 35952 6316
rect 39304 6409 39313 6443
rect 39313 6409 39347 6443
rect 39347 6409 39356 6443
rect 39304 6400 39356 6409
rect 40224 6443 40276 6452
rect 40224 6409 40233 6443
rect 40233 6409 40267 6443
rect 40267 6409 40276 6443
rect 40224 6400 40276 6409
rect 41236 6400 41288 6452
rect 44732 6400 44784 6452
rect 45192 6443 45244 6452
rect 45192 6409 45201 6443
rect 45201 6409 45235 6443
rect 45235 6409 45244 6443
rect 45192 6400 45244 6409
rect 46388 6400 46440 6452
rect 48136 6400 48188 6452
rect 38016 6307 38068 6316
rect 38016 6273 38025 6307
rect 38025 6273 38059 6307
rect 38059 6273 38068 6307
rect 38016 6264 38068 6273
rect 38568 6264 38620 6316
rect 40132 6307 40184 6316
rect 37924 6239 37976 6248
rect 37924 6205 37933 6239
rect 37933 6205 37967 6239
rect 37967 6205 37976 6239
rect 37924 6196 37976 6205
rect 39028 6196 39080 6248
rect 40132 6273 40141 6307
rect 40141 6273 40175 6307
rect 40175 6273 40184 6307
rect 40132 6264 40184 6273
rect 40316 6307 40368 6316
rect 40316 6273 40325 6307
rect 40325 6273 40359 6307
rect 40359 6273 40368 6307
rect 40316 6264 40368 6273
rect 48044 6332 48096 6384
rect 30104 6128 30156 6180
rect 32680 6128 32732 6180
rect 34244 6128 34296 6180
rect 35348 6171 35400 6180
rect 35348 6137 35357 6171
rect 35357 6137 35391 6171
rect 35391 6137 35400 6171
rect 35348 6128 35400 6137
rect 44180 6264 44232 6316
rect 44548 6307 44600 6316
rect 44548 6273 44557 6307
rect 44557 6273 44591 6307
rect 44591 6273 44600 6307
rect 44548 6264 44600 6273
rect 45560 6307 45612 6316
rect 45560 6273 45569 6307
rect 45569 6273 45603 6307
rect 45603 6273 45612 6307
rect 45560 6264 45612 6273
rect 46204 6307 46256 6316
rect 46204 6273 46213 6307
rect 46213 6273 46247 6307
rect 46247 6273 46256 6307
rect 46204 6264 46256 6273
rect 40960 6128 41012 6180
rect 42708 6128 42760 6180
rect 44088 6196 44140 6248
rect 45468 6239 45520 6248
rect 45468 6205 45477 6239
rect 45477 6205 45511 6239
rect 45511 6205 45520 6239
rect 45468 6196 45520 6205
rect 46940 6196 46992 6248
rect 48688 6400 48740 6452
rect 48320 6332 48372 6384
rect 49516 6400 49568 6452
rect 50160 6400 50212 6452
rect 49884 6375 49936 6384
rect 48780 6264 48832 6316
rect 49884 6341 49893 6375
rect 49893 6341 49927 6375
rect 49927 6341 49936 6375
rect 49884 6332 49936 6341
rect 53840 6375 53892 6384
rect 53840 6341 53849 6375
rect 53849 6341 53883 6375
rect 53883 6341 53892 6375
rect 53840 6332 53892 6341
rect 49148 6307 49200 6316
rect 49148 6273 49151 6307
rect 49151 6273 49185 6307
rect 49185 6273 49200 6307
rect 49148 6264 49200 6273
rect 50068 6264 50120 6316
rect 52276 6264 52328 6316
rect 48228 6239 48280 6248
rect 48228 6205 48237 6239
rect 48237 6205 48271 6239
rect 48271 6205 48280 6239
rect 48228 6196 48280 6205
rect 51448 6196 51500 6248
rect 53656 6239 53708 6248
rect 53656 6205 53665 6239
rect 53665 6205 53699 6239
rect 53699 6205 53708 6239
rect 53656 6196 53708 6205
rect 53932 6239 53984 6248
rect 53932 6205 53941 6239
rect 53941 6205 53975 6239
rect 53975 6205 53984 6239
rect 53932 6196 53984 6205
rect 56140 6400 56192 6452
rect 58256 6400 58308 6452
rect 58992 6400 59044 6452
rect 59544 6443 59596 6452
rect 59544 6409 59553 6443
rect 59553 6409 59587 6443
rect 59587 6409 59596 6443
rect 59544 6400 59596 6409
rect 60648 6443 60700 6452
rect 60648 6409 60657 6443
rect 60657 6409 60691 6443
rect 60691 6409 60700 6443
rect 60648 6400 60700 6409
rect 62120 6400 62172 6452
rect 65616 6400 65668 6452
rect 65708 6400 65760 6452
rect 67640 6400 67692 6452
rect 68560 6443 68612 6452
rect 68560 6409 68569 6443
rect 68569 6409 68603 6443
rect 68603 6409 68612 6443
rect 68560 6400 68612 6409
rect 71504 6400 71556 6452
rect 72056 6400 72108 6452
rect 55036 6332 55088 6384
rect 58716 6375 58768 6384
rect 54852 6196 54904 6248
rect 57888 6264 57940 6316
rect 57704 6196 57756 6248
rect 58716 6341 58725 6375
rect 58725 6341 58759 6375
rect 58759 6341 58768 6375
rect 58716 6332 58768 6341
rect 59176 6332 59228 6384
rect 67456 6332 67508 6384
rect 67732 6332 67784 6384
rect 75368 6400 75420 6452
rect 75460 6400 75512 6452
rect 76380 6400 76432 6452
rect 58900 6264 58952 6316
rect 59360 6307 59412 6316
rect 59360 6273 59369 6307
rect 59369 6273 59403 6307
rect 59403 6273 59412 6307
rect 59360 6264 59412 6273
rect 59268 6196 59320 6248
rect 26700 6060 26752 6112
rect 27436 6060 27488 6112
rect 28816 6060 28868 6112
rect 33876 6060 33928 6112
rect 34152 6060 34204 6112
rect 44272 6103 44324 6112
rect 44272 6069 44281 6103
rect 44281 6069 44315 6103
rect 44315 6069 44324 6103
rect 44272 6060 44324 6069
rect 49608 6171 49660 6180
rect 49608 6137 49617 6171
rect 49617 6137 49651 6171
rect 49651 6137 49660 6171
rect 49608 6128 49660 6137
rect 45744 6060 45796 6112
rect 46940 6060 46992 6112
rect 48320 6060 48372 6112
rect 48780 6060 48832 6112
rect 50712 6060 50764 6112
rect 51356 6060 51408 6112
rect 56968 6060 57020 6112
rect 57152 6060 57204 6112
rect 61660 6264 61712 6316
rect 61936 6264 61988 6316
rect 63592 6264 63644 6316
rect 63776 6307 63828 6316
rect 63776 6273 63785 6307
rect 63785 6273 63819 6307
rect 63819 6273 63828 6307
rect 63776 6264 63828 6273
rect 64512 6307 64564 6316
rect 64512 6273 64521 6307
rect 64521 6273 64555 6307
rect 64555 6273 64564 6307
rect 64512 6264 64564 6273
rect 64696 6307 64748 6316
rect 64696 6273 64705 6307
rect 64705 6273 64739 6307
rect 64739 6273 64748 6307
rect 64696 6264 64748 6273
rect 65156 6307 65208 6316
rect 65156 6273 65165 6307
rect 65165 6273 65199 6307
rect 65199 6273 65208 6307
rect 65156 6264 65208 6273
rect 65340 6307 65392 6316
rect 65340 6273 65349 6307
rect 65349 6273 65383 6307
rect 65383 6273 65392 6307
rect 65340 6264 65392 6273
rect 66076 6264 66128 6316
rect 60004 6196 60056 6248
rect 61016 6128 61068 6180
rect 61108 6128 61160 6180
rect 66168 6196 66220 6248
rect 64604 6128 64656 6180
rect 62120 6103 62172 6112
rect 62120 6069 62129 6103
rect 62129 6069 62163 6103
rect 62163 6069 62172 6103
rect 62120 6060 62172 6069
rect 63316 6103 63368 6112
rect 63316 6069 63325 6103
rect 63325 6069 63359 6103
rect 63359 6069 63368 6103
rect 63316 6060 63368 6069
rect 63500 6060 63552 6112
rect 65248 6060 65300 6112
rect 65892 6103 65944 6112
rect 65892 6069 65901 6103
rect 65901 6069 65935 6103
rect 65935 6069 65944 6103
rect 65892 6060 65944 6069
rect 66076 6060 66128 6112
rect 67548 6264 67600 6316
rect 70308 6307 70360 6316
rect 70308 6273 70317 6307
rect 70317 6273 70351 6307
rect 70351 6273 70360 6307
rect 70308 6264 70360 6273
rect 70768 6264 70820 6316
rect 71412 6307 71464 6316
rect 71412 6273 71421 6307
rect 71421 6273 71455 6307
rect 71455 6273 71464 6307
rect 71412 6264 71464 6273
rect 71688 6307 71740 6316
rect 71688 6273 71697 6307
rect 71697 6273 71731 6307
rect 71731 6273 71740 6307
rect 71688 6264 71740 6273
rect 74632 6332 74684 6384
rect 73528 6307 73580 6316
rect 66628 6128 66680 6180
rect 71504 6196 71556 6248
rect 73528 6273 73537 6307
rect 73537 6273 73571 6307
rect 73571 6273 73580 6307
rect 73528 6264 73580 6273
rect 74356 6264 74408 6316
rect 76012 6332 76064 6384
rect 77392 6400 77444 6452
rect 83188 6400 83240 6452
rect 94136 6443 94188 6452
rect 78772 6375 78824 6384
rect 75000 6264 75052 6316
rect 78772 6341 78781 6375
rect 78781 6341 78815 6375
rect 78815 6341 78824 6375
rect 78772 6332 78824 6341
rect 79232 6375 79284 6384
rect 79232 6341 79241 6375
rect 79241 6341 79275 6375
rect 79275 6341 79284 6375
rect 79232 6332 79284 6341
rect 79692 6332 79744 6384
rect 80704 6332 80756 6384
rect 84108 6332 84160 6384
rect 75460 6239 75512 6248
rect 75460 6205 75469 6239
rect 75469 6205 75503 6239
rect 75503 6205 75512 6239
rect 75460 6196 75512 6205
rect 68100 6060 68152 6112
rect 70400 6060 70452 6112
rect 72148 6060 72200 6112
rect 73528 6060 73580 6112
rect 73988 6060 74040 6112
rect 75460 6060 75512 6112
rect 76564 6196 76616 6248
rect 76656 6060 76708 6112
rect 83372 6264 83424 6316
rect 83740 6264 83792 6316
rect 80244 6239 80296 6248
rect 80244 6205 80253 6239
rect 80253 6205 80287 6239
rect 80287 6205 80296 6239
rect 80244 6196 80296 6205
rect 81256 6196 81308 6248
rect 81624 6196 81676 6248
rect 81992 6239 82044 6248
rect 81992 6205 82001 6239
rect 82001 6205 82035 6239
rect 82035 6205 82044 6239
rect 81992 6196 82044 6205
rect 82820 6239 82872 6248
rect 82820 6205 82829 6239
rect 82829 6205 82863 6239
rect 82863 6205 82872 6239
rect 82820 6196 82872 6205
rect 78588 6128 78640 6180
rect 87052 6332 87104 6384
rect 94136 6409 94145 6443
rect 94145 6409 94179 6443
rect 94179 6409 94188 6443
rect 94136 6400 94188 6409
rect 91836 6332 91888 6384
rect 84752 6307 84804 6316
rect 84752 6273 84761 6307
rect 84761 6273 84795 6307
rect 84795 6273 84804 6307
rect 85028 6307 85080 6316
rect 84752 6264 84804 6273
rect 85028 6273 85037 6307
rect 85037 6273 85071 6307
rect 85071 6273 85080 6307
rect 85028 6264 85080 6273
rect 85488 6264 85540 6316
rect 85764 6307 85816 6316
rect 85764 6273 85773 6307
rect 85773 6273 85807 6307
rect 85807 6273 85816 6307
rect 85764 6264 85816 6273
rect 86868 6264 86920 6316
rect 87420 6307 87472 6316
rect 87420 6273 87429 6307
rect 87429 6273 87463 6307
rect 87463 6273 87472 6307
rect 87420 6264 87472 6273
rect 88432 6264 88484 6316
rect 86132 6196 86184 6248
rect 88892 6196 88944 6248
rect 90824 6307 90876 6316
rect 90824 6273 90833 6307
rect 90833 6273 90867 6307
rect 90867 6273 90876 6307
rect 90824 6264 90876 6273
rect 91284 6264 91336 6316
rect 93032 6307 93084 6316
rect 93032 6273 93041 6307
rect 93041 6273 93075 6307
rect 93075 6273 93084 6307
rect 93032 6264 93084 6273
rect 89904 6196 89956 6248
rect 77852 6103 77904 6112
rect 77852 6069 77861 6103
rect 77861 6069 77895 6103
rect 77895 6069 77904 6103
rect 77852 6060 77904 6069
rect 81532 6060 81584 6112
rect 83464 6060 83516 6112
rect 83832 6060 83884 6112
rect 84384 6060 84436 6112
rect 85764 6060 85816 6112
rect 87604 6103 87656 6112
rect 87604 6069 87613 6103
rect 87613 6069 87647 6103
rect 87647 6069 87656 6103
rect 87604 6060 87656 6069
rect 87696 6060 87748 6112
rect 91008 6060 91060 6112
rect 91836 6060 91888 6112
rect 92756 6060 92808 6112
rect 12668 5958 12720 6010
rect 12732 5958 12784 6010
rect 12796 5958 12848 6010
rect 12860 5958 12912 6010
rect 12924 5958 12976 6010
rect 36105 5958 36157 6010
rect 36169 5958 36221 6010
rect 36233 5958 36285 6010
rect 36297 5958 36349 6010
rect 36361 5958 36413 6010
rect 59542 5958 59594 6010
rect 59606 5958 59658 6010
rect 59670 5958 59722 6010
rect 59734 5958 59786 6010
rect 59798 5958 59850 6010
rect 82979 5958 83031 6010
rect 83043 5958 83095 6010
rect 83107 5958 83159 6010
rect 83171 5958 83223 6010
rect 83235 5958 83287 6010
rect 9496 5856 9548 5908
rect 10692 5856 10744 5908
rect 19892 5899 19944 5908
rect 19892 5865 19901 5899
rect 19901 5865 19935 5899
rect 19935 5865 19944 5899
rect 19892 5856 19944 5865
rect 3976 5763 4028 5772
rect 3976 5729 3985 5763
rect 3985 5729 4019 5763
rect 4019 5729 4028 5763
rect 3976 5720 4028 5729
rect 6828 5763 6880 5772
rect 6828 5729 6837 5763
rect 6837 5729 6871 5763
rect 6871 5729 6880 5763
rect 6828 5720 6880 5729
rect 5724 5652 5776 5704
rect 18512 5720 18564 5772
rect 19708 5720 19760 5772
rect 4252 5627 4304 5636
rect 4252 5593 4261 5627
rect 4261 5593 4295 5627
rect 4295 5593 4304 5627
rect 4252 5584 4304 5593
rect 5724 5559 5776 5568
rect 5724 5525 5733 5559
rect 5733 5525 5767 5559
rect 5767 5525 5776 5559
rect 5724 5516 5776 5525
rect 13084 5584 13136 5636
rect 19616 5695 19668 5704
rect 19616 5661 19625 5695
rect 19625 5661 19659 5695
rect 19659 5661 19668 5695
rect 19616 5652 19668 5661
rect 22836 5856 22888 5908
rect 23572 5856 23624 5908
rect 23756 5788 23808 5840
rect 25688 5856 25740 5908
rect 25872 5899 25924 5908
rect 25872 5865 25881 5899
rect 25881 5865 25915 5899
rect 25915 5865 25924 5899
rect 25872 5856 25924 5865
rect 14556 5627 14608 5636
rect 14556 5593 14565 5627
rect 14565 5593 14599 5627
rect 14599 5593 14608 5627
rect 14556 5584 14608 5593
rect 19432 5584 19484 5636
rect 22100 5584 22152 5636
rect 22376 5584 22428 5636
rect 8392 5516 8444 5568
rect 9864 5559 9916 5568
rect 9864 5525 9873 5559
rect 9873 5525 9907 5559
rect 9907 5525 9916 5559
rect 9864 5516 9916 5525
rect 10784 5516 10836 5568
rect 22008 5559 22060 5568
rect 22008 5525 22017 5559
rect 22017 5525 22051 5559
rect 22051 5525 22060 5559
rect 22008 5516 22060 5525
rect 22652 5652 22704 5704
rect 22836 5695 22888 5704
rect 22836 5661 22845 5695
rect 22845 5661 22879 5695
rect 22879 5661 22888 5695
rect 22836 5652 22888 5661
rect 23296 5720 23348 5772
rect 24952 5788 25004 5840
rect 28724 5856 28776 5908
rect 40132 5856 40184 5908
rect 41604 5856 41656 5908
rect 42892 5856 42944 5908
rect 44548 5856 44600 5908
rect 46664 5856 46716 5908
rect 48044 5856 48096 5908
rect 49516 5856 49568 5908
rect 49792 5899 49844 5908
rect 49792 5865 49801 5899
rect 49801 5865 49835 5899
rect 49835 5865 49844 5899
rect 49792 5856 49844 5865
rect 50804 5899 50856 5908
rect 50804 5865 50813 5899
rect 50813 5865 50847 5899
rect 50847 5865 50856 5899
rect 50804 5856 50856 5865
rect 51448 5899 51500 5908
rect 51448 5865 51457 5899
rect 51457 5865 51491 5899
rect 51491 5865 51500 5899
rect 51448 5856 51500 5865
rect 51724 5856 51776 5908
rect 52552 5856 52604 5908
rect 53288 5856 53340 5908
rect 53748 5856 53800 5908
rect 54484 5899 54536 5908
rect 54484 5865 54493 5899
rect 54493 5865 54527 5899
rect 54527 5865 54536 5899
rect 54484 5856 54536 5865
rect 28448 5831 28500 5840
rect 28448 5797 28457 5831
rect 28457 5797 28491 5831
rect 28491 5797 28500 5831
rect 28448 5788 28500 5797
rect 24124 5720 24176 5772
rect 27068 5720 27120 5772
rect 31760 5720 31812 5772
rect 32496 5763 32548 5772
rect 32496 5729 32505 5763
rect 32505 5729 32539 5763
rect 32539 5729 32548 5763
rect 32496 5720 32548 5729
rect 35532 5788 35584 5840
rect 38108 5831 38160 5840
rect 38108 5797 38117 5831
rect 38117 5797 38151 5831
rect 38151 5797 38160 5831
rect 38108 5788 38160 5797
rect 38844 5831 38896 5840
rect 38844 5797 38853 5831
rect 38853 5797 38887 5831
rect 38887 5797 38896 5831
rect 38844 5788 38896 5797
rect 39028 5788 39080 5840
rect 40316 5788 40368 5840
rect 41236 5788 41288 5840
rect 44364 5788 44416 5840
rect 45284 5788 45336 5840
rect 49700 5788 49752 5840
rect 51356 5831 51408 5840
rect 35072 5720 35124 5772
rect 35900 5720 35952 5772
rect 36452 5720 36504 5772
rect 37464 5720 37516 5772
rect 40868 5720 40920 5772
rect 44272 5720 44324 5772
rect 45652 5720 45704 5772
rect 45744 5720 45796 5772
rect 48228 5720 48280 5772
rect 51356 5797 51365 5831
rect 51365 5797 51399 5831
rect 51399 5797 51408 5831
rect 51356 5788 51408 5797
rect 59452 5856 59504 5908
rect 60096 5899 60148 5908
rect 60096 5865 60105 5899
rect 60105 5865 60139 5899
rect 60139 5865 60148 5899
rect 60096 5856 60148 5865
rect 62120 5899 62172 5908
rect 62120 5865 62150 5899
rect 62150 5865 62172 5899
rect 62120 5856 62172 5865
rect 62304 5856 62356 5908
rect 63408 5856 63460 5908
rect 67364 5856 67416 5908
rect 68100 5899 68152 5908
rect 68100 5865 68109 5899
rect 68109 5865 68143 5899
rect 68143 5865 68152 5899
rect 68100 5856 68152 5865
rect 69204 5899 69256 5908
rect 69204 5865 69213 5899
rect 69213 5865 69247 5899
rect 69247 5865 69256 5899
rect 69204 5856 69256 5865
rect 69296 5856 69348 5908
rect 70124 5856 70176 5908
rect 70584 5856 70636 5908
rect 70952 5899 71004 5908
rect 70952 5865 70961 5899
rect 70961 5865 70995 5899
rect 70995 5865 71004 5899
rect 70952 5856 71004 5865
rect 71412 5856 71464 5908
rect 74356 5856 74408 5908
rect 74908 5856 74960 5908
rect 24216 5652 24268 5704
rect 24860 5652 24912 5704
rect 25228 5652 25280 5704
rect 25412 5695 25464 5704
rect 25412 5661 25421 5695
rect 25421 5661 25455 5695
rect 25455 5661 25464 5695
rect 25412 5652 25464 5661
rect 25688 5695 25740 5704
rect 25688 5661 25697 5695
rect 25697 5661 25731 5695
rect 25731 5661 25740 5695
rect 25688 5652 25740 5661
rect 26148 5652 26200 5704
rect 26700 5695 26752 5704
rect 26700 5661 26709 5695
rect 26709 5661 26743 5695
rect 26743 5661 26752 5695
rect 26700 5652 26752 5661
rect 38016 5652 38068 5704
rect 41236 5695 41288 5704
rect 41236 5661 41245 5695
rect 41245 5661 41279 5695
rect 41279 5661 41288 5695
rect 41236 5652 41288 5661
rect 44456 5695 44508 5704
rect 23020 5584 23072 5636
rect 23112 5627 23164 5636
rect 23112 5593 23121 5627
rect 23121 5593 23155 5627
rect 23155 5593 23164 5627
rect 23112 5584 23164 5593
rect 23480 5584 23532 5636
rect 25596 5584 25648 5636
rect 27436 5584 27488 5636
rect 29828 5584 29880 5636
rect 32772 5627 32824 5636
rect 32772 5593 32781 5627
rect 32781 5593 32815 5627
rect 32815 5593 32824 5627
rect 32772 5584 32824 5593
rect 33232 5584 33284 5636
rect 24032 5516 24084 5568
rect 24860 5516 24912 5568
rect 25136 5516 25188 5568
rect 25228 5516 25280 5568
rect 32588 5516 32640 5568
rect 32680 5516 32732 5568
rect 37464 5584 37516 5636
rect 42524 5584 42576 5636
rect 44456 5661 44465 5695
rect 44465 5661 44499 5695
rect 44499 5661 44508 5695
rect 44456 5652 44508 5661
rect 47676 5652 47728 5704
rect 48688 5695 48740 5704
rect 48688 5661 48697 5695
rect 48697 5661 48731 5695
rect 48731 5661 48740 5695
rect 48688 5652 48740 5661
rect 49516 5695 49568 5704
rect 46204 5584 46256 5636
rect 47308 5627 47360 5636
rect 47308 5593 47317 5627
rect 47317 5593 47351 5627
rect 47351 5593 47360 5627
rect 47308 5584 47360 5593
rect 49516 5661 49525 5695
rect 49525 5661 49559 5695
rect 49559 5661 49568 5695
rect 49516 5652 49568 5661
rect 49608 5695 49660 5704
rect 49608 5661 49617 5695
rect 49617 5661 49651 5695
rect 49651 5661 49660 5695
rect 49608 5652 49660 5661
rect 50252 5652 50304 5704
rect 51540 5763 51592 5772
rect 51540 5729 51549 5763
rect 51549 5729 51583 5763
rect 51583 5729 51592 5763
rect 51540 5720 51592 5729
rect 50620 5695 50672 5704
rect 50068 5584 50120 5636
rect 50620 5661 50629 5695
rect 50629 5661 50663 5695
rect 50663 5661 50672 5695
rect 50620 5652 50672 5661
rect 50712 5652 50764 5704
rect 58900 5788 58952 5840
rect 60280 5788 60332 5840
rect 55220 5720 55272 5772
rect 58808 5720 58860 5772
rect 60740 5763 60792 5772
rect 60740 5729 60749 5763
rect 60749 5729 60783 5763
rect 60783 5729 60792 5763
rect 60740 5720 60792 5729
rect 63592 5788 63644 5840
rect 63500 5720 63552 5772
rect 64696 5788 64748 5840
rect 65708 5788 65760 5840
rect 67548 5831 67600 5840
rect 67548 5797 67557 5831
rect 67557 5797 67591 5831
rect 67591 5797 67600 5831
rect 67548 5788 67600 5797
rect 75000 5788 75052 5840
rect 76012 5788 76064 5840
rect 64604 5763 64656 5772
rect 64604 5729 64613 5763
rect 64613 5729 64647 5763
rect 64647 5729 64656 5763
rect 64604 5720 64656 5729
rect 66076 5763 66128 5772
rect 66076 5729 66085 5763
rect 66085 5729 66119 5763
rect 66119 5729 66128 5763
rect 66076 5720 66128 5729
rect 66168 5720 66220 5772
rect 71964 5763 72016 5772
rect 44180 5516 44232 5568
rect 49148 5516 49200 5568
rect 50252 5516 50304 5568
rect 54392 5584 54444 5636
rect 56692 5652 56744 5704
rect 56968 5695 57020 5704
rect 56968 5661 56977 5695
rect 56977 5661 57011 5695
rect 57011 5661 57020 5695
rect 56968 5652 57020 5661
rect 57244 5652 57296 5704
rect 56140 5584 56192 5636
rect 57704 5627 57756 5636
rect 57704 5593 57713 5627
rect 57713 5593 57747 5627
rect 57747 5593 57756 5627
rect 57888 5627 57940 5636
rect 57704 5584 57756 5593
rect 57888 5593 57897 5627
rect 57897 5593 57931 5627
rect 57931 5593 57940 5627
rect 57888 5584 57940 5593
rect 58440 5652 58492 5704
rect 59452 5652 59504 5704
rect 60832 5695 60884 5704
rect 52276 5516 52328 5568
rect 54852 5516 54904 5568
rect 55864 5516 55916 5568
rect 56784 5516 56836 5568
rect 59360 5584 59412 5636
rect 60280 5584 60332 5636
rect 60832 5661 60841 5695
rect 60841 5661 60875 5695
rect 60875 5661 60884 5695
rect 60832 5652 60884 5661
rect 63684 5652 63736 5704
rect 59176 5516 59228 5568
rect 59820 5516 59872 5568
rect 60372 5516 60424 5568
rect 62396 5516 62448 5568
rect 63408 5584 63460 5636
rect 64880 5584 64932 5636
rect 64512 5516 64564 5568
rect 67732 5652 67784 5704
rect 69848 5695 69900 5704
rect 69848 5661 69857 5695
rect 69857 5661 69891 5695
rect 69891 5661 69900 5695
rect 69848 5652 69900 5661
rect 67456 5584 67508 5636
rect 71964 5729 71973 5763
rect 71973 5729 72007 5763
rect 72007 5729 72016 5763
rect 71964 5720 72016 5729
rect 73160 5763 73212 5772
rect 73160 5729 73169 5763
rect 73169 5729 73203 5763
rect 73203 5729 73212 5763
rect 73160 5720 73212 5729
rect 73252 5720 73304 5772
rect 70124 5652 70176 5704
rect 71412 5652 71464 5704
rect 71780 5695 71832 5704
rect 71780 5661 71789 5695
rect 71789 5661 71823 5695
rect 71823 5661 71832 5695
rect 71780 5652 71832 5661
rect 73344 5652 73396 5704
rect 74908 5652 74960 5704
rect 75276 5695 75328 5704
rect 75276 5661 75285 5695
rect 75285 5661 75319 5695
rect 75319 5661 75328 5695
rect 75276 5652 75328 5661
rect 75552 5695 75604 5704
rect 67640 5516 67692 5568
rect 68192 5516 68244 5568
rect 75184 5584 75236 5636
rect 75552 5661 75561 5695
rect 75561 5661 75595 5695
rect 75595 5661 75604 5695
rect 75552 5652 75604 5661
rect 76288 5856 76340 5908
rect 77852 5856 77904 5908
rect 80980 5856 81032 5908
rect 82820 5856 82872 5908
rect 83464 5899 83516 5908
rect 83464 5865 83473 5899
rect 83473 5865 83507 5899
rect 83507 5865 83516 5899
rect 83464 5856 83516 5865
rect 84752 5856 84804 5908
rect 76748 5788 76800 5840
rect 80796 5788 80848 5840
rect 82728 5788 82780 5840
rect 84292 5788 84344 5840
rect 86408 5856 86460 5908
rect 87604 5856 87656 5908
rect 89812 5856 89864 5908
rect 86132 5788 86184 5840
rect 87236 5788 87288 5840
rect 79048 5652 79100 5704
rect 79692 5695 79744 5704
rect 79692 5661 79701 5695
rect 79701 5661 79735 5695
rect 79735 5661 79744 5695
rect 79692 5652 79744 5661
rect 80704 5763 80756 5772
rect 80704 5729 80713 5763
rect 80713 5729 80747 5763
rect 80747 5729 80756 5763
rect 80704 5720 80756 5729
rect 81532 5720 81584 5772
rect 81624 5720 81676 5772
rect 86592 5720 86644 5772
rect 75460 5584 75512 5636
rect 75828 5584 75880 5636
rect 75920 5584 75972 5636
rect 78772 5584 78824 5636
rect 74080 5559 74132 5568
rect 74080 5525 74089 5559
rect 74089 5525 74123 5559
rect 74123 5525 74132 5559
rect 74080 5516 74132 5525
rect 75276 5516 75328 5568
rect 76288 5559 76340 5568
rect 76288 5525 76297 5559
rect 76297 5525 76331 5559
rect 76331 5525 76340 5559
rect 76288 5516 76340 5525
rect 76472 5559 76524 5568
rect 76472 5525 76481 5559
rect 76481 5525 76515 5559
rect 76515 5525 76524 5559
rect 76472 5516 76524 5525
rect 76932 5516 76984 5568
rect 77668 5516 77720 5568
rect 79876 5516 79928 5568
rect 79968 5516 80020 5568
rect 80060 5516 80112 5568
rect 81348 5652 81400 5704
rect 81992 5652 82044 5704
rect 86960 5695 87012 5704
rect 80336 5584 80388 5636
rect 86960 5661 86969 5695
rect 86969 5661 87003 5695
rect 87003 5661 87012 5695
rect 86960 5652 87012 5661
rect 87972 5763 88024 5772
rect 87972 5729 87981 5763
rect 87981 5729 88015 5763
rect 88015 5729 88024 5763
rect 87972 5720 88024 5729
rect 89720 5720 89772 5772
rect 87788 5652 87840 5704
rect 89352 5695 89404 5704
rect 89352 5661 89361 5695
rect 89361 5661 89395 5695
rect 89395 5661 89404 5695
rect 89352 5652 89404 5661
rect 93124 5856 93176 5908
rect 93400 5899 93452 5908
rect 93400 5865 93409 5899
rect 93409 5865 93443 5899
rect 93443 5865 93452 5899
rect 93400 5856 93452 5865
rect 93768 5856 93820 5908
rect 92756 5831 92808 5840
rect 92756 5797 92765 5831
rect 92765 5797 92799 5831
rect 92799 5797 92808 5831
rect 92756 5788 92808 5797
rect 91284 5720 91336 5772
rect 91836 5695 91888 5704
rect 91836 5661 91845 5695
rect 91845 5661 91879 5695
rect 91879 5661 91888 5695
rect 91836 5652 91888 5661
rect 93216 5695 93268 5704
rect 89904 5584 89956 5636
rect 93216 5661 93225 5695
rect 93225 5661 93259 5695
rect 93259 5661 93268 5695
rect 93216 5652 93268 5661
rect 81440 5516 81492 5568
rect 81624 5516 81676 5568
rect 86040 5516 86092 5568
rect 87144 5516 87196 5568
rect 87236 5516 87288 5568
rect 24386 5414 24438 5466
rect 24450 5414 24502 5466
rect 24514 5414 24566 5466
rect 24578 5414 24630 5466
rect 24642 5414 24694 5466
rect 47823 5414 47875 5466
rect 47887 5414 47939 5466
rect 47951 5414 48003 5466
rect 48015 5414 48067 5466
rect 48079 5414 48131 5466
rect 71260 5414 71312 5466
rect 71324 5414 71376 5466
rect 71388 5414 71440 5466
rect 71452 5414 71504 5466
rect 71516 5414 71568 5466
rect 94697 5414 94749 5466
rect 94761 5414 94813 5466
rect 94825 5414 94877 5466
rect 94889 5414 94941 5466
rect 94953 5414 95005 5466
rect 4252 5355 4304 5364
rect 4252 5321 4261 5355
rect 4261 5321 4295 5355
rect 4295 5321 4304 5355
rect 4252 5312 4304 5321
rect 8392 5312 8444 5364
rect 22376 5312 22428 5364
rect 23480 5312 23532 5364
rect 23756 5312 23808 5364
rect 24768 5312 24820 5364
rect 9588 5287 9640 5296
rect 9588 5253 9597 5287
rect 9597 5253 9631 5287
rect 9631 5253 9640 5287
rect 9588 5244 9640 5253
rect 12992 5287 13044 5296
rect 12992 5253 13001 5287
rect 13001 5253 13035 5287
rect 13035 5253 13044 5287
rect 12992 5244 13044 5253
rect 22008 5244 22060 5296
rect 4344 5219 4396 5228
rect 4344 5185 4353 5219
rect 4353 5185 4387 5219
rect 4387 5185 4396 5219
rect 4344 5176 4396 5185
rect 5724 5176 5776 5228
rect 14464 5176 14516 5228
rect 22100 5176 22152 5228
rect 22560 5219 22612 5228
rect 22560 5185 22569 5219
rect 22569 5185 22603 5219
rect 22603 5185 22612 5219
rect 22560 5176 22612 5185
rect 23572 5244 23624 5296
rect 24216 5244 24268 5296
rect 24400 5244 24452 5296
rect 26240 5244 26292 5296
rect 22836 5219 22888 5228
rect 22836 5185 22845 5219
rect 22845 5185 22879 5219
rect 22879 5185 22888 5219
rect 22836 5176 22888 5185
rect 24032 5176 24084 5228
rect 25044 5176 25096 5228
rect 13728 5108 13780 5160
rect 15476 5108 15528 5160
rect 15936 5108 15988 5160
rect 24860 5108 24912 5160
rect 26516 5108 26568 5160
rect 8484 5040 8536 5092
rect 24400 5040 24452 5092
rect 7012 4972 7064 5024
rect 23664 5015 23716 5024
rect 23664 4981 23673 5015
rect 23673 4981 23707 5015
rect 23707 4981 23716 5015
rect 23664 4972 23716 4981
rect 24216 5015 24268 5024
rect 24216 4981 24225 5015
rect 24225 4981 24259 5015
rect 24259 4981 24268 5015
rect 24216 4972 24268 4981
rect 24676 5015 24728 5024
rect 24676 4981 24685 5015
rect 24685 4981 24719 5015
rect 24719 4981 24728 5015
rect 24676 4972 24728 4981
rect 24768 4972 24820 5024
rect 28264 5287 28316 5296
rect 28264 5253 28273 5287
rect 28273 5253 28307 5287
rect 28307 5253 28316 5287
rect 28264 5244 28316 5253
rect 33232 5244 33284 5296
rect 27252 5151 27304 5160
rect 27252 5117 27261 5151
rect 27261 5117 27295 5151
rect 27295 5117 27304 5151
rect 27252 5108 27304 5117
rect 26700 5040 26752 5092
rect 31760 5219 31812 5228
rect 31760 5185 31769 5219
rect 31769 5185 31803 5219
rect 31803 5185 31812 5219
rect 32680 5219 32732 5228
rect 31760 5176 31812 5185
rect 32680 5185 32689 5219
rect 32689 5185 32723 5219
rect 32723 5185 32732 5219
rect 32680 5176 32732 5185
rect 34244 5312 34296 5364
rect 37924 5355 37976 5364
rect 37924 5321 37933 5355
rect 37933 5321 37967 5355
rect 37967 5321 37976 5355
rect 37924 5312 37976 5321
rect 40040 5312 40092 5364
rect 40868 5355 40920 5364
rect 40868 5321 40877 5355
rect 40877 5321 40911 5355
rect 40911 5321 40920 5355
rect 40868 5312 40920 5321
rect 33600 5244 33652 5296
rect 80060 5312 80112 5364
rect 42064 5244 42116 5296
rect 42708 5244 42760 5296
rect 45560 5244 45612 5296
rect 47768 5244 47820 5296
rect 49608 5287 49660 5296
rect 36452 5176 36504 5228
rect 36728 5176 36780 5228
rect 38016 5176 38068 5228
rect 42984 5219 43036 5228
rect 36912 5151 36964 5160
rect 28448 4972 28500 5024
rect 30012 5015 30064 5024
rect 30012 4981 30021 5015
rect 30021 4981 30055 5015
rect 30055 4981 30064 5015
rect 30012 4972 30064 4981
rect 30104 4972 30156 5024
rect 32772 5040 32824 5092
rect 33416 5040 33468 5092
rect 36912 5117 36921 5151
rect 36921 5117 36955 5151
rect 36955 5117 36964 5151
rect 36912 5108 36964 5117
rect 41236 5108 41288 5160
rect 41328 5108 41380 5160
rect 41788 5040 41840 5092
rect 42984 5185 42993 5219
rect 42993 5185 43027 5219
rect 43027 5185 43036 5219
rect 42984 5176 43036 5185
rect 45928 5176 45980 5228
rect 48136 5219 48188 5228
rect 48136 5185 48145 5219
rect 48145 5185 48179 5219
rect 48179 5185 48188 5219
rect 48136 5176 48188 5185
rect 49608 5253 49617 5287
rect 49617 5253 49651 5287
rect 49651 5253 49660 5287
rect 49608 5244 49660 5253
rect 50068 5219 50120 5228
rect 50068 5185 50077 5219
rect 50077 5185 50111 5219
rect 50111 5185 50120 5219
rect 50068 5176 50120 5185
rect 50160 5176 50212 5228
rect 52000 5244 52052 5296
rect 52184 5287 52236 5296
rect 52184 5253 52193 5287
rect 52193 5253 52227 5287
rect 52227 5253 52236 5287
rect 52184 5244 52236 5253
rect 53748 5244 53800 5296
rect 55128 5244 55180 5296
rect 55864 5287 55916 5296
rect 55864 5253 55873 5287
rect 55873 5253 55907 5287
rect 55907 5253 55916 5287
rect 55864 5244 55916 5253
rect 56600 5244 56652 5296
rect 57888 5244 57940 5296
rect 53380 5219 53432 5228
rect 53380 5185 53389 5219
rect 53389 5185 53423 5219
rect 53423 5185 53432 5219
rect 53380 5176 53432 5185
rect 53472 5219 53524 5228
rect 53472 5185 53481 5219
rect 53481 5185 53515 5219
rect 53515 5185 53524 5219
rect 56784 5219 56836 5228
rect 53472 5176 53524 5185
rect 56784 5185 56793 5219
rect 56793 5185 56827 5219
rect 56827 5185 56836 5219
rect 56784 5176 56836 5185
rect 43076 5151 43128 5160
rect 43076 5117 43085 5151
rect 43085 5117 43119 5151
rect 43119 5117 43128 5151
rect 43076 5108 43128 5117
rect 43996 5151 44048 5160
rect 43996 5117 44005 5151
rect 44005 5117 44039 5151
rect 44039 5117 44048 5151
rect 43996 5108 44048 5117
rect 44364 5108 44416 5160
rect 45744 5083 45796 5092
rect 34888 4972 34940 5024
rect 40316 4972 40368 5024
rect 40960 4972 41012 5024
rect 42064 4972 42116 5024
rect 42708 5015 42760 5024
rect 42708 4981 42717 5015
rect 42717 4981 42751 5015
rect 42751 4981 42760 5015
rect 42708 4972 42760 4981
rect 45744 5049 45753 5083
rect 45753 5049 45787 5083
rect 45787 5049 45796 5083
rect 45744 5040 45796 5049
rect 47124 5108 47176 5160
rect 45284 4972 45336 5024
rect 47676 5040 47728 5092
rect 48228 4972 48280 5024
rect 48688 5108 48740 5160
rect 50344 5151 50396 5160
rect 50344 5117 50353 5151
rect 50353 5117 50387 5151
rect 50387 5117 50396 5151
rect 50344 5108 50396 5117
rect 51172 5151 51224 5160
rect 51172 5117 51181 5151
rect 51181 5117 51215 5151
rect 51215 5117 51224 5151
rect 51172 5108 51224 5117
rect 49608 5040 49660 5092
rect 55220 5108 55272 5160
rect 56140 5151 56192 5160
rect 56140 5117 56149 5151
rect 56149 5117 56183 5151
rect 56183 5117 56192 5151
rect 56140 5108 56192 5117
rect 57060 5219 57112 5228
rect 57060 5185 57069 5219
rect 57069 5185 57103 5219
rect 57103 5185 57112 5219
rect 57060 5176 57112 5185
rect 57336 5176 57388 5228
rect 57704 5176 57756 5228
rect 58348 5219 58400 5228
rect 58348 5185 58357 5219
rect 58357 5185 58391 5219
rect 58391 5185 58400 5219
rect 58348 5176 58400 5185
rect 54392 5083 54444 5092
rect 49424 5015 49476 5024
rect 49424 4981 49433 5015
rect 49433 4981 49467 5015
rect 49467 4981 49476 5015
rect 49424 4972 49476 4981
rect 49792 4972 49844 5024
rect 52000 4972 52052 5024
rect 53472 4972 53524 5024
rect 54392 5049 54401 5083
rect 54401 5049 54435 5083
rect 54435 5049 54444 5083
rect 54392 5040 54444 5049
rect 57336 5040 57388 5092
rect 59452 5108 59504 5160
rect 58808 5083 58860 5092
rect 58808 5049 58817 5083
rect 58817 5049 58851 5083
rect 58851 5049 58860 5083
rect 58808 5040 58860 5049
rect 58992 5040 59044 5092
rect 56140 4972 56192 5024
rect 56692 4972 56744 5024
rect 59084 4972 59136 5024
rect 59820 4972 59872 5024
rect 62304 5244 62356 5296
rect 62396 5287 62448 5296
rect 62396 5253 62405 5287
rect 62405 5253 62439 5287
rect 62439 5253 62448 5287
rect 62396 5244 62448 5253
rect 63316 5244 63368 5296
rect 64696 5244 64748 5296
rect 65892 5244 65944 5296
rect 67732 5244 67784 5296
rect 63500 5176 63552 5228
rect 65340 5176 65392 5228
rect 70308 5244 70360 5296
rect 71872 5244 71924 5296
rect 72056 5244 72108 5296
rect 76748 5287 76800 5296
rect 71780 5176 71832 5228
rect 60464 5108 60516 5160
rect 63868 5108 63920 5160
rect 69296 5108 69348 5160
rect 60832 4972 60884 5024
rect 64420 5040 64472 5092
rect 63684 4972 63736 5024
rect 71780 5040 71832 5092
rect 72148 5108 72200 5160
rect 73804 5176 73856 5228
rect 73988 5176 74040 5228
rect 74448 5176 74500 5228
rect 75276 5219 75328 5228
rect 75276 5185 75285 5219
rect 75285 5185 75319 5219
rect 75319 5185 75328 5219
rect 76748 5253 76757 5287
rect 76757 5253 76791 5287
rect 76791 5253 76800 5287
rect 76748 5244 76800 5253
rect 81992 5312 82044 5364
rect 85396 5312 85448 5364
rect 86960 5312 87012 5364
rect 87696 5312 87748 5364
rect 90640 5355 90692 5364
rect 90640 5321 90649 5355
rect 90649 5321 90683 5355
rect 90683 5321 90692 5355
rect 90640 5312 90692 5321
rect 91008 5312 91060 5364
rect 91836 5312 91888 5364
rect 93676 5312 93728 5364
rect 94044 5312 94096 5364
rect 75276 5176 75328 5185
rect 75828 5176 75880 5228
rect 73528 5040 73580 5092
rect 75920 5108 75972 5160
rect 76288 5176 76340 5228
rect 76840 5219 76892 5228
rect 76840 5185 76849 5219
rect 76849 5185 76883 5219
rect 76883 5185 76892 5219
rect 76840 5176 76892 5185
rect 76932 5176 76984 5228
rect 77668 5219 77720 5228
rect 77668 5185 77677 5219
rect 77677 5185 77711 5219
rect 77711 5185 77720 5219
rect 77668 5176 77720 5185
rect 80612 5244 80664 5296
rect 84016 5244 84068 5296
rect 92020 5244 92072 5296
rect 78036 5108 78088 5160
rect 75460 5040 75512 5092
rect 69848 4972 69900 5024
rect 74264 5015 74316 5024
rect 74264 4981 74273 5015
rect 74273 4981 74307 5015
rect 74307 4981 74316 5015
rect 74264 4972 74316 4981
rect 75828 4972 75880 5024
rect 84936 5176 84988 5228
rect 85396 5219 85448 5228
rect 85396 5185 85405 5219
rect 85405 5185 85439 5219
rect 85439 5185 85448 5219
rect 85396 5176 85448 5185
rect 85672 5176 85724 5228
rect 86592 5176 86644 5228
rect 87696 5219 87748 5228
rect 80244 5108 80296 5160
rect 80980 5151 81032 5160
rect 80152 5015 80204 5024
rect 80152 4981 80161 5015
rect 80161 4981 80195 5015
rect 80195 4981 80204 5015
rect 80980 5117 80989 5151
rect 80989 5117 81023 5151
rect 81023 5117 81032 5151
rect 80980 5108 81032 5117
rect 81440 5108 81492 5160
rect 84568 5151 84620 5160
rect 84568 5117 84577 5151
rect 84577 5117 84611 5151
rect 84611 5117 84620 5151
rect 84568 5108 84620 5117
rect 87696 5185 87705 5219
rect 87705 5185 87739 5219
rect 87739 5185 87748 5219
rect 87696 5176 87748 5185
rect 92388 5219 92440 5228
rect 92388 5185 92397 5219
rect 92397 5185 92431 5219
rect 92431 5185 92440 5219
rect 92388 5176 92440 5185
rect 93032 5219 93084 5228
rect 93032 5185 93041 5219
rect 93041 5185 93075 5219
rect 93075 5185 93084 5219
rect 93032 5176 93084 5185
rect 80152 4972 80204 4981
rect 81440 4972 81492 5024
rect 82176 4972 82228 5024
rect 83372 4972 83424 5024
rect 84200 5015 84252 5024
rect 84200 4981 84209 5015
rect 84209 4981 84243 5015
rect 84243 4981 84252 5015
rect 84200 4972 84252 4981
rect 84660 5015 84712 5024
rect 84660 4981 84669 5015
rect 84669 4981 84703 5015
rect 84703 4981 84712 5015
rect 84660 4972 84712 4981
rect 85120 5015 85172 5024
rect 85120 4981 85129 5015
rect 85129 4981 85163 5015
rect 85163 4981 85172 5015
rect 85120 4972 85172 4981
rect 91284 5108 91336 5160
rect 87052 4972 87104 5024
rect 87880 4972 87932 5024
rect 88064 4972 88116 5024
rect 88984 5015 89036 5024
rect 88984 4981 88993 5015
rect 88993 4981 89027 5015
rect 89027 4981 89036 5015
rect 88984 4972 89036 4981
rect 89352 4972 89404 5024
rect 91008 4972 91060 5024
rect 12668 4870 12720 4922
rect 12732 4870 12784 4922
rect 12796 4870 12848 4922
rect 12860 4870 12912 4922
rect 12924 4870 12976 4922
rect 36105 4870 36157 4922
rect 36169 4870 36221 4922
rect 36233 4870 36285 4922
rect 36297 4870 36349 4922
rect 36361 4870 36413 4922
rect 59542 4870 59594 4922
rect 59606 4870 59658 4922
rect 59670 4870 59722 4922
rect 59734 4870 59786 4922
rect 59798 4870 59850 4922
rect 82979 4870 83031 4922
rect 83043 4870 83095 4922
rect 83107 4870 83159 4922
rect 83171 4870 83223 4922
rect 83235 4870 83287 4922
rect 4344 4768 4396 4820
rect 22836 4811 22888 4820
rect 6736 4675 6788 4684
rect 6736 4641 6745 4675
rect 6745 4641 6779 4675
rect 6779 4641 6788 4675
rect 6736 4632 6788 4641
rect 7012 4675 7064 4684
rect 7012 4641 7021 4675
rect 7021 4641 7055 4675
rect 7055 4641 7064 4675
rect 7012 4632 7064 4641
rect 8392 4564 8444 4616
rect 9128 4607 9180 4616
rect 9128 4573 9137 4607
rect 9137 4573 9171 4607
rect 9171 4573 9180 4607
rect 9128 4564 9180 4573
rect 9864 4564 9916 4616
rect 10600 4564 10652 4616
rect 22836 4777 22845 4811
rect 22845 4777 22879 4811
rect 22879 4777 22888 4811
rect 22836 4768 22888 4777
rect 23388 4768 23440 4820
rect 26332 4768 26384 4820
rect 26516 4811 26568 4820
rect 26516 4777 26525 4811
rect 26525 4777 26559 4811
rect 26559 4777 26568 4811
rect 26516 4768 26568 4777
rect 27252 4768 27304 4820
rect 31116 4768 31168 4820
rect 34888 4768 34940 4820
rect 24216 4700 24268 4752
rect 30104 4700 30156 4752
rect 23112 4632 23164 4684
rect 24676 4632 24728 4684
rect 24860 4632 24912 4684
rect 33600 4700 33652 4752
rect 37740 4768 37792 4820
rect 33416 4632 33468 4684
rect 14464 4564 14516 4616
rect 23664 4564 23716 4616
rect 25044 4607 25096 4616
rect 25044 4573 25053 4607
rect 25053 4573 25087 4607
rect 25087 4573 25096 4607
rect 25044 4564 25096 4573
rect 25136 4607 25188 4616
rect 25136 4573 25145 4607
rect 25145 4573 25179 4607
rect 25179 4573 25188 4607
rect 25136 4564 25188 4573
rect 25688 4564 25740 4616
rect 29828 4564 29880 4616
rect 30840 4564 30892 4616
rect 39028 4743 39080 4752
rect 39028 4709 39037 4743
rect 39037 4709 39071 4743
rect 39071 4709 39080 4743
rect 39028 4700 39080 4709
rect 41788 4768 41840 4820
rect 42984 4700 43036 4752
rect 43352 4743 43404 4752
rect 43352 4709 43361 4743
rect 43361 4709 43395 4743
rect 43395 4709 43404 4743
rect 43352 4700 43404 4709
rect 44456 4700 44508 4752
rect 44916 4700 44968 4752
rect 42708 4632 42760 4684
rect 45836 4632 45888 4684
rect 48136 4768 48188 4820
rect 49608 4768 49660 4820
rect 50344 4768 50396 4820
rect 50620 4768 50672 4820
rect 52368 4768 52420 4820
rect 53748 4811 53800 4820
rect 53748 4777 53757 4811
rect 53757 4777 53791 4811
rect 53791 4777 53800 4811
rect 53748 4768 53800 4777
rect 53932 4768 53984 4820
rect 50068 4700 50120 4752
rect 53564 4700 53616 4752
rect 56600 4768 56652 4820
rect 57060 4768 57112 4820
rect 58164 4768 58216 4820
rect 49976 4632 50028 4684
rect 40408 4607 40460 4616
rect 22560 4496 22612 4548
rect 23296 4496 23348 4548
rect 10324 4471 10376 4480
rect 10324 4437 10333 4471
rect 10333 4437 10367 4471
rect 10367 4437 10376 4471
rect 10324 4428 10376 4437
rect 10692 4428 10744 4480
rect 15384 4471 15436 4480
rect 15384 4437 15393 4471
rect 15393 4437 15427 4471
rect 15427 4437 15436 4471
rect 15384 4428 15436 4437
rect 22836 4428 22888 4480
rect 24308 4496 24360 4548
rect 31116 4496 31168 4548
rect 31392 4539 31444 4548
rect 31392 4505 31401 4539
rect 31401 4505 31435 4539
rect 31435 4505 31444 4539
rect 31392 4496 31444 4505
rect 32312 4539 32364 4548
rect 32312 4505 32321 4539
rect 32321 4505 32355 4539
rect 32355 4505 32364 4539
rect 32312 4496 32364 4505
rect 35348 4539 35400 4548
rect 26148 4428 26200 4480
rect 26332 4428 26384 4480
rect 33600 4428 33652 4480
rect 34612 4428 34664 4480
rect 35348 4505 35357 4539
rect 35357 4505 35391 4539
rect 35391 4505 35400 4539
rect 35348 4496 35400 4505
rect 40408 4573 40417 4607
rect 40417 4573 40451 4607
rect 40451 4573 40460 4607
rect 40408 4564 40460 4573
rect 41788 4564 41840 4616
rect 42524 4564 42576 4616
rect 47124 4564 47176 4616
rect 47768 4607 47820 4616
rect 47768 4573 47777 4607
rect 47777 4573 47811 4607
rect 47811 4573 47820 4607
rect 47768 4564 47820 4573
rect 52276 4632 52328 4684
rect 52000 4607 52052 4616
rect 52000 4573 52009 4607
rect 52009 4573 52043 4607
rect 52043 4573 52052 4607
rect 52000 4564 52052 4573
rect 53472 4564 53524 4616
rect 36912 4496 36964 4548
rect 37924 4496 37976 4548
rect 38476 4496 38528 4548
rect 40684 4539 40736 4548
rect 40684 4505 40693 4539
rect 40693 4505 40727 4539
rect 40727 4505 40736 4539
rect 40684 4496 40736 4505
rect 38016 4428 38068 4480
rect 40040 4428 40092 4480
rect 42156 4471 42208 4480
rect 42156 4437 42165 4471
rect 42165 4437 42199 4471
rect 42199 4437 42208 4471
rect 42156 4428 42208 4437
rect 42524 4428 42576 4480
rect 43812 4428 43864 4480
rect 45928 4428 45980 4480
rect 47400 4496 47452 4548
rect 49792 4539 49844 4548
rect 49792 4505 49801 4539
rect 49801 4505 49835 4539
rect 49835 4505 49844 4539
rect 49792 4496 49844 4505
rect 51540 4496 51592 4548
rect 53380 4496 53432 4548
rect 61292 4768 61344 4820
rect 63500 4768 63552 4820
rect 63684 4768 63736 4820
rect 71688 4768 71740 4820
rect 73252 4811 73304 4820
rect 73252 4777 73261 4811
rect 73261 4777 73295 4811
rect 73295 4777 73304 4811
rect 73252 4768 73304 4777
rect 73620 4811 73672 4820
rect 73620 4777 73629 4811
rect 73629 4777 73663 4811
rect 73663 4777 73672 4811
rect 73620 4768 73672 4777
rect 76196 4811 76248 4820
rect 76196 4777 76205 4811
rect 76205 4777 76239 4811
rect 76239 4777 76248 4811
rect 76196 4768 76248 4777
rect 77484 4768 77536 4820
rect 61200 4743 61252 4752
rect 56140 4675 56192 4684
rect 56140 4641 56149 4675
rect 56149 4641 56183 4675
rect 56183 4641 56192 4675
rect 56140 4632 56192 4641
rect 56416 4564 56468 4616
rect 47492 4471 47544 4480
rect 47492 4437 47501 4471
rect 47501 4437 47535 4471
rect 47535 4437 47544 4471
rect 47492 4428 47544 4437
rect 47584 4428 47636 4480
rect 49424 4428 49476 4480
rect 55864 4496 55916 4548
rect 56140 4496 56192 4548
rect 58348 4632 58400 4684
rect 57244 4607 57296 4616
rect 57244 4573 57253 4607
rect 57253 4573 57287 4607
rect 57287 4573 57296 4607
rect 57244 4564 57296 4573
rect 57336 4564 57388 4616
rect 61200 4709 61209 4743
rect 61209 4709 61243 4743
rect 61243 4709 61252 4743
rect 61200 4700 61252 4709
rect 64696 4700 64748 4752
rect 65340 4700 65392 4752
rect 58532 4632 58584 4684
rect 59912 4632 59964 4684
rect 58716 4607 58768 4616
rect 58716 4573 58725 4607
rect 58725 4573 58759 4607
rect 58759 4573 58768 4607
rect 58716 4564 58768 4573
rect 59084 4564 59136 4616
rect 62948 4564 63000 4616
rect 63592 4632 63644 4684
rect 64052 4675 64104 4684
rect 64052 4641 64061 4675
rect 64061 4641 64095 4675
rect 64095 4641 64104 4675
rect 64052 4632 64104 4641
rect 64420 4632 64472 4684
rect 67364 4675 67416 4684
rect 67364 4641 67373 4675
rect 67373 4641 67407 4675
rect 67407 4641 67416 4675
rect 67364 4632 67416 4641
rect 67640 4675 67692 4684
rect 67640 4641 67649 4675
rect 67649 4641 67683 4675
rect 67683 4641 67692 4675
rect 67640 4632 67692 4641
rect 73804 4700 73856 4752
rect 74448 4700 74500 4752
rect 76472 4700 76524 4752
rect 63868 4564 63920 4616
rect 72056 4632 72108 4684
rect 74264 4632 74316 4684
rect 74632 4632 74684 4684
rect 76380 4632 76432 4684
rect 78036 4700 78088 4752
rect 57704 4539 57756 4548
rect 57704 4505 57713 4539
rect 57713 4505 57747 4539
rect 57747 4505 57756 4539
rect 57704 4496 57756 4505
rect 57888 4539 57940 4548
rect 57888 4505 57897 4539
rect 57897 4505 57931 4539
rect 57931 4505 57940 4539
rect 57888 4496 57940 4505
rect 57796 4428 57848 4480
rect 66812 4496 66864 4548
rect 67732 4496 67784 4548
rect 73252 4564 73304 4616
rect 73436 4607 73488 4616
rect 73436 4573 73445 4607
rect 73445 4573 73479 4607
rect 73479 4573 73488 4607
rect 73436 4564 73488 4573
rect 73528 4607 73580 4616
rect 73528 4573 73537 4607
rect 73537 4573 73571 4607
rect 73571 4573 73580 4607
rect 76932 4607 76984 4616
rect 73528 4564 73580 4573
rect 76932 4573 76941 4607
rect 76941 4573 76975 4607
rect 76975 4573 76984 4607
rect 76932 4564 76984 4573
rect 73712 4539 73764 4548
rect 71596 4428 71648 4480
rect 73712 4505 73721 4539
rect 73721 4505 73755 4539
rect 73755 4505 73764 4539
rect 73712 4496 73764 4505
rect 74172 4539 74224 4548
rect 74172 4505 74181 4539
rect 74181 4505 74215 4539
rect 74215 4505 74224 4539
rect 74172 4496 74224 4505
rect 73528 4428 73580 4480
rect 78404 4496 78456 4548
rect 77392 4428 77444 4480
rect 78772 4496 78824 4548
rect 78680 4428 78732 4480
rect 79876 4768 79928 4820
rect 82452 4811 82504 4820
rect 82452 4777 82461 4811
rect 82461 4777 82495 4811
rect 82495 4777 82504 4811
rect 82452 4768 82504 4777
rect 79968 4632 80020 4684
rect 80704 4564 80756 4616
rect 81532 4607 81584 4616
rect 79692 4496 79744 4548
rect 81532 4573 81541 4607
rect 81541 4573 81575 4607
rect 81575 4573 81584 4607
rect 81532 4564 81584 4573
rect 82728 4564 82780 4616
rect 84292 4768 84344 4820
rect 84384 4700 84436 4752
rect 84936 4700 84988 4752
rect 85856 4700 85908 4752
rect 83372 4607 83424 4616
rect 83372 4573 83381 4607
rect 83381 4573 83415 4607
rect 83415 4573 83424 4607
rect 83372 4564 83424 4573
rect 83648 4607 83700 4616
rect 83648 4573 83657 4607
rect 83657 4573 83691 4607
rect 83691 4573 83700 4607
rect 83648 4564 83700 4573
rect 83740 4564 83792 4616
rect 86684 4632 86736 4684
rect 87052 4768 87104 4820
rect 87144 4768 87196 4820
rect 88064 4768 88116 4820
rect 84384 4607 84436 4616
rect 84384 4573 84393 4607
rect 84393 4573 84427 4607
rect 84427 4573 84436 4607
rect 84384 4564 84436 4573
rect 84660 4564 84712 4616
rect 85856 4607 85908 4616
rect 81716 4496 81768 4548
rect 83832 4496 83884 4548
rect 85856 4573 85865 4607
rect 85865 4573 85899 4607
rect 85899 4573 85908 4607
rect 85856 4564 85908 4573
rect 86592 4564 86644 4616
rect 87236 4564 87288 4616
rect 88524 4675 88576 4684
rect 88524 4641 88533 4675
rect 88533 4641 88567 4675
rect 88567 4641 88576 4675
rect 88524 4632 88576 4641
rect 87696 4607 87748 4616
rect 87696 4573 87705 4607
rect 87705 4573 87739 4607
rect 87739 4573 87748 4607
rect 87696 4564 87748 4573
rect 88616 4607 88668 4616
rect 88616 4573 88625 4607
rect 88625 4573 88659 4607
rect 88659 4573 88668 4607
rect 88616 4564 88668 4573
rect 90824 4607 90876 4616
rect 90824 4573 90833 4607
rect 90833 4573 90867 4607
rect 90867 4573 90876 4607
rect 90824 4564 90876 4573
rect 92020 4607 92072 4616
rect 92020 4573 92029 4607
rect 92029 4573 92063 4607
rect 92063 4573 92072 4607
rect 92020 4564 92072 4573
rect 88892 4496 88944 4548
rect 89628 4539 89680 4548
rect 82452 4428 82504 4480
rect 85120 4428 85172 4480
rect 87052 4428 87104 4480
rect 89352 4428 89404 4480
rect 89628 4505 89637 4539
rect 89637 4505 89671 4539
rect 89671 4505 89680 4539
rect 89628 4496 89680 4505
rect 89812 4539 89864 4548
rect 89812 4505 89821 4539
rect 89821 4505 89855 4539
rect 89855 4505 89864 4539
rect 89812 4496 89864 4505
rect 92112 4496 92164 4548
rect 90272 4428 90324 4480
rect 90916 4428 90968 4480
rect 92296 4496 92348 4548
rect 93124 4428 93176 4480
rect 93676 4471 93728 4480
rect 93676 4437 93685 4471
rect 93685 4437 93719 4471
rect 93719 4437 93728 4471
rect 93676 4428 93728 4437
rect 94228 4471 94280 4480
rect 94228 4437 94237 4471
rect 94237 4437 94271 4471
rect 94271 4437 94280 4471
rect 94228 4428 94280 4437
rect 24386 4326 24438 4378
rect 24450 4326 24502 4378
rect 24514 4326 24566 4378
rect 24578 4326 24630 4378
rect 24642 4326 24694 4378
rect 47823 4326 47875 4378
rect 47887 4326 47939 4378
rect 47951 4326 48003 4378
rect 48015 4326 48067 4378
rect 48079 4326 48131 4378
rect 71260 4326 71312 4378
rect 71324 4326 71376 4378
rect 71388 4326 71440 4378
rect 71452 4326 71504 4378
rect 71516 4326 71568 4378
rect 94697 4326 94749 4378
rect 94761 4326 94813 4378
rect 94825 4326 94877 4378
rect 94889 4326 94941 4378
rect 94953 4326 95005 4378
rect 15384 4224 15436 4276
rect 31392 4224 31444 4276
rect 35348 4224 35400 4276
rect 42156 4224 42208 4276
rect 9128 4088 9180 4140
rect 9864 4131 9916 4140
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 10692 4156 10744 4208
rect 15476 4156 15528 4208
rect 24216 4156 24268 4208
rect 25044 4156 25096 4208
rect 26148 4199 26200 4208
rect 26148 4165 26157 4199
rect 26157 4165 26191 4199
rect 26191 4165 26200 4199
rect 26148 4156 26200 4165
rect 30012 4156 30064 4208
rect 32680 4156 32732 4208
rect 33416 4199 33468 4208
rect 33416 4165 33425 4199
rect 33425 4165 33459 4199
rect 33459 4165 33468 4199
rect 33416 4156 33468 4165
rect 33600 4199 33652 4208
rect 33600 4165 33609 4199
rect 33609 4165 33643 4199
rect 33643 4165 33652 4199
rect 33600 4156 33652 4165
rect 41236 4156 41288 4208
rect 43996 4224 44048 4276
rect 51540 4224 51592 4276
rect 57704 4224 57756 4276
rect 10600 4131 10652 4140
rect 9864 4088 9916 4097
rect 10600 4097 10609 4131
rect 10609 4097 10643 4131
rect 10643 4097 10652 4131
rect 10600 4088 10652 4097
rect 14832 4131 14884 4140
rect 14832 4097 14841 4131
rect 14841 4097 14875 4131
rect 14875 4097 14884 4131
rect 14832 4088 14884 4097
rect 25688 4088 25740 4140
rect 30840 4088 30892 4140
rect 34612 4131 34664 4140
rect 34612 4097 34621 4131
rect 34621 4097 34655 4131
rect 34655 4097 34664 4131
rect 34612 4088 34664 4097
rect 38844 4088 38896 4140
rect 39948 4088 40000 4140
rect 41788 4088 41840 4140
rect 43812 4131 43864 4140
rect 43812 4097 43821 4131
rect 43821 4097 43855 4131
rect 43855 4097 43864 4131
rect 43812 4088 43864 4097
rect 50436 4088 50488 4140
rect 52184 4156 52236 4208
rect 55496 4199 55548 4208
rect 55496 4165 55505 4199
rect 55505 4165 55539 4199
rect 55539 4165 55548 4199
rect 55496 4156 55548 4165
rect 56416 4156 56468 4208
rect 59452 4224 59504 4276
rect 62212 4224 62264 4276
rect 63500 4224 63552 4276
rect 62304 4156 62356 4208
rect 51264 4088 51316 4140
rect 52276 4131 52328 4140
rect 52276 4097 52285 4131
rect 52285 4097 52319 4131
rect 52319 4097 52328 4131
rect 52276 4088 52328 4097
rect 53196 4131 53248 4140
rect 53196 4097 53205 4131
rect 53205 4097 53239 4131
rect 53239 4097 53248 4131
rect 53196 4088 53248 4097
rect 54668 4088 54720 4140
rect 13084 4063 13136 4072
rect 13084 4029 13093 4063
rect 13093 4029 13127 4063
rect 13127 4029 13136 4063
rect 13084 4020 13136 4029
rect 14556 4063 14608 4072
rect 14556 4029 14565 4063
rect 14565 4029 14599 4063
rect 14599 4029 14608 4063
rect 14556 4020 14608 4029
rect 25412 4020 25464 4072
rect 37464 4063 37516 4072
rect 37464 4029 37473 4063
rect 37473 4029 37507 4063
rect 37507 4029 37516 4063
rect 37464 4020 37516 4029
rect 37740 4063 37792 4072
rect 37740 4029 37749 4063
rect 37749 4029 37783 4063
rect 37783 4029 37792 4063
rect 37740 4020 37792 4029
rect 38476 4020 38528 4072
rect 40684 4020 40736 4072
rect 40776 4063 40828 4072
rect 40776 4029 40785 4063
rect 40785 4029 40819 4063
rect 40819 4029 40828 4063
rect 40776 4020 40828 4029
rect 48320 4020 48372 4072
rect 49148 4063 49200 4072
rect 49148 4029 49157 4063
rect 49157 4029 49191 4063
rect 49191 4029 49200 4063
rect 49148 4020 49200 4029
rect 10324 3952 10376 4004
rect 13544 3952 13596 4004
rect 47400 3952 47452 4004
rect 55128 4063 55180 4072
rect 55128 4029 55137 4063
rect 55137 4029 55171 4063
rect 55171 4029 55180 4063
rect 55128 4020 55180 4029
rect 57888 4088 57940 4140
rect 58072 4088 58124 4140
rect 62028 4131 62080 4140
rect 62028 4097 62037 4131
rect 62037 4097 62071 4131
rect 62071 4097 62080 4131
rect 62028 4088 62080 4097
rect 62580 4131 62632 4140
rect 62580 4097 62589 4131
rect 62589 4097 62623 4131
rect 62623 4097 62632 4131
rect 62580 4088 62632 4097
rect 62948 4088 63000 4140
rect 71872 4224 71924 4276
rect 73988 4224 74040 4276
rect 71596 4156 71648 4208
rect 73436 4156 73488 4208
rect 74172 4156 74224 4208
rect 75920 4267 75972 4276
rect 75920 4233 75929 4267
rect 75929 4233 75963 4267
rect 75963 4233 75972 4267
rect 75920 4224 75972 4233
rect 77300 4224 77352 4276
rect 77484 4267 77536 4276
rect 77484 4233 77493 4267
rect 77493 4233 77527 4267
rect 77527 4233 77536 4267
rect 77484 4224 77536 4233
rect 76932 4156 76984 4208
rect 79968 4224 80020 4276
rect 80244 4224 80296 4276
rect 83740 4224 83792 4276
rect 84016 4267 84068 4276
rect 84016 4233 84025 4267
rect 84025 4233 84059 4267
rect 84059 4233 84068 4267
rect 84016 4224 84068 4233
rect 84660 4224 84712 4276
rect 85120 4224 85172 4276
rect 87144 4224 87196 4276
rect 90272 4267 90324 4276
rect 90272 4233 90281 4267
rect 90281 4233 90315 4267
rect 90315 4233 90324 4267
rect 90272 4224 90324 4233
rect 91928 4224 91980 4276
rect 78404 4156 78456 4208
rect 80612 4156 80664 4208
rect 84568 4156 84620 4208
rect 88616 4156 88668 4208
rect 71228 4131 71280 4140
rect 71228 4097 71237 4131
rect 71237 4097 71271 4131
rect 71271 4097 71280 4131
rect 71228 4088 71280 4097
rect 73712 4088 73764 4140
rect 57060 4063 57112 4072
rect 55956 3952 56008 4004
rect 57060 4029 57069 4063
rect 57069 4029 57103 4063
rect 57103 4029 57112 4063
rect 57060 4020 57112 4029
rect 58716 4020 58768 4072
rect 10692 3884 10744 3936
rect 15200 3884 15252 3936
rect 37924 3884 37976 3936
rect 38108 3884 38160 3936
rect 40592 3884 40644 3936
rect 49148 3884 49200 3936
rect 51080 3884 51132 3936
rect 56232 3884 56284 3936
rect 57796 3952 57848 4004
rect 61292 4020 61344 4072
rect 64788 4020 64840 4072
rect 68652 4020 68704 4072
rect 73528 4020 73580 4072
rect 74356 4063 74408 4072
rect 74356 4029 74365 4063
rect 74365 4029 74399 4063
rect 74399 4029 74408 4063
rect 74356 4020 74408 4029
rect 74448 4020 74500 4072
rect 75184 4063 75236 4072
rect 75184 4029 75193 4063
rect 75193 4029 75227 4063
rect 75227 4029 75236 4063
rect 75184 4020 75236 4029
rect 78036 4020 78088 4072
rect 62028 3952 62080 4004
rect 57060 3884 57112 3936
rect 59360 3884 59412 3936
rect 62672 3884 62724 3936
rect 63776 3952 63828 4004
rect 64880 3952 64932 4004
rect 73712 3995 73764 4004
rect 73712 3961 73721 3995
rect 73721 3961 73755 3995
rect 73755 3961 73764 3995
rect 73712 3952 73764 3961
rect 76196 3952 76248 4004
rect 67732 3884 67784 3936
rect 73620 3927 73672 3936
rect 73620 3893 73629 3927
rect 73629 3893 73663 3927
rect 73663 3893 73672 3927
rect 73620 3884 73672 3893
rect 76380 3884 76432 3936
rect 80520 4088 80572 4140
rect 81992 4088 82044 4140
rect 83556 4088 83608 4140
rect 83832 4131 83884 4140
rect 83832 4097 83841 4131
rect 83841 4097 83875 4131
rect 83875 4097 83884 4131
rect 83832 4088 83884 4097
rect 84844 4131 84896 4140
rect 84844 4097 84853 4131
rect 84853 4097 84887 4131
rect 84887 4097 84896 4131
rect 84844 4088 84896 4097
rect 85488 4131 85540 4140
rect 85488 4097 85497 4131
rect 85497 4097 85531 4131
rect 85531 4097 85540 4131
rect 85488 4088 85540 4097
rect 86132 4088 86184 4140
rect 86960 4131 87012 4140
rect 86960 4097 86969 4131
rect 86969 4097 87003 4131
rect 87003 4097 87012 4131
rect 86960 4088 87012 4097
rect 87236 4088 87288 4140
rect 87972 4131 88024 4140
rect 87972 4097 87981 4131
rect 87981 4097 88015 4131
rect 88015 4097 88024 4131
rect 87972 4088 88024 4097
rect 89812 4156 89864 4208
rect 89996 4131 90048 4140
rect 89996 4097 90005 4131
rect 90005 4097 90039 4131
rect 90039 4097 90048 4131
rect 89996 4088 90048 4097
rect 78588 4020 78640 4072
rect 79968 4020 80020 4072
rect 80704 4020 80756 4072
rect 84200 3952 84252 4004
rect 84936 3952 84988 4004
rect 81992 3884 82044 3936
rect 89628 4020 89680 4072
rect 89076 3952 89128 4004
rect 89904 3952 89956 4004
rect 93124 4020 93176 4072
rect 88984 3927 89036 3936
rect 88984 3893 88993 3927
rect 88993 3893 89027 3927
rect 89027 3893 89036 3927
rect 88984 3884 89036 3893
rect 91008 3884 91060 3936
rect 94228 4020 94280 4072
rect 12668 3782 12720 3834
rect 12732 3782 12784 3834
rect 12796 3782 12848 3834
rect 12860 3782 12912 3834
rect 12924 3782 12976 3834
rect 36105 3782 36157 3834
rect 36169 3782 36221 3834
rect 36233 3782 36285 3834
rect 36297 3782 36349 3834
rect 36361 3782 36413 3834
rect 59542 3782 59594 3834
rect 59606 3782 59658 3834
rect 59670 3782 59722 3834
rect 59734 3782 59786 3834
rect 59798 3782 59850 3834
rect 82979 3782 83031 3834
rect 83043 3782 83095 3834
rect 83107 3782 83159 3834
rect 83171 3782 83223 3834
rect 83235 3782 83287 3834
rect 4068 3680 4120 3732
rect 10968 3680 11020 3732
rect 13544 3680 13596 3732
rect 32312 3680 32364 3732
rect 32956 3612 33008 3664
rect 38108 3612 38160 3664
rect 39948 3612 40000 3664
rect 37464 3544 37516 3596
rect 40408 3544 40460 3596
rect 40592 3680 40644 3732
rect 55496 3680 55548 3732
rect 40776 3612 40828 3664
rect 49792 3612 49844 3664
rect 51080 3655 51132 3664
rect 51080 3621 51089 3655
rect 51089 3621 51123 3655
rect 51123 3621 51132 3655
rect 54208 3655 54260 3664
rect 51080 3612 51132 3621
rect 54208 3621 54217 3655
rect 54217 3621 54251 3655
rect 54251 3621 54260 3655
rect 54208 3612 54260 3621
rect 54668 3655 54720 3664
rect 54668 3621 54677 3655
rect 54677 3621 54711 3655
rect 54711 3621 54720 3655
rect 54668 3612 54720 3621
rect 10600 3476 10652 3528
rect 15200 3519 15252 3528
rect 15200 3485 15209 3519
rect 15209 3485 15243 3519
rect 15243 3485 15252 3519
rect 15200 3476 15252 3485
rect 15476 3519 15528 3528
rect 15476 3485 15485 3519
rect 15485 3485 15519 3519
rect 15519 3485 15528 3519
rect 15476 3476 15528 3485
rect 38844 3408 38896 3460
rect 41328 3408 41380 3460
rect 24216 3340 24268 3392
rect 39028 3340 39080 3392
rect 55956 3587 56008 3596
rect 55956 3553 55965 3587
rect 55965 3553 55999 3587
rect 55999 3553 56008 3587
rect 55956 3544 56008 3553
rect 53840 3476 53892 3528
rect 52368 3408 52420 3460
rect 53380 3451 53432 3460
rect 53380 3417 53389 3451
rect 53389 3417 53423 3451
rect 53423 3417 53432 3451
rect 53380 3408 53432 3417
rect 55128 3408 55180 3460
rect 57336 3476 57388 3528
rect 58532 3680 58584 3732
rect 59268 3723 59320 3732
rect 59268 3689 59277 3723
rect 59277 3689 59311 3723
rect 59311 3689 59320 3723
rect 59268 3680 59320 3689
rect 61200 3680 61252 3732
rect 64604 3680 64656 3732
rect 67180 3680 67232 3732
rect 64696 3612 64748 3664
rect 55864 3408 55916 3460
rect 64328 3544 64380 3596
rect 62212 3476 62264 3528
rect 64604 3476 64656 3528
rect 68652 3680 68704 3732
rect 72056 3655 72108 3664
rect 72056 3621 72065 3655
rect 72065 3621 72099 3655
rect 72099 3621 72108 3655
rect 72056 3612 72108 3621
rect 73620 3612 73672 3664
rect 75920 3612 75972 3664
rect 76288 3612 76340 3664
rect 80704 3655 80756 3664
rect 80704 3621 80713 3655
rect 80713 3621 80747 3655
rect 80747 3621 80756 3655
rect 80704 3612 80756 3621
rect 84844 3612 84896 3664
rect 74448 3544 74500 3596
rect 78772 3544 78824 3596
rect 62304 3408 62356 3460
rect 65892 3408 65944 3460
rect 73804 3476 73856 3528
rect 76380 3476 76432 3528
rect 57428 3383 57480 3392
rect 57428 3349 57437 3383
rect 57437 3349 57471 3383
rect 57471 3349 57480 3383
rect 57428 3340 57480 3349
rect 68376 3340 68428 3392
rect 71228 3340 71280 3392
rect 72884 3383 72936 3392
rect 72884 3349 72893 3383
rect 72893 3349 72927 3383
rect 72927 3349 72936 3383
rect 72884 3340 72936 3349
rect 73712 3408 73764 3460
rect 73988 3383 74040 3392
rect 73988 3349 73997 3383
rect 73997 3349 74031 3383
rect 74031 3349 74040 3383
rect 73988 3340 74040 3349
rect 77852 3383 77904 3392
rect 77852 3349 77861 3383
rect 77861 3349 77895 3383
rect 77895 3349 77904 3383
rect 77852 3340 77904 3349
rect 81716 3519 81768 3528
rect 79048 3408 79100 3460
rect 79232 3408 79284 3460
rect 81716 3485 81725 3519
rect 81725 3485 81759 3519
rect 81759 3485 81768 3519
rect 81716 3476 81768 3485
rect 81992 3519 82044 3528
rect 81992 3485 82001 3519
rect 82001 3485 82035 3519
rect 82035 3485 82044 3519
rect 83648 3544 83700 3596
rect 85672 3544 85724 3596
rect 82728 3519 82780 3528
rect 81992 3476 82044 3485
rect 82728 3485 82737 3519
rect 82737 3485 82771 3519
rect 82771 3485 82780 3519
rect 82728 3476 82780 3485
rect 84936 3476 84988 3528
rect 79876 3408 79928 3460
rect 86040 3680 86092 3732
rect 88524 3680 88576 3732
rect 89996 3680 90048 3732
rect 90916 3680 90968 3732
rect 93216 3723 93268 3732
rect 93216 3689 93225 3723
rect 93225 3689 93259 3723
rect 93259 3689 93268 3723
rect 93216 3680 93268 3689
rect 87236 3612 87288 3664
rect 88984 3612 89036 3664
rect 93676 3612 93728 3664
rect 88892 3544 88944 3596
rect 89352 3587 89404 3596
rect 89352 3553 89361 3587
rect 89361 3553 89395 3587
rect 89395 3553 89404 3587
rect 89352 3544 89404 3553
rect 87052 3519 87104 3528
rect 87052 3485 87061 3519
rect 87061 3485 87095 3519
rect 87095 3485 87104 3519
rect 87052 3476 87104 3485
rect 89076 3519 89128 3528
rect 86868 3408 86920 3460
rect 89076 3485 89085 3519
rect 89085 3485 89119 3519
rect 89119 3485 89128 3519
rect 89076 3476 89128 3485
rect 91928 3519 91980 3528
rect 91928 3485 91937 3519
rect 91937 3485 91971 3519
rect 91971 3485 91980 3519
rect 91928 3476 91980 3485
rect 89904 3408 89956 3460
rect 80704 3340 80756 3392
rect 93768 3340 93820 3392
rect 24386 3238 24438 3290
rect 24450 3238 24502 3290
rect 24514 3238 24566 3290
rect 24578 3238 24630 3290
rect 24642 3238 24694 3290
rect 47823 3238 47875 3290
rect 47887 3238 47939 3290
rect 47951 3238 48003 3290
rect 48015 3238 48067 3290
rect 48079 3238 48131 3290
rect 71260 3238 71312 3290
rect 71324 3238 71376 3290
rect 71388 3238 71440 3290
rect 71452 3238 71504 3290
rect 71516 3238 71568 3290
rect 94697 3238 94749 3290
rect 94761 3238 94813 3290
rect 94825 3238 94877 3290
rect 94889 3238 94941 3290
rect 94953 3238 95005 3290
rect 37740 3136 37792 3188
rect 38844 3136 38896 3188
rect 53840 3179 53892 3188
rect 53840 3145 53849 3179
rect 53849 3145 53883 3179
rect 53883 3145 53892 3179
rect 53840 3136 53892 3145
rect 39028 3111 39080 3120
rect 39028 3077 39037 3111
rect 39037 3077 39071 3111
rect 39071 3077 39080 3111
rect 39028 3068 39080 3077
rect 53932 3068 53984 3120
rect 40408 3000 40460 3052
rect 51264 3043 51316 3052
rect 51264 3009 51273 3043
rect 51273 3009 51307 3043
rect 51307 3009 51316 3043
rect 51264 3000 51316 3009
rect 52368 3000 52420 3052
rect 55036 3136 55088 3188
rect 55864 3136 55916 3188
rect 56232 3179 56284 3188
rect 56232 3145 56241 3179
rect 56241 3145 56275 3179
rect 56275 3145 56284 3179
rect 56232 3136 56284 3145
rect 56784 3136 56836 3188
rect 57336 3136 57388 3188
rect 57428 3136 57480 3188
rect 61292 3111 61344 3120
rect 61292 3077 61301 3111
rect 61301 3077 61335 3111
rect 61335 3077 61344 3111
rect 61292 3068 61344 3077
rect 62304 3068 62356 3120
rect 64788 3136 64840 3188
rect 78588 3136 78640 3188
rect 79232 3179 79284 3188
rect 79232 3145 79241 3179
rect 79241 3145 79275 3179
rect 79275 3145 79284 3179
rect 79232 3136 79284 3145
rect 72884 3068 72936 3120
rect 74632 3068 74684 3120
rect 76288 3111 76340 3120
rect 76288 3077 76297 3111
rect 76297 3077 76331 3111
rect 76331 3077 76340 3111
rect 76288 3068 76340 3077
rect 78036 3111 78088 3120
rect 78036 3077 78045 3111
rect 78045 3077 78079 3111
rect 78079 3077 78088 3111
rect 78036 3068 78088 3077
rect 81440 3136 81492 3188
rect 81532 3179 81584 3188
rect 81532 3145 81541 3179
rect 81541 3145 81575 3179
rect 81575 3145 81584 3179
rect 81532 3136 81584 3145
rect 81992 3136 82044 3188
rect 84936 3136 84988 3188
rect 86868 3136 86920 3188
rect 90824 3136 90876 3188
rect 91008 3179 91060 3188
rect 91008 3145 91017 3179
rect 91017 3145 91051 3179
rect 91051 3145 91060 3179
rect 91008 3136 91060 3145
rect 92388 3136 92440 3188
rect 89628 3068 89680 3120
rect 55128 3000 55180 3052
rect 54392 2932 54444 2984
rect 55496 2932 55548 2984
rect 57060 2864 57112 2916
rect 77852 3000 77904 3052
rect 79876 3043 79928 3052
rect 79876 3009 79885 3043
rect 79885 3009 79919 3043
rect 79919 3009 79928 3043
rect 79876 3000 79928 3009
rect 85672 3000 85724 3052
rect 64972 2975 65024 2984
rect 64972 2941 64981 2975
rect 64981 2941 65015 2975
rect 65015 2941 65024 2975
rect 64972 2932 65024 2941
rect 78680 2932 78732 2984
rect 81716 2932 81768 2984
rect 83372 2932 83424 2984
rect 86132 2932 86184 2984
rect 89076 2932 89128 2984
rect 91008 2932 91060 2984
rect 91928 2932 91980 2984
rect 78680 2796 78732 2848
rect 12668 2694 12720 2746
rect 12732 2694 12784 2746
rect 12796 2694 12848 2746
rect 12860 2694 12912 2746
rect 12924 2694 12976 2746
rect 36105 2694 36157 2746
rect 36169 2694 36221 2746
rect 36233 2694 36285 2746
rect 36297 2694 36349 2746
rect 36361 2694 36413 2746
rect 59542 2694 59594 2746
rect 59606 2694 59658 2746
rect 59670 2694 59722 2746
rect 59734 2694 59786 2746
rect 59798 2694 59850 2746
rect 82979 2694 83031 2746
rect 83043 2694 83095 2746
rect 83107 2694 83159 2746
rect 83171 2694 83223 2746
rect 83235 2694 83287 2746
rect 37372 2592 37424 2644
rect 38844 2592 38896 2644
rect 41328 2592 41380 2644
rect 54392 2635 54444 2644
rect 54392 2601 54401 2635
rect 54401 2601 54435 2635
rect 54435 2601 54444 2635
rect 54392 2592 54444 2601
rect 64328 2635 64380 2644
rect 64328 2601 64337 2635
rect 64337 2601 64371 2635
rect 64371 2601 64380 2635
rect 64328 2592 64380 2601
rect 64972 2592 65024 2644
rect 75276 2592 75328 2644
rect 78588 2592 78640 2644
rect 78772 2635 78824 2644
rect 78772 2601 78781 2635
rect 78781 2601 78815 2635
rect 78815 2601 78824 2635
rect 78772 2592 78824 2601
rect 86868 2635 86920 2644
rect 86868 2601 86877 2635
rect 86877 2601 86911 2635
rect 86911 2601 86920 2635
rect 86868 2592 86920 2601
rect 90916 2635 90968 2644
rect 90916 2601 90925 2635
rect 90925 2601 90959 2635
rect 90959 2601 90968 2635
rect 90916 2592 90968 2601
rect 4160 2388 4212 2440
rect 13360 2431 13412 2440
rect 4436 2252 4488 2304
rect 12348 2252 12400 2304
rect 13360 2397 13369 2431
rect 13369 2397 13403 2431
rect 13403 2397 13412 2431
rect 13360 2388 13412 2397
rect 15476 2388 15528 2440
rect 28448 2431 28500 2440
rect 28448 2397 28457 2431
rect 28457 2397 28491 2431
rect 28491 2397 28500 2431
rect 28448 2388 28500 2397
rect 36084 2388 36136 2440
rect 65892 2524 65944 2576
rect 56324 2388 56376 2440
rect 68376 2431 68428 2440
rect 68376 2397 68385 2431
rect 68385 2397 68419 2431
rect 68419 2397 68428 2431
rect 68376 2388 68428 2397
rect 74816 2388 74868 2440
rect 75276 2320 75328 2372
rect 20352 2252 20404 2304
rect 28172 2252 28224 2304
rect 43996 2252 44048 2304
rect 51908 2252 51960 2304
rect 59820 2252 59872 2304
rect 67732 2252 67784 2304
rect 91468 2388 91520 2440
rect 75644 2252 75696 2304
rect 83556 2252 83608 2304
rect 24386 2150 24438 2202
rect 24450 2150 24502 2202
rect 24514 2150 24566 2202
rect 24578 2150 24630 2202
rect 24642 2150 24694 2202
rect 47823 2150 47875 2202
rect 47887 2150 47939 2202
rect 47951 2150 48003 2202
rect 48015 2150 48067 2202
rect 48079 2150 48131 2202
rect 71260 2150 71312 2202
rect 71324 2150 71376 2202
rect 71388 2150 71440 2202
rect 71452 2150 71504 2202
rect 71516 2150 71568 2202
rect 94697 2150 94749 2202
rect 94761 2150 94813 2202
rect 94825 2150 94877 2202
rect 94889 2150 94941 2202
rect 94953 2150 95005 2202
<< metal2 >>
rect 4434 19200 4490 20000
rect 12346 19200 12402 20000
rect 20258 19200 20314 20000
rect 28170 19200 28226 20000
rect 36082 19200 36138 20000
rect 43994 19200 44050 20000
rect 51906 19200 51962 20000
rect 59818 19200 59874 20000
rect 67730 19200 67786 20000
rect 75642 19200 75698 20000
rect 83554 19200 83610 20000
rect 91466 19200 91522 20000
rect 4448 17338 4476 19200
rect 12360 17354 12388 19200
rect 12360 17338 12480 17354
rect 20272 17338 20300 19200
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 4436 17332 4488 17338
rect 12360 17332 12492 17338
rect 12360 17326 12440 17332
rect 4436 17274 4488 17280
rect 12440 17274 12492 17280
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 1584 17196 1636 17202
rect 1584 17138 1636 17144
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 1596 16726 1624 17138
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 1584 16720 1636 16726
rect 1582 16688 1584 16697
rect 1636 16688 1638 16697
rect 1582 16623 1638 16632
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 2976 13394 3004 13874
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 2976 12238 3004 13330
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3436 12714 3464 13126
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 4080 12306 4108 13330
rect 4172 13326 4200 13874
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4816 13433 4844 13670
rect 5092 13530 5120 16934
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 4802 13424 4858 13433
rect 4802 13359 4858 13368
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4172 12918 4200 13262
rect 4436 13252 4488 13258
rect 4436 13194 4488 13200
rect 4448 12986 4476 13194
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 4540 12442 4568 13126
rect 5092 12850 5120 13466
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 3068 11830 3096 12038
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3056 11824 3108 11830
rect 3056 11766 3108 11772
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1596 10062 1624 11494
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1780 10810 1808 11290
rect 2332 11082 2360 11630
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2516 11150 2544 11290
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 3884 11144 3936 11150
rect 3988 11098 4016 11834
rect 3936 11092 4016 11098
rect 3884 11086 4016 11092
rect 2320 11076 2372 11082
rect 2320 11018 2372 11024
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 2332 10606 2360 11018
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 1584 10056 1636 10062
rect 1582 10024 1584 10033
rect 2228 10056 2280 10062
rect 1636 10024 1638 10033
rect 2332 10044 2360 10542
rect 2516 10062 2544 11086
rect 3896 11070 4016 11086
rect 3424 11008 3476 11014
rect 3424 10950 3476 10956
rect 3436 10198 3464 10950
rect 3988 10742 4016 11070
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 3424 10192 3476 10198
rect 3424 10134 3476 10140
rect 2280 10016 2360 10044
rect 2228 9998 2280 10004
rect 1582 9959 1638 9968
rect 2332 9654 2360 10016
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2148 8838 2176 9522
rect 2228 9036 2280 9042
rect 2332 9024 2360 9590
rect 2516 9178 2544 9998
rect 3436 9382 3464 10134
rect 3884 10056 3936 10062
rect 3988 10044 4016 10678
rect 4080 10198 4108 12242
rect 5184 12238 5212 12718
rect 5828 12646 5856 13262
rect 6564 12986 6592 17138
rect 8024 14544 8076 14550
rect 8024 14486 8076 14492
rect 8036 14414 8064 14486
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 7300 13938 7328 14350
rect 9128 14340 9180 14346
rect 9128 14282 9180 14288
rect 9140 14074 9168 14282
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 9312 14000 9364 14006
rect 9312 13942 9364 13948
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 13530 6868 13670
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6840 13326 6868 13466
rect 7300 13462 7328 13874
rect 7288 13456 7340 13462
rect 7288 13398 7340 13404
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6840 12850 6868 13262
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 7024 12782 7052 13126
rect 7012 12776 7064 12782
rect 7010 12744 7012 12753
rect 7064 12744 7066 12753
rect 7010 12679 7066 12688
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5644 12434 5672 12582
rect 5552 12406 5672 12434
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5552 12170 5580 12406
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 4540 11898 4568 12106
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 5552 11558 5580 12106
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 6012 11830 6040 12038
rect 6000 11824 6052 11830
rect 6000 11766 6052 11772
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5092 11354 5120 11494
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4540 10266 4568 10610
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 3936 10016 4016 10044
rect 3884 9998 3936 10004
rect 3896 9586 3924 9998
rect 3976 9920 4028 9926
rect 3976 9862 4028 9868
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2280 8996 2360 9024
rect 2228 8978 2280 8984
rect 2516 8974 2544 9114
rect 3252 8974 3280 9318
rect 3436 9178 3464 9318
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 2136 8832 2188 8838
rect 2136 8774 2188 8780
rect 2148 8634 2176 8774
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 3988 8430 4016 9862
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 4080 8974 4108 9046
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2240 7478 2268 8298
rect 2884 8090 2912 8298
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 2228 7472 2280 7478
rect 2228 7414 2280 7420
rect 3712 7342 3740 7822
rect 3988 7342 4016 8366
rect 4080 7478 4108 8910
rect 4264 8430 4292 8978
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4264 7750 4292 8366
rect 4356 8090 4384 9522
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4448 8566 4476 8910
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4540 8362 4568 10066
rect 4632 10062 4660 10950
rect 5000 10810 5028 11086
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4632 9654 4660 9998
rect 4816 9722 4844 10542
rect 5092 10266 5120 11290
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 5460 10538 5488 11222
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4632 9518 4660 9590
rect 5460 9586 5488 10474
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4724 8634 4752 8910
rect 5552 8838 5580 11494
rect 6012 11082 6040 11766
rect 6840 11762 6868 12038
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6932 11354 6960 11630
rect 7104 11620 7156 11626
rect 7104 11562 7156 11568
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 6012 10062 6040 11018
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6656 10130 6684 10406
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6748 9994 6776 10610
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6932 9926 6960 11154
rect 7116 10742 7144 11562
rect 7300 11082 7328 12038
rect 7392 11354 7420 13330
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7668 12918 7696 13126
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 7944 12102 7972 12718
rect 8036 12306 8064 13942
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8128 12782 8156 13466
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 8220 11830 8248 13806
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8496 13190 8524 13330
rect 9324 13326 9352 13942
rect 11348 13734 11376 14418
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8496 12782 8524 13126
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 7932 11688 7984 11694
rect 7984 11648 8156 11676
rect 8680 11665 8708 12786
rect 8852 11824 8904 11830
rect 8852 11766 8904 11772
rect 7932 11630 7984 11636
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 8036 10810 8064 10950
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5828 9178 5856 9522
rect 6932 9382 6960 9862
rect 7116 9586 7144 10474
rect 7484 10470 7512 10610
rect 8128 10470 8156 11648
rect 8666 11656 8722 11665
rect 8666 11591 8722 11600
rect 8482 11248 8538 11257
rect 8482 11183 8484 11192
rect 8536 11183 8538 11192
rect 8484 11154 8536 11160
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 7484 9654 7512 10406
rect 8128 10062 8156 10406
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7668 9586 7696 9998
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7852 9450 7880 9862
rect 8036 9654 8064 9998
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 7840 9444 7892 9450
rect 7840 9386 7892 9392
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 6288 8634 6316 8842
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 5080 8560 5132 8566
rect 5080 8502 5132 8508
rect 5724 8560 5776 8566
rect 6932 8514 6960 9318
rect 7024 9178 7052 9318
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 5724 8502 5776 8508
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3988 5778 4016 7278
rect 4264 6866 4292 7686
rect 4448 7478 4476 7686
rect 4436 7472 4488 7478
rect 4436 7414 4488 7420
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4160 6792 4212 6798
rect 4212 6740 4292 6746
rect 4160 6734 4292 6740
rect 4172 6718 4292 6734
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4080 3369 4108 3674
rect 4066 3360 4122 3369
rect 4066 3295 4122 3304
rect 4172 2446 4200 6598
rect 4264 6458 4292 6718
rect 5092 6662 5120 8502
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5276 7954 5304 8230
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5736 7818 5764 8502
rect 6748 8498 6960 8514
rect 7024 8498 7052 9114
rect 8036 9110 8064 9590
rect 8312 9518 8340 9998
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 6736 8492 6960 8498
rect 6788 8486 6960 8492
rect 7012 8492 7064 8498
rect 6736 8434 6788 8440
rect 7012 8434 7064 8440
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5736 7546 5764 7754
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5092 6458 5120 6598
rect 5184 6458 5212 6802
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5736 6254 5764 7482
rect 6840 7410 6868 8026
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6656 6390 6684 6598
rect 6644 6384 6696 6390
rect 6644 6326 6696 6332
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5736 5710 5764 6190
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 4264 5370 4292 5578
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 5736 5234 5764 5510
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 4356 4826 4384 5170
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 6748 4690 6776 6666
rect 6840 5778 6868 7346
rect 6920 6792 6972 6798
rect 7116 6780 7144 8774
rect 7668 8650 7696 8774
rect 8036 8650 8064 9046
rect 8312 8974 8340 9454
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 7484 8622 7696 8650
rect 7760 8622 8064 8650
rect 7484 8498 7512 8622
rect 7760 8514 7788 8622
rect 7576 8498 7788 8514
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7564 8492 7788 8498
rect 7616 8486 7788 8492
rect 8208 8492 8260 8498
rect 7564 8434 7616 8440
rect 7668 8022 7696 8486
rect 8208 8434 8260 8440
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 8220 7546 8248 8434
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8312 7206 8340 8910
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 6972 6752 7144 6780
rect 7564 6792 7616 6798
rect 6920 6734 6972 6740
rect 7564 6734 7616 6740
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 7576 6390 7604 6734
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 8128 6322 8156 6734
rect 8312 6730 8340 7142
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 8404 5574 8432 6258
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8404 5370 8432 5510
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 7024 4690 7052 4966
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 8404 4622 8432 5306
rect 8496 5098 8524 11018
rect 8864 10674 8892 11766
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8864 9994 8892 10610
rect 8852 9988 8904 9994
rect 8852 9930 8904 9936
rect 8956 9926 8984 12854
rect 9600 12850 9628 12922
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9692 11898 9720 12174
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9416 9602 9444 9862
rect 9232 9586 9444 9602
rect 9220 9580 9444 9586
rect 9272 9574 9444 9580
rect 9220 9522 9272 9528
rect 9232 9110 9260 9522
rect 9416 9518 9444 9574
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9220 9104 9272 9110
rect 9220 9046 9272 9052
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8588 8634 8616 8774
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 9140 8498 9168 8978
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9140 7886 9168 8434
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8588 6730 8616 7686
rect 8576 6724 8628 6730
rect 8576 6666 8628 6672
rect 8588 6118 8616 6666
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 9416 5137 9444 8978
rect 9508 7410 9536 11290
rect 9784 11218 9812 13330
rect 10152 13326 10180 13670
rect 11244 13456 11296 13462
rect 11244 13398 11296 13404
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10508 13320 10560 13326
rect 10560 13268 10732 13274
rect 10508 13262 10732 13268
rect 10520 13258 10732 13262
rect 10520 13252 10744 13258
rect 10520 13246 10692 13252
rect 10520 12782 10548 13246
rect 10692 13194 10744 13200
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 10152 10810 10180 11698
rect 11164 10810 11192 12582
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 10968 10532 11020 10538
rect 10968 10474 11020 10480
rect 10980 9926 11008 10474
rect 11072 10062 11100 10610
rect 11164 10538 11192 10746
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 9784 9042 9812 9862
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9508 5914 9536 7346
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9600 5302 9628 7414
rect 9692 7206 9720 7822
rect 10060 7410 10088 9522
rect 10520 9518 10548 9862
rect 11256 9654 11284 13398
rect 11440 13394 11468 14350
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 11440 13258 11468 13330
rect 11428 13252 11480 13258
rect 11428 13194 11480 13200
rect 11900 12986 11928 17138
rect 12668 16892 12976 16901
rect 12668 16890 12674 16892
rect 12730 16890 12754 16892
rect 12810 16890 12834 16892
rect 12890 16890 12914 16892
rect 12970 16890 12976 16892
rect 12730 16838 12732 16890
rect 12912 16838 12914 16890
rect 12668 16836 12674 16838
rect 12730 16836 12754 16838
rect 12810 16836 12834 16838
rect 12890 16836 12914 16838
rect 12970 16836 12976 16838
rect 12668 16827 12976 16836
rect 20352 16652 20404 16658
rect 20352 16594 20404 16600
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 19628 16182 19656 16390
rect 19616 16176 19668 16182
rect 19616 16118 19668 16124
rect 20364 16046 20392 16594
rect 15384 16040 15436 16046
rect 20352 16040 20404 16046
rect 15384 15982 15436 15988
rect 20350 16008 20352 16017
rect 20404 16008 20406 16017
rect 12668 15804 12976 15813
rect 12668 15802 12674 15804
rect 12730 15802 12754 15804
rect 12810 15802 12834 15804
rect 12890 15802 12914 15804
rect 12970 15802 12976 15804
rect 12730 15750 12732 15802
rect 12912 15750 12914 15802
rect 12668 15748 12674 15750
rect 12730 15748 12754 15750
rect 12810 15748 12834 15750
rect 12890 15748 12914 15750
rect 12970 15748 12976 15750
rect 12668 15739 12976 15748
rect 13910 15056 13966 15065
rect 13910 14991 13966 15000
rect 12714 14920 12770 14929
rect 12532 14884 12584 14890
rect 12714 14855 12716 14864
rect 12532 14826 12584 14832
rect 12768 14855 12770 14864
rect 12716 14826 12768 14832
rect 12544 14414 12572 14826
rect 12668 14716 12976 14725
rect 12668 14714 12674 14716
rect 12730 14714 12754 14716
rect 12810 14714 12834 14716
rect 12890 14714 12914 14716
rect 12970 14714 12976 14716
rect 12730 14662 12732 14714
rect 12912 14662 12914 14714
rect 12668 14660 12674 14662
rect 12730 14660 12754 14662
rect 12810 14660 12834 14662
rect 12890 14660 12914 14662
rect 12970 14660 12976 14662
rect 12668 14651 12976 14660
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 13082 14376 13138 14385
rect 12440 14340 12492 14346
rect 13082 14311 13084 14320
rect 12440 14282 12492 14288
rect 13136 14311 13138 14320
rect 13084 14282 13136 14288
rect 12452 13938 12480 14282
rect 13174 14104 13230 14113
rect 13174 14039 13230 14048
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 11980 13864 12032 13870
rect 11978 13832 11980 13841
rect 12032 13832 12034 13841
rect 11978 13767 12034 13776
rect 12668 13628 12976 13637
rect 12668 13626 12674 13628
rect 12730 13626 12754 13628
rect 12810 13626 12834 13628
rect 12890 13626 12914 13628
rect 12970 13626 12976 13628
rect 12730 13574 12732 13626
rect 12912 13574 12914 13626
rect 12668 13572 12674 13574
rect 12730 13572 12754 13574
rect 12810 13572 12834 13574
rect 12890 13572 12914 13574
rect 12970 13572 12976 13574
rect 12668 13563 12976 13572
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11900 11354 11928 11494
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11808 10266 11836 11086
rect 11886 10704 11942 10713
rect 11886 10639 11942 10648
rect 11900 10538 11928 10639
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10520 8974 10548 9454
rect 11256 9042 11284 9590
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 10508 8968 10560 8974
rect 10876 8968 10928 8974
rect 10508 8910 10560 8916
rect 10796 8928 10876 8956
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 6866 9720 7142
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9692 6322 9720 6802
rect 9876 6322 9904 6802
rect 10152 6662 10180 7822
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10704 6934 10732 7346
rect 10796 7206 10824 8928
rect 10876 8910 10928 8916
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10796 6798 10824 7142
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10508 6724 10560 6730
rect 10508 6666 10560 6672
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10152 6322 10180 6598
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10428 6118 10456 6598
rect 10520 6458 10548 6666
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10796 6322 10824 6734
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10416 6112 10468 6118
rect 10336 6060 10416 6066
rect 10336 6054 10468 6060
rect 10336 6038 10456 6054
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 9402 5128 9458 5137
rect 8484 5092 8536 5098
rect 9402 5063 9458 5072
rect 8484 5034 8536 5040
rect 9876 4622 9904 5510
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9140 4146 9168 4558
rect 9876 4146 9904 4558
rect 10336 4486 10364 6038
rect 10612 4622 10640 6258
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10704 5914 10732 6190
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10796 5574 10824 6122
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 10336 4010 10364 4422
rect 10612 4146 10640 4558
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10704 4214 10732 4422
rect 10692 4208 10744 4214
rect 10888 4185 10916 8366
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11348 7886 11376 8298
rect 11716 8090 11744 9522
rect 11900 9466 11928 10474
rect 11992 10062 12020 12038
rect 12544 11286 12572 12582
rect 12668 12540 12976 12549
rect 12668 12538 12674 12540
rect 12730 12538 12754 12540
rect 12810 12538 12834 12540
rect 12890 12538 12914 12540
rect 12970 12538 12976 12540
rect 12730 12486 12732 12538
rect 12912 12486 12914 12538
rect 12668 12484 12674 12486
rect 12730 12484 12754 12486
rect 12810 12484 12834 12486
rect 12890 12484 12914 12486
rect 12970 12484 12976 12486
rect 12668 12475 12976 12484
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 13004 11937 13032 12106
rect 12990 11928 13046 11937
rect 12990 11863 13046 11872
rect 13188 11694 13216 14039
rect 13924 13938 13952 14991
rect 15016 14816 15068 14822
rect 15016 14758 15068 14764
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 14016 13870 14044 14214
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14016 13462 14044 13806
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 14004 13456 14056 13462
rect 14004 13398 14056 13404
rect 13268 13184 13320 13190
rect 13268 13126 13320 13132
rect 13280 12986 13308 13126
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13372 11762 13400 13398
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13832 12306 13860 12582
rect 13924 12442 13952 12786
rect 14016 12646 14044 13262
rect 14292 12918 14320 13262
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 12668 11452 12976 11461
rect 12668 11450 12674 11452
rect 12730 11450 12754 11452
rect 12810 11450 12834 11452
rect 12890 11450 12914 11452
rect 12970 11450 12976 11452
rect 12730 11398 12732 11450
rect 12912 11398 12914 11450
rect 12668 11396 12674 11398
rect 12730 11396 12754 11398
rect 12810 11396 12834 11398
rect 12890 11396 12914 11398
rect 12970 11396 12976 11398
rect 12668 11387 12976 11396
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 12268 10810 12296 11154
rect 12544 11082 12572 11222
rect 12532 11076 12584 11082
rect 12532 11018 12584 11024
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 12084 9518 12112 10610
rect 12164 10600 12216 10606
rect 12268 10588 12296 10746
rect 13004 10742 13032 11494
rect 13372 11218 13400 11698
rect 13464 11354 13492 12106
rect 13924 11762 13952 12378
rect 14004 12164 14056 12170
rect 14004 12106 14056 12112
rect 14016 11898 14044 12106
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14004 11892 14056 11898
rect 14004 11834 14056 11840
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 12992 10736 13044 10742
rect 12992 10678 13044 10684
rect 12216 10560 12296 10588
rect 12532 10600 12584 10606
rect 12164 10542 12216 10548
rect 12532 10542 12584 10548
rect 12544 10130 12572 10542
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 12668 10364 12976 10373
rect 12668 10362 12674 10364
rect 12730 10362 12754 10364
rect 12810 10362 12834 10364
rect 12890 10362 12914 10364
rect 12970 10362 12976 10364
rect 12730 10310 12732 10362
rect 12912 10310 12914 10362
rect 12668 10308 12674 10310
rect 12730 10308 12754 10310
rect 12810 10308 12834 10310
rect 12890 10308 12914 10310
rect 12970 10308 12976 10310
rect 12668 10299 12976 10308
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12072 9512 12124 9518
rect 11900 9450 12020 9466
rect 12072 9454 12124 9460
rect 11900 9444 12032 9450
rect 11900 9438 11980 9444
rect 11980 9386 12032 9392
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 8634 11928 9318
rect 12544 9042 12572 10066
rect 13004 9654 13032 10406
rect 13556 10130 13584 11630
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13648 10470 13676 10950
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 12668 9276 12976 9285
rect 12668 9274 12674 9276
rect 12730 9274 12754 9276
rect 12810 9274 12834 9276
rect 12890 9274 12914 9276
rect 12970 9274 12976 9276
rect 12730 9222 12732 9274
rect 12912 9222 12914 9274
rect 12668 9220 12674 9222
rect 12730 9220 12754 9222
rect 12810 9220 12834 9222
rect 12890 9220 12914 9222
rect 12970 9220 12976 9222
rect 12668 9211 12976 9220
rect 13464 9110 13492 9522
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11716 7886 11744 8026
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 12360 7818 12388 8434
rect 12544 8090 12572 8978
rect 12668 8188 12976 8197
rect 12668 8186 12674 8188
rect 12730 8186 12754 8188
rect 12810 8186 12834 8188
rect 12890 8186 12914 8188
rect 12970 8186 12976 8188
rect 12730 8134 12732 8186
rect 12912 8134 12914 8186
rect 12668 8132 12674 8134
rect 12730 8132 12754 8134
rect 12810 8132 12834 8134
rect 12890 8132 12914 8134
rect 12970 8132 12976 8134
rect 12668 8123 12976 8132
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 13464 7993 13492 9046
rect 13556 9042 13584 9862
rect 13648 9654 13676 10406
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13832 8974 13860 9998
rect 13924 9994 13952 11698
rect 14384 11286 14412 12038
rect 14476 11626 14504 13806
rect 14568 13394 14596 14418
rect 15028 13977 15056 14758
rect 15396 14550 15424 15982
rect 20350 15943 20406 15952
rect 20364 15917 20392 15943
rect 16946 15600 17002 15609
rect 16946 15535 17002 15544
rect 19616 15564 19668 15570
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15384 14544 15436 14550
rect 15384 14486 15436 14492
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15108 14408 15160 14414
rect 15108 14350 15160 14356
rect 15014 13968 15070 13977
rect 15120 13938 15148 14350
rect 15014 13903 15070 13912
rect 15108 13932 15160 13938
rect 15028 13870 15056 13903
rect 15108 13874 15160 13880
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 15016 13388 15068 13394
rect 15016 13330 15068 13336
rect 15028 12918 15056 13330
rect 15016 12912 15068 12918
rect 15016 12854 15068 12860
rect 15120 12782 15148 13874
rect 15212 13802 15240 14418
rect 15568 14272 15620 14278
rect 15568 14214 15620 14220
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 15580 13258 15608 14214
rect 15764 13734 15792 14894
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 15856 12850 15884 13806
rect 16132 13394 16160 14758
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 16224 14006 16252 14214
rect 16212 14000 16264 14006
rect 16212 13942 16264 13948
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15120 12442 15148 12718
rect 16316 12646 16344 15098
rect 16960 14006 16988 15535
rect 19616 15506 19668 15512
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15764 12306 15792 12378
rect 16120 12368 16172 12374
rect 16120 12310 16172 12316
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 16132 12238 16160 12310
rect 16120 12232 16172 12238
rect 15396 12170 15608 12186
rect 16120 12174 16172 12180
rect 15396 12164 15620 12170
rect 15396 12158 15568 12164
rect 15396 11937 15424 12158
rect 15568 12106 15620 12112
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15382 11928 15438 11937
rect 15382 11863 15438 11872
rect 15396 11830 15424 11863
rect 15384 11824 15436 11830
rect 15384 11766 15436 11772
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 14464 11620 14516 11626
rect 14464 11562 14516 11568
rect 14844 11354 14872 11630
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14096 11280 14148 11286
rect 14096 11222 14148 11228
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14108 10674 14136 11222
rect 15212 11150 15240 11630
rect 15488 11150 15516 12038
rect 16132 11694 16160 12174
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 14832 10736 14884 10742
rect 14832 10678 14884 10684
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 13556 8022 13584 8842
rect 14200 8566 14228 9522
rect 14648 9512 14700 9518
rect 14554 9480 14610 9489
rect 14648 9454 14700 9460
rect 14554 9415 14556 9424
rect 14608 9415 14610 9424
rect 14556 9386 14608 9392
rect 14660 9178 14688 9454
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14844 9110 14872 10678
rect 14924 9716 14976 9722
rect 14924 9658 14976 9664
rect 14936 9110 14964 9658
rect 14832 9104 14884 9110
rect 14832 9046 14884 9052
rect 14924 9104 14976 9110
rect 14924 9046 14976 9052
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 13728 8492 13780 8498
rect 13648 8452 13728 8480
rect 13544 8016 13596 8022
rect 13450 7984 13506 7993
rect 13544 7958 13596 7964
rect 13450 7919 13506 7928
rect 13174 7848 13230 7857
rect 12348 7812 12400 7818
rect 13174 7783 13176 7792
rect 12348 7754 12400 7760
rect 13228 7783 13230 7792
rect 13176 7754 13228 7760
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10692 4150 10744 4156
rect 10874 4176 10930 4185
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 10612 3534 10640 4082
rect 10704 3942 10732 4150
rect 10874 4111 10930 4120
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10980 3738 11008 7142
rect 12360 7002 12388 7754
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 12668 7100 12976 7109
rect 12668 7098 12674 7100
rect 12730 7098 12754 7100
rect 12810 7098 12834 7100
rect 12890 7098 12914 7100
rect 12970 7098 12976 7100
rect 12730 7046 12732 7098
rect 12912 7046 12914 7098
rect 12668 7044 12674 7046
rect 12730 7044 12754 7046
rect 12810 7044 12834 7046
rect 12890 7044 12914 7046
rect 12970 7044 12976 7046
rect 12668 7035 12976 7044
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12636 6186 12664 6734
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12668 6012 12976 6021
rect 12668 6010 12674 6012
rect 12730 6010 12754 6012
rect 12810 6010 12834 6012
rect 12890 6010 12914 6012
rect 12970 6010 12976 6012
rect 12730 5958 12732 6010
rect 12912 5958 12914 6010
rect 12668 5956 12674 5958
rect 12730 5956 12754 5958
rect 12810 5956 12834 5958
rect 12890 5956 12914 5958
rect 12970 5956 12976 5958
rect 12668 5947 12976 5956
rect 13004 5302 13032 7414
rect 13648 6662 13676 8452
rect 13728 8434 13780 8440
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13740 7478 13768 7754
rect 13728 7472 13780 7478
rect 13728 7414 13780 7420
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13740 7002 13768 7278
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13084 5636 13136 5642
rect 13084 5578 13136 5584
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 12668 4924 12976 4933
rect 12668 4922 12674 4924
rect 12730 4922 12754 4924
rect 12810 4922 12834 4924
rect 12890 4922 12914 4924
rect 12970 4922 12976 4924
rect 12730 4870 12732 4922
rect 12912 4870 12914 4922
rect 12668 4868 12674 4870
rect 12730 4868 12754 4870
rect 12810 4868 12834 4870
rect 12890 4868 12914 4870
rect 12970 4868 12976 4870
rect 12668 4859 12976 4868
rect 13096 4078 13124 5578
rect 13740 5166 13768 6938
rect 14844 6322 14872 9046
rect 15028 8634 15056 10950
rect 15212 10810 15240 11086
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15106 10296 15162 10305
rect 15106 10231 15162 10240
rect 15120 10130 15148 10231
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15120 9042 15148 10066
rect 15396 9926 15424 10746
rect 15476 10736 15528 10742
rect 15580 10724 15608 11086
rect 15528 10696 15608 10724
rect 15476 10678 15528 10684
rect 15948 10606 15976 11154
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16500 10674 16528 11018
rect 16776 10742 16804 13262
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16868 12918 16896 13126
rect 16856 12912 16908 12918
rect 16856 12854 16908 12860
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16868 12170 16896 12582
rect 16960 12306 16988 13942
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17420 13326 17448 13670
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17512 13258 17540 13670
rect 19352 13410 19380 15438
rect 19628 15094 19656 15506
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 19616 15088 19668 15094
rect 19616 15030 19668 15036
rect 20088 14006 20116 15302
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20076 14000 20128 14006
rect 20076 13942 20128 13948
rect 19628 13802 20116 13818
rect 19628 13796 20128 13802
rect 19628 13790 20076 13796
rect 19628 13734 19656 13790
rect 20076 13738 20128 13744
rect 19616 13728 19668 13734
rect 19616 13670 19668 13676
rect 19708 13728 19760 13734
rect 20456 13705 20484 14010
rect 19708 13670 19760 13676
rect 20442 13696 20498 13705
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 19260 13382 19380 13410
rect 19260 13326 19288 13382
rect 19444 13326 19472 13466
rect 19248 13320 19300 13326
rect 19248 13262 19300 13268
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19720 13258 19748 13670
rect 20442 13631 20498 13640
rect 17500 13252 17552 13258
rect 17500 13194 17552 13200
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19708 13252 19760 13258
rect 19708 13194 19760 13200
rect 17960 13184 18012 13190
rect 17960 13126 18012 13132
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 17512 11762 17540 12582
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17144 11150 17172 11698
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 16764 10736 16816 10742
rect 16764 10678 16816 10684
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 15028 6798 15056 8570
rect 15108 8356 15160 8362
rect 15108 8298 15160 8304
rect 15120 8022 15148 8298
rect 15108 8016 15160 8022
rect 15108 7958 15160 7964
rect 15304 6798 15332 8774
rect 15856 8566 15884 8774
rect 15844 8560 15896 8566
rect 15844 8502 15896 8508
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15028 6458 15056 6734
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 14556 5636 14608 5642
rect 14556 5578 14608 5584
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 14476 4622 14504 5170
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14568 4078 14596 5578
rect 14844 4146 14872 6258
rect 15948 5166 15976 10542
rect 16132 9654 16160 10542
rect 16776 10538 16804 10678
rect 16764 10532 16816 10538
rect 16764 10474 16816 10480
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16120 9648 16172 9654
rect 16120 9590 16172 9596
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16040 9178 16068 9522
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 16040 8566 16068 9114
rect 16132 8974 16160 9454
rect 16224 9178 16252 9522
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 16316 8294 16344 9522
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16316 7478 16344 8230
rect 16304 7472 16356 7478
rect 16304 7414 16356 7420
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15396 4282 15424 4422
rect 15384 4276 15436 4282
rect 15384 4218 15436 4224
rect 15488 4214 15516 5102
rect 16408 4593 16436 9862
rect 17880 9722 17908 11018
rect 17972 10606 18000 13126
rect 19156 12708 19208 12714
rect 19156 12650 19208 12656
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18616 12306 18644 12582
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 18236 12164 18288 12170
rect 18236 12106 18288 12112
rect 18052 11824 18104 11830
rect 18052 11766 18104 11772
rect 18064 11694 18092 11766
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 18248 10810 18276 12106
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18432 11830 18460 12038
rect 18420 11824 18472 11830
rect 18420 11766 18472 11772
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 18340 10690 18368 11086
rect 18156 10674 18368 10690
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 18156 10668 18380 10674
rect 18156 10662 18328 10668
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 18064 10198 18092 10610
rect 18156 10470 18184 10662
rect 18328 10610 18380 10616
rect 18432 10554 18460 11086
rect 19064 11008 19116 11014
rect 19064 10950 19116 10956
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18248 10526 18460 10554
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 18052 10192 18104 10198
rect 18052 10134 18104 10140
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16960 9178 16988 9454
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 16534 9036 16586 9042
rect 16672 9036 16724 9042
rect 16586 8996 16672 9024
rect 16534 8978 16586 8984
rect 16672 8978 16724 8984
rect 16776 8974 16804 9046
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16672 8900 16724 8906
rect 16672 8842 16724 8848
rect 16684 8401 16712 8842
rect 16868 8634 16896 8910
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16670 8392 16726 8401
rect 16670 8327 16726 8336
rect 16960 7750 16988 8978
rect 17052 8634 17080 9590
rect 17972 9586 18000 10066
rect 18064 9994 18092 10134
rect 18052 9988 18104 9994
rect 18052 9930 18104 9936
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17130 8664 17186 8673
rect 17040 8628 17092 8634
rect 17130 8599 17186 8608
rect 17040 8570 17092 8576
rect 17144 8566 17172 8599
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17236 8362 17264 9114
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 17328 8090 17356 8910
rect 17406 8528 17462 8537
rect 17604 8498 17632 8978
rect 17682 8800 17738 8809
rect 17682 8735 17738 8744
rect 17696 8498 17724 8735
rect 17406 8463 17462 8472
rect 17500 8492 17552 8498
rect 17420 8430 17448 8463
rect 17500 8434 17552 8440
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17684 8492 17736 8498
rect 17788 8480 17816 9114
rect 18052 9104 18104 9110
rect 18052 9046 18104 9052
rect 18064 8974 18092 9046
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17788 8452 17908 8480
rect 17684 8434 17736 8440
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17512 8090 17540 8434
rect 17880 8412 17908 8452
rect 17960 8424 18012 8430
rect 17590 8392 17646 8401
rect 17880 8384 17960 8412
rect 17960 8366 18012 8372
rect 17590 8327 17592 8336
rect 17644 8327 17646 8336
rect 17592 8298 17644 8304
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16960 6934 16988 7686
rect 17328 7478 17356 8026
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17316 7472 17368 7478
rect 17316 7414 17368 7420
rect 16948 6928 17000 6934
rect 16948 6870 17000 6876
rect 17328 6798 17356 7414
rect 17972 6934 18000 7890
rect 18156 7886 18184 10406
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18248 7410 18276 10526
rect 18616 10146 18644 10542
rect 18800 10282 18828 10746
rect 19076 10674 19104 10950
rect 19064 10668 19116 10674
rect 19064 10610 19116 10616
rect 18708 10266 18828 10282
rect 18696 10260 18828 10266
rect 18748 10254 18828 10260
rect 18696 10202 18748 10208
rect 19064 10192 19116 10198
rect 18616 10118 18736 10146
rect 19064 10134 19116 10140
rect 18328 9920 18380 9926
rect 18604 9920 18656 9926
rect 18328 9862 18380 9868
rect 18432 9880 18604 9908
rect 18340 9450 18368 9862
rect 18432 9722 18460 9880
rect 18604 9862 18656 9868
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18328 9444 18380 9450
rect 18328 9386 18380 9392
rect 18432 9178 18460 9658
rect 18420 9172 18472 9178
rect 18420 9114 18472 9120
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18328 8900 18380 8906
rect 18328 8842 18380 8848
rect 18340 8809 18368 8842
rect 18420 8832 18472 8838
rect 18326 8800 18382 8809
rect 18524 8820 18552 9114
rect 18708 9081 18736 10118
rect 19076 9926 19104 10134
rect 19168 10130 19196 12650
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19260 11762 19288 12310
rect 19352 12306 19380 13194
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 19616 12640 19668 12646
rect 19616 12582 19668 12588
rect 19628 12434 19656 12582
rect 20456 12442 20484 12786
rect 20444 12436 20496 12442
rect 19628 12406 19748 12434
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19338 11520 19394 11529
rect 19338 11455 19394 11464
rect 19352 11286 19380 11455
rect 19340 11280 19392 11286
rect 19340 11222 19392 11228
rect 19432 11280 19484 11286
rect 19484 11240 19564 11268
rect 19432 11222 19484 11228
rect 19340 11144 19392 11150
rect 19338 11112 19340 11121
rect 19536 11132 19564 11240
rect 19616 11144 19668 11150
rect 19392 11112 19394 11121
rect 19536 11104 19616 11132
rect 19616 11086 19668 11092
rect 19338 11047 19394 11056
rect 19294 11008 19346 11014
rect 19432 11008 19484 11014
rect 19346 10976 19394 10985
rect 19294 10950 19338 10956
rect 19306 10934 19338 10950
rect 19432 10950 19484 10956
rect 19338 10911 19394 10920
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 19076 9518 19104 9862
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 18694 9072 18750 9081
rect 19168 9042 19196 10066
rect 19260 9654 19288 10406
rect 19444 9674 19472 10950
rect 19720 10674 19748 12406
rect 20444 12378 20496 12384
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 19890 11384 19946 11393
rect 19890 11319 19946 11328
rect 19800 11008 19852 11014
rect 19798 10976 19800 10985
rect 19852 10976 19854 10985
rect 19798 10911 19854 10920
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 19720 10062 19748 10610
rect 19904 10606 19932 11319
rect 19996 11150 20024 11494
rect 20180 11354 20208 11494
rect 20548 11354 20576 17138
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20640 16114 20668 16526
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20640 15502 20668 16050
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 20732 15094 20760 15846
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20824 14414 20852 15302
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 20640 13546 20668 14214
rect 20640 13518 20760 13546
rect 20732 13462 20760 13518
rect 20720 13456 20772 13462
rect 20720 13398 20772 13404
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20812 11212 20864 11218
rect 20812 11154 20864 11160
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19996 10606 20024 11086
rect 19892 10600 19944 10606
rect 19892 10542 19944 10548
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19996 10130 20024 10542
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19708 10056 19760 10062
rect 20732 10033 20760 10202
rect 19708 9998 19760 10004
rect 20718 10024 20774 10033
rect 20718 9959 20774 9968
rect 19706 9752 19762 9761
rect 19706 9687 19762 9696
rect 20720 9716 20772 9722
rect 19248 9648 19300 9654
rect 19248 9590 19300 9596
rect 19352 9646 19472 9674
rect 18694 9007 18750 9016
rect 19156 9036 19208 9042
rect 19156 8978 19208 8984
rect 18696 8900 18748 8906
rect 18696 8842 18748 8848
rect 18472 8792 18552 8820
rect 18420 8774 18472 8780
rect 18326 8735 18382 8744
rect 18708 8498 18736 8842
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18340 7546 18368 8366
rect 19260 8294 19288 9590
rect 19352 9518 19380 9646
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19720 9178 19748 9687
rect 20720 9658 20772 9664
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 19708 9172 19760 9178
rect 19708 9114 19760 9120
rect 19892 9172 19944 9178
rect 19892 9114 19944 9120
rect 19904 9081 19932 9114
rect 19890 9072 19946 9081
rect 19536 9030 19840 9058
rect 19536 8906 19564 9030
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19524 8900 19576 8906
rect 19524 8842 19576 8848
rect 19628 8498 19656 8910
rect 19720 8838 19748 8910
rect 19812 8906 19840 9030
rect 19890 9007 19946 9016
rect 19800 8900 19852 8906
rect 19800 8842 19852 8848
rect 19708 8832 19760 8838
rect 19708 8774 19760 8780
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19904 8294 19932 9007
rect 20088 8401 20116 9522
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20272 8566 20300 8774
rect 20442 8664 20498 8673
rect 20548 8634 20576 8978
rect 20732 8974 20760 9658
rect 20824 9518 20852 11154
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20628 8968 20680 8974
rect 20626 8936 20628 8945
rect 20720 8968 20772 8974
rect 20680 8936 20682 8945
rect 20720 8910 20772 8916
rect 20626 8871 20682 8880
rect 20442 8599 20498 8608
rect 20536 8628 20588 8634
rect 20260 8560 20312 8566
rect 20260 8502 20312 8508
rect 20456 8498 20484 8599
rect 20536 8570 20588 8576
rect 20732 8537 20760 8910
rect 20718 8528 20774 8537
rect 20444 8492 20496 8498
rect 20718 8463 20774 8472
rect 20444 8434 20496 8440
rect 20074 8392 20130 8401
rect 20074 8327 20130 8336
rect 19260 8266 19380 8294
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18616 7410 18644 7686
rect 18708 7546 18736 7822
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18892 7478 18920 8026
rect 18880 7472 18932 7478
rect 18880 7414 18932 7420
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18248 6934 18276 7346
rect 19352 7206 19380 8266
rect 19892 8288 19944 8294
rect 19892 8230 19944 8236
rect 20088 7478 20116 8327
rect 20732 7954 20760 8463
rect 20916 7954 20944 17478
rect 24386 17436 24694 17445
rect 24386 17434 24392 17436
rect 24448 17434 24472 17436
rect 24528 17434 24552 17436
rect 24608 17434 24632 17436
rect 24688 17434 24694 17436
rect 24448 17382 24450 17434
rect 24630 17382 24632 17434
rect 24386 17380 24392 17382
rect 24448 17380 24472 17382
rect 24528 17380 24552 17382
rect 24608 17380 24632 17382
rect 24688 17380 24694 17382
rect 24386 17371 24694 17380
rect 28184 17338 28212 19200
rect 36096 17898 36124 19200
rect 36004 17870 36124 17898
rect 28172 17332 28224 17338
rect 28172 17274 28224 17280
rect 34336 17264 34388 17270
rect 34336 17206 34388 17212
rect 28448 17196 28500 17202
rect 28448 17138 28500 17144
rect 24308 16720 24360 16726
rect 24308 16662 24360 16668
rect 22100 15972 22152 15978
rect 22100 15914 22152 15920
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21100 13190 21128 13466
rect 21284 13394 21312 13874
rect 22112 13682 22140 15914
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22376 14816 22428 14822
rect 22376 14758 22428 14764
rect 22192 13864 22244 13870
rect 22192 13806 22244 13812
rect 21928 13654 22140 13682
rect 21928 13530 21956 13654
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 22008 13524 22060 13530
rect 22008 13466 22060 13472
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 21272 13388 21324 13394
rect 21272 13330 21324 13336
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 21284 12850 21312 13330
rect 21456 13252 21508 13258
rect 21456 13194 21508 13200
rect 21468 12986 21496 13194
rect 21456 12980 21508 12986
rect 21456 12922 21508 12928
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 20996 11008 21048 11014
rect 20996 10950 21048 10956
rect 21008 10742 21036 10950
rect 21284 10742 21312 12786
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21652 11694 21680 12174
rect 22020 11778 22048 13466
rect 22112 13394 22140 13466
rect 22100 13388 22152 13394
rect 22100 13330 22152 13336
rect 22204 13326 22232 13806
rect 22192 13320 22244 13326
rect 22098 13288 22154 13297
rect 22192 13262 22244 13268
rect 22098 13223 22154 13232
rect 22112 12442 22140 13223
rect 22388 12918 22416 14758
rect 22572 13870 22600 15098
rect 22664 14074 22692 15438
rect 22744 15360 22796 15366
rect 22744 15302 22796 15308
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 22756 14346 22784 15302
rect 23676 14958 23704 15302
rect 23664 14952 23716 14958
rect 23664 14894 23716 14900
rect 23756 14544 23808 14550
rect 23676 14492 23756 14498
rect 23676 14486 23808 14492
rect 23676 14470 23796 14486
rect 22744 14340 22796 14346
rect 22744 14282 22796 14288
rect 22652 14068 22704 14074
rect 22652 14010 22704 14016
rect 23676 14006 23704 14470
rect 24214 14104 24270 14113
rect 24214 14039 24270 14048
rect 23664 14000 23716 14006
rect 23664 13942 23716 13948
rect 22560 13864 22612 13870
rect 22560 13806 22612 13812
rect 24228 13818 24256 14039
rect 24320 14006 24348 16662
rect 24386 16348 24694 16357
rect 24386 16346 24392 16348
rect 24448 16346 24472 16348
rect 24528 16346 24552 16348
rect 24608 16346 24632 16348
rect 24688 16346 24694 16348
rect 24448 16294 24450 16346
rect 24630 16294 24632 16346
rect 24386 16292 24392 16294
rect 24448 16292 24472 16294
rect 24528 16292 24552 16294
rect 24608 16292 24632 16294
rect 24688 16292 24694 16294
rect 24386 16283 24694 16292
rect 27712 15904 27764 15910
rect 27712 15846 27764 15852
rect 27620 15496 27672 15502
rect 27620 15438 27672 15444
rect 24768 15360 24820 15366
rect 24768 15302 24820 15308
rect 24386 15260 24694 15269
rect 24386 15258 24392 15260
rect 24448 15258 24472 15260
rect 24528 15258 24552 15260
rect 24608 15258 24632 15260
rect 24688 15258 24694 15260
rect 24448 15206 24450 15258
rect 24630 15206 24632 15258
rect 24386 15204 24392 15206
rect 24448 15204 24472 15206
rect 24528 15204 24552 15206
rect 24608 15204 24632 15206
rect 24688 15204 24694 15206
rect 24386 15195 24694 15204
rect 24780 15094 24808 15302
rect 24768 15088 24820 15094
rect 24768 15030 24820 15036
rect 24860 15088 24912 15094
rect 24860 15030 24912 15036
rect 24584 15020 24636 15026
rect 24584 14962 24636 14968
rect 24400 14884 24452 14890
rect 24400 14826 24452 14832
rect 24412 14618 24440 14826
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24400 14612 24452 14618
rect 24400 14554 24452 14560
rect 24504 14414 24532 14758
rect 24596 14618 24624 14962
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 24780 14414 24808 15030
rect 24492 14408 24544 14414
rect 24492 14350 24544 14356
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 24872 14346 24900 15030
rect 25872 14952 25924 14958
rect 25872 14894 25924 14900
rect 25594 14784 25650 14793
rect 25594 14719 25650 14728
rect 25044 14612 25096 14618
rect 25044 14554 25096 14560
rect 24860 14340 24912 14346
rect 24860 14282 24912 14288
rect 24386 14172 24694 14181
rect 24386 14170 24392 14172
rect 24448 14170 24472 14172
rect 24528 14170 24552 14172
rect 24608 14170 24632 14172
rect 24688 14170 24694 14172
rect 24448 14118 24450 14170
rect 24630 14118 24632 14170
rect 24386 14116 24392 14118
rect 24448 14116 24472 14118
rect 24528 14116 24552 14118
rect 24608 14116 24632 14118
rect 24688 14116 24694 14118
rect 24386 14107 24694 14116
rect 24766 14104 24822 14113
rect 24766 14039 24822 14048
rect 24308 14000 24360 14006
rect 24780 13954 24808 14039
rect 24308 13942 24360 13948
rect 24412 13926 24808 13954
rect 25056 13938 25084 14554
rect 25608 14414 25636 14719
rect 25596 14408 25648 14414
rect 25596 14350 25648 14356
rect 25596 14272 25648 14278
rect 25596 14214 25648 14220
rect 25608 14006 25636 14214
rect 25884 14090 25912 14894
rect 26792 14816 26844 14822
rect 26792 14758 26844 14764
rect 26884 14816 26936 14822
rect 26884 14758 26936 14764
rect 26240 14272 26292 14278
rect 26240 14214 26292 14220
rect 25700 14074 25912 14090
rect 25688 14068 25912 14074
rect 25740 14062 25912 14068
rect 25688 14010 25740 14016
rect 25596 14000 25648 14006
rect 25596 13942 25648 13948
rect 25044 13932 25096 13938
rect 24412 13818 24440 13926
rect 25044 13874 25096 13880
rect 24228 13790 24440 13818
rect 25320 13796 25372 13802
rect 25320 13738 25372 13744
rect 25332 13530 25360 13738
rect 25320 13524 25372 13530
rect 25320 13466 25372 13472
rect 25884 13410 25912 14062
rect 26148 14068 26200 14074
rect 26148 14010 26200 14016
rect 26160 13954 26188 14010
rect 25976 13926 26188 13954
rect 25976 13870 26004 13926
rect 25964 13864 26016 13870
rect 25964 13806 26016 13812
rect 25884 13382 26004 13410
rect 25976 13326 26004 13382
rect 25964 13320 26016 13326
rect 25964 13262 26016 13268
rect 23204 13252 23256 13258
rect 23204 13194 23256 13200
rect 23216 12918 23244 13194
rect 24386 13084 24694 13093
rect 24386 13082 24392 13084
rect 24448 13082 24472 13084
rect 24528 13082 24552 13084
rect 24608 13082 24632 13084
rect 24688 13082 24694 13084
rect 24448 13030 24450 13082
rect 24630 13030 24632 13082
rect 24386 13028 24392 13030
rect 24448 13028 24472 13030
rect 24528 13028 24552 13030
rect 24608 13028 24632 13030
rect 24688 13028 24694 13030
rect 24386 13019 24694 13028
rect 26148 12980 26200 12986
rect 26148 12922 26200 12928
rect 22376 12912 22428 12918
rect 22376 12854 22428 12860
rect 23204 12912 23256 12918
rect 23204 12854 23256 12860
rect 25136 12912 25188 12918
rect 25320 12912 25372 12918
rect 25188 12872 25320 12900
rect 25136 12854 25188 12860
rect 25320 12854 25372 12860
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 22204 12442 22232 12718
rect 22284 12640 22336 12646
rect 22284 12582 22336 12588
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22192 12436 22244 12442
rect 22192 12378 22244 12384
rect 22296 12306 22324 12582
rect 22744 12436 22796 12442
rect 22744 12378 22796 12384
rect 22756 12322 22784 12378
rect 22284 12300 22336 12306
rect 22756 12294 22876 12322
rect 22284 12242 22336 12248
rect 22744 12096 22796 12102
rect 22744 12038 22796 12044
rect 22560 11824 22612 11830
rect 21928 11762 22048 11778
rect 21916 11756 22048 11762
rect 21968 11750 22048 11756
rect 22558 11792 22560 11801
rect 22612 11792 22614 11801
rect 22558 11727 22614 11736
rect 21916 11698 21968 11704
rect 21640 11688 21692 11694
rect 21640 11630 21692 11636
rect 22756 11150 22784 12038
rect 22848 11830 22876 12294
rect 23216 12102 23244 12854
rect 26160 12434 26188 12922
rect 26252 12850 26280 14214
rect 26804 13462 26832 14758
rect 26896 14482 26924 14758
rect 27160 14544 27212 14550
rect 27212 14492 27384 14498
rect 27160 14486 27384 14492
rect 26884 14476 26936 14482
rect 27172 14470 27384 14486
rect 26884 14418 26936 14424
rect 27160 14408 27212 14414
rect 27160 14350 27212 14356
rect 26792 13456 26844 13462
rect 26792 13398 26844 13404
rect 26332 13252 26384 13258
rect 26332 13194 26384 13200
rect 26240 12844 26292 12850
rect 26240 12786 26292 12792
rect 26068 12406 26188 12434
rect 24032 12368 24084 12374
rect 24030 12336 24032 12345
rect 24084 12336 24086 12345
rect 24030 12271 24086 12280
rect 23204 12096 23256 12102
rect 23204 12038 23256 12044
rect 25412 12096 25464 12102
rect 25412 12038 25464 12044
rect 25872 12096 25924 12102
rect 25872 12038 25924 12044
rect 24386 11996 24694 12005
rect 24386 11994 24392 11996
rect 24448 11994 24472 11996
rect 24528 11994 24552 11996
rect 24608 11994 24632 11996
rect 24688 11994 24694 11996
rect 24448 11942 24450 11994
rect 24630 11942 24632 11994
rect 24386 11940 24392 11942
rect 24448 11940 24472 11942
rect 24528 11940 24552 11942
rect 24608 11940 24632 11942
rect 24688 11940 24694 11942
rect 24386 11931 24694 11940
rect 25424 11937 25452 12038
rect 25410 11928 25466 11937
rect 25410 11863 25466 11872
rect 22836 11824 22888 11830
rect 22836 11766 22888 11772
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 22756 10742 22784 11086
rect 20996 10736 21048 10742
rect 20996 10678 21048 10684
rect 21272 10736 21324 10742
rect 21272 10678 21324 10684
rect 22744 10736 22796 10742
rect 22744 10678 22796 10684
rect 22558 10432 22614 10441
rect 22558 10367 22614 10376
rect 22572 10266 22600 10367
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22006 10160 22062 10169
rect 22006 10095 22008 10104
rect 22060 10095 22062 10104
rect 22008 10066 22060 10072
rect 22572 10062 22600 10202
rect 22560 10056 22612 10062
rect 22560 9998 22612 10004
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22468 9988 22520 9994
rect 22468 9930 22520 9936
rect 20996 9648 21048 9654
rect 20996 9590 21048 9596
rect 21180 9648 21232 9654
rect 21180 9590 21232 9596
rect 21008 9518 21036 9590
rect 20996 9512 21048 9518
rect 20996 9454 21048 9460
rect 21192 9178 21220 9590
rect 21824 9512 21876 9518
rect 21824 9454 21876 9460
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 21836 9178 21864 9454
rect 21916 9376 21968 9382
rect 21914 9344 21916 9353
rect 21968 9344 21970 9353
rect 21914 9279 21970 9288
rect 22112 9178 22140 9454
rect 22190 9344 22246 9353
rect 22190 9279 22246 9288
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21824 9172 21876 9178
rect 21824 9114 21876 9120
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 21638 8800 21694 8809
rect 21638 8735 21694 8744
rect 21456 8560 21508 8566
rect 21454 8528 21456 8537
rect 21508 8528 21510 8537
rect 21454 8463 21510 8472
rect 21652 8090 21680 8735
rect 21836 8430 21864 9114
rect 22204 9042 22232 9279
rect 22100 9036 22152 9042
rect 22100 8978 22152 8984
rect 22192 9036 22244 9042
rect 22192 8978 22244 8984
rect 22112 8922 22140 8978
rect 22376 8968 22428 8974
rect 21916 8900 21968 8906
rect 22112 8894 22232 8922
rect 22376 8910 22428 8916
rect 21916 8842 21968 8848
rect 21824 8424 21876 8430
rect 21928 8401 21956 8842
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 21824 8366 21876 8372
rect 21914 8392 21970 8401
rect 21836 8090 21864 8366
rect 21914 8327 21970 8336
rect 21640 8084 21692 8090
rect 21640 8026 21692 8032
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 20076 7472 20128 7478
rect 20076 7414 20128 7420
rect 20272 7410 20300 7822
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 20916 7002 20944 7890
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 20996 7472 21048 7478
rect 20994 7440 20996 7449
rect 21048 7440 21050 7449
rect 21284 7410 21312 7822
rect 21836 7546 21864 8026
rect 21928 7954 21956 8026
rect 21916 7948 21968 7954
rect 21916 7890 21968 7896
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 20994 7375 21050 7384
rect 21272 7404 21324 7410
rect 21272 7346 21324 7352
rect 20904 6996 20956 7002
rect 20904 6938 20956 6944
rect 17960 6928 18012 6934
rect 17960 6870 18012 6876
rect 18236 6928 18288 6934
rect 18236 6870 18288 6876
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17972 6730 18000 6870
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 17972 6458 18000 6666
rect 18248 6662 18276 6870
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 18236 6656 18288 6662
rect 18236 6598 18288 6604
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 17972 6254 18000 6394
rect 19248 6384 19300 6390
rect 19248 6326 19300 6332
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 19260 6186 19288 6326
rect 19248 6180 19300 6186
rect 19248 6122 19300 6128
rect 18512 6112 18564 6118
rect 18512 6054 18564 6060
rect 18524 5778 18552 6054
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 19444 5642 19472 6394
rect 20456 6322 20484 6802
rect 20548 6458 20576 6802
rect 22112 6730 22140 8434
rect 22204 7818 22232 8894
rect 22388 8566 22416 8910
rect 22376 8560 22428 8566
rect 22376 8502 22428 8508
rect 22192 7812 22244 7818
rect 22192 7754 22244 7760
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22296 7002 22324 7414
rect 22480 7342 22508 9930
rect 22664 9722 22692 9998
rect 22848 9994 22876 11766
rect 25044 11688 25096 11694
rect 25044 11630 25096 11636
rect 22926 11112 22982 11121
rect 22926 11047 22928 11056
rect 22980 11047 22982 11056
rect 24306 11112 24362 11121
rect 24306 11047 24362 11056
rect 22928 11018 22980 11024
rect 23940 11008 23992 11014
rect 23940 10950 23992 10956
rect 23952 10577 23980 10950
rect 24320 10810 24348 11047
rect 24768 11008 24820 11014
rect 24768 10950 24820 10956
rect 24386 10908 24694 10917
rect 24386 10906 24392 10908
rect 24448 10906 24472 10908
rect 24528 10906 24552 10908
rect 24608 10906 24632 10908
rect 24688 10906 24694 10908
rect 24448 10854 24450 10906
rect 24630 10854 24632 10906
rect 24386 10852 24392 10854
rect 24448 10852 24472 10854
rect 24528 10852 24552 10854
rect 24608 10852 24632 10854
rect 24688 10852 24694 10854
rect 24386 10843 24694 10852
rect 24308 10804 24360 10810
rect 24308 10746 24360 10752
rect 24492 10804 24544 10810
rect 24492 10746 24544 10752
rect 23938 10568 23994 10577
rect 24504 10538 24532 10746
rect 24780 10554 24808 10950
rect 24952 10736 25004 10742
rect 24952 10678 25004 10684
rect 24964 10606 24992 10678
rect 24860 10600 24912 10606
rect 24780 10548 24860 10554
rect 24780 10542 24912 10548
rect 24952 10600 25004 10606
rect 24952 10542 25004 10548
rect 23938 10503 23994 10512
rect 24492 10532 24544 10538
rect 24780 10526 24900 10542
rect 24492 10474 24544 10480
rect 23756 10464 23808 10470
rect 23756 10406 23808 10412
rect 23768 10266 23796 10406
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 24596 10084 24900 10112
rect 22836 9988 22888 9994
rect 22836 9930 22888 9936
rect 24596 9926 24624 10084
rect 24688 9994 24808 10010
rect 24676 9988 24808 9994
rect 24728 9982 24808 9988
rect 24676 9930 24728 9936
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 24584 9920 24636 9926
rect 24584 9862 24636 9868
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 23400 9654 23428 9862
rect 24386 9820 24694 9829
rect 24386 9818 24392 9820
rect 24448 9818 24472 9820
rect 24528 9818 24552 9820
rect 24608 9818 24632 9820
rect 24688 9818 24694 9820
rect 24448 9766 24450 9818
rect 24630 9766 24632 9818
rect 24386 9764 24392 9766
rect 24448 9764 24472 9766
rect 24528 9764 24552 9766
rect 24608 9764 24632 9766
rect 24688 9764 24694 9766
rect 23570 9752 23626 9761
rect 24386 9755 24694 9764
rect 23570 9687 23626 9696
rect 23388 9648 23440 9654
rect 23386 9616 23388 9625
rect 23440 9616 23442 9625
rect 23386 9551 23442 9560
rect 23584 9489 23612 9687
rect 23386 9480 23442 9489
rect 22928 9444 22980 9450
rect 23386 9415 23442 9424
rect 23570 9480 23626 9489
rect 23570 9415 23626 9424
rect 22928 9386 22980 9392
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22560 8968 22612 8974
rect 22664 8945 22692 9318
rect 22560 8910 22612 8916
rect 22650 8936 22706 8945
rect 22572 8809 22600 8910
rect 22650 8871 22706 8880
rect 22664 8838 22692 8871
rect 22652 8832 22704 8838
rect 22558 8800 22614 8809
rect 22652 8774 22704 8780
rect 22558 8735 22614 8744
rect 22572 8498 22600 8735
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 22940 8430 22968 9386
rect 23400 9382 23428 9415
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 23202 9208 23258 9217
rect 23202 9143 23258 9152
rect 22928 8424 22980 8430
rect 22928 8366 22980 8372
rect 22928 7744 22980 7750
rect 22928 7686 22980 7692
rect 22468 7336 22520 7342
rect 22468 7278 22520 7284
rect 22480 7206 22508 7278
rect 22468 7200 22520 7206
rect 22468 7142 22520 7148
rect 22284 6996 22336 7002
rect 22284 6938 22336 6944
rect 22192 6928 22244 6934
rect 22192 6870 22244 6876
rect 22100 6724 22152 6730
rect 22100 6666 22152 6672
rect 22204 6458 22232 6870
rect 22744 6724 22796 6730
rect 22744 6666 22796 6672
rect 22756 6458 22784 6666
rect 22940 6662 22968 7686
rect 23112 7336 23164 7342
rect 23110 7304 23112 7313
rect 23164 7304 23166 7313
rect 23110 7239 23166 7248
rect 23020 6792 23072 6798
rect 23020 6734 23072 6740
rect 22928 6656 22980 6662
rect 22928 6598 22980 6604
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 22192 6452 22244 6458
rect 22192 6394 22244 6400
rect 22744 6452 22796 6458
rect 22744 6394 22796 6400
rect 20904 6384 20956 6390
rect 22652 6384 22704 6390
rect 20956 6332 21220 6338
rect 20904 6326 21220 6332
rect 22652 6326 22704 6332
rect 20916 6322 21220 6326
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 20444 6316 20496 6322
rect 20916 6316 21232 6322
rect 20916 6310 21180 6316
rect 20444 6258 20496 6264
rect 21180 6258 21232 6264
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19628 5710 19656 6054
rect 19720 5778 19748 6258
rect 19890 5944 19946 5953
rect 19890 5879 19892 5888
rect 19944 5879 19946 5888
rect 19892 5850 19944 5856
rect 22664 5794 22692 6326
rect 22756 6186 22784 6394
rect 22744 6180 22796 6186
rect 22744 6122 22796 6128
rect 22836 6112 22888 6118
rect 22836 6054 22888 6060
rect 22848 5914 22876 6054
rect 22836 5908 22888 5914
rect 22836 5850 22888 5856
rect 22940 5817 22968 6598
rect 23032 6254 23060 6734
rect 23216 6322 23244 9143
rect 24386 8732 24694 8741
rect 24386 8730 24392 8732
rect 24448 8730 24472 8732
rect 24528 8730 24552 8732
rect 24608 8730 24632 8732
rect 24688 8730 24694 8732
rect 24448 8678 24450 8730
rect 24630 8678 24632 8730
rect 24386 8676 24392 8678
rect 24448 8676 24472 8678
rect 24528 8676 24552 8678
rect 24608 8676 24632 8678
rect 24688 8676 24694 8678
rect 24386 8667 24694 8676
rect 23754 8528 23810 8537
rect 23754 8463 23756 8472
rect 23808 8463 23810 8472
rect 23756 8434 23808 8440
rect 23296 8424 23348 8430
rect 23296 8366 23348 8372
rect 23308 7750 23336 8366
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 24386 7644 24694 7653
rect 24386 7642 24392 7644
rect 24448 7642 24472 7644
rect 24528 7642 24552 7644
rect 24608 7642 24632 7644
rect 24688 7642 24694 7644
rect 24448 7590 24450 7642
rect 24630 7590 24632 7642
rect 24386 7588 24392 7590
rect 24448 7588 24472 7590
rect 24528 7588 24552 7590
rect 24608 7588 24632 7590
rect 24688 7588 24694 7590
rect 24386 7579 24694 7588
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 23388 7336 23440 7342
rect 23388 7278 23440 7284
rect 23400 7206 23428 7278
rect 23676 7206 23704 7346
rect 23388 7200 23440 7206
rect 23664 7200 23716 7206
rect 23388 7142 23440 7148
rect 23662 7168 23664 7177
rect 24216 7200 24268 7206
rect 23716 7168 23718 7177
rect 24216 7142 24268 7148
rect 23662 7103 23718 7112
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 23204 6316 23256 6322
rect 23204 6258 23256 6264
rect 23020 6248 23072 6254
rect 23020 6190 23072 6196
rect 22926 5808 22982 5817
rect 19708 5772 19760 5778
rect 19708 5714 19760 5720
rect 22480 5766 22876 5794
rect 19616 5704 19668 5710
rect 22480 5658 22508 5766
rect 22848 5710 22876 5766
rect 22926 5743 22982 5752
rect 22652 5704 22704 5710
rect 19616 5646 19668 5652
rect 22388 5642 22508 5658
rect 19432 5636 19484 5642
rect 19432 5578 19484 5584
rect 22100 5636 22152 5642
rect 22100 5578 22152 5584
rect 22376 5636 22508 5642
rect 22428 5630 22508 5636
rect 22650 5672 22652 5681
rect 22836 5704 22888 5710
rect 22704 5672 22706 5681
rect 22836 5646 22888 5652
rect 22650 5607 22706 5616
rect 22376 5578 22428 5584
rect 22008 5568 22060 5574
rect 22008 5510 22060 5516
rect 22020 5302 22048 5510
rect 22008 5296 22060 5302
rect 22008 5238 22060 5244
rect 22112 5234 22140 5578
rect 22388 5370 22416 5578
rect 22376 5364 22428 5370
rect 22376 5306 22428 5312
rect 22848 5234 22876 5646
rect 23032 5642 23060 6190
rect 23296 5772 23348 5778
rect 23296 5714 23348 5720
rect 23020 5636 23072 5642
rect 23020 5578 23072 5584
rect 23112 5636 23164 5642
rect 23112 5578 23164 5584
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22560 5228 22612 5234
rect 22560 5170 22612 5176
rect 22836 5228 22888 5234
rect 22836 5170 22888 5176
rect 16394 4584 16450 4593
rect 22572 4554 22600 5170
rect 22848 4826 22876 5170
rect 22836 4820 22888 4826
rect 22836 4762 22888 4768
rect 16394 4519 16450 4528
rect 22560 4548 22612 4554
rect 22560 4490 22612 4496
rect 22848 4486 22876 4762
rect 23124 4690 23152 5578
rect 23112 4684 23164 4690
rect 23112 4626 23164 4632
rect 23308 4554 23336 5714
rect 23400 4826 23428 6598
rect 23768 6118 23796 6734
rect 24124 6656 24176 6662
rect 24124 6598 24176 6604
rect 23756 6112 23808 6118
rect 23756 6054 23808 6060
rect 23572 5908 23624 5914
rect 23572 5850 23624 5856
rect 23480 5636 23532 5642
rect 23480 5578 23532 5584
rect 23492 5370 23520 5578
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 23584 5302 23612 5850
rect 23756 5840 23808 5846
rect 23756 5782 23808 5788
rect 23768 5370 23796 5782
rect 24136 5778 24164 6598
rect 24228 6254 24256 7142
rect 24780 7018 24808 9982
rect 24872 9654 24900 10084
rect 24860 9648 24912 9654
rect 24860 9590 24912 9596
rect 24872 8566 24900 9590
rect 25056 9042 25084 11630
rect 25884 11286 25912 12038
rect 26068 11694 26096 12406
rect 26252 12374 26280 12786
rect 26344 12782 26372 13194
rect 27172 12782 27200 14350
rect 27356 14346 27384 14470
rect 27344 14340 27396 14346
rect 27344 14282 27396 14288
rect 27632 14278 27660 15438
rect 27724 14890 27752 15846
rect 28080 15700 28132 15706
rect 28080 15642 28132 15648
rect 27804 15632 27856 15638
rect 27804 15574 27856 15580
rect 27816 15094 27844 15574
rect 28092 15162 28120 15642
rect 28080 15156 28132 15162
rect 28080 15098 28132 15104
rect 27804 15088 27856 15094
rect 27804 15030 27856 15036
rect 27712 14884 27764 14890
rect 27712 14826 27764 14832
rect 27620 14272 27672 14278
rect 27620 14214 27672 14220
rect 27632 13530 27660 14214
rect 27896 13932 27948 13938
rect 27896 13874 27948 13880
rect 27436 13524 27488 13530
rect 27436 13466 27488 13472
rect 27620 13524 27672 13530
rect 27620 13466 27672 13472
rect 27448 13190 27476 13466
rect 27712 13320 27764 13326
rect 27712 13262 27764 13268
rect 27436 13184 27488 13190
rect 27436 13126 27488 13132
rect 27344 12844 27396 12850
rect 27344 12786 27396 12792
rect 26332 12776 26384 12782
rect 26332 12718 26384 12724
rect 27160 12776 27212 12782
rect 27160 12718 27212 12724
rect 27252 12640 27304 12646
rect 27252 12582 27304 12588
rect 26424 12436 26476 12442
rect 26424 12378 26476 12384
rect 26240 12368 26292 12374
rect 26240 12310 26292 12316
rect 26252 11830 26280 12310
rect 26436 12238 26464 12378
rect 27160 12368 27212 12374
rect 27066 12336 27122 12345
rect 27160 12310 27212 12316
rect 27066 12271 27122 12280
rect 27080 12238 27108 12271
rect 26424 12232 26476 12238
rect 26424 12174 26476 12180
rect 27068 12232 27120 12238
rect 27068 12174 27120 12180
rect 27172 12170 27200 12310
rect 27264 12238 27292 12582
rect 27356 12434 27384 12786
rect 27620 12640 27672 12646
rect 27620 12582 27672 12588
rect 27356 12406 27568 12434
rect 27252 12232 27304 12238
rect 27252 12174 27304 12180
rect 26884 12164 26936 12170
rect 26884 12106 26936 12112
rect 27160 12164 27212 12170
rect 27160 12106 27212 12112
rect 26896 11880 26924 12106
rect 26976 11892 27028 11898
rect 26896 11852 26976 11880
rect 26976 11834 27028 11840
rect 26240 11824 26292 11830
rect 26240 11766 26292 11772
rect 27172 11762 27200 12106
rect 27434 11928 27490 11937
rect 27434 11863 27490 11872
rect 27160 11756 27212 11762
rect 27160 11698 27212 11704
rect 27448 11694 27476 11863
rect 26056 11688 26108 11694
rect 26056 11630 26108 11636
rect 26608 11688 26660 11694
rect 26608 11630 26660 11636
rect 27436 11688 27488 11694
rect 27436 11630 27488 11636
rect 25872 11280 25924 11286
rect 25872 11222 25924 11228
rect 25872 11144 25924 11150
rect 25872 11086 25924 11092
rect 25136 10736 25188 10742
rect 25136 10678 25188 10684
rect 25044 9036 25096 9042
rect 25044 8978 25096 8984
rect 24860 8560 24912 8566
rect 24860 8502 24912 8508
rect 24872 7954 24900 8502
rect 24860 7948 24912 7954
rect 24860 7890 24912 7896
rect 25148 7410 25176 10678
rect 25884 10470 25912 11086
rect 26240 11008 26292 11014
rect 26240 10950 26292 10956
rect 25872 10464 25924 10470
rect 25872 10406 25924 10412
rect 25780 10124 25832 10130
rect 25884 10112 25912 10406
rect 25832 10084 25912 10112
rect 25780 10066 25832 10072
rect 25320 9920 25372 9926
rect 25320 9862 25372 9868
rect 25332 9518 25360 9862
rect 25884 9722 25912 10084
rect 26056 9920 26108 9926
rect 26056 9862 26108 9868
rect 25872 9716 25924 9722
rect 25872 9658 25924 9664
rect 25884 9602 25912 9658
rect 25792 9574 25912 9602
rect 25320 9512 25372 9518
rect 25320 9454 25372 9460
rect 25332 9110 25360 9454
rect 25320 9104 25372 9110
rect 25320 9046 25372 9052
rect 25792 9042 25820 9574
rect 26068 9518 26096 9862
rect 26252 9722 26280 10950
rect 26240 9716 26292 9722
rect 26240 9658 26292 9664
rect 26056 9512 26108 9518
rect 26620 9489 26648 11630
rect 27448 11218 27476 11630
rect 27436 11212 27488 11218
rect 27436 11154 27488 11160
rect 27540 11150 27568 12406
rect 27632 11354 27660 12582
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 27528 11144 27580 11150
rect 27528 11086 27580 11092
rect 26700 11076 26752 11082
rect 26700 11018 26752 11024
rect 26712 10470 26740 11018
rect 27540 10826 27568 11086
rect 27448 10798 27568 10826
rect 27448 10674 27476 10798
rect 27528 10736 27580 10742
rect 27526 10704 27528 10713
rect 27580 10704 27582 10713
rect 27436 10668 27488 10674
rect 27724 10674 27752 13262
rect 27908 12345 27936 13874
rect 28264 13864 28316 13870
rect 28264 13806 28316 13812
rect 28276 13025 28304 13806
rect 28460 13530 28488 17138
rect 32220 16992 32272 16998
rect 32220 16934 32272 16940
rect 31852 16652 31904 16658
rect 31852 16594 31904 16600
rect 29368 16516 29420 16522
rect 29368 16458 29420 16464
rect 28540 15360 28592 15366
rect 28540 15302 28592 15308
rect 28908 15360 28960 15366
rect 28908 15302 28960 15308
rect 28552 14414 28580 15302
rect 28920 15094 28948 15302
rect 28908 15088 28960 15094
rect 28908 15030 28960 15036
rect 28724 14612 28776 14618
rect 28724 14554 28776 14560
rect 28736 14464 28764 14554
rect 28816 14476 28868 14482
rect 28736 14436 28816 14464
rect 28816 14418 28868 14424
rect 28540 14408 28592 14414
rect 28540 14350 28592 14356
rect 28540 13728 28592 13734
rect 28540 13670 28592 13676
rect 28552 13530 28580 13670
rect 28448 13524 28500 13530
rect 28448 13466 28500 13472
rect 28540 13524 28592 13530
rect 28540 13466 28592 13472
rect 29092 13184 29144 13190
rect 29092 13126 29144 13132
rect 28262 13016 28318 13025
rect 28262 12951 28318 12960
rect 29104 12866 29132 13126
rect 29104 12838 29316 12866
rect 29288 12782 29316 12838
rect 29276 12776 29328 12782
rect 29276 12718 29328 12724
rect 27894 12336 27950 12345
rect 27894 12271 27950 12280
rect 28356 12232 28408 12238
rect 28356 12174 28408 12180
rect 28998 12200 29054 12209
rect 27896 12096 27948 12102
rect 27896 12038 27948 12044
rect 27804 11688 27856 11694
rect 27804 11630 27856 11636
rect 27816 11121 27844 11630
rect 27908 11626 27936 12038
rect 27896 11620 27948 11626
rect 27896 11562 27948 11568
rect 28078 11384 28134 11393
rect 28368 11354 28396 12174
rect 28998 12135 29054 12144
rect 28816 11824 28868 11830
rect 28868 11784 28948 11812
rect 28816 11766 28868 11772
rect 28920 11694 28948 11784
rect 29012 11762 29040 12135
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 29380 11694 29408 16458
rect 31392 16176 31444 16182
rect 31392 16118 31444 16124
rect 29552 16108 29604 16114
rect 29552 16050 29604 16056
rect 30104 16108 30156 16114
rect 30104 16050 30156 16056
rect 29564 15910 29592 16050
rect 29736 15972 29788 15978
rect 29736 15914 29788 15920
rect 29552 15904 29604 15910
rect 29552 15846 29604 15852
rect 29564 15337 29592 15846
rect 29550 15328 29606 15337
rect 29550 15263 29606 15272
rect 29644 14952 29696 14958
rect 29644 14894 29696 14900
rect 29656 14657 29684 14894
rect 29642 14648 29698 14657
rect 29642 14583 29698 14592
rect 29458 14512 29514 14521
rect 29458 14447 29514 14456
rect 29472 13530 29500 14447
rect 29644 13728 29696 13734
rect 29644 13670 29696 13676
rect 29656 13569 29684 13670
rect 29642 13560 29698 13569
rect 29460 13524 29512 13530
rect 29642 13495 29698 13504
rect 29460 13466 29512 13472
rect 29552 13456 29604 13462
rect 29552 13398 29604 13404
rect 29564 12850 29592 13398
rect 29748 13326 29776 15914
rect 30116 15706 30144 16050
rect 31404 15706 31432 16118
rect 30104 15700 30156 15706
rect 30104 15642 30156 15648
rect 31392 15700 31444 15706
rect 31392 15642 31444 15648
rect 30116 15026 30144 15642
rect 30472 15496 30524 15502
rect 30472 15438 30524 15444
rect 30104 15020 30156 15026
rect 30104 14962 30156 14968
rect 29920 14952 29972 14958
rect 29920 14894 29972 14900
rect 29826 14240 29882 14249
rect 29826 14175 29882 14184
rect 29840 13870 29868 14175
rect 29828 13864 29880 13870
rect 29828 13806 29880 13812
rect 29736 13320 29788 13326
rect 29736 13262 29788 13268
rect 29644 13184 29696 13190
rect 29644 13126 29696 13132
rect 29552 12844 29604 12850
rect 29552 12786 29604 12792
rect 29460 11756 29512 11762
rect 29460 11698 29512 11704
rect 28816 11688 28868 11694
rect 28816 11630 28868 11636
rect 28908 11688 28960 11694
rect 28908 11630 28960 11636
rect 29184 11688 29236 11694
rect 29184 11630 29236 11636
rect 29368 11688 29420 11694
rect 29368 11630 29420 11636
rect 28632 11552 28684 11558
rect 28630 11520 28632 11529
rect 28684 11520 28686 11529
rect 28630 11455 28686 11464
rect 28078 11319 28134 11328
rect 28356 11348 28408 11354
rect 27802 11112 27858 11121
rect 27802 11047 27858 11056
rect 27986 11112 28042 11121
rect 27986 11047 28042 11056
rect 27526 10639 27582 10648
rect 27712 10668 27764 10674
rect 27436 10610 27488 10616
rect 27712 10610 27764 10616
rect 26700 10464 26752 10470
rect 27528 10464 27580 10470
rect 26700 10406 26752 10412
rect 27066 10432 27122 10441
rect 26056 9454 26108 9460
rect 26606 9480 26662 9489
rect 26606 9415 26608 9424
rect 26660 9415 26662 9424
rect 26608 9386 26660 9392
rect 26712 9330 26740 10406
rect 27528 10406 27580 10412
rect 27066 10367 27122 10376
rect 26792 10192 26844 10198
rect 26792 10134 26844 10140
rect 26804 9625 26832 10134
rect 27080 10033 27108 10367
rect 27436 10056 27488 10062
rect 27066 10024 27122 10033
rect 27436 9998 27488 10004
rect 27066 9959 27122 9968
rect 26790 9616 26846 9625
rect 26790 9551 26846 9560
rect 27068 9580 27120 9586
rect 27068 9522 27120 9528
rect 26528 9302 26740 9330
rect 25780 9036 25832 9042
rect 25780 8978 25832 8984
rect 26528 8906 26556 9302
rect 27080 9110 27108 9522
rect 27448 9178 27476 9998
rect 27540 9518 27568 10406
rect 27724 9654 27752 10610
rect 28000 10577 28028 11047
rect 27986 10568 28042 10577
rect 27986 10503 28042 10512
rect 28000 9994 28028 10503
rect 28092 10470 28120 11319
rect 28356 11290 28408 11296
rect 28828 11286 28856 11630
rect 29196 11529 29224 11630
rect 29182 11520 29238 11529
rect 29182 11455 29238 11464
rect 28816 11280 28868 11286
rect 28816 11222 28868 11228
rect 28906 11248 28962 11257
rect 29380 11218 29408 11630
rect 28906 11183 28962 11192
rect 29368 11212 29420 11218
rect 28920 10810 28948 11183
rect 29368 11154 29420 11160
rect 29092 11076 29144 11082
rect 29092 11018 29144 11024
rect 29000 11008 29052 11014
rect 29000 10950 29052 10956
rect 28908 10804 28960 10810
rect 28908 10746 28960 10752
rect 29012 10742 29040 10950
rect 29000 10736 29052 10742
rect 29000 10678 29052 10684
rect 28080 10464 28132 10470
rect 28080 10406 28132 10412
rect 27988 9988 28040 9994
rect 27988 9930 28040 9936
rect 27712 9648 27764 9654
rect 27712 9590 27764 9596
rect 27528 9512 27580 9518
rect 27528 9454 27580 9460
rect 27526 9208 27582 9217
rect 27436 9172 27488 9178
rect 27526 9143 27528 9152
rect 27436 9114 27488 9120
rect 27580 9143 27582 9152
rect 27528 9114 27580 9120
rect 27068 9104 27120 9110
rect 27068 9046 27120 9052
rect 26516 8900 26568 8906
rect 26516 8842 26568 8848
rect 26148 8288 26200 8294
rect 26148 8230 26200 8236
rect 26160 7478 26188 8230
rect 26528 7954 26556 8842
rect 27080 8838 27108 9046
rect 27068 8832 27120 8838
rect 27068 8774 27120 8780
rect 27724 8634 27752 9590
rect 27712 8628 27764 8634
rect 27712 8570 27764 8576
rect 27526 8392 27582 8401
rect 27526 8327 27582 8336
rect 26240 7948 26292 7954
rect 26240 7890 26292 7896
rect 26516 7948 26568 7954
rect 26516 7890 26568 7896
rect 27160 7948 27212 7954
rect 27160 7890 27212 7896
rect 27252 7948 27304 7954
rect 27252 7890 27304 7896
rect 26252 7478 26280 7890
rect 26148 7472 26200 7478
rect 26148 7414 26200 7420
rect 26240 7472 26292 7478
rect 26240 7414 26292 7420
rect 25136 7404 25188 7410
rect 25136 7346 25188 7352
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 24780 6990 24992 7018
rect 25148 7002 25176 7142
rect 24860 6860 24912 6866
rect 24860 6802 24912 6808
rect 24386 6556 24694 6565
rect 24386 6554 24392 6556
rect 24448 6554 24472 6556
rect 24528 6554 24552 6556
rect 24608 6554 24632 6556
rect 24688 6554 24694 6556
rect 24448 6502 24450 6554
rect 24630 6502 24632 6554
rect 24386 6500 24392 6502
rect 24448 6500 24472 6502
rect 24528 6500 24552 6502
rect 24608 6500 24632 6502
rect 24688 6500 24694 6502
rect 24386 6491 24694 6500
rect 24766 6352 24822 6361
rect 24766 6287 24822 6296
rect 24780 6254 24808 6287
rect 24216 6248 24268 6254
rect 24216 6190 24268 6196
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24308 6112 24360 6118
rect 24308 6054 24360 6060
rect 24124 5772 24176 5778
rect 24124 5714 24176 5720
rect 24216 5704 24268 5710
rect 24216 5646 24268 5652
rect 24032 5568 24084 5574
rect 24032 5510 24084 5516
rect 23756 5364 23808 5370
rect 23756 5306 23808 5312
rect 23572 5296 23624 5302
rect 23572 5238 23624 5244
rect 24044 5234 24072 5510
rect 24228 5302 24256 5646
rect 24216 5296 24268 5302
rect 24216 5238 24268 5244
rect 24032 5228 24084 5234
rect 24032 5170 24084 5176
rect 24228 5030 24256 5238
rect 23664 5024 23716 5030
rect 23664 4966 23716 4972
rect 24216 5024 24268 5030
rect 24216 4966 24268 4972
rect 23388 4820 23440 4826
rect 23388 4762 23440 4768
rect 23676 4622 23704 4966
rect 24228 4758 24256 4966
rect 24216 4752 24268 4758
rect 24216 4694 24268 4700
rect 23664 4616 23716 4622
rect 23664 4558 23716 4564
rect 23296 4548 23348 4554
rect 23296 4490 23348 4496
rect 22836 4480 22888 4486
rect 22836 4422 22888 4428
rect 24228 4214 24256 4694
rect 24320 4554 24348 6054
rect 24872 5710 24900 6802
rect 24964 6474 24992 6990
rect 25136 6996 25188 7002
rect 25136 6938 25188 6944
rect 26146 6896 26202 6905
rect 26146 6831 26202 6840
rect 25594 6760 25650 6769
rect 25594 6695 25596 6704
rect 25648 6695 25650 6704
rect 25596 6666 25648 6672
rect 24964 6446 25268 6474
rect 24952 5840 25004 5846
rect 24952 5782 25004 5788
rect 24860 5704 24912 5710
rect 24964 5681 24992 5782
rect 24860 5646 24912 5652
rect 24950 5672 25006 5681
rect 24872 5574 24900 5646
rect 24950 5607 25006 5616
rect 24860 5568 24912 5574
rect 24860 5510 24912 5516
rect 24386 5468 24694 5477
rect 24386 5466 24392 5468
rect 24448 5466 24472 5468
rect 24528 5466 24552 5468
rect 24608 5466 24632 5468
rect 24688 5466 24694 5468
rect 24448 5414 24450 5466
rect 24630 5414 24632 5466
rect 24386 5412 24392 5414
rect 24448 5412 24472 5414
rect 24528 5412 24552 5414
rect 24608 5412 24632 5414
rect 24688 5412 24694 5414
rect 24386 5403 24694 5412
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 24400 5296 24452 5302
rect 24400 5238 24452 5244
rect 24412 5098 24440 5238
rect 24400 5092 24452 5098
rect 24400 5034 24452 5040
rect 24780 5030 24808 5306
rect 25056 5234 25084 6446
rect 25240 6390 25268 6446
rect 25228 6384 25280 6390
rect 25228 6326 25280 6332
rect 25596 6384 25648 6390
rect 25596 6326 25648 6332
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 25148 5953 25176 6190
rect 25134 5944 25190 5953
rect 25134 5879 25190 5888
rect 25228 5704 25280 5710
rect 25228 5646 25280 5652
rect 25412 5704 25464 5710
rect 25412 5646 25464 5652
rect 25240 5574 25268 5646
rect 25136 5568 25188 5574
rect 25136 5510 25188 5516
rect 25228 5568 25280 5574
rect 25228 5510 25280 5516
rect 25044 5228 25096 5234
rect 25044 5170 25096 5176
rect 24860 5160 24912 5166
rect 24860 5102 24912 5108
rect 24676 5024 24728 5030
rect 24674 4992 24676 5001
rect 24768 5024 24820 5030
rect 24728 4992 24730 5001
rect 24768 4966 24820 4972
rect 24674 4927 24730 4936
rect 24688 4690 24716 4927
rect 24872 4690 24900 5102
rect 24676 4684 24728 4690
rect 24676 4626 24728 4632
rect 24860 4684 24912 4690
rect 24860 4626 24912 4632
rect 25148 4622 25176 5510
rect 25044 4616 25096 4622
rect 25044 4558 25096 4564
rect 25136 4616 25188 4622
rect 25136 4558 25188 4564
rect 24308 4548 24360 4554
rect 24308 4490 24360 4496
rect 24386 4380 24694 4389
rect 24386 4378 24392 4380
rect 24448 4378 24472 4380
rect 24528 4378 24552 4380
rect 24608 4378 24632 4380
rect 24688 4378 24694 4380
rect 24448 4326 24450 4378
rect 24630 4326 24632 4378
rect 24386 4324 24392 4326
rect 24448 4324 24472 4326
rect 24528 4324 24552 4326
rect 24608 4324 24632 4326
rect 24688 4324 24694 4326
rect 24386 4315 24694 4324
rect 25056 4214 25084 4558
rect 15476 4208 15528 4214
rect 15476 4150 15528 4156
rect 24216 4208 24268 4214
rect 24216 4150 24268 4156
rect 25044 4208 25096 4214
rect 25044 4150 25096 4156
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 13544 4004 13596 4010
rect 13544 3946 13596 3952
rect 12668 3836 12976 3845
rect 12668 3834 12674 3836
rect 12730 3834 12754 3836
rect 12810 3834 12834 3836
rect 12890 3834 12914 3836
rect 12970 3834 12976 3836
rect 12730 3782 12732 3834
rect 12912 3782 12914 3834
rect 12668 3780 12674 3782
rect 12730 3780 12754 3782
rect 12810 3780 12834 3782
rect 12890 3780 12914 3782
rect 12970 3780 12976 3782
rect 12668 3771 12976 3780
rect 13556 3738 13584 3946
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 13556 2774 13584 3674
rect 15212 3534 15240 3878
rect 15488 3534 15516 4150
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 12668 2748 12976 2757
rect 12668 2746 12674 2748
rect 12730 2746 12754 2748
rect 12810 2746 12834 2748
rect 12890 2746 12914 2748
rect 12970 2746 12976 2748
rect 12730 2694 12732 2746
rect 12912 2694 12914 2746
rect 12668 2692 12674 2694
rect 12730 2692 12754 2694
rect 12810 2692 12834 2694
rect 12890 2692 12914 2694
rect 12970 2692 12976 2694
rect 12668 2683 12976 2692
rect 13372 2746 13584 2774
rect 13372 2446 13400 2746
rect 15488 2446 15516 3470
rect 24228 3398 24256 4150
rect 25424 4078 25452 5646
rect 25608 5642 25636 6326
rect 25872 6248 25924 6254
rect 25872 6190 25924 6196
rect 25884 5914 25912 6190
rect 25688 5908 25740 5914
rect 25688 5850 25740 5856
rect 25872 5908 25924 5914
rect 25872 5850 25924 5856
rect 25700 5710 25728 5850
rect 26160 5710 26188 6831
rect 26252 6730 26280 7414
rect 27172 7342 27200 7890
rect 26608 7336 26660 7342
rect 26608 7278 26660 7284
rect 27160 7336 27212 7342
rect 27160 7278 27212 7284
rect 26620 6882 26648 7278
rect 27264 7206 27292 7890
rect 27540 7546 27568 8327
rect 28000 8022 28028 9930
rect 29012 9926 29040 10678
rect 29104 10198 29132 11018
rect 29092 10192 29144 10198
rect 29092 10134 29144 10140
rect 29000 9920 29052 9926
rect 29000 9862 29052 9868
rect 29012 9761 29040 9862
rect 28998 9752 29054 9761
rect 28998 9687 29054 9696
rect 29000 9376 29052 9382
rect 29000 9318 29052 9324
rect 29012 9178 29040 9318
rect 29380 9178 29408 11154
rect 29472 11150 29500 11698
rect 29460 11144 29512 11150
rect 29460 11086 29512 11092
rect 29656 10674 29684 13126
rect 29644 10668 29696 10674
rect 29644 10610 29696 10616
rect 29656 10130 29684 10610
rect 29748 10538 29776 13262
rect 29826 12880 29882 12889
rect 29826 12815 29882 12824
rect 29840 12782 29868 12815
rect 29828 12776 29880 12782
rect 29828 12718 29880 12724
rect 29932 12442 29960 14894
rect 30484 14414 30512 15438
rect 31404 15026 31432 15642
rect 31392 15020 31444 15026
rect 31392 14962 31444 14968
rect 31484 15020 31536 15026
rect 31484 14962 31536 14968
rect 30748 14952 30800 14958
rect 30748 14894 30800 14900
rect 30656 14476 30708 14482
rect 30656 14418 30708 14424
rect 30472 14408 30524 14414
rect 30472 14350 30524 14356
rect 30012 14272 30064 14278
rect 30012 14214 30064 14220
rect 30196 14272 30248 14278
rect 30196 14214 30248 14220
rect 30024 13258 30052 14214
rect 30208 14006 30236 14214
rect 30288 14068 30340 14074
rect 30288 14010 30340 14016
rect 30196 14000 30248 14006
rect 30196 13942 30248 13948
rect 30104 13932 30156 13938
rect 30104 13874 30156 13880
rect 30116 13734 30144 13874
rect 30300 13818 30328 14010
rect 30300 13802 30512 13818
rect 30196 13796 30248 13802
rect 30300 13796 30524 13802
rect 30300 13790 30472 13796
rect 30196 13738 30248 13744
rect 30472 13738 30524 13744
rect 30104 13728 30156 13734
rect 30104 13670 30156 13676
rect 30208 13530 30236 13738
rect 30668 13734 30696 14418
rect 30760 14090 30788 14894
rect 31392 14272 31444 14278
rect 31392 14214 31444 14220
rect 30760 14062 30880 14090
rect 30748 13864 30800 13870
rect 30748 13806 30800 13812
rect 30656 13728 30708 13734
rect 30656 13670 30708 13676
rect 30196 13524 30248 13530
rect 30196 13466 30248 13472
rect 30564 13388 30616 13394
rect 30564 13330 30616 13336
rect 30012 13252 30064 13258
rect 30012 13194 30064 13200
rect 30472 13252 30524 13258
rect 30472 13194 30524 13200
rect 30484 12986 30512 13194
rect 30576 12986 30604 13330
rect 30472 12980 30524 12986
rect 30472 12922 30524 12928
rect 30564 12980 30616 12986
rect 30564 12922 30616 12928
rect 30116 12850 30512 12866
rect 30104 12844 30524 12850
rect 30156 12838 30472 12844
rect 30104 12786 30156 12792
rect 30472 12786 30524 12792
rect 30760 12442 30788 13806
rect 30852 12646 30880 14062
rect 30932 13864 30984 13870
rect 30932 13806 30984 13812
rect 30944 13569 30972 13806
rect 31024 13728 31076 13734
rect 31024 13670 31076 13676
rect 30930 13560 30986 13569
rect 31036 13530 31064 13670
rect 30930 13495 30986 13504
rect 31024 13524 31076 13530
rect 31024 13466 31076 13472
rect 31114 13152 31170 13161
rect 31114 13087 31170 13096
rect 30840 12640 30892 12646
rect 30840 12582 30892 12588
rect 29920 12436 29972 12442
rect 29920 12378 29972 12384
rect 30748 12436 30800 12442
rect 30748 12378 30800 12384
rect 30656 12368 30708 12374
rect 30656 12310 30708 12316
rect 30288 12300 30340 12306
rect 30288 12242 30340 12248
rect 30196 12232 30248 12238
rect 30196 12174 30248 12180
rect 30208 11937 30236 12174
rect 30194 11928 30250 11937
rect 30194 11863 30250 11872
rect 30010 11656 30066 11665
rect 30010 11591 30066 11600
rect 30024 11354 30052 11591
rect 30012 11348 30064 11354
rect 30012 11290 30064 11296
rect 30024 11014 30052 11290
rect 30300 11082 30328 12242
rect 30668 11830 30696 12310
rect 31128 12306 31156 13087
rect 31404 12850 31432 14214
rect 31496 13938 31524 14962
rect 31758 14648 31814 14657
rect 31758 14583 31814 14592
rect 31772 13938 31800 14583
rect 31864 14482 31892 16594
rect 32232 16454 32260 16934
rect 32220 16448 32272 16454
rect 32220 16390 32272 16396
rect 32864 16448 32916 16454
rect 32864 16390 32916 16396
rect 32232 15502 32260 16390
rect 32876 16250 32904 16390
rect 32864 16244 32916 16250
rect 32864 16186 32916 16192
rect 32876 15978 32904 16186
rect 32864 15972 32916 15978
rect 32864 15914 32916 15920
rect 32772 15904 32824 15910
rect 32772 15846 32824 15852
rect 32220 15496 32272 15502
rect 32220 15438 32272 15444
rect 32784 15434 32812 15846
rect 32876 15502 32904 15914
rect 34060 15904 34112 15910
rect 34060 15846 34112 15852
rect 32864 15496 32916 15502
rect 32864 15438 32916 15444
rect 32404 15428 32456 15434
rect 32404 15370 32456 15376
rect 32588 15428 32640 15434
rect 32588 15370 32640 15376
rect 32772 15428 32824 15434
rect 32772 15370 32824 15376
rect 32036 14884 32088 14890
rect 32036 14826 32088 14832
rect 32048 14482 32076 14826
rect 31852 14476 31904 14482
rect 31852 14418 31904 14424
rect 32036 14476 32088 14482
rect 32036 14418 32088 14424
rect 31484 13932 31536 13938
rect 31484 13874 31536 13880
rect 31760 13932 31812 13938
rect 31760 13874 31812 13880
rect 31496 13530 31524 13874
rect 31772 13530 31800 13874
rect 31484 13524 31536 13530
rect 31484 13466 31536 13472
rect 31760 13524 31812 13530
rect 31760 13466 31812 13472
rect 31484 13252 31536 13258
rect 31484 13194 31536 13200
rect 31300 12844 31352 12850
rect 31300 12786 31352 12792
rect 31392 12844 31444 12850
rect 31392 12786 31444 12792
rect 31312 12646 31340 12786
rect 31496 12782 31524 13194
rect 31484 12776 31536 12782
rect 31484 12718 31536 12724
rect 31668 12776 31720 12782
rect 31668 12718 31720 12724
rect 31392 12708 31444 12714
rect 31392 12650 31444 12656
rect 31300 12640 31352 12646
rect 31300 12582 31352 12588
rect 31404 12374 31432 12650
rect 31392 12368 31444 12374
rect 31392 12310 31444 12316
rect 31116 12300 31168 12306
rect 31116 12242 31168 12248
rect 31128 11830 31156 12242
rect 31300 12232 31352 12238
rect 31300 12174 31352 12180
rect 30656 11824 30708 11830
rect 30656 11766 30708 11772
rect 31116 11824 31168 11830
rect 31116 11766 31168 11772
rect 31312 11286 31340 12174
rect 31576 11756 31628 11762
rect 31576 11698 31628 11704
rect 31484 11620 31536 11626
rect 31484 11562 31536 11568
rect 31496 11354 31524 11562
rect 31588 11558 31616 11698
rect 31576 11552 31628 11558
rect 31576 11494 31628 11500
rect 31484 11348 31536 11354
rect 31484 11290 31536 11296
rect 30472 11280 30524 11286
rect 30472 11222 30524 11228
rect 31300 11280 31352 11286
rect 31300 11222 31352 11228
rect 30288 11076 30340 11082
rect 30288 11018 30340 11024
rect 30380 11076 30432 11082
rect 30380 11018 30432 11024
rect 30012 11008 30064 11014
rect 30012 10950 30064 10956
rect 30288 10668 30340 10674
rect 30288 10610 30340 10616
rect 29736 10532 29788 10538
rect 29736 10474 29788 10480
rect 29826 10432 29882 10441
rect 29826 10367 29882 10376
rect 29644 10124 29696 10130
rect 29644 10066 29696 10072
rect 29840 10062 29868 10367
rect 29828 10056 29880 10062
rect 29828 9998 29880 10004
rect 29920 10056 29972 10062
rect 29920 9998 29972 10004
rect 29458 9752 29514 9761
rect 29458 9687 29514 9696
rect 29000 9172 29052 9178
rect 29000 9114 29052 9120
rect 29368 9172 29420 9178
rect 29368 9114 29420 9120
rect 28540 9036 28592 9042
rect 28540 8978 28592 8984
rect 28448 8968 28500 8974
rect 28448 8910 28500 8916
rect 27988 8016 28040 8022
rect 27988 7958 28040 7964
rect 28460 7886 28488 8910
rect 28552 8634 28580 8978
rect 28724 8832 28776 8838
rect 28776 8780 29040 8786
rect 28724 8774 29040 8780
rect 28736 8758 29040 8774
rect 28540 8628 28592 8634
rect 28540 8570 28592 8576
rect 28632 8084 28684 8090
rect 28632 8026 28684 8032
rect 28448 7880 28500 7886
rect 28448 7822 28500 7828
rect 27712 7812 27764 7818
rect 27712 7754 27764 7760
rect 27528 7540 27580 7546
rect 27528 7482 27580 7488
rect 27724 7410 27752 7754
rect 28460 7546 28488 7822
rect 28448 7540 28500 7546
rect 28448 7482 28500 7488
rect 27712 7404 27764 7410
rect 27712 7346 27764 7352
rect 28644 7274 28672 8026
rect 29012 8022 29040 8758
rect 29472 8362 29500 9687
rect 29932 9518 29960 9998
rect 30196 9648 30248 9654
rect 30194 9616 30196 9625
rect 30248 9616 30250 9625
rect 30194 9551 30250 9560
rect 29920 9512 29972 9518
rect 30300 9489 30328 10610
rect 30392 10266 30420 11018
rect 30484 10985 30512 11222
rect 31680 10985 31708 12718
rect 31772 12238 31800 13466
rect 31864 12434 31892 14418
rect 32416 14006 32444 15370
rect 32404 14000 32456 14006
rect 32404 13942 32456 13948
rect 32220 13184 32272 13190
rect 32220 13126 32272 13132
rect 31864 12406 32076 12434
rect 31760 12232 31812 12238
rect 31760 12174 31812 12180
rect 31772 11070 31984 11098
rect 31772 11014 31800 11070
rect 31760 11008 31812 11014
rect 30470 10976 30526 10985
rect 30470 10911 30526 10920
rect 31666 10976 31722 10985
rect 31760 10950 31812 10956
rect 31852 11008 31904 11014
rect 31852 10950 31904 10956
rect 31666 10911 31722 10920
rect 31208 10804 31260 10810
rect 31208 10746 31260 10752
rect 31220 10470 31248 10746
rect 31300 10736 31352 10742
rect 31300 10678 31352 10684
rect 31312 10588 31340 10678
rect 31864 10674 31892 10950
rect 31956 10674 31984 11070
rect 31852 10668 31904 10674
rect 31852 10610 31904 10616
rect 31944 10668 31996 10674
rect 31944 10610 31996 10616
rect 31484 10600 31536 10606
rect 31312 10560 31484 10588
rect 31484 10542 31536 10548
rect 31864 10538 31892 10610
rect 31852 10532 31904 10538
rect 31852 10474 31904 10480
rect 31208 10464 31260 10470
rect 31208 10406 31260 10412
rect 30380 10260 30432 10266
rect 30380 10202 30432 10208
rect 30656 9512 30708 9518
rect 29920 9454 29972 9460
rect 30286 9480 30342 9489
rect 29736 9104 29788 9110
rect 29736 9046 29788 9052
rect 29644 8832 29696 8838
rect 29644 8774 29696 8780
rect 29460 8356 29512 8362
rect 29460 8298 29512 8304
rect 29000 8016 29052 8022
rect 29000 7958 29052 7964
rect 28724 7744 28776 7750
rect 28724 7686 28776 7692
rect 28908 7744 28960 7750
rect 28908 7686 28960 7692
rect 28736 7342 28764 7686
rect 28724 7336 28776 7342
rect 28776 7284 28856 7290
rect 28724 7278 28856 7284
rect 28632 7268 28684 7274
rect 28632 7210 28684 7216
rect 28736 7262 28856 7278
rect 28736 7213 28764 7262
rect 27252 7200 27304 7206
rect 27252 7142 27304 7148
rect 28080 7200 28132 7206
rect 28080 7142 28132 7148
rect 28092 7002 28120 7142
rect 28080 6996 28132 7002
rect 28080 6938 28132 6944
rect 28448 6996 28500 7002
rect 28448 6938 28500 6944
rect 26700 6928 26752 6934
rect 26344 6866 26648 6882
rect 26332 6860 26648 6866
rect 26384 6854 26648 6860
rect 26332 6802 26384 6808
rect 26620 6746 26648 6854
rect 26698 6896 26700 6905
rect 26752 6896 26754 6905
rect 28460 6866 28488 6938
rect 26698 6831 26754 6840
rect 28448 6860 28500 6866
rect 28448 6802 28500 6808
rect 26240 6724 26292 6730
rect 26620 6718 26740 6746
rect 26240 6666 26292 6672
rect 26424 6384 26476 6390
rect 26422 6352 26424 6361
rect 26476 6352 26478 6361
rect 26422 6287 26478 6296
rect 26516 6316 26568 6322
rect 26516 6258 26568 6264
rect 26240 6180 26292 6186
rect 26240 6122 26292 6128
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 26148 5704 26200 5710
rect 26148 5646 26200 5652
rect 25596 5636 25648 5642
rect 25596 5578 25648 5584
rect 25700 4622 25728 5646
rect 26252 5302 26280 6122
rect 26240 5296 26292 5302
rect 26528 5250 26556 6258
rect 26712 6118 26740 6718
rect 28172 6724 28224 6730
rect 28172 6666 28224 6672
rect 28184 6458 28212 6666
rect 28172 6452 28224 6458
rect 28172 6394 28224 6400
rect 26700 6112 26752 6118
rect 26700 6054 26752 6060
rect 27436 6112 27488 6118
rect 27436 6054 27488 6060
rect 26712 5710 26740 6054
rect 27066 5808 27122 5817
rect 27066 5743 27068 5752
rect 27120 5743 27122 5752
rect 27068 5714 27120 5720
rect 26700 5704 26752 5710
rect 26700 5646 26752 5652
rect 26240 5238 26292 5244
rect 26436 5222 26556 5250
rect 26436 5001 26464 5222
rect 26516 5160 26568 5166
rect 26712 5114 26740 5646
rect 27448 5642 27476 6054
rect 28460 5846 28488 6802
rect 28724 6656 28776 6662
rect 28724 6598 28776 6604
rect 28736 5914 28764 6598
rect 28828 6118 28856 7262
rect 28920 7206 28948 7686
rect 28908 7200 28960 7206
rect 28908 7142 28960 7148
rect 29472 6866 29500 8298
rect 29656 7478 29684 8774
rect 29748 8430 29776 9046
rect 29932 9042 29960 9454
rect 30656 9454 30708 9460
rect 30286 9415 30342 9424
rect 29920 9036 29972 9042
rect 29920 8978 29972 8984
rect 29828 8560 29880 8566
rect 29828 8502 29880 8508
rect 29736 8424 29788 8430
rect 29736 8366 29788 8372
rect 29840 7818 29868 8502
rect 29932 8498 29960 8978
rect 30012 8832 30064 8838
rect 30012 8774 30064 8780
rect 29920 8492 29972 8498
rect 29920 8434 29972 8440
rect 29920 8356 29972 8362
rect 30024 8344 30052 8774
rect 30668 8566 30696 9454
rect 31484 9444 31536 9450
rect 31484 9386 31536 9392
rect 31496 9110 31524 9386
rect 31668 9376 31720 9382
rect 31668 9318 31720 9324
rect 31680 9178 31708 9318
rect 31668 9172 31720 9178
rect 31668 9114 31720 9120
rect 31484 9104 31536 9110
rect 31484 9046 31536 9052
rect 31484 8900 31536 8906
rect 31484 8842 31536 8848
rect 31760 8900 31812 8906
rect 32048 8888 32076 12406
rect 32126 12336 32182 12345
rect 32126 12271 32182 12280
rect 32140 12238 32168 12271
rect 32232 12238 32260 13126
rect 32416 12918 32444 13942
rect 32600 13938 32628 15370
rect 32680 15360 32732 15366
rect 33140 15360 33192 15366
rect 32680 15302 32732 15308
rect 33060 15320 33140 15348
rect 32588 13932 32640 13938
rect 32588 13874 32640 13880
rect 32692 13394 32720 15302
rect 32956 15020 33008 15026
rect 32956 14962 33008 14968
rect 32772 14952 32824 14958
rect 32772 14894 32824 14900
rect 32784 14482 32812 14894
rect 32772 14476 32824 14482
rect 32772 14418 32824 14424
rect 32968 14346 32996 14962
rect 33060 14822 33088 15320
rect 33140 15302 33192 15308
rect 33324 15156 33376 15162
rect 33324 15098 33376 15104
rect 33232 14952 33284 14958
rect 33232 14894 33284 14900
rect 33048 14816 33100 14822
rect 33048 14758 33100 14764
rect 33244 14634 33272 14894
rect 33060 14606 33272 14634
rect 32956 14340 33008 14346
rect 32956 14282 33008 14288
rect 32772 13524 32824 13530
rect 32772 13466 32824 13472
rect 32864 13524 32916 13530
rect 32864 13466 32916 13472
rect 32784 13394 32812 13466
rect 32680 13388 32732 13394
rect 32680 13330 32732 13336
rect 32772 13388 32824 13394
rect 32772 13330 32824 13336
rect 32496 13320 32548 13326
rect 32876 13274 32904 13466
rect 32496 13262 32548 13268
rect 32404 12912 32456 12918
rect 32404 12854 32456 12860
rect 32508 12434 32536 13262
rect 32784 13246 32904 13274
rect 32586 12880 32642 12889
rect 32586 12815 32588 12824
rect 32640 12815 32642 12824
rect 32588 12786 32640 12792
rect 32508 12406 32628 12434
rect 32404 12300 32456 12306
rect 32404 12242 32456 12248
rect 32128 12232 32180 12238
rect 32128 12174 32180 12180
rect 32220 12232 32272 12238
rect 32220 12174 32272 12180
rect 32416 12170 32444 12242
rect 32404 12164 32456 12170
rect 32404 12106 32456 12112
rect 32402 12064 32458 12073
rect 32402 11999 32458 12008
rect 32416 10305 32444 11999
rect 32496 11892 32548 11898
rect 32496 11834 32548 11840
rect 32508 11286 32536 11834
rect 32496 11280 32548 11286
rect 32496 11222 32548 11228
rect 32496 11144 32548 11150
rect 32496 11086 32548 11092
rect 32402 10296 32458 10305
rect 32402 10231 32458 10240
rect 32508 10130 32536 11086
rect 32496 10124 32548 10130
rect 32496 10066 32548 10072
rect 32508 9586 32536 10066
rect 32496 9580 32548 9586
rect 32496 9522 32548 9528
rect 32508 9042 32536 9522
rect 32600 9489 32628 12406
rect 32678 11248 32734 11257
rect 32678 11183 32734 11192
rect 32692 10606 32720 11183
rect 32784 10674 32812 13246
rect 32864 13184 32916 13190
rect 32864 13126 32916 13132
rect 32876 12918 32904 13126
rect 32864 12912 32916 12918
rect 32864 12854 32916 12860
rect 33060 12170 33088 14606
rect 33336 14498 33364 15098
rect 33244 14470 33364 14498
rect 33140 13728 33192 13734
rect 33244 13716 33272 14470
rect 33968 14340 34020 14346
rect 33968 14282 34020 14288
rect 33980 13870 34008 14282
rect 34072 13870 34100 15846
rect 34244 14272 34296 14278
rect 34244 14214 34296 14220
rect 34256 14006 34284 14214
rect 34244 14000 34296 14006
rect 34244 13942 34296 13948
rect 33968 13864 34020 13870
rect 33968 13806 34020 13812
rect 34060 13864 34112 13870
rect 34060 13806 34112 13812
rect 33192 13688 33272 13716
rect 33324 13728 33376 13734
rect 33140 13670 33192 13676
rect 33324 13670 33376 13676
rect 33416 13728 33468 13734
rect 33416 13670 33468 13676
rect 33336 12918 33364 13670
rect 33428 13530 33456 13670
rect 33416 13524 33468 13530
rect 33416 13466 33468 13472
rect 33980 13258 34008 13806
rect 33968 13252 34020 13258
rect 33968 13194 34020 13200
rect 33324 12912 33376 12918
rect 33324 12854 33376 12860
rect 33600 12640 33652 12646
rect 33600 12582 33652 12588
rect 33968 12640 34020 12646
rect 33968 12582 34020 12588
rect 33048 12164 33100 12170
rect 33048 12106 33100 12112
rect 32864 12096 32916 12102
rect 32864 12038 32916 12044
rect 32772 10668 32824 10674
rect 32772 10610 32824 10616
rect 32680 10600 32732 10606
rect 32680 10542 32732 10548
rect 32876 10146 32904 12038
rect 33508 11688 33560 11694
rect 33508 11630 33560 11636
rect 33416 11552 33468 11558
rect 33414 11520 33416 11529
rect 33468 11520 33470 11529
rect 33414 11455 33470 11464
rect 33048 11076 33100 11082
rect 33048 11018 33100 11024
rect 32954 10568 33010 10577
rect 32954 10503 32956 10512
rect 33008 10503 33010 10512
rect 32956 10474 33008 10480
rect 33060 10470 33088 11018
rect 33520 10742 33548 11630
rect 33508 10736 33560 10742
rect 33508 10678 33560 10684
rect 33048 10464 33100 10470
rect 33048 10406 33100 10412
rect 33140 10192 33192 10198
rect 32876 10118 32996 10146
rect 33192 10140 33364 10146
rect 33140 10134 33364 10140
rect 33152 10118 33364 10134
rect 32772 9988 32824 9994
rect 32824 9948 32904 9976
rect 32772 9930 32824 9936
rect 32586 9480 32642 9489
rect 32586 9415 32642 9424
rect 32496 9036 32548 9042
rect 32496 8978 32548 8984
rect 31812 8860 32076 8888
rect 31760 8842 31812 8848
rect 31496 8566 31524 8842
rect 31668 8832 31720 8838
rect 31720 8780 31892 8786
rect 31668 8774 31892 8780
rect 31680 8758 31892 8774
rect 30656 8560 30708 8566
rect 30656 8502 30708 8508
rect 31484 8560 31536 8566
rect 31484 8502 31536 8508
rect 31864 8362 31892 8758
rect 32508 8498 32536 8978
rect 32876 8974 32904 9948
rect 32864 8968 32916 8974
rect 32864 8910 32916 8916
rect 32496 8492 32548 8498
rect 32496 8434 32548 8440
rect 29972 8316 30052 8344
rect 31852 8356 31904 8362
rect 29920 8298 29972 8304
rect 31852 8298 31904 8304
rect 32404 8356 32456 8362
rect 32404 8298 32456 8304
rect 31668 8288 31720 8294
rect 31668 8230 31720 8236
rect 30472 7880 30524 7886
rect 30472 7822 30524 7828
rect 29828 7812 29880 7818
rect 29828 7754 29880 7760
rect 29644 7472 29696 7478
rect 29644 7414 29696 7420
rect 29460 6860 29512 6866
rect 29460 6802 29512 6808
rect 29736 6656 29788 6662
rect 29736 6598 29788 6604
rect 29748 6390 29776 6598
rect 29736 6384 29788 6390
rect 29736 6326 29788 6332
rect 28816 6112 28868 6118
rect 28816 6054 28868 6060
rect 28724 5908 28776 5914
rect 28724 5850 28776 5856
rect 28448 5840 28500 5846
rect 28448 5782 28500 5788
rect 29840 5642 29868 7754
rect 30196 7336 30248 7342
rect 30196 7278 30248 7284
rect 30208 6866 30236 7278
rect 30196 6860 30248 6866
rect 30196 6802 30248 6808
rect 30104 6792 30156 6798
rect 30104 6734 30156 6740
rect 30116 6186 30144 6734
rect 30208 6322 30236 6802
rect 30484 6730 30512 7822
rect 30748 7540 30800 7546
rect 30748 7482 30800 7488
rect 30472 6724 30524 6730
rect 30472 6666 30524 6672
rect 30484 6497 30512 6666
rect 30470 6488 30526 6497
rect 30470 6423 30526 6432
rect 30196 6316 30248 6322
rect 30196 6258 30248 6264
rect 30760 6254 30788 7482
rect 31680 7274 31708 8230
rect 32416 7478 32444 8298
rect 32772 8288 32824 8294
rect 32772 8230 32824 8236
rect 31760 7472 31812 7478
rect 31760 7414 31812 7420
rect 32404 7472 32456 7478
rect 32404 7414 32456 7420
rect 31668 7268 31720 7274
rect 31668 7210 31720 7216
rect 31208 6928 31260 6934
rect 31206 6896 31208 6905
rect 31772 6914 31800 7414
rect 32784 7206 32812 8230
rect 32864 7336 32916 7342
rect 32864 7278 32916 7284
rect 32772 7200 32824 7206
rect 32772 7142 32824 7148
rect 32876 6934 32904 7278
rect 31260 6896 31262 6905
rect 31206 6831 31262 6840
rect 31680 6886 31800 6914
rect 32864 6928 32916 6934
rect 31680 6730 31708 6886
rect 32864 6870 32916 6876
rect 31668 6724 31720 6730
rect 31668 6666 31720 6672
rect 32312 6452 32364 6458
rect 32312 6394 32364 6400
rect 32324 6361 32352 6394
rect 32310 6352 32366 6361
rect 32876 6322 32904 6870
rect 32310 6287 32366 6296
rect 32496 6316 32548 6322
rect 32496 6258 32548 6264
rect 32864 6316 32916 6322
rect 32864 6258 32916 6264
rect 30748 6248 30800 6254
rect 30748 6190 30800 6196
rect 30104 6180 30156 6186
rect 30104 6122 30156 6128
rect 32508 5778 32536 6258
rect 32680 6180 32732 6186
rect 32680 6122 32732 6128
rect 31760 5772 31812 5778
rect 31760 5714 31812 5720
rect 32496 5772 32548 5778
rect 32496 5714 32548 5720
rect 27436 5636 27488 5642
rect 27436 5578 27488 5584
rect 29828 5636 29880 5642
rect 29828 5578 29880 5584
rect 28264 5296 28316 5302
rect 28262 5264 28264 5273
rect 28316 5264 28318 5273
rect 28262 5199 28318 5208
rect 26568 5108 26740 5114
rect 26516 5102 26740 5108
rect 27252 5160 27304 5166
rect 27252 5102 27304 5108
rect 26528 5098 26740 5102
rect 26528 5092 26752 5098
rect 26528 5086 26700 5092
rect 26422 4992 26478 5001
rect 26422 4927 26478 4936
rect 26528 4826 26556 5086
rect 26700 5034 26752 5040
rect 27264 4826 27292 5102
rect 28448 5024 28500 5030
rect 28448 4966 28500 4972
rect 26332 4820 26384 4826
rect 26332 4762 26384 4768
rect 26516 4820 26568 4826
rect 26516 4762 26568 4768
rect 27252 4820 27304 4826
rect 27252 4762 27304 4768
rect 25688 4616 25740 4622
rect 25688 4558 25740 4564
rect 25700 4146 25728 4558
rect 26344 4486 26372 4762
rect 26148 4480 26200 4486
rect 26148 4422 26200 4428
rect 26332 4480 26384 4486
rect 26332 4422 26384 4428
rect 26160 4214 26188 4422
rect 26148 4208 26200 4214
rect 26148 4150 26200 4156
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 25412 4072 25464 4078
rect 25412 4014 25464 4020
rect 24216 3392 24268 3398
rect 24216 3334 24268 3340
rect 24386 3292 24694 3301
rect 24386 3290 24392 3292
rect 24448 3290 24472 3292
rect 24528 3290 24552 3292
rect 24608 3290 24632 3292
rect 24688 3290 24694 3292
rect 24448 3238 24450 3290
rect 24630 3238 24632 3290
rect 24386 3236 24392 3238
rect 24448 3236 24472 3238
rect 24528 3236 24552 3238
rect 24608 3236 24632 3238
rect 24688 3236 24694 3238
rect 24386 3227 24694 3236
rect 28460 2446 28488 4966
rect 29840 4622 29868 5578
rect 31772 5234 31800 5714
rect 32692 5574 32720 6122
rect 32770 5672 32826 5681
rect 32770 5607 32772 5616
rect 32824 5607 32826 5616
rect 32772 5578 32824 5584
rect 32588 5568 32640 5574
rect 32588 5510 32640 5516
rect 32680 5568 32732 5574
rect 32680 5510 32732 5516
rect 32600 5352 32628 5510
rect 32600 5324 32812 5352
rect 31760 5228 31812 5234
rect 31760 5170 31812 5176
rect 32680 5228 32732 5234
rect 32680 5170 32732 5176
rect 30012 5024 30064 5030
rect 30012 4966 30064 4972
rect 30104 5024 30156 5030
rect 30104 4966 30156 4972
rect 29828 4616 29880 4622
rect 29828 4558 29880 4564
rect 30024 4214 30052 4966
rect 30116 4758 30144 4966
rect 31116 4820 31168 4826
rect 31116 4762 31168 4768
rect 30104 4752 30156 4758
rect 30104 4694 30156 4700
rect 30840 4616 30892 4622
rect 30840 4558 30892 4564
rect 30012 4208 30064 4214
rect 30012 4150 30064 4156
rect 30852 4146 30880 4558
rect 31128 4554 31156 4762
rect 31116 4548 31168 4554
rect 31116 4490 31168 4496
rect 31392 4548 31444 4554
rect 31392 4490 31444 4496
rect 32312 4548 32364 4554
rect 32312 4490 32364 4496
rect 31404 4282 31432 4490
rect 31392 4276 31444 4282
rect 31392 4218 31444 4224
rect 30840 4140 30892 4146
rect 30840 4082 30892 4088
rect 32324 3738 32352 4490
rect 32692 4214 32720 5170
rect 32784 5098 32812 5324
rect 32772 5092 32824 5098
rect 32772 5034 32824 5040
rect 32680 4208 32732 4214
rect 32680 4150 32732 4156
rect 32312 3732 32364 3738
rect 32312 3674 32364 3680
rect 32968 3670 32996 10118
rect 33140 10056 33192 10062
rect 33192 10004 33272 10010
rect 33140 9998 33272 10004
rect 33152 9982 33272 9998
rect 33140 9920 33192 9926
rect 33140 9862 33192 9868
rect 33152 9722 33180 9862
rect 33140 9716 33192 9722
rect 33140 9658 33192 9664
rect 33048 9376 33100 9382
rect 33048 9318 33100 9324
rect 33060 9217 33088 9318
rect 33046 9208 33102 9217
rect 33046 9143 33102 9152
rect 33244 9110 33272 9982
rect 33336 9489 33364 10118
rect 33416 9988 33468 9994
rect 33468 9948 33548 9976
rect 33416 9930 33468 9936
rect 33520 9654 33548 9948
rect 33508 9648 33560 9654
rect 33508 9590 33560 9596
rect 33322 9480 33378 9489
rect 33322 9415 33378 9424
rect 33324 9376 33376 9382
rect 33324 9318 33376 9324
rect 33232 9104 33284 9110
rect 33232 9046 33284 9052
rect 33336 8838 33364 9318
rect 33520 9058 33548 9590
rect 33428 9030 33548 9058
rect 33324 8832 33376 8838
rect 33324 8774 33376 8780
rect 33046 8528 33102 8537
rect 33046 8463 33102 8472
rect 33324 8492 33376 8498
rect 33060 7954 33088 8463
rect 33324 8434 33376 8440
rect 33336 8090 33364 8434
rect 33428 8362 33456 9030
rect 33508 8968 33560 8974
rect 33508 8910 33560 8916
rect 33416 8356 33468 8362
rect 33416 8298 33468 8304
rect 33140 8084 33192 8090
rect 33140 8026 33192 8032
rect 33324 8084 33376 8090
rect 33324 8026 33376 8032
rect 33152 7954 33180 8026
rect 33048 7948 33100 7954
rect 33048 7890 33100 7896
rect 33140 7948 33192 7954
rect 33140 7890 33192 7896
rect 33520 7818 33548 8910
rect 33612 7886 33640 12582
rect 33784 12232 33836 12238
rect 33784 12174 33836 12180
rect 33796 11830 33824 12174
rect 33784 11824 33836 11830
rect 33784 11766 33836 11772
rect 33980 11762 34008 12582
rect 34256 12238 34284 13942
rect 34244 12232 34296 12238
rect 34244 12174 34296 12180
rect 33968 11756 34020 11762
rect 33968 11698 34020 11704
rect 34348 11082 34376 17206
rect 34888 17128 34940 17134
rect 34888 17070 34940 17076
rect 34796 15972 34848 15978
rect 34796 15914 34848 15920
rect 34520 15904 34572 15910
rect 34520 15846 34572 15852
rect 34532 15366 34560 15846
rect 34808 15502 34836 15914
rect 34796 15496 34848 15502
rect 34900 15473 34928 17070
rect 36004 16590 36032 17870
rect 44008 17338 44036 19200
rect 47823 17436 48131 17445
rect 47823 17434 47829 17436
rect 47885 17434 47909 17436
rect 47965 17434 47989 17436
rect 48045 17434 48069 17436
rect 48125 17434 48131 17436
rect 47885 17382 47887 17434
rect 48067 17382 48069 17434
rect 47823 17380 47829 17382
rect 47885 17380 47909 17382
rect 47965 17380 47989 17382
rect 48045 17380 48069 17382
rect 48125 17380 48131 17382
rect 47823 17371 48131 17380
rect 51920 17338 51948 19200
rect 59832 17338 59860 19200
rect 67744 17338 67772 19200
rect 69664 17536 69716 17542
rect 69664 17478 69716 17484
rect 43996 17332 44048 17338
rect 43996 17274 44048 17280
rect 50344 17332 50396 17338
rect 50344 17274 50396 17280
rect 51908 17332 51960 17338
rect 51908 17274 51960 17280
rect 59820 17332 59872 17338
rect 59820 17274 59872 17280
rect 67732 17332 67784 17338
rect 67732 17274 67784 17280
rect 44008 17202 44036 17274
rect 49516 17264 49568 17270
rect 49516 17206 49568 17212
rect 43996 17196 44048 17202
rect 43996 17138 44048 17144
rect 36912 17128 36964 17134
rect 36912 17070 36964 17076
rect 46204 17128 46256 17134
rect 46204 17070 46256 17076
rect 36105 16892 36413 16901
rect 36105 16890 36111 16892
rect 36167 16890 36191 16892
rect 36247 16890 36271 16892
rect 36327 16890 36351 16892
rect 36407 16890 36413 16892
rect 36167 16838 36169 16890
rect 36349 16838 36351 16890
rect 36105 16836 36111 16838
rect 36167 16836 36191 16838
rect 36247 16836 36271 16838
rect 36327 16836 36351 16838
rect 36407 16836 36413 16838
rect 36105 16827 36413 16836
rect 36924 16794 36952 17070
rect 38660 16992 38712 16998
rect 38660 16934 38712 16940
rect 40592 16992 40644 16998
rect 40592 16934 40644 16940
rect 46020 16992 46072 16998
rect 46020 16934 46072 16940
rect 38672 16794 38700 16934
rect 36912 16788 36964 16794
rect 36912 16730 36964 16736
rect 38660 16788 38712 16794
rect 38660 16730 38712 16736
rect 35992 16584 36044 16590
rect 35992 16526 36044 16532
rect 35808 15904 35860 15910
rect 35808 15846 35860 15852
rect 34980 15700 35032 15706
rect 34980 15642 35032 15648
rect 34796 15438 34848 15444
rect 34886 15464 34942 15473
rect 34520 15360 34572 15366
rect 34808 15348 34836 15438
rect 34886 15399 34942 15408
rect 34992 15366 35020 15642
rect 35346 15464 35402 15473
rect 35346 15399 35402 15408
rect 34980 15360 35032 15366
rect 34520 15302 34572 15308
rect 34702 15328 34758 15337
rect 34808 15320 34928 15348
rect 34702 15263 34758 15272
rect 34716 14958 34744 15263
rect 34796 15020 34848 15026
rect 34796 14962 34848 14968
rect 34704 14952 34756 14958
rect 34704 14894 34756 14900
rect 34520 11348 34572 11354
rect 34520 11290 34572 11296
rect 34336 11076 34388 11082
rect 34336 11018 34388 11024
rect 33692 10668 33744 10674
rect 33692 10610 33744 10616
rect 33704 10538 33732 10610
rect 33692 10532 33744 10538
rect 33692 10474 33744 10480
rect 33704 10266 33732 10474
rect 34348 10266 34376 11018
rect 34532 10606 34560 11290
rect 34808 11082 34836 14962
rect 34900 14414 34928 15320
rect 34980 15302 35032 15308
rect 34992 15026 35020 15302
rect 34980 15020 35032 15026
rect 34980 14962 35032 14968
rect 35072 14952 35124 14958
rect 35072 14894 35124 14900
rect 35084 14793 35112 14894
rect 35070 14784 35126 14793
rect 35070 14719 35126 14728
rect 35070 14512 35126 14521
rect 35070 14447 35126 14456
rect 34888 14408 34940 14414
rect 34888 14350 34940 14356
rect 35084 14278 35112 14447
rect 35072 14272 35124 14278
rect 35072 14214 35124 14220
rect 35072 13864 35124 13870
rect 35072 13806 35124 13812
rect 34980 12844 35032 12850
rect 34980 12786 35032 12792
rect 34992 12442 35020 12786
rect 34980 12436 35032 12442
rect 34980 12378 35032 12384
rect 34980 12096 35032 12102
rect 34980 12038 35032 12044
rect 34992 11762 35020 12038
rect 34980 11756 35032 11762
rect 34980 11698 35032 11704
rect 34796 11076 34848 11082
rect 34796 11018 34848 11024
rect 34520 10600 34572 10606
rect 34520 10542 34572 10548
rect 35084 10441 35112 13806
rect 35256 11144 35308 11150
rect 35256 11086 35308 11092
rect 35070 10432 35126 10441
rect 35070 10367 35126 10376
rect 33692 10260 33744 10266
rect 34336 10260 34388 10266
rect 33692 10202 33744 10208
rect 34256 10220 34336 10248
rect 33692 9648 33744 9654
rect 34256 9602 34284 10220
rect 34336 10202 34388 10208
rect 35084 10198 35112 10367
rect 35164 10260 35216 10266
rect 35164 10202 35216 10208
rect 35072 10192 35124 10198
rect 35072 10134 35124 10140
rect 35176 9994 35204 10202
rect 35164 9988 35216 9994
rect 35164 9930 35216 9936
rect 34612 9920 34664 9926
rect 34518 9888 34574 9897
rect 34612 9862 34664 9868
rect 34518 9823 34574 9832
rect 33744 9596 34284 9602
rect 33692 9590 34284 9596
rect 33704 9574 34284 9590
rect 34532 9518 34560 9823
rect 34520 9512 34572 9518
rect 34520 9454 34572 9460
rect 33690 9208 33746 9217
rect 33690 9143 33746 9152
rect 33704 8974 33732 9143
rect 33692 8968 33744 8974
rect 33692 8910 33744 8916
rect 33968 8968 34020 8974
rect 33968 8910 34020 8916
rect 34336 8968 34388 8974
rect 34336 8910 34388 8916
rect 34518 8936 34574 8945
rect 33876 8832 33928 8838
rect 33876 8774 33928 8780
rect 33888 8634 33916 8774
rect 33876 8628 33928 8634
rect 33876 8570 33928 8576
rect 33980 8430 34008 8910
rect 34152 8832 34204 8838
rect 34152 8774 34204 8780
rect 33876 8424 33928 8430
rect 33874 8392 33876 8401
rect 33968 8424 34020 8430
rect 33928 8392 33930 8401
rect 33968 8366 34020 8372
rect 33874 8327 33930 8336
rect 33600 7880 33652 7886
rect 33600 7822 33652 7828
rect 33508 7812 33560 7818
rect 33508 7754 33560 7760
rect 33138 7712 33194 7721
rect 33520 7698 33548 7754
rect 33520 7670 33640 7698
rect 33138 7647 33194 7656
rect 33152 7478 33180 7647
rect 33612 7478 33640 7670
rect 33140 7472 33192 7478
rect 33140 7414 33192 7420
rect 33600 7472 33652 7478
rect 33600 7414 33652 7420
rect 33140 6860 33192 6866
rect 33140 6802 33192 6808
rect 33416 6860 33468 6866
rect 33416 6802 33468 6808
rect 33048 6724 33100 6730
rect 33048 6666 33100 6672
rect 33060 6633 33088 6666
rect 33046 6624 33102 6633
rect 33046 6559 33102 6568
rect 33152 6390 33180 6802
rect 33324 6792 33376 6798
rect 33324 6734 33376 6740
rect 33336 6458 33364 6734
rect 33428 6662 33456 6802
rect 33416 6656 33468 6662
rect 33416 6598 33468 6604
rect 33324 6452 33376 6458
rect 33324 6394 33376 6400
rect 33140 6384 33192 6390
rect 33140 6326 33192 6332
rect 33232 6384 33284 6390
rect 33232 6326 33284 6332
rect 33244 5642 33272 6326
rect 33232 5636 33284 5642
rect 33232 5578 33284 5584
rect 33244 5302 33272 5578
rect 33232 5296 33284 5302
rect 33232 5238 33284 5244
rect 33428 5098 33456 6598
rect 33612 6390 33640 7414
rect 33784 7200 33836 7206
rect 33784 7142 33836 7148
rect 33876 7200 33928 7206
rect 33876 7142 33928 7148
rect 33796 6798 33824 7142
rect 33784 6792 33836 6798
rect 33784 6734 33836 6740
rect 33888 6730 33916 7142
rect 34060 6996 34112 7002
rect 34060 6938 34112 6944
rect 33876 6724 33928 6730
rect 33876 6666 33928 6672
rect 33600 6384 33652 6390
rect 33600 6326 33652 6332
rect 33888 6118 33916 6666
rect 33876 6112 33928 6118
rect 34072 6100 34100 6938
rect 34164 6934 34192 8774
rect 34348 8673 34376 8910
rect 34518 8871 34520 8880
rect 34572 8871 34574 8880
rect 34520 8842 34572 8848
rect 34334 8664 34390 8673
rect 34334 8599 34390 8608
rect 34520 8560 34572 8566
rect 34624 8548 34652 9862
rect 35268 9674 35296 11086
rect 35176 9646 35296 9674
rect 35360 9654 35388 15399
rect 35532 15360 35584 15366
rect 35820 15337 35848 15846
rect 36105 15804 36413 15813
rect 36105 15802 36111 15804
rect 36167 15802 36191 15804
rect 36247 15802 36271 15804
rect 36327 15802 36351 15804
rect 36407 15802 36413 15804
rect 36167 15750 36169 15802
rect 36349 15750 36351 15802
rect 36105 15748 36111 15750
rect 36167 15748 36191 15750
rect 36247 15748 36271 15750
rect 36327 15748 36351 15750
rect 36407 15748 36413 15750
rect 36105 15739 36413 15748
rect 35898 15600 35954 15609
rect 35898 15535 35954 15544
rect 35532 15302 35584 15308
rect 35806 15328 35862 15337
rect 35440 14272 35492 14278
rect 35440 14214 35492 14220
rect 35452 14006 35480 14214
rect 35440 14000 35492 14006
rect 35440 13942 35492 13948
rect 35440 13320 35492 13326
rect 35440 13262 35492 13268
rect 35452 12102 35480 13262
rect 35544 12889 35572 15302
rect 35806 15263 35862 15272
rect 35624 14000 35676 14006
rect 35624 13942 35676 13948
rect 35636 13705 35664 13942
rect 35622 13696 35678 13705
rect 35622 13631 35678 13640
rect 35912 13530 35940 15535
rect 37096 15496 37148 15502
rect 37096 15438 37148 15444
rect 36268 15360 36320 15366
rect 36268 15302 36320 15308
rect 36280 15094 36308 15302
rect 35992 15088 36044 15094
rect 35992 15030 36044 15036
rect 36268 15088 36320 15094
rect 36268 15030 36320 15036
rect 36004 14906 36032 15030
rect 36004 14878 36124 14906
rect 36096 14822 36124 14878
rect 35992 14816 36044 14822
rect 35992 14758 36044 14764
rect 36084 14816 36136 14822
rect 36084 14758 36136 14764
rect 36004 14618 36032 14758
rect 36105 14716 36413 14725
rect 36105 14714 36111 14716
rect 36167 14714 36191 14716
rect 36247 14714 36271 14716
rect 36327 14714 36351 14716
rect 36407 14714 36413 14716
rect 36167 14662 36169 14714
rect 36349 14662 36351 14714
rect 36105 14660 36111 14662
rect 36167 14660 36191 14662
rect 36247 14660 36271 14662
rect 36327 14660 36351 14662
rect 36407 14660 36413 14662
rect 36105 14651 36413 14660
rect 35992 14612 36044 14618
rect 35992 14554 36044 14560
rect 37108 14414 37136 15438
rect 37740 15360 37792 15366
rect 37740 15302 37792 15308
rect 38108 15360 38160 15366
rect 38108 15302 38160 15308
rect 37280 15020 37332 15026
rect 37332 14980 37412 15008
rect 37280 14962 37332 14968
rect 37384 14414 37412 14980
rect 37096 14408 37148 14414
rect 37096 14350 37148 14356
rect 37372 14408 37424 14414
rect 37372 14350 37424 14356
rect 37108 14249 37136 14350
rect 37094 14240 37150 14249
rect 37094 14175 37150 14184
rect 37384 14074 37412 14350
rect 37372 14068 37424 14074
rect 37372 14010 37424 14016
rect 36728 14000 36780 14006
rect 36728 13942 36780 13948
rect 35992 13728 36044 13734
rect 35992 13670 36044 13676
rect 36452 13728 36504 13734
rect 36740 13705 36768 13942
rect 37464 13932 37516 13938
rect 37464 13874 37516 13880
rect 37280 13864 37332 13870
rect 37280 13806 37332 13812
rect 36452 13670 36504 13676
rect 36726 13696 36782 13705
rect 35900 13524 35952 13530
rect 35900 13466 35952 13472
rect 36004 13394 36032 13670
rect 36105 13628 36413 13637
rect 36105 13626 36111 13628
rect 36167 13626 36191 13628
rect 36247 13626 36271 13628
rect 36327 13626 36351 13628
rect 36407 13626 36413 13628
rect 36167 13574 36169 13626
rect 36349 13574 36351 13626
rect 36105 13572 36111 13574
rect 36167 13572 36191 13574
rect 36247 13572 36271 13574
rect 36327 13572 36351 13574
rect 36407 13572 36413 13574
rect 36105 13563 36413 13572
rect 36464 13462 36492 13670
rect 36726 13631 36782 13640
rect 37292 13530 37320 13806
rect 37280 13524 37332 13530
rect 37280 13466 37332 13472
rect 36452 13456 36504 13462
rect 36452 13398 36504 13404
rect 36636 13456 36688 13462
rect 36636 13398 36688 13404
rect 35992 13388 36044 13394
rect 35992 13330 36044 13336
rect 36452 13320 36504 13326
rect 36452 13262 36504 13268
rect 35716 13252 35768 13258
rect 35716 13194 35768 13200
rect 35624 13184 35676 13190
rect 35624 13126 35676 13132
rect 35530 12880 35586 12889
rect 35530 12815 35532 12824
rect 35584 12815 35586 12824
rect 35532 12786 35584 12792
rect 35544 12755 35572 12786
rect 35636 12782 35664 13126
rect 35624 12776 35676 12782
rect 35624 12718 35676 12724
rect 35728 12594 35756 13194
rect 35636 12566 35756 12594
rect 35440 12096 35492 12102
rect 35440 12038 35492 12044
rect 35440 11688 35492 11694
rect 35440 11630 35492 11636
rect 35452 9674 35480 11630
rect 35636 11082 35664 12566
rect 36105 12540 36413 12549
rect 36105 12538 36111 12540
rect 36167 12538 36191 12540
rect 36247 12538 36271 12540
rect 36327 12538 36351 12540
rect 36407 12538 36413 12540
rect 36167 12486 36169 12538
rect 36349 12486 36351 12538
rect 36105 12484 36111 12486
rect 36167 12484 36191 12486
rect 36247 12484 36271 12486
rect 36327 12484 36351 12486
rect 36407 12484 36413 12486
rect 36105 12475 36413 12484
rect 36464 12442 36492 13262
rect 36452 12436 36504 12442
rect 36452 12378 36504 12384
rect 36360 11892 36412 11898
rect 36360 11834 36412 11840
rect 36372 11694 36400 11834
rect 36464 11762 36492 12378
rect 36648 12306 36676 13398
rect 37292 12782 37320 13466
rect 37476 13161 37504 13874
rect 37462 13152 37518 13161
rect 37462 13087 37518 13096
rect 37004 12776 37056 12782
rect 37004 12718 37056 12724
rect 37280 12776 37332 12782
rect 37280 12718 37332 12724
rect 36912 12640 36964 12646
rect 36912 12582 36964 12588
rect 36636 12300 36688 12306
rect 36636 12242 36688 12248
rect 36544 12164 36596 12170
rect 36544 12106 36596 12112
rect 36556 11898 36584 12106
rect 36544 11892 36596 11898
rect 36544 11834 36596 11840
rect 36648 11762 36676 12242
rect 36924 12209 36952 12582
rect 37016 12306 37044 12718
rect 37004 12300 37056 12306
rect 37004 12242 37056 12248
rect 37292 12238 37320 12718
rect 37280 12232 37332 12238
rect 36910 12200 36966 12209
rect 37280 12174 37332 12180
rect 36910 12135 36966 12144
rect 36728 12096 36780 12102
rect 36728 12038 36780 12044
rect 36740 11898 36768 12038
rect 36728 11892 36780 11898
rect 36728 11834 36780 11840
rect 36452 11756 36504 11762
rect 36452 11698 36504 11704
rect 36636 11756 36688 11762
rect 36636 11698 36688 11704
rect 36360 11688 36412 11694
rect 36360 11630 36412 11636
rect 35716 11552 35768 11558
rect 35714 11520 35716 11529
rect 35768 11520 35770 11529
rect 35714 11455 35770 11464
rect 36105 11452 36413 11461
rect 36105 11450 36111 11452
rect 36167 11450 36191 11452
rect 36247 11450 36271 11452
rect 36327 11450 36351 11452
rect 36407 11450 36413 11452
rect 36167 11398 36169 11450
rect 36349 11398 36351 11450
rect 36105 11396 36111 11398
rect 36167 11396 36191 11398
rect 36247 11396 36271 11398
rect 36327 11396 36351 11398
rect 36407 11396 36413 11398
rect 36105 11387 36413 11396
rect 36544 11212 36596 11218
rect 36820 11212 36872 11218
rect 36596 11172 36820 11200
rect 36544 11154 36596 11160
rect 36820 11154 36872 11160
rect 36924 11121 36952 12135
rect 37004 12096 37056 12102
rect 37004 12038 37056 12044
rect 37016 11665 37044 12038
rect 37188 11824 37240 11830
rect 37188 11766 37240 11772
rect 37002 11656 37058 11665
rect 37002 11591 37058 11600
rect 37200 11354 37228 11766
rect 37096 11348 37148 11354
rect 37096 11290 37148 11296
rect 37188 11348 37240 11354
rect 37188 11290 37240 11296
rect 36910 11112 36966 11121
rect 35624 11076 35676 11082
rect 36910 11047 36966 11056
rect 35624 11018 35676 11024
rect 35636 10742 35664 11018
rect 36542 10976 36598 10985
rect 36542 10911 36598 10920
rect 35624 10736 35676 10742
rect 35624 10678 35676 10684
rect 35716 10600 35768 10606
rect 35716 10542 35768 10548
rect 35728 10470 35756 10542
rect 35716 10464 35768 10470
rect 36556 10441 36584 10911
rect 36636 10668 36688 10674
rect 36636 10610 36688 10616
rect 35716 10406 35768 10412
rect 36542 10432 36598 10441
rect 36105 10364 36413 10373
rect 36542 10367 36598 10376
rect 36105 10362 36111 10364
rect 36167 10362 36191 10364
rect 36247 10362 36271 10364
rect 36327 10362 36351 10364
rect 36407 10362 36413 10364
rect 36167 10310 36169 10362
rect 36349 10310 36351 10362
rect 36105 10308 36111 10310
rect 36167 10308 36191 10310
rect 36247 10308 36271 10310
rect 36327 10308 36351 10310
rect 36407 10308 36413 10310
rect 36105 10299 36413 10308
rect 36544 10260 36596 10266
rect 36544 10202 36596 10208
rect 36452 10192 36504 10198
rect 36452 10134 36504 10140
rect 35716 10124 35768 10130
rect 35716 10066 35768 10072
rect 35728 9722 35756 10066
rect 35992 9920 36044 9926
rect 35992 9862 36044 9868
rect 35716 9716 35768 9722
rect 35348 9648 35400 9654
rect 34704 9444 34756 9450
rect 34704 9386 34756 9392
rect 34572 8520 34652 8548
rect 34520 8502 34572 8508
rect 34426 7848 34482 7857
rect 34532 7818 34560 8502
rect 34426 7783 34482 7792
rect 34520 7812 34572 7818
rect 34152 6928 34204 6934
rect 34152 6870 34204 6876
rect 34244 6724 34296 6730
rect 34244 6666 34296 6672
rect 34256 6186 34284 6666
rect 34244 6180 34296 6186
rect 34244 6122 34296 6128
rect 34152 6112 34204 6118
rect 34072 6072 34152 6100
rect 33876 6054 33928 6060
rect 34152 6054 34204 6060
rect 34256 5370 34284 6122
rect 34244 5364 34296 5370
rect 34244 5306 34296 5312
rect 33600 5296 33652 5302
rect 33600 5238 33652 5244
rect 33416 5092 33468 5098
rect 33416 5034 33468 5040
rect 33612 4758 33640 5238
rect 33600 4752 33652 4758
rect 34440 4729 34468 7783
rect 34520 7754 34572 7760
rect 34532 6730 34560 7754
rect 34716 7041 34744 9386
rect 35176 9382 35204 9646
rect 35452 9646 35664 9674
rect 36004 9674 36032 9862
rect 36464 9722 36492 10134
rect 36556 10062 36584 10202
rect 36544 10056 36596 10062
rect 36544 9998 36596 10004
rect 36648 9897 36676 10610
rect 36820 10532 36872 10538
rect 36820 10474 36872 10480
rect 36728 10056 36780 10062
rect 36832 10044 36860 10474
rect 36780 10016 36860 10044
rect 36728 9998 36780 10004
rect 36634 9888 36690 9897
rect 36634 9823 36690 9832
rect 36818 9752 36874 9761
rect 35716 9658 35768 9664
rect 35348 9590 35400 9596
rect 35164 9376 35216 9382
rect 34886 9344 34942 9353
rect 35216 9336 35296 9364
rect 35164 9318 35216 9324
rect 34886 9279 34942 9288
rect 34900 8838 34928 9279
rect 35070 9208 35126 9217
rect 35070 9143 35126 9152
rect 34888 8832 34940 8838
rect 34888 8774 34940 8780
rect 34888 7880 34940 7886
rect 34888 7822 34940 7828
rect 34702 7032 34758 7041
rect 34702 6967 34758 6976
rect 34900 6866 34928 7822
rect 34888 6860 34940 6866
rect 34888 6802 34940 6808
rect 34704 6792 34756 6798
rect 34704 6734 34756 6740
rect 34520 6724 34572 6730
rect 34520 6666 34572 6672
rect 34716 6497 34744 6734
rect 34888 6656 34940 6662
rect 34888 6598 34940 6604
rect 34702 6488 34758 6497
rect 34702 6423 34758 6432
rect 34716 6322 34744 6423
rect 34900 6390 34928 6598
rect 34888 6384 34940 6390
rect 34888 6326 34940 6332
rect 34704 6316 34756 6322
rect 34704 6258 34756 6264
rect 35084 5778 35112 9143
rect 35164 8900 35216 8906
rect 35164 8842 35216 8848
rect 35176 8809 35204 8842
rect 35162 8800 35218 8809
rect 35162 8735 35218 8744
rect 35162 7848 35218 7857
rect 35162 7783 35218 7792
rect 35176 7002 35204 7783
rect 35268 7002 35296 9336
rect 35164 6996 35216 7002
rect 35164 6938 35216 6944
rect 35256 6996 35308 7002
rect 35256 6938 35308 6944
rect 35360 6186 35388 9590
rect 35636 9450 35664 9646
rect 35820 9646 36032 9674
rect 36452 9716 36504 9722
rect 36818 9687 36874 9696
rect 36452 9658 36504 9664
rect 35532 9444 35584 9450
rect 35452 9404 35532 9432
rect 35452 9330 35480 9404
rect 35532 9386 35584 9392
rect 35624 9444 35676 9450
rect 35624 9386 35676 9392
rect 35452 9302 35572 9330
rect 35544 9024 35572 9302
rect 35714 9208 35770 9217
rect 35820 9194 35848 9646
rect 36832 9586 36860 9687
rect 36544 9580 36596 9586
rect 36544 9522 36596 9528
rect 36820 9580 36872 9586
rect 36820 9522 36872 9528
rect 36452 9512 36504 9518
rect 36096 9460 36452 9466
rect 36096 9454 36504 9460
rect 36096 9450 36492 9454
rect 36556 9450 36584 9522
rect 36084 9444 36492 9450
rect 36136 9438 36492 9444
rect 36544 9444 36596 9450
rect 36084 9386 36136 9392
rect 36544 9386 36596 9392
rect 36268 9376 36320 9382
rect 36320 9336 36492 9364
rect 36268 9318 36320 9324
rect 36105 9276 36413 9285
rect 36105 9274 36111 9276
rect 36167 9274 36191 9276
rect 36247 9274 36271 9276
rect 36327 9274 36351 9276
rect 36407 9274 36413 9276
rect 36167 9222 36169 9274
rect 36349 9222 36351 9274
rect 36105 9220 36111 9222
rect 36167 9220 36191 9222
rect 36247 9220 36271 9222
rect 36327 9220 36351 9222
rect 36407 9220 36413 9222
rect 36105 9211 36413 9220
rect 35770 9166 35848 9194
rect 35714 9143 35770 9152
rect 35544 8996 35756 9024
rect 35624 8900 35676 8906
rect 35624 8842 35676 8848
rect 35530 8800 35586 8809
rect 35530 8735 35586 8744
rect 35348 6180 35400 6186
rect 35348 6122 35400 6128
rect 35544 5846 35572 8735
rect 35636 7818 35664 8842
rect 35728 8786 35756 8996
rect 35728 8758 35848 8786
rect 35716 8628 35768 8634
rect 35716 8570 35768 8576
rect 35728 8090 35756 8570
rect 35820 8430 35848 8758
rect 36464 8634 36492 9336
rect 36832 8906 36860 9522
rect 36820 8900 36872 8906
rect 36820 8842 36872 8848
rect 36728 8832 36780 8838
rect 36728 8774 36780 8780
rect 36268 8628 36320 8634
rect 36268 8570 36320 8576
rect 36452 8628 36504 8634
rect 36452 8570 36504 8576
rect 35808 8424 35860 8430
rect 35808 8366 35860 8372
rect 36280 8294 36308 8570
rect 36360 8492 36412 8498
rect 36360 8434 36412 8440
rect 36372 8378 36400 8434
rect 36372 8350 36492 8378
rect 35808 8288 35860 8294
rect 35808 8230 35860 8236
rect 35900 8288 35952 8294
rect 35900 8230 35952 8236
rect 36268 8288 36320 8294
rect 36268 8230 36320 8236
rect 36464 8242 36492 8350
rect 36542 8256 36598 8265
rect 35820 8090 35848 8230
rect 35716 8084 35768 8090
rect 35716 8026 35768 8032
rect 35808 8084 35860 8090
rect 35808 8026 35860 8032
rect 35624 7812 35676 7818
rect 35624 7754 35676 7760
rect 35636 6730 35664 7754
rect 35912 7410 35940 8230
rect 36464 8214 36542 8242
rect 36105 8188 36413 8197
rect 36105 8186 36111 8188
rect 36167 8186 36191 8188
rect 36247 8186 36271 8188
rect 36327 8186 36351 8188
rect 36407 8186 36413 8188
rect 36167 8134 36169 8186
rect 36349 8134 36351 8186
rect 36105 8132 36111 8134
rect 36167 8132 36191 8134
rect 36247 8132 36271 8134
rect 36327 8132 36351 8134
rect 36407 8132 36413 8134
rect 36105 8123 36413 8132
rect 35808 7404 35860 7410
rect 35808 7346 35860 7352
rect 35900 7404 35952 7410
rect 35900 7346 35952 7352
rect 35820 7206 35848 7346
rect 35808 7200 35860 7206
rect 35808 7142 35860 7148
rect 36105 7100 36413 7109
rect 36105 7098 36111 7100
rect 36167 7098 36191 7100
rect 36247 7098 36271 7100
rect 36327 7098 36351 7100
rect 36407 7098 36413 7100
rect 36167 7046 36169 7098
rect 36349 7046 36351 7098
rect 36105 7044 36111 7046
rect 36167 7044 36191 7046
rect 36247 7044 36271 7046
rect 36327 7044 36351 7046
rect 36407 7044 36413 7046
rect 35898 7032 35954 7041
rect 36105 7035 36413 7044
rect 35898 6967 35954 6976
rect 35912 6916 35940 6967
rect 36176 6928 36228 6934
rect 35912 6888 36176 6916
rect 36176 6870 36228 6876
rect 35808 6860 35860 6866
rect 35808 6802 35860 6808
rect 35624 6724 35676 6730
rect 35624 6666 35676 6672
rect 35820 6361 35848 6802
rect 35806 6352 35862 6361
rect 35806 6287 35862 6296
rect 35900 6316 35952 6322
rect 35900 6258 35952 6264
rect 35624 6248 35676 6254
rect 35622 6216 35624 6225
rect 35676 6216 35678 6225
rect 35622 6151 35678 6160
rect 35532 5840 35584 5846
rect 35532 5782 35584 5788
rect 35912 5778 35940 6258
rect 36105 6012 36413 6021
rect 36105 6010 36111 6012
rect 36167 6010 36191 6012
rect 36247 6010 36271 6012
rect 36327 6010 36351 6012
rect 36407 6010 36413 6012
rect 36167 5958 36169 6010
rect 36349 5958 36351 6010
rect 36105 5956 36111 5958
rect 36167 5956 36191 5958
rect 36247 5956 36271 5958
rect 36327 5956 36351 5958
rect 36407 5956 36413 5958
rect 36105 5947 36413 5956
rect 36464 5778 36492 8214
rect 36542 8191 36598 8200
rect 36544 7744 36596 7750
rect 36544 7686 36596 7692
rect 36636 7744 36688 7750
rect 36636 7686 36688 7692
rect 36556 7546 36584 7686
rect 36544 7540 36596 7546
rect 36544 7482 36596 7488
rect 36648 7342 36676 7686
rect 36740 7410 36768 8774
rect 36728 7404 36780 7410
rect 36728 7346 36780 7352
rect 36636 7336 36688 7342
rect 36636 7278 36688 7284
rect 36544 7268 36596 7274
rect 36544 7210 36596 7216
rect 35072 5772 35124 5778
rect 35072 5714 35124 5720
rect 35900 5772 35952 5778
rect 35900 5714 35952 5720
rect 36452 5772 36504 5778
rect 36452 5714 36504 5720
rect 36556 5681 36584 7210
rect 36728 6656 36780 6662
rect 36726 6624 36728 6633
rect 36780 6624 36782 6633
rect 36726 6559 36782 6568
rect 36542 5672 36598 5681
rect 36542 5607 36598 5616
rect 36924 5386 36952 11047
rect 37108 10538 37136 11290
rect 37096 10532 37148 10538
rect 37096 10474 37148 10480
rect 37292 10470 37320 12174
rect 37476 11830 37504 13087
rect 37752 12850 37780 15302
rect 38014 13016 38070 13025
rect 38014 12951 38070 12960
rect 37740 12844 37792 12850
rect 37740 12786 37792 12792
rect 37464 11824 37516 11830
rect 37464 11766 37516 11772
rect 37752 11626 37780 12786
rect 37832 12436 37884 12442
rect 37832 12378 37884 12384
rect 37844 12345 37872 12378
rect 37830 12336 37886 12345
rect 37830 12271 37886 12280
rect 37740 11620 37792 11626
rect 37740 11562 37792 11568
rect 37464 11552 37516 11558
rect 37464 11494 37516 11500
rect 37476 11014 37504 11494
rect 38028 11218 38056 12951
rect 38120 11880 38148 15302
rect 38672 15026 38700 16730
rect 40132 16652 40184 16658
rect 40132 16594 40184 16600
rect 39580 16448 39632 16454
rect 39580 16390 39632 16396
rect 39592 16250 39620 16390
rect 39580 16244 39632 16250
rect 39580 16186 39632 16192
rect 39764 16176 39816 16182
rect 39764 16118 39816 16124
rect 38844 15904 38896 15910
rect 38844 15846 38896 15852
rect 38752 15564 38804 15570
rect 38752 15506 38804 15512
rect 38764 15162 38792 15506
rect 38752 15156 38804 15162
rect 38752 15098 38804 15104
rect 38660 15020 38712 15026
rect 38660 14962 38712 14968
rect 38856 14414 38884 15846
rect 39776 15706 39804 16118
rect 39764 15700 39816 15706
rect 39764 15642 39816 15648
rect 39304 15564 39356 15570
rect 39304 15506 39356 15512
rect 39316 15026 39344 15506
rect 39304 15020 39356 15026
rect 39304 14962 39356 14968
rect 40144 14414 40172 16594
rect 40316 16040 40368 16046
rect 40316 15982 40368 15988
rect 40328 15502 40356 15982
rect 40316 15496 40368 15502
rect 40368 15456 40448 15484
rect 40316 15438 40368 15444
rect 40420 15026 40448 15456
rect 40316 15020 40368 15026
rect 40316 14962 40368 14968
rect 40408 15020 40460 15026
rect 40408 14962 40460 14968
rect 40224 14816 40276 14822
rect 40224 14758 40276 14764
rect 38844 14408 38896 14414
rect 38844 14350 38896 14356
rect 40132 14408 40184 14414
rect 40132 14350 40184 14356
rect 38568 14340 38620 14346
rect 38568 14282 38620 14288
rect 38580 14006 38608 14282
rect 38568 14000 38620 14006
rect 38568 13942 38620 13948
rect 38476 13932 38528 13938
rect 38476 13874 38528 13880
rect 38200 13864 38252 13870
rect 38200 13806 38252 13812
rect 38212 12170 38240 13806
rect 38488 13530 38516 13874
rect 38660 13796 38712 13802
rect 38660 13738 38712 13744
rect 38476 13524 38528 13530
rect 38476 13466 38528 13472
rect 38488 13326 38516 13466
rect 38292 13320 38344 13326
rect 38292 13262 38344 13268
rect 38476 13320 38528 13326
rect 38476 13262 38528 13268
rect 38304 12434 38332 13262
rect 38672 12918 38700 13738
rect 38856 13734 38884 14350
rect 39120 14340 39172 14346
rect 39120 14282 39172 14288
rect 39132 14006 39160 14282
rect 40236 14006 40264 14758
rect 40328 14362 40356 14962
rect 40604 14521 40632 16934
rect 42340 16652 42392 16658
rect 42340 16594 42392 16600
rect 42432 16652 42484 16658
rect 42432 16594 42484 16600
rect 45836 16652 45888 16658
rect 45836 16594 45888 16600
rect 42352 16561 42380 16594
rect 42338 16552 42394 16561
rect 40776 16516 40828 16522
rect 40776 16458 40828 16464
rect 42260 16510 42338 16538
rect 40788 16182 40816 16458
rect 41604 16244 41656 16250
rect 41604 16186 41656 16192
rect 40776 16176 40828 16182
rect 40776 16118 40828 16124
rect 40868 16108 40920 16114
rect 40868 16050 40920 16056
rect 40776 16040 40828 16046
rect 40774 16008 40776 16017
rect 40828 16008 40830 16017
rect 40774 15943 40830 15952
rect 40774 15600 40830 15609
rect 40880 15586 40908 16050
rect 40960 16040 41012 16046
rect 40960 15982 41012 15988
rect 40830 15558 40908 15586
rect 40774 15535 40830 15544
rect 40788 15502 40816 15535
rect 40776 15496 40828 15502
rect 40776 15438 40828 15444
rect 40868 15496 40920 15502
rect 40868 15438 40920 15444
rect 40880 15366 40908 15438
rect 40868 15360 40920 15366
rect 40868 15302 40920 15308
rect 40972 14929 41000 15982
rect 41616 15434 41644 16186
rect 41880 15972 41932 15978
rect 41880 15914 41932 15920
rect 41892 15434 41920 15914
rect 41604 15428 41656 15434
rect 41604 15370 41656 15376
rect 41880 15428 41932 15434
rect 41880 15370 41932 15376
rect 41144 15360 41196 15366
rect 41144 15302 41196 15308
rect 41696 15360 41748 15366
rect 41696 15302 41748 15308
rect 40958 14920 41014 14929
rect 40958 14855 41014 14864
rect 40590 14512 40646 14521
rect 40590 14447 40592 14456
rect 40644 14447 40646 14456
rect 40684 14476 40736 14482
rect 40592 14418 40644 14424
rect 40684 14418 40736 14424
rect 40696 14362 40724 14418
rect 40328 14334 40724 14362
rect 39120 14000 39172 14006
rect 39120 13942 39172 13948
rect 40224 14000 40276 14006
rect 40224 13942 40276 13948
rect 38844 13728 38896 13734
rect 38844 13670 38896 13676
rect 40328 13326 40356 14334
rect 40500 14000 40552 14006
rect 40500 13942 40552 13948
rect 40316 13320 40368 13326
rect 40316 13262 40368 13268
rect 39396 13252 39448 13258
rect 39396 13194 39448 13200
rect 38660 12912 38712 12918
rect 38660 12854 38712 12860
rect 39408 12782 39436 13194
rect 39948 13184 40000 13190
rect 39948 13126 40000 13132
rect 40132 13184 40184 13190
rect 40132 13126 40184 13132
rect 39960 12850 39988 13126
rect 40144 12918 40172 13126
rect 40132 12912 40184 12918
rect 40132 12854 40184 12860
rect 39948 12844 40000 12850
rect 39948 12786 40000 12792
rect 39304 12776 39356 12782
rect 39304 12718 39356 12724
rect 39396 12776 39448 12782
rect 39396 12718 39448 12724
rect 39212 12640 39264 12646
rect 39212 12582 39264 12588
rect 39316 12594 39344 12718
rect 40040 12708 40092 12714
rect 40040 12650 40092 12656
rect 39026 12472 39082 12481
rect 38304 12406 38424 12434
rect 39026 12407 39082 12416
rect 38200 12164 38252 12170
rect 38200 12106 38252 12112
rect 38120 11852 38240 11880
rect 38212 11626 38240 11852
rect 38396 11694 38424 12406
rect 38934 12200 38990 12209
rect 38934 12135 38936 12144
rect 38988 12135 38990 12144
rect 38936 12106 38988 12112
rect 38658 11928 38714 11937
rect 38658 11863 38714 11872
rect 38384 11688 38436 11694
rect 38384 11630 38436 11636
rect 38200 11620 38252 11626
rect 38200 11562 38252 11568
rect 38292 11620 38344 11626
rect 38292 11562 38344 11568
rect 38304 11336 38332 11562
rect 38212 11308 38332 11336
rect 37556 11212 37608 11218
rect 37556 11154 37608 11160
rect 38016 11212 38068 11218
rect 38016 11154 38068 11160
rect 37372 11008 37424 11014
rect 37372 10950 37424 10956
rect 37464 11008 37516 11014
rect 37464 10950 37516 10956
rect 37384 10674 37412 10950
rect 37476 10810 37504 10950
rect 37568 10810 37596 11154
rect 38212 11082 38240 11308
rect 38396 11234 38424 11630
rect 38304 11218 38424 11234
rect 38672 11218 38700 11863
rect 39040 11830 39068 12407
rect 39224 12306 39252 12582
rect 39316 12566 39528 12594
rect 39500 12306 39528 12566
rect 39212 12300 39264 12306
rect 39212 12242 39264 12248
rect 39488 12300 39540 12306
rect 39488 12242 39540 12248
rect 38844 11824 38896 11830
rect 38844 11766 38896 11772
rect 39028 11824 39080 11830
rect 39028 11766 39080 11772
rect 38856 11665 38884 11766
rect 39580 11688 39632 11694
rect 38842 11656 38898 11665
rect 39580 11630 39632 11636
rect 39764 11688 39816 11694
rect 39764 11630 39816 11636
rect 38842 11591 38898 11600
rect 39592 11529 39620 11630
rect 39578 11520 39634 11529
rect 39578 11455 39634 11464
rect 38750 11384 38806 11393
rect 38750 11319 38806 11328
rect 39120 11348 39172 11354
rect 38292 11212 38424 11218
rect 38344 11206 38424 11212
rect 38660 11212 38712 11218
rect 38292 11154 38344 11160
rect 38660 11154 38712 11160
rect 38200 11076 38252 11082
rect 38200 11018 38252 11024
rect 38304 11014 38332 11154
rect 38292 11008 38344 11014
rect 38292 10950 38344 10956
rect 38384 11008 38436 11014
rect 38384 10950 38436 10956
rect 38396 10826 38424 10950
rect 37464 10804 37516 10810
rect 37464 10746 37516 10752
rect 37556 10804 37608 10810
rect 37556 10746 37608 10752
rect 38212 10798 38424 10826
rect 37738 10704 37794 10713
rect 37372 10668 37424 10674
rect 38212 10674 38240 10798
rect 37738 10639 37794 10648
rect 38200 10668 38252 10674
rect 37372 10610 37424 10616
rect 37384 10470 37412 10610
rect 37280 10464 37332 10470
rect 37280 10406 37332 10412
rect 37372 10464 37424 10470
rect 37372 10406 37424 10412
rect 37004 9648 37056 9654
rect 37004 9590 37056 9596
rect 37016 7002 37044 9590
rect 37188 8832 37240 8838
rect 37188 8774 37240 8780
rect 37094 8664 37150 8673
rect 37094 8599 37096 8608
rect 37148 8599 37150 8608
rect 37096 8570 37148 8576
rect 37200 8566 37228 8774
rect 37188 8560 37240 8566
rect 37188 8502 37240 8508
rect 37004 6996 37056 7002
rect 37004 6938 37056 6944
rect 37292 6866 37320 10406
rect 37752 9897 37780 10639
rect 38200 10610 38252 10616
rect 38292 10668 38344 10674
rect 38292 10610 38344 10616
rect 37738 9888 37794 9897
rect 37738 9823 37794 9832
rect 37752 9586 37780 9823
rect 38304 9602 38332 10610
rect 38568 10056 38620 10062
rect 38568 9998 38620 10004
rect 38384 9716 38436 9722
rect 38384 9658 38436 9664
rect 37464 9580 37516 9586
rect 37464 9522 37516 9528
rect 37740 9580 37792 9586
rect 37740 9522 37792 9528
rect 38212 9574 38332 9602
rect 37372 9512 37424 9518
rect 37372 9454 37424 9460
rect 37384 6934 37412 9454
rect 37476 8106 37504 9522
rect 37556 8968 37608 8974
rect 37556 8910 37608 8916
rect 37568 8566 37596 8910
rect 37556 8560 37608 8566
rect 37556 8502 37608 8508
rect 37568 8294 37596 8502
rect 37648 8492 37700 8498
rect 37648 8434 37700 8440
rect 37556 8288 37608 8294
rect 37556 8230 37608 8236
rect 37476 8078 37596 8106
rect 37464 7812 37516 7818
rect 37464 7754 37516 7760
rect 37372 6928 37424 6934
rect 37372 6870 37424 6876
rect 37280 6860 37332 6866
rect 37280 6802 37332 6808
rect 37476 5778 37504 7754
rect 37568 6361 37596 8078
rect 37660 7206 37688 8434
rect 37752 7886 37780 9522
rect 37924 9444 37976 9450
rect 37924 9386 37976 9392
rect 37832 8356 37884 8362
rect 37832 8298 37884 8304
rect 37844 8265 37872 8298
rect 37830 8256 37886 8265
rect 37830 8191 37886 8200
rect 37740 7880 37792 7886
rect 37740 7822 37792 7828
rect 37648 7200 37700 7206
rect 37648 7142 37700 7148
rect 37832 7200 37884 7206
rect 37832 7142 37884 7148
rect 37844 7002 37872 7142
rect 37832 6996 37884 7002
rect 37832 6938 37884 6944
rect 37554 6352 37610 6361
rect 37554 6287 37610 6296
rect 37936 6254 37964 9386
rect 38212 9382 38240 9574
rect 38396 9382 38424 9658
rect 38580 9518 38608 9998
rect 38568 9512 38620 9518
rect 38568 9454 38620 9460
rect 38200 9376 38252 9382
rect 38384 9376 38436 9382
rect 38200 9318 38252 9324
rect 38304 9336 38384 9364
rect 38108 8968 38160 8974
rect 38108 8910 38160 8916
rect 38120 8537 38148 8910
rect 38106 8528 38162 8537
rect 38028 8486 38106 8514
rect 38028 6934 38056 8486
rect 38106 8463 38162 8472
rect 38108 7404 38160 7410
rect 38108 7346 38160 7352
rect 38016 6928 38068 6934
rect 38120 6905 38148 7346
rect 38016 6870 38068 6876
rect 38106 6896 38162 6905
rect 38028 6780 38056 6870
rect 38106 6831 38162 6840
rect 38028 6752 38148 6780
rect 38016 6316 38068 6322
rect 38016 6258 38068 6264
rect 37924 6248 37976 6254
rect 37924 6190 37976 6196
rect 37464 5772 37516 5778
rect 37464 5714 37516 5720
rect 37476 5642 37504 5714
rect 38028 5710 38056 6258
rect 38120 5846 38148 6752
rect 38108 5840 38160 5846
rect 38108 5782 38160 5788
rect 38016 5704 38068 5710
rect 38016 5646 38068 5652
rect 37464 5636 37516 5642
rect 37464 5578 37516 5584
rect 36740 5358 36952 5386
rect 37924 5364 37976 5370
rect 36740 5250 36768 5358
rect 37924 5306 37976 5312
rect 36464 5234 36768 5250
rect 36452 5228 36780 5234
rect 36504 5222 36728 5228
rect 36452 5170 36504 5176
rect 36728 5170 36780 5176
rect 36740 5139 36768 5170
rect 36912 5160 36964 5166
rect 36912 5102 36964 5108
rect 34888 5024 34940 5030
rect 34888 4966 34940 4972
rect 34900 4826 34928 4966
rect 36105 4924 36413 4933
rect 36105 4922 36111 4924
rect 36167 4922 36191 4924
rect 36247 4922 36271 4924
rect 36327 4922 36351 4924
rect 36407 4922 36413 4924
rect 36167 4870 36169 4922
rect 36349 4870 36351 4922
rect 36105 4868 36111 4870
rect 36167 4868 36191 4870
rect 36247 4868 36271 4870
rect 36327 4868 36351 4870
rect 36407 4868 36413 4870
rect 36105 4859 36413 4868
rect 34888 4820 34940 4826
rect 34888 4762 34940 4768
rect 33600 4694 33652 4700
rect 34426 4720 34482 4729
rect 33416 4684 33468 4690
rect 34426 4655 34482 4664
rect 33416 4626 33468 4632
rect 33428 4214 33456 4626
rect 36924 4554 36952 5102
rect 37740 4820 37792 4826
rect 37740 4762 37792 4768
rect 35348 4548 35400 4554
rect 35348 4490 35400 4496
rect 36912 4548 36964 4554
rect 36912 4490 36964 4496
rect 33600 4480 33652 4486
rect 33600 4422 33652 4428
rect 34612 4480 34664 4486
rect 34612 4422 34664 4428
rect 33612 4214 33640 4422
rect 33416 4208 33468 4214
rect 33416 4150 33468 4156
rect 33600 4208 33652 4214
rect 33600 4150 33652 4156
rect 34624 4146 34652 4422
rect 35360 4282 35388 4490
rect 35348 4276 35400 4282
rect 35348 4218 35400 4224
rect 34612 4140 34664 4146
rect 34612 4082 34664 4088
rect 37752 4078 37780 4762
rect 37936 4554 37964 5306
rect 38016 5228 38068 5234
rect 38016 5170 38068 5176
rect 37924 4548 37976 4554
rect 37924 4490 37976 4496
rect 37464 4072 37516 4078
rect 37464 4014 37516 4020
rect 37740 4072 37792 4078
rect 37740 4014 37792 4020
rect 36105 3836 36413 3845
rect 36105 3834 36111 3836
rect 36167 3834 36191 3836
rect 36247 3834 36271 3836
rect 36327 3834 36351 3836
rect 36407 3834 36413 3836
rect 36167 3782 36169 3834
rect 36349 3782 36351 3834
rect 36105 3780 36111 3782
rect 36167 3780 36191 3782
rect 36247 3780 36271 3782
rect 36327 3780 36351 3782
rect 36407 3780 36413 3782
rect 36105 3771 36413 3780
rect 32956 3664 33008 3670
rect 32956 3606 33008 3612
rect 37476 3602 37504 4014
rect 37464 3596 37516 3602
rect 37464 3538 37516 3544
rect 37476 2774 37504 3538
rect 37752 3194 37780 4014
rect 37936 3942 37964 4490
rect 38028 4486 38056 5170
rect 38212 4593 38240 9318
rect 38304 7206 38332 9336
rect 38384 9318 38436 9324
rect 38474 9072 38530 9081
rect 38474 9007 38530 9016
rect 38384 8968 38436 8974
rect 38384 8910 38436 8916
rect 38396 8634 38424 8910
rect 38384 8628 38436 8634
rect 38384 8570 38436 8576
rect 38292 7200 38344 7206
rect 38292 7142 38344 7148
rect 38488 6866 38516 9007
rect 38672 8922 38700 11154
rect 38764 10674 38792 11319
rect 39120 11290 39172 11296
rect 38844 11144 38896 11150
rect 38844 11086 38896 11092
rect 38856 10674 38884 11086
rect 38752 10668 38804 10674
rect 38752 10610 38804 10616
rect 38844 10668 38896 10674
rect 38844 10610 38896 10616
rect 39028 9648 39080 9654
rect 39028 9590 39080 9596
rect 38752 9580 38804 9586
rect 38752 9522 38804 9528
rect 38764 9081 38792 9522
rect 38936 9512 38988 9518
rect 38936 9454 38988 9460
rect 38948 9382 38976 9454
rect 38936 9376 38988 9382
rect 38842 9344 38898 9353
rect 38936 9318 38988 9324
rect 38842 9279 38898 9288
rect 38856 9110 38884 9279
rect 38844 9104 38896 9110
rect 38750 9072 38806 9081
rect 38844 9046 38896 9052
rect 38934 9072 38990 9081
rect 38750 9007 38806 9016
rect 38934 9007 38990 9016
rect 38842 8936 38898 8945
rect 38672 8894 38792 8922
rect 38660 8832 38712 8838
rect 38660 8774 38712 8780
rect 38672 8498 38700 8774
rect 38660 8492 38712 8498
rect 38660 8434 38712 8440
rect 38764 8294 38792 8894
rect 38842 8871 38898 8880
rect 38856 8838 38884 8871
rect 38844 8832 38896 8838
rect 38844 8774 38896 8780
rect 38752 8288 38804 8294
rect 38752 8230 38804 8236
rect 38844 7404 38896 7410
rect 38844 7346 38896 7352
rect 38856 7206 38884 7346
rect 38844 7200 38896 7206
rect 38844 7142 38896 7148
rect 38856 6866 38884 7142
rect 38476 6860 38528 6866
rect 38476 6802 38528 6808
rect 38844 6860 38896 6866
rect 38844 6802 38896 6808
rect 38568 6316 38620 6322
rect 38568 6258 38620 6264
rect 38580 6225 38608 6258
rect 38566 6216 38622 6225
rect 38566 6151 38622 6160
rect 38856 5846 38884 6802
rect 38948 6662 38976 9007
rect 39040 8974 39068 9590
rect 39028 8968 39080 8974
rect 39028 8910 39080 8916
rect 39132 7750 39160 11290
rect 39776 11150 39804 11630
rect 39764 11144 39816 11150
rect 39764 11086 39816 11092
rect 39776 11014 39804 11086
rect 39764 11008 39816 11014
rect 39764 10950 39816 10956
rect 40052 10674 40080 12650
rect 40512 12442 40540 13942
rect 40972 13938 41000 14855
rect 40960 13932 41012 13938
rect 40960 13874 41012 13880
rect 40590 12608 40646 12617
rect 40590 12543 40646 12552
rect 40500 12436 40552 12442
rect 40500 12378 40552 12384
rect 40604 11830 40632 12543
rect 40592 11824 40644 11830
rect 40592 11766 40644 11772
rect 40224 11756 40276 11762
rect 40224 11698 40276 11704
rect 40236 11529 40264 11698
rect 40222 11520 40278 11529
rect 40222 11455 40278 11464
rect 40500 11144 40552 11150
rect 40130 11112 40186 11121
rect 40500 11086 40552 11092
rect 40130 11047 40186 11056
rect 40144 10742 40172 11047
rect 40512 10985 40540 11086
rect 40498 10976 40554 10985
rect 40498 10911 40554 10920
rect 41156 10742 41184 15302
rect 41328 14952 41380 14958
rect 41328 14894 41380 14900
rect 41236 14884 41288 14890
rect 41236 14826 41288 14832
rect 41248 14657 41276 14826
rect 41234 14648 41290 14657
rect 41234 14583 41290 14592
rect 41340 14482 41368 14894
rect 41604 14816 41656 14822
rect 41604 14758 41656 14764
rect 41328 14476 41380 14482
rect 41328 14418 41380 14424
rect 41616 14346 41644 14758
rect 41604 14340 41656 14346
rect 41604 14282 41656 14288
rect 41418 14240 41474 14249
rect 41418 14175 41474 14184
rect 41432 14074 41460 14175
rect 41420 14068 41472 14074
rect 41420 14010 41472 14016
rect 41708 12850 41736 15302
rect 41880 14544 41932 14550
rect 41880 14486 41932 14492
rect 41892 14278 41920 14486
rect 41880 14272 41932 14278
rect 41880 14214 41932 14220
rect 42260 14113 42288 16510
rect 42338 16487 42394 16496
rect 42340 15360 42392 15366
rect 42340 15302 42392 15308
rect 42246 14104 42302 14113
rect 42246 14039 42302 14048
rect 41788 13932 41840 13938
rect 41788 13874 41840 13880
rect 41800 13161 41828 13874
rect 42260 13734 42288 14039
rect 42248 13728 42300 13734
rect 42248 13670 42300 13676
rect 41786 13152 41842 13161
rect 41786 13087 41842 13096
rect 41696 12844 41748 12850
rect 41696 12786 41748 12792
rect 42352 12782 42380 15302
rect 42444 15065 42472 16594
rect 43720 16448 43772 16454
rect 43720 16390 43772 16396
rect 44824 16448 44876 16454
rect 44824 16390 44876 16396
rect 42800 16108 42852 16114
rect 42800 16050 42852 16056
rect 42430 15056 42486 15065
rect 42430 14991 42486 15000
rect 42444 13938 42472 14991
rect 42708 14952 42760 14958
rect 42708 14894 42760 14900
rect 42720 14822 42748 14894
rect 42708 14816 42760 14822
rect 42708 14758 42760 14764
rect 42720 14618 42748 14758
rect 42708 14612 42760 14618
rect 42708 14554 42760 14560
rect 42708 14272 42760 14278
rect 42708 14214 42760 14220
rect 42432 13932 42484 13938
rect 42432 13874 42484 13880
rect 42432 13524 42484 13530
rect 42432 13466 42484 13472
rect 42444 13326 42472 13466
rect 42524 13456 42576 13462
rect 42524 13398 42576 13404
rect 42432 13320 42484 13326
rect 42432 13262 42484 13268
rect 41604 12776 41656 12782
rect 41604 12718 41656 12724
rect 42340 12776 42392 12782
rect 42340 12718 42392 12724
rect 41616 12073 41644 12718
rect 41696 12640 41748 12646
rect 41696 12582 41748 12588
rect 41788 12640 41840 12646
rect 41788 12582 41840 12588
rect 41602 12064 41658 12073
rect 41602 11999 41658 12008
rect 41420 11756 41472 11762
rect 41420 11698 41472 11704
rect 41432 11665 41460 11698
rect 41604 11688 41656 11694
rect 41418 11656 41474 11665
rect 41604 11630 41656 11636
rect 41418 11591 41474 11600
rect 40132 10736 40184 10742
rect 40132 10678 40184 10684
rect 41144 10736 41196 10742
rect 41144 10678 41196 10684
rect 40040 10668 40092 10674
rect 40040 10610 40092 10616
rect 39672 10600 39724 10606
rect 39672 10542 39724 10548
rect 39764 10600 39816 10606
rect 39764 10542 39816 10548
rect 39302 9752 39358 9761
rect 39302 9687 39358 9696
rect 39316 9042 39344 9687
rect 39396 9512 39448 9518
rect 39396 9454 39448 9460
rect 39304 9036 39356 9042
rect 39304 8978 39356 8984
rect 39120 7744 39172 7750
rect 39120 7686 39172 7692
rect 39028 7336 39080 7342
rect 39028 7278 39080 7284
rect 39040 7002 39068 7278
rect 39408 7274 39436 9454
rect 39684 9081 39712 10542
rect 39776 9994 39804 10542
rect 41142 10296 41198 10305
rect 41142 10231 41198 10240
rect 40224 10192 40276 10198
rect 40224 10134 40276 10140
rect 39948 10056 40000 10062
rect 40236 10010 40264 10134
rect 41156 10062 41184 10231
rect 39948 9998 40000 10004
rect 39764 9988 39816 9994
rect 39764 9930 39816 9936
rect 39856 9920 39908 9926
rect 39856 9862 39908 9868
rect 39960 9874 39988 9998
rect 40144 9982 40264 10010
rect 40316 10056 40368 10062
rect 40316 9998 40368 10004
rect 41144 10056 41196 10062
rect 41144 9998 41196 10004
rect 40144 9874 40172 9982
rect 40328 9926 40356 9998
rect 40592 9988 40644 9994
rect 40592 9930 40644 9936
rect 39670 9072 39726 9081
rect 39670 9007 39726 9016
rect 39764 9036 39816 9042
rect 39764 8978 39816 8984
rect 39776 8362 39804 8978
rect 39764 8356 39816 8362
rect 39764 8298 39816 8304
rect 39868 7546 39896 9862
rect 39960 9846 40172 9874
rect 40224 9920 40276 9926
rect 40224 9862 40276 9868
rect 40316 9920 40368 9926
rect 40316 9862 40368 9868
rect 40236 9722 40264 9862
rect 40224 9716 40276 9722
rect 40224 9658 40276 9664
rect 40222 9480 40278 9489
rect 40040 9444 40092 9450
rect 40222 9415 40224 9424
rect 40040 9386 40092 9392
rect 40276 9415 40278 9424
rect 40224 9386 40276 9392
rect 40052 8022 40080 9386
rect 40328 8498 40356 9862
rect 40604 9654 40632 9930
rect 41156 9897 41184 9998
rect 41236 9988 41288 9994
rect 41236 9930 41288 9936
rect 41142 9888 41198 9897
rect 41248 9874 41276 9930
rect 41326 9888 41382 9897
rect 41248 9846 41326 9874
rect 41142 9823 41198 9832
rect 41326 9823 41382 9832
rect 40592 9648 40644 9654
rect 40592 9590 40644 9596
rect 41052 9512 41104 9518
rect 41236 9512 41288 9518
rect 41052 9454 41104 9460
rect 41234 9480 41236 9489
rect 41288 9480 41290 9489
rect 40500 8968 40552 8974
rect 40500 8910 40552 8916
rect 40684 8968 40736 8974
rect 40684 8910 40736 8916
rect 40512 8673 40540 8910
rect 40498 8664 40554 8673
rect 40498 8599 40554 8608
rect 40512 8498 40540 8599
rect 40316 8492 40368 8498
rect 40316 8434 40368 8440
rect 40500 8492 40552 8498
rect 40500 8434 40552 8440
rect 40696 8430 40724 8910
rect 40960 8832 41012 8838
rect 40960 8774 41012 8780
rect 40774 8528 40830 8537
rect 40774 8463 40776 8472
rect 40828 8463 40830 8472
rect 40776 8434 40828 8440
rect 40408 8424 40460 8430
rect 40408 8366 40460 8372
rect 40684 8424 40736 8430
rect 40684 8366 40736 8372
rect 40420 8129 40448 8366
rect 40696 8294 40724 8366
rect 40684 8288 40736 8294
rect 40684 8230 40736 8236
rect 40406 8120 40462 8129
rect 40406 8055 40462 8064
rect 40696 8022 40724 8230
rect 40040 8016 40092 8022
rect 40040 7958 40092 7964
rect 40684 8016 40736 8022
rect 40684 7958 40736 7964
rect 40132 7948 40184 7954
rect 40132 7890 40184 7896
rect 40776 7948 40828 7954
rect 40776 7890 40828 7896
rect 40040 7880 40092 7886
rect 40040 7822 40092 7828
rect 39856 7540 39908 7546
rect 39856 7482 39908 7488
rect 39396 7268 39448 7274
rect 39396 7210 39448 7216
rect 39868 7206 39896 7482
rect 39856 7200 39908 7206
rect 39856 7142 39908 7148
rect 39028 6996 39080 7002
rect 39028 6938 39080 6944
rect 40052 6866 40080 7822
rect 40144 7410 40172 7890
rect 40132 7404 40184 7410
rect 40132 7346 40184 7352
rect 40592 7336 40644 7342
rect 40592 7278 40644 7284
rect 40132 7268 40184 7274
rect 40132 7210 40184 7216
rect 40040 6860 40092 6866
rect 40040 6802 40092 6808
rect 39028 6792 39080 6798
rect 39028 6734 39080 6740
rect 38936 6656 38988 6662
rect 38936 6598 38988 6604
rect 39040 6254 39068 6734
rect 39304 6656 39356 6662
rect 39304 6598 39356 6604
rect 39316 6458 39344 6598
rect 39304 6452 39356 6458
rect 39304 6394 39356 6400
rect 39028 6248 39080 6254
rect 39028 6190 39080 6196
rect 39040 5846 39068 6190
rect 38844 5840 38896 5846
rect 38844 5782 38896 5788
rect 39028 5840 39080 5846
rect 39028 5782 39080 5788
rect 39040 4758 39068 5782
rect 40052 5370 40080 6802
rect 40144 6322 40172 7210
rect 40604 7177 40632 7278
rect 40590 7168 40646 7177
rect 40590 7103 40646 7112
rect 40788 7002 40816 7890
rect 40972 7818 41000 8774
rect 41064 8498 41092 9454
rect 41234 9415 41290 9424
rect 41234 9208 41290 9217
rect 41234 9143 41236 9152
rect 41288 9143 41290 9152
rect 41328 9172 41380 9178
rect 41236 9114 41288 9120
rect 41328 9114 41380 9120
rect 41340 8566 41368 9114
rect 41432 8838 41460 11591
rect 41616 11393 41644 11630
rect 41602 11384 41658 11393
rect 41708 11370 41736 12582
rect 41800 12170 41828 12582
rect 42352 12345 42380 12718
rect 42338 12336 42394 12345
rect 42338 12271 42394 12280
rect 42536 12238 42564 13398
rect 42616 12436 42668 12442
rect 42616 12378 42668 12384
rect 42628 12238 42656 12378
rect 42720 12306 42748 14214
rect 42812 13938 42840 16050
rect 42892 15904 42944 15910
rect 42892 15846 42944 15852
rect 42800 13932 42852 13938
rect 42800 13874 42852 13880
rect 42904 13297 42932 15846
rect 43732 15502 43760 16390
rect 44836 16250 44864 16390
rect 44824 16244 44876 16250
rect 44824 16186 44876 16192
rect 44638 16144 44694 16153
rect 44272 16108 44324 16114
rect 44638 16079 44694 16088
rect 44272 16050 44324 16056
rect 44284 15910 44312 16050
rect 44364 16040 44416 16046
rect 44364 15982 44416 15988
rect 43812 15904 43864 15910
rect 43812 15846 43864 15852
rect 44272 15904 44324 15910
rect 44272 15846 44324 15852
rect 43720 15496 43772 15502
rect 43720 15438 43772 15444
rect 43076 15428 43128 15434
rect 43076 15370 43128 15376
rect 42890 13288 42946 13297
rect 42890 13223 42892 13232
rect 42944 13223 42946 13232
rect 42892 13194 42944 13200
rect 42904 13163 42932 13194
rect 43088 12850 43116 15370
rect 43444 15020 43496 15026
rect 43444 14962 43496 14968
rect 43168 13252 43220 13258
rect 43168 13194 43220 13200
rect 43076 12844 43128 12850
rect 43076 12786 43128 12792
rect 42892 12776 42944 12782
rect 42892 12718 42944 12724
rect 42708 12300 42760 12306
rect 42708 12242 42760 12248
rect 42524 12232 42576 12238
rect 42524 12174 42576 12180
rect 42616 12232 42668 12238
rect 42616 12174 42668 12180
rect 41788 12164 41840 12170
rect 41788 12106 41840 12112
rect 41972 11892 42024 11898
rect 41972 11834 42024 11840
rect 41984 11558 42012 11834
rect 41972 11552 42024 11558
rect 41972 11494 42024 11500
rect 41786 11384 41842 11393
rect 41708 11354 41786 11370
rect 41602 11319 41658 11328
rect 41696 11348 41786 11354
rect 41748 11342 41786 11348
rect 41984 11354 42012 11494
rect 41786 11319 41842 11328
rect 41972 11348 42024 11354
rect 41696 11290 41748 11296
rect 41708 11259 41736 11290
rect 41800 11150 41828 11319
rect 41972 11290 42024 11296
rect 41788 11144 41840 11150
rect 41788 11086 41840 11092
rect 41984 11082 42012 11290
rect 42156 11144 42208 11150
rect 42156 11086 42208 11092
rect 41972 11076 42024 11082
rect 41972 11018 42024 11024
rect 42168 10985 42196 11086
rect 42154 10976 42210 10985
rect 42154 10911 42210 10920
rect 41786 10840 41842 10849
rect 41786 10775 41842 10784
rect 41604 10736 41656 10742
rect 41524 10696 41604 10724
rect 41524 9586 41552 10696
rect 41604 10678 41656 10684
rect 41800 10198 41828 10775
rect 41880 10600 41932 10606
rect 41880 10542 41932 10548
rect 41892 10470 41920 10542
rect 41880 10464 41932 10470
rect 41880 10406 41932 10412
rect 41972 10464 42024 10470
rect 41972 10406 42024 10412
rect 41880 10260 41932 10266
rect 41880 10202 41932 10208
rect 41788 10192 41840 10198
rect 41788 10134 41840 10140
rect 41788 9988 41840 9994
rect 41788 9930 41840 9936
rect 41800 9722 41828 9930
rect 41788 9716 41840 9722
rect 41788 9658 41840 9664
rect 41512 9580 41564 9586
rect 41512 9522 41564 9528
rect 41524 9110 41552 9522
rect 41800 9382 41828 9658
rect 41892 9654 41920 10202
rect 41984 10062 42012 10406
rect 42062 10296 42118 10305
rect 42062 10231 42064 10240
rect 42116 10231 42118 10240
rect 42064 10202 42116 10208
rect 41972 10056 42024 10062
rect 41972 9998 42024 10004
rect 41984 9926 42012 9998
rect 41972 9920 42024 9926
rect 41972 9862 42024 9868
rect 41880 9648 41932 9654
rect 41880 9590 41932 9596
rect 42168 9586 42196 10911
rect 42536 10810 42564 12174
rect 42616 11892 42668 11898
rect 42616 11834 42668 11840
rect 42628 11801 42656 11834
rect 42614 11792 42670 11801
rect 42614 11727 42670 11736
rect 42904 11694 42932 12718
rect 43180 12714 43208 13194
rect 43168 12708 43220 12714
rect 43168 12650 43220 12656
rect 43260 12708 43312 12714
rect 43260 12650 43312 12656
rect 42892 11688 42944 11694
rect 42892 11630 42944 11636
rect 42890 11520 42946 11529
rect 42890 11455 42946 11464
rect 42904 11354 42932 11455
rect 42892 11348 42944 11354
rect 42892 11290 42944 11296
rect 42800 11076 42852 11082
rect 42800 11018 42852 11024
rect 42708 11008 42760 11014
rect 42708 10950 42760 10956
rect 42524 10804 42576 10810
rect 42524 10746 42576 10752
rect 42432 10668 42484 10674
rect 42432 10610 42484 10616
rect 42444 10198 42472 10610
rect 42720 10606 42748 10950
rect 42812 10674 42840 11018
rect 42800 10668 42852 10674
rect 42800 10610 42852 10616
rect 42904 10606 42932 11290
rect 43272 10606 43300 12650
rect 43456 12442 43484 14962
rect 43824 14657 43852 15846
rect 44086 15736 44142 15745
rect 44086 15671 44142 15680
rect 43810 14648 43866 14657
rect 43810 14583 43866 14592
rect 43824 14414 43852 14583
rect 43812 14408 43864 14414
rect 43812 14350 43864 14356
rect 44100 14006 44128 15671
rect 44284 15638 44312 15846
rect 44376 15706 44404 15982
rect 44364 15700 44416 15706
rect 44364 15642 44416 15648
rect 44272 15632 44324 15638
rect 44272 15574 44324 15580
rect 44088 14000 44140 14006
rect 44088 13942 44140 13948
rect 43996 12844 44048 12850
rect 43996 12786 44048 12792
rect 44272 12844 44324 12850
rect 44272 12786 44324 12792
rect 44008 12646 44036 12786
rect 43904 12640 43956 12646
rect 43904 12582 43956 12588
rect 43996 12640 44048 12646
rect 43996 12582 44048 12588
rect 43444 12436 43496 12442
rect 43444 12378 43496 12384
rect 43812 12232 43864 12238
rect 43812 12174 43864 12180
rect 43720 12096 43772 12102
rect 43720 12038 43772 12044
rect 43732 11898 43760 12038
rect 43720 11892 43772 11898
rect 43720 11834 43772 11840
rect 43824 11150 43852 12174
rect 43916 12073 43944 12582
rect 43996 12232 44048 12238
rect 43996 12174 44048 12180
rect 43902 12064 43958 12073
rect 43902 11999 43958 12008
rect 43916 11354 43944 11999
rect 44008 11393 44036 12174
rect 44088 11824 44140 11830
rect 44088 11766 44140 11772
rect 44100 11694 44128 11766
rect 44088 11688 44140 11694
rect 44088 11630 44140 11636
rect 43994 11384 44050 11393
rect 43904 11348 43956 11354
rect 43994 11319 44050 11328
rect 43904 11290 43956 11296
rect 44008 11218 44036 11319
rect 43996 11212 44048 11218
rect 43996 11154 44048 11160
rect 43812 11144 43864 11150
rect 43812 11086 43864 11092
rect 44284 10810 44312 12786
rect 44546 12200 44602 12209
rect 44546 12135 44548 12144
rect 44600 12135 44602 12144
rect 44548 12106 44600 12112
rect 44364 11892 44416 11898
rect 44416 11852 44496 11880
rect 44364 11834 44416 11840
rect 44364 11688 44416 11694
rect 44364 11630 44416 11636
rect 44272 10804 44324 10810
rect 44272 10746 44324 10752
rect 42708 10600 42760 10606
rect 42708 10542 42760 10548
rect 42892 10600 42944 10606
rect 42892 10542 42944 10548
rect 43260 10600 43312 10606
rect 43260 10542 43312 10548
rect 43904 10600 43956 10606
rect 43904 10542 43956 10548
rect 43916 10266 43944 10542
rect 44376 10305 44404 11630
rect 44468 11286 44496 11852
rect 44456 11280 44508 11286
rect 44456 11222 44508 11228
rect 44652 11218 44680 16079
rect 45468 15904 45520 15910
rect 45468 15846 45520 15852
rect 45480 15706 45508 15846
rect 45468 15700 45520 15706
rect 45468 15642 45520 15648
rect 45744 15496 45796 15502
rect 45744 15438 45796 15444
rect 45652 15360 45704 15366
rect 45652 15302 45704 15308
rect 44732 14816 44784 14822
rect 44732 14758 44784 14764
rect 44744 13190 44772 14758
rect 45468 14408 45520 14414
rect 45468 14350 45520 14356
rect 44916 14272 44968 14278
rect 44916 14214 44968 14220
rect 45192 14272 45244 14278
rect 45192 14214 45244 14220
rect 44824 13864 44876 13870
rect 44824 13806 44876 13812
rect 44732 13184 44784 13190
rect 44732 13126 44784 13132
rect 44744 12918 44772 13126
rect 44732 12912 44784 12918
rect 44732 12854 44784 12860
rect 44836 12850 44864 13806
rect 44824 12844 44876 12850
rect 44824 12786 44876 12792
rect 44640 11212 44692 11218
rect 44640 11154 44692 11160
rect 44928 10742 44956 14214
rect 45204 13394 45232 14214
rect 45192 13388 45244 13394
rect 45192 13330 45244 13336
rect 45480 12986 45508 14350
rect 45664 14006 45692 15302
rect 45756 14414 45784 15438
rect 45744 14408 45796 14414
rect 45744 14350 45796 14356
rect 45652 14000 45704 14006
rect 45652 13942 45704 13948
rect 45744 13864 45796 13870
rect 45848 13852 45876 16594
rect 46032 16114 46060 16934
rect 46216 16794 46244 17070
rect 46480 16992 46532 16998
rect 46480 16934 46532 16940
rect 47032 16992 47084 16998
rect 47032 16934 47084 16940
rect 46204 16788 46256 16794
rect 46204 16730 46256 16736
rect 46388 16652 46440 16658
rect 46388 16594 46440 16600
rect 46110 16552 46166 16561
rect 46110 16487 46166 16496
rect 46020 16108 46072 16114
rect 46020 16050 46072 16056
rect 46032 15978 46060 16050
rect 46020 15972 46072 15978
rect 46020 15914 46072 15920
rect 46020 15088 46072 15094
rect 46020 15030 46072 15036
rect 46032 14958 46060 15030
rect 46020 14952 46072 14958
rect 46020 14894 46072 14900
rect 46124 13870 46152 16487
rect 46400 16250 46428 16594
rect 46388 16244 46440 16250
rect 46388 16186 46440 16192
rect 46400 16028 46428 16186
rect 46492 16182 46520 16934
rect 47044 16726 47072 16934
rect 47032 16720 47084 16726
rect 47032 16662 47084 16668
rect 46572 16652 46624 16658
rect 46572 16594 46624 16600
rect 46480 16176 46532 16182
rect 46480 16118 46532 16124
rect 46400 16000 46520 16028
rect 46204 15972 46256 15978
rect 46204 15914 46256 15920
rect 46216 15570 46244 15914
rect 46492 15570 46520 16000
rect 46204 15564 46256 15570
rect 46204 15506 46256 15512
rect 46480 15564 46532 15570
rect 46480 15506 46532 15512
rect 46296 14952 46348 14958
rect 46296 14894 46348 14900
rect 45796 13824 45876 13852
rect 46112 13864 46164 13870
rect 45744 13806 45796 13812
rect 46112 13806 46164 13812
rect 45756 13705 45784 13806
rect 45742 13696 45798 13705
rect 45742 13631 45798 13640
rect 45468 12980 45520 12986
rect 45468 12922 45520 12928
rect 45928 12980 45980 12986
rect 45928 12922 45980 12928
rect 45284 12368 45336 12374
rect 45284 12310 45336 12316
rect 45560 12368 45612 12374
rect 45560 12310 45612 12316
rect 45296 12220 45324 12310
rect 45296 12192 45508 12220
rect 45480 12102 45508 12192
rect 45468 12096 45520 12102
rect 45468 12038 45520 12044
rect 45192 11620 45244 11626
rect 45192 11562 45244 11568
rect 44916 10736 44968 10742
rect 44916 10678 44968 10684
rect 44456 10668 44508 10674
rect 44456 10610 44508 10616
rect 44362 10296 44418 10305
rect 43904 10260 43956 10266
rect 44468 10266 44496 10610
rect 45204 10606 45232 11562
rect 45480 11354 45508 12038
rect 45572 11626 45600 12310
rect 45652 12096 45704 12102
rect 45652 12038 45704 12044
rect 45664 11830 45692 12038
rect 45652 11824 45704 11830
rect 45652 11766 45704 11772
rect 45560 11620 45612 11626
rect 45560 11562 45612 11568
rect 45744 11552 45796 11558
rect 45744 11494 45796 11500
rect 45468 11348 45520 11354
rect 45468 11290 45520 11296
rect 45756 11150 45784 11494
rect 45744 11144 45796 11150
rect 45744 11086 45796 11092
rect 45192 10600 45244 10606
rect 45192 10542 45244 10548
rect 45192 10464 45244 10470
rect 45192 10406 45244 10412
rect 44362 10231 44418 10240
rect 44456 10260 44508 10266
rect 43904 10202 43956 10208
rect 42432 10192 42484 10198
rect 42432 10134 42484 10140
rect 43352 10124 43404 10130
rect 43352 10066 43404 10072
rect 42616 10056 42668 10062
rect 42616 9998 42668 10004
rect 42628 9926 42656 9998
rect 42616 9920 42668 9926
rect 42616 9862 42668 9868
rect 42708 9920 42760 9926
rect 42708 9862 42760 9868
rect 42720 9761 42748 9862
rect 42706 9752 42762 9761
rect 42706 9687 42762 9696
rect 42156 9580 42208 9586
rect 42156 9522 42208 9528
rect 42800 9580 42852 9586
rect 42800 9522 42852 9528
rect 42064 9512 42116 9518
rect 42064 9454 42116 9460
rect 41788 9376 41840 9382
rect 41788 9318 41840 9324
rect 41602 9208 41658 9217
rect 41602 9143 41658 9152
rect 41616 9110 41644 9143
rect 41512 9104 41564 9110
rect 41512 9046 41564 9052
rect 41604 9104 41656 9110
rect 41604 9046 41656 9052
rect 41604 8900 41656 8906
rect 41604 8842 41656 8848
rect 41420 8832 41472 8838
rect 41420 8774 41472 8780
rect 41328 8560 41380 8566
rect 41328 8502 41380 8508
rect 41052 8492 41104 8498
rect 41052 8434 41104 8440
rect 41616 8430 41644 8842
rect 42076 8430 42104 9454
rect 42430 8664 42486 8673
rect 42430 8599 42432 8608
rect 42484 8599 42486 8608
rect 42432 8570 42484 8576
rect 41604 8424 41656 8430
rect 41604 8366 41656 8372
rect 42064 8424 42116 8430
rect 42064 8366 42116 8372
rect 41604 7880 41656 7886
rect 41604 7822 41656 7828
rect 40960 7812 41012 7818
rect 40960 7754 41012 7760
rect 41328 7744 41380 7750
rect 41328 7686 41380 7692
rect 40868 7336 40920 7342
rect 40868 7278 40920 7284
rect 40960 7336 41012 7342
rect 40960 7278 41012 7284
rect 41236 7336 41288 7342
rect 41236 7278 41288 7284
rect 40776 6996 40828 7002
rect 40776 6938 40828 6944
rect 40880 6934 40908 7278
rect 40224 6928 40276 6934
rect 40224 6870 40276 6876
rect 40868 6928 40920 6934
rect 40868 6870 40920 6876
rect 40236 6458 40264 6870
rect 40776 6792 40828 6798
rect 40776 6734 40828 6740
rect 40316 6724 40368 6730
rect 40316 6666 40368 6672
rect 40224 6452 40276 6458
rect 40224 6394 40276 6400
rect 40328 6322 40356 6666
rect 40132 6316 40184 6322
rect 40132 6258 40184 6264
rect 40316 6316 40368 6322
rect 40316 6258 40368 6264
rect 40144 5914 40172 6258
rect 40132 5908 40184 5914
rect 40132 5850 40184 5856
rect 40328 5846 40356 6258
rect 40316 5840 40368 5846
rect 40316 5782 40368 5788
rect 40040 5364 40092 5370
rect 40040 5306 40092 5312
rect 39028 4752 39080 4758
rect 39028 4694 39080 4700
rect 38198 4584 38254 4593
rect 38198 4519 38254 4528
rect 38476 4548 38528 4554
rect 38476 4490 38528 4496
rect 38016 4480 38068 4486
rect 38016 4422 38068 4428
rect 38488 4078 38516 4490
rect 40052 4486 40080 5306
rect 40328 5030 40356 5782
rect 40316 5024 40368 5030
rect 40316 4966 40368 4972
rect 40408 4616 40460 4622
rect 40408 4558 40460 4564
rect 40040 4480 40092 4486
rect 40040 4422 40092 4428
rect 38844 4140 38896 4146
rect 38844 4082 38896 4088
rect 39948 4140 40000 4146
rect 39948 4082 40000 4088
rect 38476 4072 38528 4078
rect 38476 4014 38528 4020
rect 37924 3936 37976 3942
rect 37924 3878 37976 3884
rect 38108 3936 38160 3942
rect 38108 3878 38160 3884
rect 38120 3670 38148 3878
rect 38108 3664 38160 3670
rect 38108 3606 38160 3612
rect 38856 3466 38884 4082
rect 39960 3670 39988 4082
rect 39948 3664 40000 3670
rect 39948 3606 40000 3612
rect 40420 3602 40448 4558
rect 40684 4548 40736 4554
rect 40684 4490 40736 4496
rect 40696 4078 40724 4490
rect 40788 4078 40816 6734
rect 40868 6724 40920 6730
rect 40868 6666 40920 6672
rect 40880 5778 40908 6666
rect 40972 6186 41000 7278
rect 41144 7200 41196 7206
rect 41144 7142 41196 7148
rect 41156 6798 41184 7142
rect 41248 6934 41276 7278
rect 41236 6928 41288 6934
rect 41236 6870 41288 6876
rect 41144 6792 41196 6798
rect 41144 6734 41196 6740
rect 41248 6458 41276 6870
rect 41236 6452 41288 6458
rect 41236 6394 41288 6400
rect 40960 6180 41012 6186
rect 40960 6122 41012 6128
rect 40868 5772 40920 5778
rect 40868 5714 40920 5720
rect 40880 5370 40908 5714
rect 40868 5364 40920 5370
rect 40868 5306 40920 5312
rect 40972 5030 41000 6122
rect 41236 5840 41288 5846
rect 41340 5794 41368 7686
rect 41616 7546 41644 7822
rect 42444 7546 42472 8570
rect 42812 8514 42840 9522
rect 42892 9172 42944 9178
rect 42892 9114 42944 9120
rect 42536 8486 42840 8514
rect 42904 8498 42932 9114
rect 42892 8492 42944 8498
rect 42536 7886 42564 8486
rect 42892 8434 42944 8440
rect 43168 8492 43220 8498
rect 43168 8434 43220 8440
rect 42708 8424 42760 8430
rect 42760 8372 42932 8378
rect 42708 8366 42932 8372
rect 42720 8350 42932 8366
rect 42904 8294 42932 8350
rect 42892 8288 42944 8294
rect 42892 8230 42944 8236
rect 42616 8016 42668 8022
rect 42616 7958 42668 7964
rect 42524 7880 42576 7886
rect 42524 7822 42576 7828
rect 42628 7721 42656 7958
rect 42904 7954 42932 8230
rect 43076 8084 43128 8090
rect 43076 8026 43128 8032
rect 42892 7948 42944 7954
rect 42892 7890 42944 7896
rect 42984 7880 43036 7886
rect 42984 7822 43036 7828
rect 42892 7744 42944 7750
rect 42614 7712 42670 7721
rect 42892 7686 42944 7692
rect 42614 7647 42670 7656
rect 41604 7540 41656 7546
rect 41604 7482 41656 7488
rect 42432 7540 42484 7546
rect 42432 7482 42484 7488
rect 41512 7472 41564 7478
rect 41512 7414 41564 7420
rect 41524 7002 41552 7414
rect 42444 7410 42472 7482
rect 42432 7404 42484 7410
rect 42432 7346 42484 7352
rect 41604 7336 41656 7342
rect 41604 7278 41656 7284
rect 41512 6996 41564 7002
rect 41512 6938 41564 6944
rect 41616 5914 41644 7278
rect 41880 7268 41932 7274
rect 41880 7210 41932 7216
rect 42064 7268 42116 7274
rect 42064 7210 42116 7216
rect 41892 7177 41920 7210
rect 41972 7200 42024 7206
rect 41878 7168 41934 7177
rect 41972 7142 42024 7148
rect 41878 7103 41934 7112
rect 41984 6866 42012 7142
rect 41972 6860 42024 6866
rect 41972 6802 42024 6808
rect 41604 5908 41656 5914
rect 41604 5850 41656 5856
rect 41288 5788 41368 5794
rect 41236 5782 41368 5788
rect 41248 5766 41368 5782
rect 41236 5704 41288 5710
rect 41236 5646 41288 5652
rect 41248 5166 41276 5646
rect 41340 5166 41368 5766
rect 42076 5302 42104 7210
rect 42904 6866 42932 7686
rect 42996 7546 43024 7822
rect 42984 7540 43036 7546
rect 42984 7482 43036 7488
rect 43088 7478 43116 8026
rect 43076 7472 43128 7478
rect 43076 7414 43128 7420
rect 43076 7336 43128 7342
rect 43076 7278 43128 7284
rect 43088 6934 43116 7278
rect 43076 6928 43128 6934
rect 43076 6870 43128 6876
rect 42892 6860 42944 6866
rect 42892 6802 42944 6808
rect 43088 6798 43116 6870
rect 43076 6792 43128 6798
rect 42430 6760 42486 6769
rect 43076 6734 43128 6740
rect 43180 6730 43208 8434
rect 43364 6730 43392 10066
rect 44376 10062 44404 10231
rect 44456 10202 44508 10208
rect 43536 10056 43588 10062
rect 43536 9998 43588 10004
rect 43812 10056 43864 10062
rect 43812 9998 43864 10004
rect 44364 10056 44416 10062
rect 44364 9998 44416 10004
rect 43548 9586 43576 9998
rect 43824 9586 43852 9998
rect 43904 9920 43956 9926
rect 43904 9862 43956 9868
rect 43916 9586 43944 9862
rect 44272 9716 44324 9722
rect 44272 9658 44324 9664
rect 43536 9580 43588 9586
rect 43536 9522 43588 9528
rect 43812 9580 43864 9586
rect 43812 9522 43864 9528
rect 43904 9580 43956 9586
rect 43904 9522 43956 9528
rect 43824 9178 43852 9522
rect 43812 9172 43864 9178
rect 43812 9114 43864 9120
rect 43536 9104 43588 9110
rect 43442 9072 43498 9081
rect 43536 9046 43588 9052
rect 43442 9007 43444 9016
rect 43496 9007 43498 9016
rect 43444 8978 43496 8984
rect 43548 8430 43576 9046
rect 44284 9042 44312 9658
rect 44364 9580 44416 9586
rect 44364 9522 44416 9528
rect 44272 9036 44324 9042
rect 44272 8978 44324 8984
rect 43812 8968 43864 8974
rect 44376 8922 44404 9522
rect 44468 8974 44496 10202
rect 44916 10192 44968 10198
rect 44916 10134 44968 10140
rect 44548 10124 44600 10130
rect 44732 10124 44784 10130
rect 44600 10084 44732 10112
rect 44548 10066 44600 10072
rect 44732 10066 44784 10072
rect 44824 10056 44876 10062
rect 44824 9998 44876 10004
rect 44836 9897 44864 9998
rect 44928 9994 44956 10134
rect 44916 9988 44968 9994
rect 44916 9930 44968 9936
rect 44822 9888 44878 9897
rect 44822 9823 44878 9832
rect 44640 9648 44692 9654
rect 44640 9590 44692 9596
rect 43812 8910 43864 8916
rect 43444 8424 43496 8430
rect 43444 8366 43496 8372
rect 43536 8424 43588 8430
rect 43536 8366 43588 8372
rect 43456 7342 43484 8366
rect 43824 7886 43852 8910
rect 44100 8894 44404 8922
rect 44456 8968 44508 8974
rect 44456 8910 44508 8916
rect 44100 8430 44128 8894
rect 44364 8832 44416 8838
rect 44652 8820 44680 9590
rect 44732 8968 44784 8974
rect 44732 8910 44784 8916
rect 44416 8792 44680 8820
rect 44364 8774 44416 8780
rect 44180 8628 44232 8634
rect 44180 8570 44232 8576
rect 44088 8424 44140 8430
rect 44088 8366 44140 8372
rect 43812 7880 43864 7886
rect 43812 7822 43864 7828
rect 44100 7750 44128 8366
rect 44192 7750 44220 8570
rect 44088 7744 44140 7750
rect 44088 7686 44140 7692
rect 44180 7744 44232 7750
rect 44180 7686 44232 7692
rect 44100 7478 44128 7686
rect 44088 7472 44140 7478
rect 44088 7414 44140 7420
rect 43444 7336 43496 7342
rect 43444 7278 43496 7284
rect 43456 6866 43484 7278
rect 43444 6860 43496 6866
rect 43444 6802 43496 6808
rect 42430 6695 42486 6704
rect 43168 6724 43220 6730
rect 42444 6662 42472 6695
rect 43168 6666 43220 6672
rect 43352 6724 43404 6730
rect 43352 6666 43404 6672
rect 42432 6656 42484 6662
rect 42432 6598 42484 6604
rect 42892 6656 42944 6662
rect 42892 6598 42944 6604
rect 42708 6180 42760 6186
rect 42708 6122 42760 6128
rect 42524 5636 42576 5642
rect 42524 5578 42576 5584
rect 42064 5296 42116 5302
rect 42064 5238 42116 5244
rect 41236 5160 41288 5166
rect 41236 5102 41288 5108
rect 41328 5160 41380 5166
rect 41328 5102 41380 5108
rect 40960 5024 41012 5030
rect 40960 4966 41012 4972
rect 41248 4214 41276 5102
rect 41788 5092 41840 5098
rect 41788 5034 41840 5040
rect 41800 4826 41828 5034
rect 42076 5030 42104 5238
rect 42064 5024 42116 5030
rect 42064 4966 42116 4972
rect 41788 4820 41840 4826
rect 41788 4762 41840 4768
rect 42536 4622 42564 5578
rect 42720 5302 42748 6122
rect 42904 5914 42932 6598
rect 42892 5908 42944 5914
rect 42892 5850 42944 5856
rect 43074 5400 43130 5409
rect 43074 5335 43130 5344
rect 42708 5296 42760 5302
rect 42708 5238 42760 5244
rect 42984 5228 43036 5234
rect 42984 5170 43036 5176
rect 42708 5024 42760 5030
rect 42996 5001 43024 5170
rect 43088 5166 43116 5335
rect 43076 5160 43128 5166
rect 43076 5102 43128 5108
rect 42708 4966 42760 4972
rect 42982 4992 43038 5001
rect 42720 4690 42748 4966
rect 42982 4927 43038 4936
rect 42996 4758 43024 4927
rect 43364 4758 43392 6666
rect 44100 6254 44128 7414
rect 44192 6322 44220 7686
rect 44364 7540 44416 7546
rect 44364 7482 44416 7488
rect 44180 6316 44232 6322
rect 44180 6258 44232 6264
rect 44088 6248 44140 6254
rect 44088 6190 44140 6196
rect 44272 6112 44324 6118
rect 44272 6054 44324 6060
rect 44284 5778 44312 6054
rect 44376 5846 44404 7482
rect 44652 6866 44680 8792
rect 44640 6860 44692 6866
rect 44640 6802 44692 6808
rect 44640 6724 44692 6730
rect 44640 6666 44692 6672
rect 44652 6610 44680 6666
rect 44560 6582 44680 6610
rect 44560 6322 44588 6582
rect 44744 6458 44772 8910
rect 44928 8838 44956 9930
rect 45204 9897 45232 10406
rect 45190 9888 45246 9897
rect 45190 9823 45246 9832
rect 45006 9616 45062 9625
rect 45006 9551 45062 9560
rect 45020 9450 45048 9551
rect 45098 9480 45154 9489
rect 45008 9444 45060 9450
rect 45098 9415 45154 9424
rect 45008 9386 45060 9392
rect 45112 9178 45140 9415
rect 45100 9172 45152 9178
rect 45100 9114 45152 9120
rect 45204 8974 45232 9823
rect 45560 9376 45612 9382
rect 45560 9318 45612 9324
rect 45192 8968 45244 8974
rect 45192 8910 45244 8916
rect 45468 8968 45520 8974
rect 45468 8910 45520 8916
rect 44916 8832 44968 8838
rect 44916 8774 44968 8780
rect 44928 8498 44956 8774
rect 45204 8634 45232 8910
rect 45480 8838 45508 8910
rect 45468 8832 45520 8838
rect 45468 8774 45520 8780
rect 45192 8628 45244 8634
rect 45192 8570 45244 8576
rect 45376 8628 45428 8634
rect 45376 8570 45428 8576
rect 44916 8492 44968 8498
rect 44916 8434 44968 8440
rect 44928 7546 44956 8434
rect 45388 7954 45416 8570
rect 45466 8120 45522 8129
rect 45572 8106 45600 9318
rect 45652 8968 45704 8974
rect 45652 8910 45704 8916
rect 45664 8430 45692 8910
rect 45652 8424 45704 8430
rect 45652 8366 45704 8372
rect 45744 8288 45796 8294
rect 45744 8230 45796 8236
rect 45522 8078 45600 8106
rect 45650 8120 45706 8129
rect 45466 8055 45522 8064
rect 45650 8055 45652 8064
rect 45376 7948 45428 7954
rect 45376 7890 45428 7896
rect 45190 7848 45246 7857
rect 45190 7783 45246 7792
rect 44916 7540 44968 7546
rect 44916 7482 44968 7488
rect 44916 7200 44968 7206
rect 44916 7142 44968 7148
rect 44928 6866 44956 7142
rect 44916 6860 44968 6866
rect 44916 6802 44968 6808
rect 44928 6662 44956 6802
rect 44916 6656 44968 6662
rect 44916 6598 44968 6604
rect 44732 6452 44784 6458
rect 44732 6394 44784 6400
rect 44548 6316 44600 6322
rect 44548 6258 44600 6264
rect 44560 5914 44588 6258
rect 44548 5908 44600 5914
rect 44548 5850 44600 5856
rect 44364 5840 44416 5846
rect 44364 5782 44416 5788
rect 44272 5772 44324 5778
rect 44272 5714 44324 5720
rect 44456 5704 44508 5710
rect 44456 5646 44508 5652
rect 44180 5568 44232 5574
rect 44180 5510 44232 5516
rect 44192 5409 44220 5510
rect 44178 5400 44234 5409
rect 44178 5335 44234 5344
rect 43996 5160 44048 5166
rect 44364 5160 44416 5166
rect 44048 5120 44364 5148
rect 43996 5102 44048 5108
rect 44364 5102 44416 5108
rect 42984 4752 43036 4758
rect 42984 4694 43036 4700
rect 43352 4752 43404 4758
rect 43352 4694 43404 4700
rect 42708 4684 42760 4690
rect 42708 4626 42760 4632
rect 41788 4616 41840 4622
rect 41788 4558 41840 4564
rect 42524 4616 42576 4622
rect 42524 4558 42576 4564
rect 41236 4208 41288 4214
rect 41236 4150 41288 4156
rect 41800 4146 41828 4558
rect 42536 4486 42564 4558
rect 42156 4480 42208 4486
rect 42156 4422 42208 4428
rect 42524 4480 42576 4486
rect 42524 4422 42576 4428
rect 43812 4480 43864 4486
rect 43812 4422 43864 4428
rect 42168 4282 42196 4422
rect 42156 4276 42208 4282
rect 42156 4218 42208 4224
rect 43824 4146 43852 4422
rect 44008 4282 44036 5102
rect 44468 4758 44496 5646
rect 44928 4758 44956 6598
rect 45204 6458 45232 7783
rect 45480 7546 45508 8055
rect 45704 8055 45706 8064
rect 45652 8026 45704 8032
rect 45652 7880 45704 7886
rect 45756 7868 45784 8230
rect 45836 7948 45888 7954
rect 45836 7890 45888 7896
rect 45704 7840 45784 7868
rect 45652 7822 45704 7828
rect 45468 7540 45520 7546
rect 45468 7482 45520 7488
rect 45480 7206 45508 7482
rect 45560 7268 45612 7274
rect 45560 7210 45612 7216
rect 45468 7200 45520 7206
rect 45468 7142 45520 7148
rect 45284 6792 45336 6798
rect 45284 6734 45336 6740
rect 45192 6452 45244 6458
rect 45192 6394 45244 6400
rect 45296 5846 45324 6734
rect 45468 6656 45520 6662
rect 45468 6598 45520 6604
rect 45480 6254 45508 6598
rect 45572 6322 45600 7210
rect 45756 7206 45784 7840
rect 45744 7200 45796 7206
rect 45744 7142 45796 7148
rect 45756 7002 45784 7142
rect 45744 6996 45796 7002
rect 45744 6938 45796 6944
rect 45560 6316 45612 6322
rect 45560 6258 45612 6264
rect 45468 6248 45520 6254
rect 45468 6190 45520 6196
rect 45284 5840 45336 5846
rect 45284 5782 45336 5788
rect 45296 5030 45324 5782
rect 45572 5302 45600 6258
rect 45756 6202 45784 6938
rect 45848 6866 45876 7890
rect 45836 6860 45888 6866
rect 45836 6802 45888 6808
rect 45664 6174 45784 6202
rect 45664 5778 45692 6174
rect 45744 6112 45796 6118
rect 45744 6054 45796 6060
rect 45756 5778 45784 6054
rect 45652 5772 45704 5778
rect 45652 5714 45704 5720
rect 45744 5772 45796 5778
rect 45744 5714 45796 5720
rect 45560 5296 45612 5302
rect 45560 5238 45612 5244
rect 45756 5098 45784 5714
rect 45940 5234 45968 12922
rect 46308 12306 46336 14894
rect 46492 14006 46520 15506
rect 46480 14000 46532 14006
rect 46480 13942 46532 13948
rect 46492 13258 46520 13942
rect 46480 13252 46532 13258
rect 46480 13194 46532 13200
rect 46492 12986 46520 13194
rect 46480 12980 46532 12986
rect 46480 12922 46532 12928
rect 46296 12300 46348 12306
rect 46296 12242 46348 12248
rect 46020 12232 46072 12238
rect 46020 12174 46072 12180
rect 46032 11694 46060 12174
rect 46584 11830 46612 16594
rect 47136 16522 47440 16538
rect 47124 16516 47452 16522
rect 47176 16510 47400 16516
rect 47124 16458 47176 16464
rect 47400 16458 47452 16464
rect 48872 16448 48924 16454
rect 48872 16390 48924 16396
rect 47823 16348 48131 16357
rect 47823 16346 47829 16348
rect 47885 16346 47909 16348
rect 47965 16346 47989 16348
rect 48045 16346 48069 16348
rect 48125 16346 48131 16348
rect 47885 16294 47887 16346
rect 48067 16294 48069 16346
rect 47823 16292 47829 16294
rect 47885 16292 47909 16294
rect 47965 16292 47989 16294
rect 48045 16292 48069 16294
rect 48125 16292 48131 16294
rect 47823 16283 48131 16292
rect 47032 16108 47084 16114
rect 47032 16050 47084 16056
rect 47044 15910 47072 16050
rect 48688 16040 48740 16046
rect 48688 15982 48740 15988
rect 47032 15904 47084 15910
rect 47032 15846 47084 15852
rect 47124 15904 47176 15910
rect 47124 15846 47176 15852
rect 46664 15496 46716 15502
rect 46664 15438 46716 15444
rect 46676 14618 46704 15438
rect 46940 15428 46992 15434
rect 46940 15370 46992 15376
rect 46664 14612 46716 14618
rect 46664 14554 46716 14560
rect 46848 14340 46900 14346
rect 46848 14282 46900 14288
rect 46860 13530 46888 14282
rect 46848 13524 46900 13530
rect 46848 13466 46900 13472
rect 46756 13184 46808 13190
rect 46756 13126 46808 13132
rect 46768 12850 46796 13126
rect 46952 12986 46980 15370
rect 47136 15026 47164 15846
rect 47950 15736 48006 15745
rect 47950 15671 48006 15680
rect 47964 15638 47992 15671
rect 47952 15632 48004 15638
rect 47952 15574 48004 15580
rect 48700 15502 48728 15982
rect 48884 15910 48912 16390
rect 49056 16108 49108 16114
rect 49056 16050 49108 16056
rect 48780 15904 48832 15910
rect 48780 15846 48832 15852
rect 48872 15904 48924 15910
rect 48872 15846 48924 15852
rect 48688 15496 48740 15502
rect 48792 15473 48820 15846
rect 48688 15438 48740 15444
rect 48778 15464 48834 15473
rect 48504 15360 48556 15366
rect 48504 15302 48556 15308
rect 47823 15260 48131 15269
rect 47823 15258 47829 15260
rect 47885 15258 47909 15260
rect 47965 15258 47989 15260
rect 48045 15258 48069 15260
rect 48125 15258 48131 15260
rect 47885 15206 47887 15258
rect 48067 15206 48069 15258
rect 47823 15204 47829 15206
rect 47885 15204 47909 15206
rect 47965 15204 47989 15206
rect 48045 15204 48069 15206
rect 48125 15204 48131 15206
rect 47823 15195 48131 15204
rect 47124 15020 47176 15026
rect 47124 14962 47176 14968
rect 47216 15020 47268 15026
rect 47216 14962 47268 14968
rect 47136 14618 47164 14962
rect 47124 14612 47176 14618
rect 47124 14554 47176 14560
rect 47032 14340 47084 14346
rect 47032 14282 47084 14288
rect 47044 14249 47072 14282
rect 47030 14240 47086 14249
rect 47030 14175 47086 14184
rect 47228 14074 47256 14962
rect 48320 14952 48372 14958
rect 48320 14894 48372 14900
rect 48332 14385 48360 14894
rect 48318 14376 48374 14385
rect 48318 14311 48374 14320
rect 47308 14272 47360 14278
rect 47308 14214 47360 14220
rect 48320 14272 48372 14278
rect 48320 14214 48372 14220
rect 47320 14074 47348 14214
rect 47823 14172 48131 14181
rect 47823 14170 47829 14172
rect 47885 14170 47909 14172
rect 47965 14170 47989 14172
rect 48045 14170 48069 14172
rect 48125 14170 48131 14172
rect 47885 14118 47887 14170
rect 48067 14118 48069 14170
rect 47823 14116 47829 14118
rect 47885 14116 47909 14118
rect 47965 14116 47989 14118
rect 48045 14116 48069 14118
rect 48125 14116 48131 14118
rect 47823 14107 48131 14116
rect 47216 14068 47268 14074
rect 47216 14010 47268 14016
rect 47308 14068 47360 14074
rect 47308 14010 47360 14016
rect 48332 14006 48360 14214
rect 48320 14000 48372 14006
rect 48320 13942 48372 13948
rect 47676 13252 47728 13258
rect 47676 13194 47728 13200
rect 46940 12980 46992 12986
rect 46940 12922 46992 12928
rect 46756 12844 46808 12850
rect 46756 12786 46808 12792
rect 47032 12776 47084 12782
rect 47032 12718 47084 12724
rect 47044 12646 47072 12718
rect 47032 12640 47084 12646
rect 47032 12582 47084 12588
rect 47584 12436 47636 12442
rect 47584 12378 47636 12384
rect 46756 12300 46808 12306
rect 46756 12242 46808 12248
rect 46768 12073 46796 12242
rect 47124 12164 47176 12170
rect 47124 12106 47176 12112
rect 46754 12064 46810 12073
rect 46754 11999 46810 12008
rect 46572 11824 46624 11830
rect 46572 11766 46624 11772
rect 46020 11688 46072 11694
rect 46020 11630 46072 11636
rect 46296 11688 46348 11694
rect 46296 11630 46348 11636
rect 46308 10062 46336 11630
rect 46768 11150 46796 11999
rect 46848 11756 46900 11762
rect 46848 11698 46900 11704
rect 46860 11558 46888 11698
rect 46848 11552 46900 11558
rect 46848 11494 46900 11500
rect 46756 11144 46808 11150
rect 46756 11086 46808 11092
rect 47030 10840 47086 10849
rect 47030 10775 47086 10784
rect 47044 10266 47072 10775
rect 47032 10260 47084 10266
rect 47032 10202 47084 10208
rect 46112 10056 46164 10062
rect 46112 9998 46164 10004
rect 46296 10056 46348 10062
rect 46296 9998 46348 10004
rect 46124 9602 46152 9998
rect 46308 9722 46336 9998
rect 46572 9988 46624 9994
rect 46572 9930 46624 9936
rect 46584 9897 46612 9930
rect 46570 9888 46626 9897
rect 46570 9823 46626 9832
rect 46296 9716 46348 9722
rect 46296 9658 46348 9664
rect 47136 9654 47164 12106
rect 47596 11694 47624 12378
rect 47584 11688 47636 11694
rect 47584 11630 47636 11636
rect 47596 10266 47624 11630
rect 47688 10577 47716 13194
rect 47823 13084 48131 13093
rect 47823 13082 47829 13084
rect 47885 13082 47909 13084
rect 47965 13082 47989 13084
rect 48045 13082 48069 13084
rect 48125 13082 48131 13084
rect 47885 13030 47887 13082
rect 48067 13030 48069 13082
rect 47823 13028 47829 13030
rect 47885 13028 47909 13030
rect 47965 13028 47989 13030
rect 48045 13028 48069 13030
rect 48125 13028 48131 13030
rect 47823 13019 48131 13028
rect 48136 12844 48188 12850
rect 48136 12786 48188 12792
rect 48148 12306 48176 12786
rect 48226 12744 48282 12753
rect 48226 12679 48282 12688
rect 48240 12434 48268 12679
rect 48240 12406 48360 12434
rect 48136 12300 48188 12306
rect 48136 12242 48188 12248
rect 47823 11996 48131 12005
rect 47823 11994 47829 11996
rect 47885 11994 47909 11996
rect 47965 11994 47989 11996
rect 48045 11994 48069 11996
rect 48125 11994 48131 11996
rect 47885 11942 47887 11994
rect 48067 11942 48069 11994
rect 47823 11940 47829 11942
rect 47885 11940 47909 11942
rect 47965 11940 47989 11942
rect 48045 11940 48069 11942
rect 48125 11940 48131 11942
rect 47823 11931 48131 11940
rect 47823 10908 48131 10917
rect 47823 10906 47829 10908
rect 47885 10906 47909 10908
rect 47965 10906 47989 10908
rect 48045 10906 48069 10908
rect 48125 10906 48131 10908
rect 47885 10854 47887 10906
rect 48067 10854 48069 10906
rect 47823 10852 47829 10854
rect 47885 10852 47909 10854
rect 47965 10852 47989 10854
rect 48045 10852 48069 10854
rect 48125 10852 48131 10854
rect 47823 10843 48131 10852
rect 48332 10810 48360 12406
rect 48516 12238 48544 15302
rect 48700 15094 48728 15438
rect 48778 15399 48834 15408
rect 48792 15094 48820 15399
rect 48688 15088 48740 15094
rect 48688 15030 48740 15036
rect 48780 15088 48832 15094
rect 48780 15030 48832 15036
rect 48780 14000 48832 14006
rect 48780 13942 48832 13948
rect 48792 13734 48820 13942
rect 48780 13728 48832 13734
rect 48780 13670 48832 13676
rect 48792 13326 48820 13670
rect 48780 13320 48832 13326
rect 48780 13262 48832 13268
rect 49068 13258 49096 16050
rect 49528 15502 49556 17206
rect 50356 16794 50384 17274
rect 57060 17264 57112 17270
rect 57060 17206 57112 17212
rect 65892 17264 65944 17270
rect 65892 17206 65944 17212
rect 52276 17196 52328 17202
rect 52276 17138 52328 17144
rect 50344 16788 50396 16794
rect 50344 16730 50396 16736
rect 50528 16788 50580 16794
rect 50528 16730 50580 16736
rect 50356 16114 50384 16730
rect 50344 16108 50396 16114
rect 50344 16050 50396 16056
rect 50436 16108 50488 16114
rect 50436 16050 50488 16056
rect 49148 15496 49200 15502
rect 49148 15438 49200 15444
rect 49516 15496 49568 15502
rect 49516 15438 49568 15444
rect 49160 15026 49188 15438
rect 49700 15360 49752 15366
rect 49700 15302 49752 15308
rect 49712 15094 49740 15302
rect 49700 15088 49752 15094
rect 49700 15030 49752 15036
rect 49148 15020 49200 15026
rect 49148 14962 49200 14968
rect 49332 14544 49384 14550
rect 49332 14486 49384 14492
rect 49240 14408 49292 14414
rect 49240 14350 49292 14356
rect 49252 13326 49280 14350
rect 49344 13938 49372 14486
rect 49712 14278 49740 15030
rect 50356 14929 50384 16050
rect 50448 15638 50476 16050
rect 50540 16046 50568 16730
rect 51816 16516 51868 16522
rect 51816 16458 51868 16464
rect 51172 16448 51224 16454
rect 51172 16390 51224 16396
rect 50528 16040 50580 16046
rect 50528 15982 50580 15988
rect 50436 15632 50488 15638
rect 50436 15574 50488 15580
rect 50540 15366 50568 15982
rect 51184 15502 51212 16390
rect 51448 16176 51500 16182
rect 51448 16118 51500 16124
rect 51172 15496 51224 15502
rect 51172 15438 51224 15444
rect 50528 15360 50580 15366
rect 50528 15302 50580 15308
rect 50712 15088 50764 15094
rect 50712 15030 50764 15036
rect 50342 14920 50398 14929
rect 50342 14855 50398 14864
rect 50724 14618 50752 15030
rect 50896 14816 50948 14822
rect 50896 14758 50948 14764
rect 50908 14618 50936 14758
rect 50712 14612 50764 14618
rect 50712 14554 50764 14560
rect 50896 14612 50948 14618
rect 50896 14554 50948 14560
rect 50620 14408 50672 14414
rect 50620 14350 50672 14356
rect 49700 14272 49752 14278
rect 49700 14214 49752 14220
rect 50068 14272 50120 14278
rect 50068 14214 50120 14220
rect 50252 14272 50304 14278
rect 50252 14214 50304 14220
rect 49516 14000 49568 14006
rect 49516 13942 49568 13948
rect 49332 13932 49384 13938
rect 49332 13874 49384 13880
rect 49332 13524 49384 13530
rect 49332 13466 49384 13472
rect 49240 13320 49292 13326
rect 49240 13262 49292 13268
rect 49056 13252 49108 13258
rect 49056 13194 49108 13200
rect 48964 13184 49016 13190
rect 48964 13126 49016 13132
rect 48976 12850 49004 13126
rect 49344 12850 49372 13466
rect 48964 12844 49016 12850
rect 48964 12786 49016 12792
rect 49332 12844 49384 12850
rect 49332 12786 49384 12792
rect 48504 12232 48556 12238
rect 48504 12174 48556 12180
rect 48780 12164 48832 12170
rect 48780 12106 48832 12112
rect 49240 12164 49292 12170
rect 49240 12106 49292 12112
rect 48792 11150 48820 12106
rect 48962 11248 49018 11257
rect 48962 11183 48964 11192
rect 49016 11183 49018 11192
rect 48964 11154 49016 11160
rect 48780 11144 48832 11150
rect 48780 11086 48832 11092
rect 49252 11014 49280 12106
rect 49344 11778 49372 12786
rect 49528 12238 49556 13942
rect 49712 13734 49740 14214
rect 50080 14006 50108 14214
rect 50068 14000 50120 14006
rect 50068 13942 50120 13948
rect 49792 13796 49844 13802
rect 49792 13738 49844 13744
rect 49700 13728 49752 13734
rect 49700 13670 49752 13676
rect 49608 13456 49660 13462
rect 49608 13398 49660 13404
rect 49620 12442 49648 13398
rect 49700 12776 49752 12782
rect 49700 12718 49752 12724
rect 49712 12442 49740 12718
rect 49608 12436 49660 12442
rect 49608 12378 49660 12384
rect 49700 12436 49752 12442
rect 49804 12434 49832 13738
rect 49976 12776 50028 12782
rect 49976 12718 50028 12724
rect 49804 12406 49924 12434
rect 49700 12378 49752 12384
rect 49516 12232 49568 12238
rect 49516 12174 49568 12180
rect 49344 11750 49464 11778
rect 49332 11688 49384 11694
rect 49332 11630 49384 11636
rect 49240 11008 49292 11014
rect 49240 10950 49292 10956
rect 48410 10840 48466 10849
rect 48320 10804 48372 10810
rect 48410 10775 48466 10784
rect 48320 10746 48372 10752
rect 48424 10742 48452 10775
rect 48412 10736 48464 10742
rect 48412 10678 48464 10684
rect 48504 10668 48556 10674
rect 48504 10610 48556 10616
rect 47674 10568 47730 10577
rect 47674 10503 47730 10512
rect 48320 10464 48372 10470
rect 48320 10406 48372 10412
rect 47584 10260 47636 10266
rect 47584 10202 47636 10208
rect 47823 9820 48131 9829
rect 47823 9818 47829 9820
rect 47885 9818 47909 9820
rect 47965 9818 47989 9820
rect 48045 9818 48069 9820
rect 48125 9818 48131 9820
rect 47885 9766 47887 9818
rect 48067 9766 48069 9818
rect 47823 9764 47829 9766
rect 47885 9764 47909 9766
rect 47965 9764 47989 9766
rect 48045 9764 48069 9766
rect 48125 9764 48131 9766
rect 47823 9755 48131 9764
rect 48332 9654 48360 10406
rect 48516 9654 48544 10610
rect 48780 10532 48832 10538
rect 48780 10474 48832 10480
rect 48792 10198 48820 10474
rect 48780 10192 48832 10198
rect 48780 10134 48832 10140
rect 49252 10146 49280 10950
rect 49344 10577 49372 11630
rect 49330 10568 49386 10577
rect 49330 10503 49386 10512
rect 49252 10118 49372 10146
rect 48780 10056 48832 10062
rect 48780 9998 48832 10004
rect 49240 10056 49292 10062
rect 49240 9998 49292 10004
rect 48792 9722 48820 9998
rect 48780 9716 48832 9722
rect 48780 9658 48832 9664
rect 47124 9648 47176 9654
rect 46124 9574 46428 9602
rect 47124 9590 47176 9596
rect 48320 9648 48372 9654
rect 48320 9590 48372 9596
rect 48504 9648 48556 9654
rect 48504 9590 48556 9596
rect 46204 9512 46256 9518
rect 46204 9454 46256 9460
rect 46296 9512 46348 9518
rect 46296 9454 46348 9460
rect 46216 9178 46244 9454
rect 46308 9178 46336 9454
rect 46204 9172 46256 9178
rect 46204 9114 46256 9120
rect 46296 9172 46348 9178
rect 46296 9114 46348 9120
rect 46204 8968 46256 8974
rect 46308 8956 46336 9114
rect 46400 8974 46428 9574
rect 46572 9512 46624 9518
rect 46572 9454 46624 9460
rect 48228 9512 48280 9518
rect 48228 9454 48280 9460
rect 48688 9512 48740 9518
rect 48688 9454 48740 9460
rect 46584 9353 46612 9454
rect 47492 9444 47544 9450
rect 47492 9386 47544 9392
rect 46570 9344 46626 9353
rect 46626 9302 46704 9330
rect 46570 9279 46626 9288
rect 46256 8928 46336 8956
rect 46388 8968 46440 8974
rect 46204 8910 46256 8916
rect 46388 8910 46440 8916
rect 46400 6458 46428 8910
rect 46572 8832 46624 8838
rect 46570 8800 46572 8809
rect 46624 8800 46626 8809
rect 46570 8735 46626 8744
rect 46584 8566 46612 8597
rect 46572 8560 46624 8566
rect 46570 8528 46572 8537
rect 46624 8528 46626 8537
rect 46570 8463 46626 8472
rect 46584 8362 46612 8463
rect 46572 8356 46624 8362
rect 46572 8298 46624 8304
rect 46570 7576 46626 7585
rect 46570 7511 46572 7520
rect 46624 7511 46626 7520
rect 46572 7482 46624 7488
rect 46584 7410 46612 7482
rect 46572 7404 46624 7410
rect 46572 7346 46624 7352
rect 46388 6452 46440 6458
rect 46388 6394 46440 6400
rect 46204 6316 46256 6322
rect 46204 6258 46256 6264
rect 46216 5642 46244 6258
rect 46676 5914 46704 9302
rect 46754 9072 46810 9081
rect 46754 9007 46810 9016
rect 46768 8838 46796 9007
rect 47400 8968 47452 8974
rect 47400 8910 47452 8916
rect 46756 8832 46808 8838
rect 46756 8774 46808 8780
rect 47214 8800 47270 8809
rect 47214 8735 47270 8744
rect 46848 8492 46900 8498
rect 46848 8434 46900 8440
rect 46756 8288 46808 8294
rect 46756 8230 46808 8236
rect 46768 7698 46796 8230
rect 46860 7818 46888 8434
rect 47032 8424 47084 8430
rect 47032 8366 47084 8372
rect 47044 8022 47072 8366
rect 47228 8090 47256 8735
rect 47412 8634 47440 8910
rect 47400 8628 47452 8634
rect 47400 8570 47452 8576
rect 47308 8424 47360 8430
rect 47308 8366 47360 8372
rect 47216 8084 47268 8090
rect 47216 8026 47268 8032
rect 47032 8016 47084 8022
rect 47032 7958 47084 7964
rect 47216 7948 47268 7954
rect 47216 7890 47268 7896
rect 47032 7880 47084 7886
rect 47032 7822 47084 7828
rect 46848 7812 46900 7818
rect 46848 7754 46900 7760
rect 47044 7698 47072 7822
rect 47228 7818 47256 7890
rect 47216 7812 47268 7818
rect 47216 7754 47268 7760
rect 46768 7670 47072 7698
rect 47320 7546 47348 8366
rect 47398 8120 47454 8129
rect 47398 8055 47454 8064
rect 47412 8022 47440 8055
rect 47400 8016 47452 8022
rect 47400 7958 47452 7964
rect 47308 7540 47360 7546
rect 47308 7482 47360 7488
rect 47320 7342 47348 7482
rect 47308 7336 47360 7342
rect 47308 7278 47360 7284
rect 47308 6656 47360 6662
rect 47308 6598 47360 6604
rect 46940 6248 46992 6254
rect 46940 6190 46992 6196
rect 46952 6118 46980 6190
rect 46940 6112 46992 6118
rect 46940 6054 46992 6060
rect 46664 5908 46716 5914
rect 46664 5850 46716 5856
rect 47320 5681 47348 6598
rect 47306 5672 47362 5681
rect 46204 5636 46256 5642
rect 47306 5607 47308 5616
rect 46204 5578 46256 5584
rect 47360 5607 47362 5616
rect 47308 5578 47360 5584
rect 45928 5228 45980 5234
rect 45928 5170 45980 5176
rect 45744 5092 45796 5098
rect 45744 5034 45796 5040
rect 45284 5024 45336 5030
rect 45284 4966 45336 4972
rect 44456 4752 44508 4758
rect 44456 4694 44508 4700
rect 44916 4752 44968 4758
rect 44916 4694 44968 4700
rect 45836 4684 45888 4690
rect 45836 4626 45888 4632
rect 45848 4593 45876 4626
rect 45834 4584 45890 4593
rect 45834 4519 45890 4528
rect 45940 4486 45968 5170
rect 47124 5160 47176 5166
rect 47504 5137 47532 9386
rect 47582 9072 47638 9081
rect 47582 9007 47638 9016
rect 47596 8906 47624 9007
rect 47584 8900 47636 8906
rect 47584 8842 47636 8848
rect 47823 8732 48131 8741
rect 47823 8730 47829 8732
rect 47885 8730 47909 8732
rect 47965 8730 47989 8732
rect 48045 8730 48069 8732
rect 48125 8730 48131 8732
rect 47885 8678 47887 8730
rect 48067 8678 48069 8730
rect 47823 8676 47829 8678
rect 47885 8676 47909 8678
rect 47965 8676 47989 8678
rect 48045 8676 48069 8678
rect 48125 8676 48131 8678
rect 47823 8667 48131 8676
rect 48240 8090 48268 9454
rect 48700 8430 48728 9454
rect 48872 9376 48924 9382
rect 48870 9344 48872 9353
rect 49056 9376 49108 9382
rect 48924 9344 48926 9353
rect 49056 9318 49108 9324
rect 48870 9279 48926 9288
rect 48778 9072 48834 9081
rect 49068 9042 49096 9318
rect 48778 9007 48834 9016
rect 49056 9036 49108 9042
rect 48688 8424 48740 8430
rect 48688 8366 48740 8372
rect 48320 8356 48372 8362
rect 48320 8298 48372 8304
rect 48228 8084 48280 8090
rect 48228 8026 48280 8032
rect 48332 7886 48360 8298
rect 48228 7880 48280 7886
rect 48228 7822 48280 7828
rect 48320 7880 48372 7886
rect 48320 7822 48372 7828
rect 47823 7644 48131 7653
rect 47823 7642 47829 7644
rect 47885 7642 47909 7644
rect 47965 7642 47989 7644
rect 48045 7642 48069 7644
rect 48125 7642 48131 7644
rect 47885 7590 47887 7642
rect 48067 7590 48069 7642
rect 47823 7588 47829 7590
rect 47885 7588 47909 7590
rect 47965 7588 47989 7590
rect 48045 7588 48069 7590
rect 48125 7588 48131 7590
rect 47823 7579 48131 7588
rect 48240 7274 48268 7822
rect 48700 7274 48728 8366
rect 48228 7268 48280 7274
rect 48228 7210 48280 7216
rect 48688 7268 48740 7274
rect 48688 7210 48740 7216
rect 48792 6866 48820 9007
rect 49056 8978 49108 8984
rect 48872 8288 48924 8294
rect 48872 8230 48924 8236
rect 48884 7750 48912 8230
rect 49252 8090 49280 9998
rect 49344 9926 49372 10118
rect 49436 9994 49464 11750
rect 49620 11626 49648 12378
rect 49896 11665 49924 12406
rect 49882 11656 49938 11665
rect 49608 11620 49660 11626
rect 49882 11591 49938 11600
rect 49608 11562 49660 11568
rect 49698 11248 49754 11257
rect 49698 11183 49754 11192
rect 49712 11150 49740 11183
rect 49608 11144 49660 11150
rect 49608 11086 49660 11092
rect 49700 11144 49752 11150
rect 49700 11086 49752 11092
rect 49514 10976 49570 10985
rect 49514 10911 49570 10920
rect 49528 10062 49556 10911
rect 49620 10130 49648 11086
rect 49700 11008 49752 11014
rect 49700 10950 49752 10956
rect 49712 10606 49740 10950
rect 49700 10600 49752 10606
rect 49700 10542 49752 10548
rect 49712 10266 49740 10542
rect 49884 10464 49936 10470
rect 49884 10406 49936 10412
rect 49700 10260 49752 10266
rect 49700 10202 49752 10208
rect 49896 10198 49924 10406
rect 49884 10192 49936 10198
rect 49884 10134 49936 10140
rect 49608 10124 49660 10130
rect 49608 10066 49660 10072
rect 49516 10056 49568 10062
rect 49516 9998 49568 10004
rect 49792 10056 49844 10062
rect 49792 9998 49844 10004
rect 49424 9988 49476 9994
rect 49424 9930 49476 9936
rect 49332 9920 49384 9926
rect 49332 9862 49384 9868
rect 49608 9648 49660 9654
rect 49608 9590 49660 9596
rect 49332 9580 49384 9586
rect 49332 9522 49384 9528
rect 49240 8084 49292 8090
rect 49240 8026 49292 8032
rect 49344 7954 49372 9522
rect 49424 9444 49476 9450
rect 49424 9386 49476 9392
rect 49436 9178 49464 9386
rect 49620 9353 49648 9590
rect 49700 9512 49752 9518
rect 49700 9454 49752 9460
rect 49606 9344 49662 9353
rect 49606 9279 49662 9288
rect 49424 9172 49476 9178
rect 49424 9114 49476 9120
rect 49424 8832 49476 8838
rect 49424 8774 49476 8780
rect 49436 8498 49464 8774
rect 49516 8628 49568 8634
rect 49516 8570 49568 8576
rect 49424 8492 49476 8498
rect 49424 8434 49476 8440
rect 49528 8401 49556 8570
rect 49620 8498 49648 9279
rect 49608 8492 49660 8498
rect 49608 8434 49660 8440
rect 49514 8392 49570 8401
rect 49514 8327 49570 8336
rect 49712 8090 49740 9454
rect 49804 8974 49832 9998
rect 49988 9654 50016 12718
rect 50264 12434 50292 14214
rect 50344 13864 50396 13870
rect 50344 13806 50396 13812
rect 50356 13326 50384 13806
rect 50436 13728 50488 13734
rect 50436 13670 50488 13676
rect 50344 13320 50396 13326
rect 50344 13262 50396 13268
rect 50448 13172 50476 13670
rect 50356 13144 50476 13172
rect 50356 12986 50384 13144
rect 50344 12980 50396 12986
rect 50344 12922 50396 12928
rect 50356 12646 50384 12922
rect 50344 12640 50396 12646
rect 50344 12582 50396 12588
rect 50172 12406 50292 12434
rect 50172 12170 50200 12406
rect 50356 12238 50384 12582
rect 50344 12232 50396 12238
rect 50344 12174 50396 12180
rect 50160 12164 50212 12170
rect 50160 12106 50212 12112
rect 50068 12096 50120 12102
rect 50068 12038 50120 12044
rect 50080 11150 50108 12038
rect 50172 11762 50200 12106
rect 50344 12096 50396 12102
rect 50344 12038 50396 12044
rect 50252 11824 50304 11830
rect 50252 11766 50304 11772
rect 50160 11756 50212 11762
rect 50160 11698 50212 11704
rect 50068 11144 50120 11150
rect 50068 11086 50120 11092
rect 50158 10840 50214 10849
rect 50068 10804 50120 10810
rect 50158 10775 50160 10784
rect 50068 10746 50120 10752
rect 50212 10775 50214 10784
rect 50160 10746 50212 10752
rect 50080 10470 50108 10746
rect 50068 10464 50120 10470
rect 50068 10406 50120 10412
rect 50264 10062 50292 11766
rect 50356 11098 50384 12038
rect 50528 11688 50580 11694
rect 50528 11630 50580 11636
rect 50436 11552 50488 11558
rect 50436 11494 50488 11500
rect 50448 11218 50476 11494
rect 50436 11212 50488 11218
rect 50436 11154 50488 11160
rect 50356 11070 50476 11098
rect 50540 11082 50568 11630
rect 50632 11257 50660 14350
rect 51184 13546 51212 15438
rect 51460 15434 51488 16118
rect 51448 15428 51500 15434
rect 51448 15370 51500 15376
rect 51724 14816 51776 14822
rect 51724 14758 51776 14764
rect 51448 14612 51500 14618
rect 51448 14554 51500 14560
rect 51540 14612 51592 14618
rect 51540 14554 51592 14560
rect 51354 14376 51410 14385
rect 51354 14311 51410 14320
rect 51000 13518 51212 13546
rect 51000 12730 51028 13518
rect 51264 13184 51316 13190
rect 51264 13126 51316 13132
rect 51172 12776 51224 12782
rect 51000 12702 51120 12730
rect 51172 12718 51224 12724
rect 51092 12434 51120 12702
rect 51046 12406 51120 12434
rect 51046 12220 51074 12406
rect 51046 12192 51120 12220
rect 50896 12164 50948 12170
rect 50896 12106 50948 12112
rect 50618 11248 50674 11257
rect 50618 11183 50674 11192
rect 50632 11150 50660 11183
rect 50620 11144 50672 11150
rect 50620 11086 50672 11092
rect 50712 11144 50764 11150
rect 50712 11086 50764 11092
rect 50344 10668 50396 10674
rect 50344 10610 50396 10616
rect 50252 10056 50304 10062
rect 50252 9998 50304 10004
rect 50356 9722 50384 10610
rect 50448 10606 50476 11070
rect 50528 11076 50580 11082
rect 50528 11018 50580 11024
rect 50436 10600 50488 10606
rect 50436 10542 50488 10548
rect 50344 9716 50396 9722
rect 50344 9658 50396 9664
rect 49976 9648 50028 9654
rect 49976 9590 50028 9596
rect 49792 8968 49844 8974
rect 49792 8910 49844 8916
rect 49976 8424 50028 8430
rect 49976 8366 50028 8372
rect 49988 8090 50016 8366
rect 49700 8084 49752 8090
rect 49700 8026 49752 8032
rect 49976 8084 50028 8090
rect 49976 8026 50028 8032
rect 49332 7948 49384 7954
rect 49332 7890 49384 7896
rect 49700 7948 49752 7954
rect 49700 7890 49752 7896
rect 48872 7744 48924 7750
rect 48872 7686 48924 7692
rect 49148 7404 49200 7410
rect 49148 7346 49200 7352
rect 49160 7177 49188 7346
rect 49344 7342 49372 7890
rect 49712 7478 49740 7890
rect 50448 7818 50476 10542
rect 50632 9178 50660 11086
rect 50724 10985 50752 11086
rect 50908 11082 50936 12106
rect 50896 11076 50948 11082
rect 50896 11018 50948 11024
rect 50804 11008 50856 11014
rect 50710 10976 50766 10985
rect 50804 10950 50856 10956
rect 50710 10911 50766 10920
rect 50816 10742 50844 10950
rect 50804 10736 50856 10742
rect 50804 10678 50856 10684
rect 50712 10600 50764 10606
rect 50712 10542 50764 10548
rect 50724 10266 50752 10542
rect 50712 10260 50764 10266
rect 50712 10202 50764 10208
rect 50804 10260 50856 10266
rect 50804 10202 50856 10208
rect 50816 9994 50844 10202
rect 50804 9988 50856 9994
rect 50804 9930 50856 9936
rect 50620 9172 50672 9178
rect 50672 9132 50752 9160
rect 50620 9114 50672 9120
rect 50724 9042 50752 9132
rect 50712 9036 50764 9042
rect 50712 8978 50764 8984
rect 50620 8968 50672 8974
rect 50620 8910 50672 8916
rect 50632 8634 50660 8910
rect 50620 8628 50672 8634
rect 50620 8570 50672 8576
rect 51092 7993 51120 12192
rect 51184 11937 51212 12718
rect 51276 12238 51304 13126
rect 51264 12232 51316 12238
rect 51368 12209 51396 14311
rect 51460 13870 51488 14554
rect 51552 14414 51580 14554
rect 51540 14408 51592 14414
rect 51540 14350 51592 14356
rect 51448 13864 51500 13870
rect 51448 13806 51500 13812
rect 51632 13728 51684 13734
rect 51632 13670 51684 13676
rect 51540 13388 51592 13394
rect 51540 13330 51592 13336
rect 51552 12628 51580 13330
rect 51644 12782 51672 13670
rect 51736 13462 51764 14758
rect 51828 14346 51856 16458
rect 52288 16250 52316 17138
rect 55128 17060 55180 17066
rect 55128 17002 55180 17008
rect 55140 16794 55168 17002
rect 56692 16992 56744 16998
rect 56692 16934 56744 16940
rect 55128 16788 55180 16794
rect 55128 16730 55180 16736
rect 54944 16720 54996 16726
rect 54944 16662 54996 16668
rect 53564 16652 53616 16658
rect 53564 16594 53616 16600
rect 52368 16448 52420 16454
rect 52368 16390 52420 16396
rect 52092 16244 52144 16250
rect 52092 16186 52144 16192
rect 52276 16244 52328 16250
rect 52276 16186 52328 16192
rect 52104 14958 52132 16186
rect 52380 16114 52408 16390
rect 53576 16182 53604 16594
rect 54852 16516 54904 16522
rect 54852 16458 54904 16464
rect 53564 16176 53616 16182
rect 53564 16118 53616 16124
rect 52368 16108 52420 16114
rect 52368 16050 52420 16056
rect 52380 16017 52408 16050
rect 52366 16008 52422 16017
rect 52366 15943 52422 15952
rect 53012 15904 53064 15910
rect 53012 15846 53064 15852
rect 53024 15434 53052 15846
rect 53012 15428 53064 15434
rect 53012 15370 53064 15376
rect 53104 15088 53156 15094
rect 53104 15030 53156 15036
rect 52092 14952 52144 14958
rect 52092 14894 52144 14900
rect 52000 14816 52052 14822
rect 52000 14758 52052 14764
rect 51816 14340 51868 14346
rect 51816 14282 51868 14288
rect 51724 13456 51776 13462
rect 51724 13398 51776 13404
rect 51736 12850 51764 13398
rect 52012 12986 52040 14758
rect 53116 14550 53144 15030
rect 53104 14544 53156 14550
rect 53104 14486 53156 14492
rect 53576 13938 53604 16118
rect 53656 16108 53708 16114
rect 53656 16050 53708 16056
rect 54208 16108 54260 16114
rect 54208 16050 54260 16056
rect 53668 15502 53696 16050
rect 53656 15496 53708 15502
rect 53656 15438 53708 15444
rect 53668 14396 53696 15438
rect 53748 15360 53800 15366
rect 53748 15302 53800 15308
rect 53760 15094 53788 15302
rect 53748 15088 53800 15094
rect 53748 15030 53800 15036
rect 53838 15056 53894 15065
rect 53838 14991 53894 15000
rect 53748 14408 53800 14414
rect 53668 14368 53748 14396
rect 53748 14350 53800 14356
rect 53760 13938 53788 14350
rect 52368 13932 52420 13938
rect 52368 13874 52420 13880
rect 53564 13932 53616 13938
rect 53564 13874 53616 13880
rect 53748 13932 53800 13938
rect 53748 13874 53800 13880
rect 52276 13796 52328 13802
rect 52276 13738 52328 13744
rect 52184 13728 52236 13734
rect 52184 13670 52236 13676
rect 52092 13252 52144 13258
rect 52092 13194 52144 13200
rect 52104 13161 52132 13194
rect 52196 13190 52224 13670
rect 52184 13184 52236 13190
rect 52090 13152 52146 13161
rect 52184 13126 52236 13132
rect 52090 13087 52146 13096
rect 52000 12980 52052 12986
rect 52000 12922 52052 12928
rect 52012 12850 52040 12922
rect 51724 12844 51776 12850
rect 51724 12786 51776 12792
rect 52000 12844 52052 12850
rect 52000 12786 52052 12792
rect 52196 12782 52224 13126
rect 51632 12776 51684 12782
rect 51632 12718 51684 12724
rect 52184 12776 52236 12782
rect 52184 12718 52236 12724
rect 51552 12600 51764 12628
rect 51552 12406 51672 12434
rect 51552 12374 51580 12406
rect 51540 12368 51592 12374
rect 51540 12310 51592 12316
rect 51644 12238 51672 12406
rect 51736 12374 51764 12600
rect 51724 12368 51776 12374
rect 51724 12310 51776 12316
rect 51632 12232 51684 12238
rect 51264 12174 51316 12180
rect 51354 12200 51410 12209
rect 51632 12174 51684 12180
rect 51354 12135 51410 12144
rect 51170 11928 51226 11937
rect 51170 11863 51226 11872
rect 51264 11688 51316 11694
rect 51184 11636 51264 11642
rect 51184 11630 51316 11636
rect 51184 11614 51304 11630
rect 51184 11558 51212 11614
rect 51172 11552 51224 11558
rect 51172 11494 51224 11500
rect 51264 11552 51316 11558
rect 51264 11494 51316 11500
rect 51276 11150 51304 11494
rect 51736 11150 51764 12310
rect 52184 12300 52236 12306
rect 52184 12242 52236 12248
rect 52000 12096 52052 12102
rect 52000 12038 52052 12044
rect 51908 11756 51960 11762
rect 51908 11698 51960 11704
rect 51816 11348 51868 11354
rect 51816 11290 51868 11296
rect 51264 11144 51316 11150
rect 51264 11086 51316 11092
rect 51724 11144 51776 11150
rect 51724 11086 51776 11092
rect 51356 11076 51408 11082
rect 51356 11018 51408 11024
rect 51264 9988 51316 9994
rect 51264 9930 51316 9936
rect 51276 9466 51304 9930
rect 51368 9654 51396 11018
rect 51828 11014 51856 11290
rect 51920 11218 51948 11698
rect 52012 11354 52040 12038
rect 52196 11762 52224 12242
rect 52288 11830 52316 13738
rect 52380 13530 52408 13874
rect 53656 13728 53708 13734
rect 53656 13670 53708 13676
rect 52368 13524 52420 13530
rect 52368 13466 52420 13472
rect 53668 13258 53696 13670
rect 53656 13252 53708 13258
rect 53656 13194 53708 13200
rect 53760 12986 53788 13874
rect 53852 13802 53880 14991
rect 54220 14618 54248 16050
rect 54864 15366 54892 16458
rect 54484 15360 54536 15366
rect 54484 15302 54536 15308
rect 54852 15360 54904 15366
rect 54852 15302 54904 15308
rect 54208 14612 54260 14618
rect 54208 14554 54260 14560
rect 54496 14278 54524 15302
rect 54864 14346 54892 15302
rect 54956 15094 54984 16662
rect 54944 15088 54996 15094
rect 54944 15030 54996 15036
rect 54944 14408 54996 14414
rect 54944 14350 54996 14356
rect 54852 14340 54904 14346
rect 54852 14282 54904 14288
rect 54484 14272 54536 14278
rect 54484 14214 54536 14220
rect 54208 13864 54260 13870
rect 54208 13806 54260 13812
rect 53840 13796 53892 13802
rect 53840 13738 53892 13744
rect 53748 12980 53800 12986
rect 53748 12922 53800 12928
rect 54220 12434 54248 13806
rect 54220 12406 54340 12434
rect 52828 12232 52880 12238
rect 52828 12174 52880 12180
rect 52920 12232 52972 12238
rect 52920 12174 52972 12180
rect 53288 12232 53340 12238
rect 53288 12174 53340 12180
rect 52368 12096 52420 12102
rect 52368 12038 52420 12044
rect 52276 11824 52328 11830
rect 52276 11766 52328 11772
rect 52380 11762 52408 12038
rect 52840 11898 52868 12174
rect 52828 11892 52880 11898
rect 52828 11834 52880 11840
rect 52932 11762 52960 12174
rect 52184 11756 52236 11762
rect 52184 11698 52236 11704
rect 52368 11756 52420 11762
rect 52368 11698 52420 11704
rect 52920 11756 52972 11762
rect 52920 11698 52972 11704
rect 53012 11756 53064 11762
rect 53012 11698 53064 11704
rect 52276 11688 52328 11694
rect 52276 11630 52328 11636
rect 52288 11558 52316 11630
rect 52932 11626 52960 11698
rect 52920 11620 52972 11626
rect 52920 11562 52972 11568
rect 53024 11558 53052 11698
rect 52276 11552 52328 11558
rect 52276 11494 52328 11500
rect 53012 11552 53064 11558
rect 53012 11494 53064 11500
rect 52000 11348 52052 11354
rect 52000 11290 52052 11296
rect 52368 11280 52420 11286
rect 52368 11222 52420 11228
rect 51908 11212 51960 11218
rect 51908 11154 51960 11160
rect 51816 11008 51868 11014
rect 51816 10950 51868 10956
rect 52184 10464 52236 10470
rect 52184 10406 52236 10412
rect 52276 10464 52328 10470
rect 52276 10406 52328 10412
rect 51356 9648 51408 9654
rect 51356 9590 51408 9596
rect 52196 9586 52224 10406
rect 52288 10130 52316 10406
rect 52276 10124 52328 10130
rect 52276 10066 52328 10072
rect 52380 9738 52408 11222
rect 53024 11082 53052 11494
rect 52736 11076 52788 11082
rect 52736 11018 52788 11024
rect 53012 11076 53064 11082
rect 53012 11018 53064 11024
rect 52552 9988 52604 9994
rect 52552 9930 52604 9936
rect 52564 9897 52592 9930
rect 52550 9888 52606 9897
rect 52550 9823 52606 9832
rect 52380 9710 52500 9738
rect 52472 9586 52500 9710
rect 51448 9580 51500 9586
rect 51448 9522 51500 9528
rect 52184 9580 52236 9586
rect 52184 9522 52236 9528
rect 52276 9580 52328 9586
rect 52276 9522 52328 9528
rect 52460 9580 52512 9586
rect 52460 9522 52512 9528
rect 51356 9512 51408 9518
rect 51276 9460 51356 9466
rect 51276 9454 51408 9460
rect 51276 9438 51396 9454
rect 51368 8906 51396 9438
rect 51460 8974 51488 9522
rect 52288 9160 52316 9522
rect 52104 9132 52316 9160
rect 51448 8968 51500 8974
rect 51448 8910 51500 8916
rect 51356 8900 51408 8906
rect 51356 8842 51408 8848
rect 51632 8832 51684 8838
rect 51632 8774 51684 8780
rect 51644 8566 51672 8774
rect 52104 8566 52132 9132
rect 52460 9104 52512 9110
rect 52380 9052 52460 9058
rect 52380 9046 52512 9052
rect 52380 9030 52500 9046
rect 52276 8968 52328 8974
rect 52276 8910 52328 8916
rect 51632 8560 51684 8566
rect 51632 8502 51684 8508
rect 52092 8560 52144 8566
rect 52092 8502 52144 8508
rect 52184 8560 52236 8566
rect 52184 8502 52236 8508
rect 51448 8288 51500 8294
rect 51448 8230 51500 8236
rect 51078 7984 51134 7993
rect 51078 7919 51134 7928
rect 50436 7812 50488 7818
rect 50436 7754 50488 7760
rect 50988 7812 51040 7818
rect 50988 7754 51040 7760
rect 50344 7540 50396 7546
rect 50344 7482 50396 7488
rect 49700 7472 49752 7478
rect 49700 7414 49752 7420
rect 49516 7404 49568 7410
rect 49516 7346 49568 7352
rect 49332 7336 49384 7342
rect 49332 7278 49384 7284
rect 49146 7168 49202 7177
rect 49146 7103 49202 7112
rect 48780 6860 48832 6866
rect 48780 6802 48832 6808
rect 49528 6798 49556 7346
rect 49608 6996 49660 7002
rect 49608 6938 49660 6944
rect 49516 6792 49568 6798
rect 49516 6734 49568 6740
rect 49620 6746 49648 6938
rect 50356 6905 50384 7482
rect 50342 6896 50398 6905
rect 50068 6860 50120 6866
rect 51000 6866 51028 7754
rect 51092 7585 51120 7919
rect 51460 7886 51488 8230
rect 52196 8090 52224 8502
rect 52184 8084 52236 8090
rect 52012 8044 52184 8072
rect 51172 7880 51224 7886
rect 51170 7848 51172 7857
rect 51448 7880 51500 7886
rect 51224 7848 51226 7857
rect 51448 7822 51500 7828
rect 51722 7848 51778 7857
rect 51170 7783 51226 7792
rect 51356 7812 51408 7818
rect 51722 7783 51778 7792
rect 51816 7812 51868 7818
rect 51356 7754 51408 7760
rect 51078 7576 51134 7585
rect 51368 7546 51396 7754
rect 51078 7511 51134 7520
rect 51356 7540 51408 7546
rect 51356 7482 51408 7488
rect 51632 7336 51684 7342
rect 51632 7278 51684 7284
rect 50342 6831 50344 6840
rect 50068 6802 50120 6808
rect 50396 6831 50398 6840
rect 50988 6860 51040 6866
rect 50344 6802 50396 6808
rect 50988 6802 51040 6808
rect 49148 6724 49200 6730
rect 49148 6666 49200 6672
rect 47823 6556 48131 6565
rect 47823 6554 47829 6556
rect 47885 6554 47909 6556
rect 47965 6554 47989 6556
rect 48045 6554 48069 6556
rect 48125 6554 48131 6556
rect 47885 6502 47887 6554
rect 48067 6502 48069 6554
rect 47823 6500 47829 6502
rect 47885 6500 47909 6502
rect 47965 6500 47989 6502
rect 48045 6500 48069 6502
rect 48125 6500 48131 6502
rect 47823 6491 48131 6500
rect 48226 6488 48282 6497
rect 48136 6452 48188 6458
rect 48188 6432 48226 6440
rect 48188 6423 48282 6432
rect 48688 6452 48740 6458
rect 48188 6412 48268 6423
rect 48136 6394 48188 6400
rect 48688 6394 48740 6400
rect 48044 6384 48096 6390
rect 48320 6384 48372 6390
rect 48044 6326 48096 6332
rect 48240 6344 48320 6372
rect 48056 5914 48084 6326
rect 48240 6254 48268 6344
rect 48320 6326 48372 6332
rect 48228 6248 48280 6254
rect 48228 6190 48280 6196
rect 48044 5908 48096 5914
rect 48044 5850 48096 5856
rect 48240 5778 48268 6190
rect 48320 6112 48372 6118
rect 48320 6054 48372 6060
rect 48332 5817 48360 6054
rect 48318 5808 48374 5817
rect 48228 5772 48280 5778
rect 48318 5743 48374 5752
rect 48228 5714 48280 5720
rect 48700 5710 48728 6394
rect 49160 6322 49188 6666
rect 49528 6458 49556 6734
rect 49620 6718 49924 6746
rect 49700 6656 49752 6662
rect 49700 6598 49752 6604
rect 49516 6452 49568 6458
rect 49516 6394 49568 6400
rect 48780 6316 48832 6322
rect 48780 6258 48832 6264
rect 49148 6316 49200 6322
rect 49148 6258 49200 6264
rect 48792 6118 48820 6258
rect 48780 6112 48832 6118
rect 48780 6054 48832 6060
rect 47676 5704 47728 5710
rect 47676 5646 47728 5652
rect 48688 5704 48740 5710
rect 48688 5646 48740 5652
rect 47124 5102 47176 5108
rect 47490 5128 47546 5137
rect 47136 4622 47164 5102
rect 47688 5098 47716 5646
rect 47823 5468 48131 5477
rect 47823 5466 47829 5468
rect 47885 5466 47909 5468
rect 47965 5466 47989 5468
rect 48045 5466 48069 5468
rect 48125 5466 48131 5468
rect 47885 5414 47887 5466
rect 48067 5414 48069 5466
rect 47823 5412 47829 5414
rect 47885 5412 47909 5414
rect 47965 5412 47989 5414
rect 48045 5412 48069 5414
rect 48125 5412 48131 5414
rect 47823 5403 48131 5412
rect 47768 5296 47820 5302
rect 47768 5238 47820 5244
rect 47490 5063 47546 5072
rect 47676 5092 47728 5098
rect 47676 5034 47728 5040
rect 47582 4992 47638 5001
rect 47582 4927 47638 4936
rect 47124 4616 47176 4622
rect 47124 4558 47176 4564
rect 47490 4584 47546 4593
rect 47400 4548 47452 4554
rect 47490 4519 47546 4528
rect 47400 4490 47452 4496
rect 45928 4480 45980 4486
rect 45928 4422 45980 4428
rect 43996 4276 44048 4282
rect 43996 4218 44048 4224
rect 41788 4140 41840 4146
rect 41788 4082 41840 4088
rect 43812 4140 43864 4146
rect 43812 4082 43864 4088
rect 40684 4072 40736 4078
rect 40684 4014 40736 4020
rect 40776 4072 40828 4078
rect 40776 4014 40828 4020
rect 40592 3936 40644 3942
rect 40592 3878 40644 3884
rect 40604 3738 40632 3878
rect 40592 3732 40644 3738
rect 40592 3674 40644 3680
rect 40788 3670 40816 4014
rect 47412 4010 47440 4490
rect 47504 4486 47532 4519
rect 47596 4486 47624 4927
rect 47780 4622 47808 5238
rect 48136 5228 48188 5234
rect 48136 5170 48188 5176
rect 48148 4826 48176 5170
rect 48700 5166 48728 5646
rect 49160 5574 49188 6258
rect 49608 6180 49660 6186
rect 49608 6122 49660 6128
rect 49514 5944 49570 5953
rect 49514 5879 49516 5888
rect 49568 5879 49570 5888
rect 49516 5850 49568 5856
rect 49620 5710 49648 6122
rect 49712 5846 49740 6598
rect 49896 6390 49924 6718
rect 49884 6384 49936 6390
rect 49884 6326 49936 6332
rect 50080 6322 50108 6802
rect 51644 6662 51672 7278
rect 51632 6656 51684 6662
rect 51632 6598 51684 6604
rect 51736 6497 51764 7783
rect 51816 7754 51868 7760
rect 51828 7274 51856 7754
rect 51908 7744 51960 7750
rect 51908 7686 51960 7692
rect 51816 7268 51868 7274
rect 51816 7210 51868 7216
rect 51920 6934 51948 7686
rect 51908 6928 51960 6934
rect 51908 6870 51960 6876
rect 51722 6488 51778 6497
rect 50160 6452 50212 6458
rect 51722 6423 51778 6432
rect 50160 6394 50212 6400
rect 50068 6316 50120 6322
rect 50068 6258 50120 6264
rect 49974 6080 50030 6089
rect 49974 6015 50030 6024
rect 49792 5908 49844 5914
rect 49792 5850 49844 5856
rect 49700 5840 49752 5846
rect 49700 5782 49752 5788
rect 49516 5704 49568 5710
rect 49516 5646 49568 5652
rect 49608 5704 49660 5710
rect 49608 5646 49660 5652
rect 49148 5568 49200 5574
rect 49148 5510 49200 5516
rect 49528 5386 49556 5646
rect 49528 5358 49648 5386
rect 49620 5302 49648 5358
rect 49608 5296 49660 5302
rect 49608 5238 49660 5244
rect 48688 5160 48740 5166
rect 48688 5102 48740 5108
rect 49620 5098 49648 5238
rect 49608 5092 49660 5098
rect 49608 5034 49660 5040
rect 48228 5024 48280 5030
rect 49424 5024 49476 5030
rect 48280 4984 48360 5012
rect 48228 4966 48280 4972
rect 48136 4820 48188 4826
rect 48136 4762 48188 4768
rect 47768 4616 47820 4622
rect 47768 4558 47820 4564
rect 47492 4480 47544 4486
rect 47492 4422 47544 4428
rect 47584 4480 47636 4486
rect 47584 4422 47636 4428
rect 47823 4380 48131 4389
rect 47823 4378 47829 4380
rect 47885 4378 47909 4380
rect 47965 4378 47989 4380
rect 48045 4378 48069 4380
rect 48125 4378 48131 4380
rect 47885 4326 47887 4378
rect 48067 4326 48069 4378
rect 47823 4324 47829 4326
rect 47885 4324 47909 4326
rect 47965 4324 47989 4326
rect 48045 4324 48069 4326
rect 48125 4324 48131 4326
rect 47823 4315 48131 4324
rect 48332 4078 48360 4984
rect 49424 4966 49476 4972
rect 49436 4486 49464 4966
rect 49620 4826 49648 5034
rect 49804 5030 49832 5850
rect 49792 5024 49844 5030
rect 49792 4966 49844 4972
rect 49608 4820 49660 4826
rect 49608 4762 49660 4768
rect 49988 4690 50016 6015
rect 50068 5636 50120 5642
rect 50068 5578 50120 5584
rect 50080 5234 50108 5578
rect 50172 5234 50200 6394
rect 51448 6248 51500 6254
rect 51448 6190 51500 6196
rect 50712 6112 50764 6118
rect 50712 6054 50764 6060
rect 51356 6112 51408 6118
rect 51356 6054 51408 6060
rect 50724 5710 50752 6054
rect 50802 5944 50858 5953
rect 50802 5879 50804 5888
rect 50856 5879 50858 5888
rect 50804 5850 50856 5856
rect 51368 5846 51396 6054
rect 51460 5914 51488 6190
rect 51736 5914 51764 6423
rect 51448 5908 51500 5914
rect 51448 5850 51500 5856
rect 51724 5908 51776 5914
rect 51724 5850 51776 5856
rect 51356 5840 51408 5846
rect 51356 5782 51408 5788
rect 51540 5772 51592 5778
rect 51540 5714 51592 5720
rect 50252 5704 50304 5710
rect 50252 5646 50304 5652
rect 50620 5704 50672 5710
rect 50620 5646 50672 5652
rect 50712 5704 50764 5710
rect 50712 5646 50764 5652
rect 50264 5574 50292 5646
rect 50252 5568 50304 5574
rect 50252 5510 50304 5516
rect 50068 5228 50120 5234
rect 50068 5170 50120 5176
rect 50160 5228 50212 5234
rect 50160 5170 50212 5176
rect 50080 4758 50108 5170
rect 50344 5160 50396 5166
rect 50632 5137 50660 5646
rect 51172 5160 51224 5166
rect 50344 5102 50396 5108
rect 50618 5128 50674 5137
rect 50356 4826 50384 5102
rect 51172 5102 51224 5108
rect 50618 5063 50674 5072
rect 50632 4826 50660 5063
rect 51184 5001 51212 5102
rect 51552 5001 51580 5714
rect 52012 5302 52040 8044
rect 52184 8026 52236 8032
rect 52092 7744 52144 7750
rect 52092 7686 52144 7692
rect 52104 7410 52132 7686
rect 52288 7546 52316 8910
rect 52380 8430 52408 9030
rect 52368 8424 52420 8430
rect 52368 8366 52420 8372
rect 52276 7540 52328 7546
rect 52276 7482 52328 7488
rect 52092 7404 52144 7410
rect 52092 7346 52144 7352
rect 52184 7336 52236 7342
rect 52288 7324 52316 7482
rect 52236 7296 52316 7324
rect 52184 7278 52236 7284
rect 52092 7268 52144 7274
rect 52092 7210 52144 7216
rect 52000 5296 52052 5302
rect 52000 5238 52052 5244
rect 52000 5024 52052 5030
rect 51170 4992 51226 5001
rect 51170 4927 51226 4936
rect 51538 4992 51594 5001
rect 52104 5012 52132 7210
rect 52276 6316 52328 6322
rect 52276 6258 52328 6264
rect 52288 5574 52316 6258
rect 52276 5568 52328 5574
rect 52276 5510 52328 5516
rect 52184 5296 52236 5302
rect 52184 5238 52236 5244
rect 52052 4984 52132 5012
rect 52000 4966 52052 4972
rect 51538 4927 51594 4936
rect 50344 4820 50396 4826
rect 50344 4762 50396 4768
rect 50620 4820 50672 4826
rect 50620 4762 50672 4768
rect 50068 4752 50120 4758
rect 50068 4694 50120 4700
rect 49976 4684 50028 4690
rect 49976 4626 50028 4632
rect 49792 4548 49844 4554
rect 49792 4490 49844 4496
rect 49424 4480 49476 4486
rect 49424 4422 49476 4428
rect 48320 4072 48372 4078
rect 48320 4014 48372 4020
rect 49148 4072 49200 4078
rect 49148 4014 49200 4020
rect 47400 4004 47452 4010
rect 47400 3946 47452 3952
rect 49160 3942 49188 4014
rect 49148 3936 49200 3942
rect 49148 3878 49200 3884
rect 49804 3670 49832 4490
rect 50356 4128 50384 4762
rect 51552 4554 51580 4927
rect 52012 4622 52040 4966
rect 52000 4616 52052 4622
rect 51998 4584 52000 4593
rect 52052 4584 52054 4593
rect 51540 4548 51592 4554
rect 51998 4519 52054 4528
rect 51540 4490 51592 4496
rect 51552 4282 51580 4490
rect 51540 4276 51592 4282
rect 51540 4218 51592 4224
rect 52196 4214 52224 5238
rect 52288 4690 52316 5510
rect 52380 4826 52408 8366
rect 52564 5914 52592 9823
rect 52644 8424 52696 8430
rect 52644 8366 52696 8372
rect 52656 7954 52684 8366
rect 52748 7954 52776 11018
rect 53024 9994 53052 11018
rect 53300 10849 53328 12174
rect 54312 12170 54340 12406
rect 54208 12164 54260 12170
rect 54208 12106 54260 12112
rect 54300 12164 54352 12170
rect 54300 12106 54352 12112
rect 53748 11892 53800 11898
rect 53748 11834 53800 11840
rect 53656 11552 53708 11558
rect 53656 11494 53708 11500
rect 53668 11286 53696 11494
rect 53472 11280 53524 11286
rect 53392 11240 53472 11268
rect 53286 10840 53342 10849
rect 53286 10775 53342 10784
rect 53300 10674 53328 10775
rect 53288 10668 53340 10674
rect 53288 10610 53340 10616
rect 53104 10600 53156 10606
rect 53104 10542 53156 10548
rect 53012 9988 53064 9994
rect 53012 9930 53064 9936
rect 53116 9654 53144 10542
rect 53300 10418 53328 10610
rect 53392 10538 53420 11240
rect 53472 11222 53524 11228
rect 53656 11280 53708 11286
rect 53656 11222 53708 11228
rect 53564 11212 53616 11218
rect 53564 11154 53616 11160
rect 53576 11014 53604 11154
rect 53564 11008 53616 11014
rect 53564 10950 53616 10956
rect 53576 10674 53604 10950
rect 53654 10840 53710 10849
rect 53654 10775 53710 10784
rect 53472 10668 53524 10674
rect 53472 10610 53524 10616
rect 53564 10668 53616 10674
rect 53564 10610 53616 10616
rect 53380 10532 53432 10538
rect 53380 10474 53432 10480
rect 53208 10390 53328 10418
rect 53104 9648 53156 9654
rect 53104 9590 53156 9596
rect 53208 8616 53236 10390
rect 53286 10296 53342 10305
rect 53286 10231 53288 10240
rect 53340 10231 53342 10240
rect 53288 10202 53340 10208
rect 53392 10146 53420 10474
rect 53484 10266 53512 10610
rect 53668 10266 53696 10775
rect 53760 10674 53788 11834
rect 54220 11014 54248 12106
rect 54312 11830 54340 12106
rect 54496 12102 54524 14214
rect 54864 13977 54892 14282
rect 54850 13968 54906 13977
rect 54956 13938 54984 14350
rect 54850 13903 54906 13912
rect 54944 13932 54996 13938
rect 54864 12782 54892 13903
rect 54944 13874 54996 13880
rect 55140 13818 55168 16730
rect 55956 16652 56008 16658
rect 55956 16594 56008 16600
rect 55220 16448 55272 16454
rect 55220 16390 55272 16396
rect 55232 14958 55260 16390
rect 55864 16176 55916 16182
rect 55864 16118 55916 16124
rect 55312 15972 55364 15978
rect 55312 15914 55364 15920
rect 55220 14952 55272 14958
rect 55220 14894 55272 14900
rect 54956 13790 55168 13818
rect 54852 12776 54904 12782
rect 54852 12718 54904 12724
rect 54484 12096 54536 12102
rect 54484 12038 54536 12044
rect 54300 11824 54352 11830
rect 54300 11766 54352 11772
rect 54864 11762 54892 12718
rect 54852 11756 54904 11762
rect 54852 11698 54904 11704
rect 54668 11280 54720 11286
rect 54666 11248 54668 11257
rect 54760 11280 54812 11286
rect 54720 11248 54722 11257
rect 54392 11212 54444 11218
rect 54444 11172 54616 11200
rect 54760 11222 54812 11228
rect 54666 11183 54722 11192
rect 54392 11154 54444 11160
rect 54588 11098 54616 11172
rect 54668 11144 54720 11150
rect 54588 11092 54668 11098
rect 54588 11086 54720 11092
rect 54392 11076 54444 11082
rect 54588 11070 54708 11086
rect 54392 11018 54444 11024
rect 54208 11008 54260 11014
rect 53838 10976 53894 10985
rect 54208 10950 54260 10956
rect 53838 10911 53894 10920
rect 53748 10668 53800 10674
rect 53748 10610 53800 10616
rect 53472 10260 53524 10266
rect 53472 10202 53524 10208
rect 53656 10260 53708 10266
rect 53656 10202 53708 10208
rect 53288 10124 53340 10130
rect 53392 10118 53604 10146
rect 53288 10066 53340 10072
rect 53300 9586 53328 10066
rect 53380 10056 53432 10062
rect 53380 9998 53432 10004
rect 53288 9580 53340 9586
rect 53288 9522 53340 9528
rect 53208 8588 53328 8616
rect 53196 8492 53248 8498
rect 53196 8434 53248 8440
rect 53208 8090 53236 8434
rect 53196 8084 53248 8090
rect 53196 8026 53248 8032
rect 52644 7948 52696 7954
rect 52644 7890 52696 7896
rect 52736 7948 52788 7954
rect 52736 7890 52788 7896
rect 53196 7880 53248 7886
rect 53196 7822 53248 7828
rect 52920 7744 52972 7750
rect 52920 7686 52972 7692
rect 52932 6730 52960 7686
rect 52920 6724 52972 6730
rect 52920 6666 52972 6672
rect 52552 5908 52604 5914
rect 52552 5850 52604 5856
rect 52368 4820 52420 4826
rect 52368 4762 52420 4768
rect 52276 4684 52328 4690
rect 52276 4626 52328 4632
rect 52184 4208 52236 4214
rect 52184 4150 52236 4156
rect 52288 4146 52316 4626
rect 53208 4146 53236 7822
rect 53300 7002 53328 8588
rect 53392 8022 53420 9998
rect 53472 8424 53524 8430
rect 53576 8412 53604 10118
rect 53656 10124 53708 10130
rect 53656 10066 53708 10072
rect 53668 8634 53696 10066
rect 53748 10056 53800 10062
rect 53748 9998 53800 10004
rect 53760 8634 53788 9998
rect 53852 9654 53880 10911
rect 54220 10742 54248 10950
rect 54404 10742 54432 11018
rect 54024 10736 54076 10742
rect 54024 10678 54076 10684
rect 54208 10736 54260 10742
rect 54208 10678 54260 10684
rect 54392 10736 54444 10742
rect 54392 10678 54444 10684
rect 54036 10266 54064 10678
rect 54208 10532 54260 10538
rect 54404 10520 54432 10678
rect 54484 10668 54536 10674
rect 54484 10610 54536 10616
rect 54260 10492 54432 10520
rect 54208 10474 54260 10480
rect 54496 10305 54524 10610
rect 54576 10600 54628 10606
rect 54576 10542 54628 10548
rect 54482 10296 54538 10305
rect 54024 10260 54076 10266
rect 54588 10266 54616 10542
rect 54482 10231 54538 10240
rect 54576 10260 54628 10266
rect 54024 10202 54076 10208
rect 54576 10202 54628 10208
rect 54484 9920 54536 9926
rect 54484 9862 54536 9868
rect 53840 9648 53892 9654
rect 53840 9590 53892 9596
rect 53656 8628 53708 8634
rect 53656 8570 53708 8576
rect 53748 8628 53800 8634
rect 53748 8570 53800 8576
rect 53932 8492 53984 8498
rect 53932 8434 53984 8440
rect 53576 8384 53788 8412
rect 53472 8366 53524 8372
rect 53380 8016 53432 8022
rect 53380 7958 53432 7964
rect 53288 6996 53340 7002
rect 53288 6938 53340 6944
rect 53300 5914 53328 6938
rect 53484 6866 53512 8366
rect 53564 7404 53616 7410
rect 53564 7346 53616 7352
rect 53472 6860 53524 6866
rect 53472 6802 53524 6808
rect 53576 6662 53604 7346
rect 53656 7200 53708 7206
rect 53656 7142 53708 7148
rect 53668 6798 53696 7142
rect 53656 6792 53708 6798
rect 53656 6734 53708 6740
rect 53564 6656 53616 6662
rect 53564 6598 53616 6604
rect 53656 6248 53708 6254
rect 53654 6216 53656 6225
rect 53708 6216 53710 6225
rect 53654 6151 53710 6160
rect 53288 5908 53340 5914
rect 53288 5850 53340 5856
rect 53668 5273 53696 6151
rect 53760 5914 53788 8384
rect 53944 7818 53972 8434
rect 53932 7812 53984 7818
rect 53932 7754 53984 7760
rect 54208 7336 54260 7342
rect 54208 7278 54260 7284
rect 54220 7177 54248 7278
rect 54206 7168 54262 7177
rect 54206 7103 54262 7112
rect 53840 6384 53892 6390
rect 53838 6352 53840 6361
rect 53892 6352 53894 6361
rect 53838 6287 53894 6296
rect 53748 5908 53800 5914
rect 53748 5850 53800 5856
rect 53748 5296 53800 5302
rect 53654 5264 53710 5273
rect 53380 5228 53432 5234
rect 53380 5170 53432 5176
rect 53472 5228 53524 5234
rect 53524 5188 53604 5216
rect 53748 5238 53800 5244
rect 53654 5199 53710 5208
rect 53472 5170 53524 5176
rect 53392 4554 53420 5170
rect 53472 5024 53524 5030
rect 53472 4966 53524 4972
rect 53484 4622 53512 4966
rect 53576 4758 53604 5188
rect 53760 4826 53788 5238
rect 53748 4820 53800 4826
rect 53748 4762 53800 4768
rect 53564 4752 53616 4758
rect 53564 4694 53616 4700
rect 53472 4616 53524 4622
rect 53472 4558 53524 4564
rect 53380 4548 53432 4554
rect 53380 4490 53432 4496
rect 50436 4140 50488 4146
rect 50356 4100 50436 4128
rect 50436 4082 50488 4088
rect 51264 4140 51316 4146
rect 51264 4082 51316 4088
rect 52276 4140 52328 4146
rect 52276 4082 52328 4088
rect 53196 4140 53248 4146
rect 53196 4082 53248 4088
rect 51080 3936 51132 3942
rect 51080 3878 51132 3884
rect 51092 3670 51120 3878
rect 40776 3664 40828 3670
rect 40776 3606 40828 3612
rect 49792 3664 49844 3670
rect 49792 3606 49844 3612
rect 51080 3664 51132 3670
rect 51080 3606 51132 3612
rect 40408 3596 40460 3602
rect 40408 3538 40460 3544
rect 38844 3460 38896 3466
rect 38844 3402 38896 3408
rect 38856 3194 38884 3402
rect 39028 3392 39080 3398
rect 39028 3334 39080 3340
rect 37740 3188 37792 3194
rect 37740 3130 37792 3136
rect 38844 3188 38896 3194
rect 38844 3130 38896 3136
rect 36105 2748 36413 2757
rect 36105 2746 36111 2748
rect 36167 2746 36191 2748
rect 36247 2746 36271 2748
rect 36327 2746 36351 2748
rect 36407 2746 36413 2748
rect 36167 2694 36169 2746
rect 36349 2694 36351 2746
rect 36105 2692 36111 2694
rect 36167 2692 36191 2694
rect 36247 2692 36271 2694
rect 36327 2692 36351 2694
rect 36407 2692 36413 2694
rect 36105 2683 36413 2692
rect 37384 2746 37504 2774
rect 37384 2650 37412 2746
rect 38856 2650 38884 3130
rect 39040 3126 39068 3334
rect 39028 3120 39080 3126
rect 39028 3062 39080 3068
rect 40420 3058 40448 3538
rect 41328 3460 41380 3466
rect 41328 3402 41380 3408
rect 40408 3052 40460 3058
rect 40408 2994 40460 3000
rect 41340 2650 41368 3402
rect 47823 3292 48131 3301
rect 47823 3290 47829 3292
rect 47885 3290 47909 3292
rect 47965 3290 47989 3292
rect 48045 3290 48069 3292
rect 48125 3290 48131 3292
rect 47885 3238 47887 3290
rect 48067 3238 48069 3290
rect 47823 3236 47829 3238
rect 47885 3236 47909 3238
rect 47965 3236 47989 3238
rect 48045 3236 48069 3238
rect 48125 3236 48131 3238
rect 47823 3227 48131 3236
rect 51276 3058 51304 4082
rect 52368 3460 52420 3466
rect 52368 3402 52420 3408
rect 53380 3460 53432 3466
rect 53484 3448 53512 4558
rect 53852 3618 53880 6287
rect 53932 6248 53984 6254
rect 53932 6190 53984 6196
rect 53944 4826 53972 6190
rect 53932 4820 53984 4826
rect 53932 4762 53984 4768
rect 54220 3670 54248 7103
rect 54496 5914 54524 9862
rect 54588 6089 54616 10202
rect 54772 10198 54800 11222
rect 54956 11098 54984 13790
rect 55232 13716 55260 14894
rect 55324 13938 55352 15914
rect 55496 15088 55548 15094
rect 55496 15030 55548 15036
rect 55508 14822 55536 15030
rect 55588 14952 55640 14958
rect 55588 14894 55640 14900
rect 55496 14816 55548 14822
rect 55496 14758 55548 14764
rect 55600 14414 55628 14894
rect 55772 14476 55824 14482
rect 55772 14418 55824 14424
rect 55588 14408 55640 14414
rect 55588 14350 55640 14356
rect 55784 14074 55812 14418
rect 55772 14068 55824 14074
rect 55772 14010 55824 14016
rect 55312 13932 55364 13938
rect 55312 13874 55364 13880
rect 55140 13688 55260 13716
rect 55036 12980 55088 12986
rect 55036 12922 55088 12928
rect 55048 12850 55076 12922
rect 55036 12844 55088 12850
rect 55036 12786 55088 12792
rect 55048 11762 55076 12786
rect 55036 11756 55088 11762
rect 55036 11698 55088 11704
rect 55140 11150 55168 13688
rect 55876 13190 55904 16118
rect 55968 15910 55996 16594
rect 56704 16114 56732 16934
rect 57072 16794 57100 17206
rect 59360 17128 59412 17134
rect 59360 17070 59412 17076
rect 61844 17128 61896 17134
rect 61844 17070 61896 17076
rect 63592 17128 63644 17134
rect 63592 17070 63644 17076
rect 65800 17128 65852 17134
rect 65800 17070 65852 17076
rect 57980 17060 58032 17066
rect 57980 17002 58032 17008
rect 57060 16788 57112 16794
rect 57060 16730 57112 16736
rect 56784 16652 56836 16658
rect 56784 16594 56836 16600
rect 56416 16108 56468 16114
rect 56416 16050 56468 16056
rect 56692 16108 56744 16114
rect 56692 16050 56744 16056
rect 56324 16040 56376 16046
rect 56324 15982 56376 15988
rect 55956 15904 56008 15910
rect 55956 15846 56008 15852
rect 55968 14414 55996 15846
rect 56048 15360 56100 15366
rect 56048 15302 56100 15308
rect 55956 14408 56008 14414
rect 55956 14350 56008 14356
rect 55864 13184 55916 13190
rect 55864 13126 55916 13132
rect 55678 13016 55734 13025
rect 55678 12951 55734 12960
rect 55404 12708 55456 12714
rect 55456 12668 55536 12696
rect 55404 12650 55456 12656
rect 55220 12096 55272 12102
rect 55220 12038 55272 12044
rect 55128 11144 55180 11150
rect 54956 11070 55076 11098
rect 55128 11086 55180 11092
rect 54944 11008 54996 11014
rect 54944 10950 54996 10956
rect 54956 10674 54984 10950
rect 54944 10668 54996 10674
rect 54944 10610 54996 10616
rect 54760 10192 54812 10198
rect 54760 10134 54812 10140
rect 54852 10192 54904 10198
rect 54852 10134 54904 10140
rect 54864 9926 54892 10134
rect 54852 9920 54904 9926
rect 54852 9862 54904 9868
rect 54944 8968 54996 8974
rect 54944 8910 54996 8916
rect 54852 7880 54904 7886
rect 54956 7868 54984 8910
rect 54904 7840 54984 7868
rect 54852 7822 54904 7828
rect 54956 7342 54984 7840
rect 54852 7336 54904 7342
rect 54852 7278 54904 7284
rect 54944 7336 54996 7342
rect 54944 7278 54996 7284
rect 54864 7002 54892 7278
rect 54852 6996 54904 7002
rect 54852 6938 54904 6944
rect 55048 6390 55076 11070
rect 55232 9178 55260 12038
rect 55508 10606 55536 12668
rect 55692 12617 55720 12951
rect 55678 12608 55734 12617
rect 55678 12543 55734 12552
rect 55876 12434 55904 13126
rect 55968 12986 55996 14350
rect 56060 14006 56088 15302
rect 56336 14482 56364 15982
rect 56428 15502 56456 16050
rect 56600 15904 56652 15910
rect 56600 15846 56652 15852
rect 56416 15496 56468 15502
rect 56416 15438 56468 15444
rect 56612 15026 56640 15846
rect 56704 15434 56732 16050
rect 56692 15428 56744 15434
rect 56692 15370 56744 15376
rect 56600 15020 56652 15026
rect 56600 14962 56652 14968
rect 56704 14958 56732 15370
rect 56692 14952 56744 14958
rect 56692 14894 56744 14900
rect 56324 14476 56376 14482
rect 56324 14418 56376 14424
rect 56232 14340 56284 14346
rect 56232 14282 56284 14288
rect 56048 14000 56100 14006
rect 56048 13942 56100 13948
rect 56244 13394 56272 14282
rect 56692 14000 56744 14006
rect 56692 13942 56744 13948
rect 56704 13870 56732 13942
rect 56692 13864 56744 13870
rect 56692 13806 56744 13812
rect 56600 13524 56652 13530
rect 56600 13466 56652 13472
rect 56232 13388 56284 13394
rect 56232 13330 56284 13336
rect 56322 13288 56378 13297
rect 56322 13223 56378 13232
rect 55956 12980 56008 12986
rect 55956 12922 56008 12928
rect 56232 12776 56284 12782
rect 56336 12764 56364 13223
rect 56612 12918 56640 13466
rect 56600 12912 56652 12918
rect 56600 12854 56652 12860
rect 56284 12736 56364 12764
rect 56232 12718 56284 12724
rect 56416 12708 56468 12714
rect 56416 12650 56468 12656
rect 55784 12406 55904 12434
rect 56138 12472 56194 12481
rect 56138 12407 56194 12416
rect 55784 12170 55812 12406
rect 56152 12374 56180 12407
rect 56428 12374 56456 12650
rect 56140 12368 56192 12374
rect 56140 12310 56192 12316
rect 56416 12368 56468 12374
rect 56416 12310 56468 12316
rect 55956 12300 56008 12306
rect 55956 12242 56008 12248
rect 55772 12164 55824 12170
rect 55772 12106 55824 12112
rect 55784 10674 55812 12106
rect 55968 11286 55996 12242
rect 56600 12096 56652 12102
rect 56598 12064 56600 12073
rect 56652 12064 56654 12073
rect 56598 11999 56654 12008
rect 56690 11792 56746 11801
rect 56690 11727 56692 11736
rect 56744 11727 56746 11736
rect 56692 11698 56744 11704
rect 56324 11688 56376 11694
rect 56324 11630 56376 11636
rect 56506 11656 56562 11665
rect 56140 11552 56192 11558
rect 56140 11494 56192 11500
rect 55956 11280 56008 11286
rect 55956 11222 56008 11228
rect 56152 11150 56180 11494
rect 56336 11150 56364 11630
rect 56506 11591 56508 11600
rect 56560 11591 56562 11600
rect 56508 11562 56560 11568
rect 56048 11144 56100 11150
rect 56048 11086 56100 11092
rect 56140 11144 56192 11150
rect 56140 11086 56192 11092
rect 56324 11144 56376 11150
rect 56796 11121 56824 16594
rect 56966 15600 57022 15609
rect 56966 15535 57022 15544
rect 56980 14958 57008 15535
rect 57072 15502 57100 16730
rect 57336 16652 57388 16658
rect 57336 16594 57388 16600
rect 57060 15496 57112 15502
rect 57060 15438 57112 15444
rect 56968 14952 57020 14958
rect 56968 14894 57020 14900
rect 57244 14340 57296 14346
rect 57244 14282 57296 14288
rect 57152 13864 57204 13870
rect 57072 13824 57152 13852
rect 56968 13728 57020 13734
rect 56968 13670 57020 13676
rect 56980 13274 57008 13670
rect 56888 13246 57008 13274
rect 56888 12782 56916 13246
rect 56968 13184 57020 13190
rect 56968 13126 57020 13132
rect 56876 12776 56928 12782
rect 56876 12718 56928 12724
rect 56324 11086 56376 11092
rect 56782 11112 56838 11121
rect 55772 10668 55824 10674
rect 55772 10610 55824 10616
rect 55496 10600 55548 10606
rect 55496 10542 55548 10548
rect 55312 10464 55364 10470
rect 55312 10406 55364 10412
rect 55402 10432 55458 10441
rect 55220 9172 55272 9178
rect 55220 9114 55272 9120
rect 55220 8424 55272 8430
rect 55220 8366 55272 8372
rect 55232 6905 55260 8366
rect 55324 7954 55352 10406
rect 55402 10367 55458 10376
rect 55416 8537 55444 10367
rect 55680 10056 55732 10062
rect 55680 9998 55732 10004
rect 55864 10056 55916 10062
rect 55864 9998 55916 10004
rect 55496 9920 55548 9926
rect 55496 9862 55548 9868
rect 55508 8945 55536 9862
rect 55494 8936 55550 8945
rect 55494 8871 55550 8880
rect 55402 8528 55458 8537
rect 55402 8463 55458 8472
rect 55496 8424 55548 8430
rect 55496 8366 55548 8372
rect 55508 8090 55536 8366
rect 55496 8084 55548 8090
rect 55496 8026 55548 8032
rect 55312 7948 55364 7954
rect 55312 7890 55364 7896
rect 55692 7886 55720 9998
rect 55772 9512 55824 9518
rect 55772 9454 55824 9460
rect 55784 9042 55812 9454
rect 55876 9382 55904 9998
rect 56060 9674 56088 11086
rect 56508 11076 56560 11082
rect 56782 11047 56838 11056
rect 56508 11018 56560 11024
rect 56520 10674 56548 11018
rect 56600 10736 56652 10742
rect 56600 10678 56652 10684
rect 56508 10668 56560 10674
rect 56508 10610 56560 10616
rect 56324 10532 56376 10538
rect 56324 10474 56376 10480
rect 56060 9646 56180 9674
rect 56048 9512 56100 9518
rect 56046 9480 56048 9489
rect 56100 9480 56102 9489
rect 56046 9415 56102 9424
rect 55864 9376 55916 9382
rect 55864 9318 55916 9324
rect 55772 9036 55824 9042
rect 55772 8978 55824 8984
rect 55876 8430 55904 9318
rect 55864 8424 55916 8430
rect 55864 8366 55916 8372
rect 55680 7880 55732 7886
rect 55680 7822 55732 7828
rect 55956 7812 56008 7818
rect 55956 7754 56008 7760
rect 55864 7744 55916 7750
rect 55864 7686 55916 7692
rect 55876 7478 55904 7686
rect 55864 7472 55916 7478
rect 55864 7414 55916 7420
rect 55968 7274 55996 7754
rect 55956 7268 56008 7274
rect 55956 7210 56008 7216
rect 55218 6896 55274 6905
rect 55218 6831 55274 6840
rect 55036 6384 55088 6390
rect 55036 6326 55088 6332
rect 54852 6248 54904 6254
rect 54852 6190 54904 6196
rect 54574 6080 54630 6089
rect 54574 6015 54630 6024
rect 54484 5908 54536 5914
rect 54484 5850 54536 5856
rect 54392 5636 54444 5642
rect 54392 5578 54444 5584
rect 54404 5098 54432 5578
rect 54864 5574 54892 6190
rect 55048 5930 55076 6326
rect 55048 5902 55168 5930
rect 54852 5568 54904 5574
rect 54852 5510 54904 5516
rect 55140 5302 55168 5902
rect 55220 5772 55272 5778
rect 55220 5714 55272 5720
rect 55128 5296 55180 5302
rect 55128 5238 55180 5244
rect 54392 5092 54444 5098
rect 54392 5034 54444 5040
rect 55140 4162 55168 5238
rect 55232 5166 55260 5714
rect 55864 5568 55916 5574
rect 55864 5510 55916 5516
rect 55876 5302 55904 5510
rect 56060 5409 56088 9415
rect 56152 9178 56180 9646
rect 56140 9172 56192 9178
rect 56140 9114 56192 9120
rect 56140 6452 56192 6458
rect 56140 6394 56192 6400
rect 56152 5642 56180 6394
rect 56140 5636 56192 5642
rect 56140 5578 56192 5584
rect 56046 5400 56102 5409
rect 56046 5335 56102 5344
rect 55864 5296 55916 5302
rect 55864 5238 55916 5244
rect 56152 5166 56180 5578
rect 55220 5160 55272 5166
rect 55220 5102 55272 5108
rect 56140 5160 56192 5166
rect 56192 5108 56272 5114
rect 56140 5102 56272 5108
rect 56152 5086 56272 5102
rect 56140 5024 56192 5030
rect 56140 4966 56192 4972
rect 56152 4690 56180 4966
rect 56140 4684 56192 4690
rect 56140 4626 56192 4632
rect 55864 4548 55916 4554
rect 56140 4548 56192 4554
rect 55916 4508 56140 4536
rect 55864 4490 55916 4496
rect 56140 4490 56192 4496
rect 54668 4140 54720 4146
rect 54668 4082 54720 4088
rect 55048 4134 55168 4162
rect 55496 4208 55548 4214
rect 55496 4150 55548 4156
rect 54680 3670 54708 4082
rect 54208 3664 54260 3670
rect 53852 3590 53972 3618
rect 54208 3606 54260 3612
rect 54668 3664 54720 3670
rect 54668 3606 54720 3612
rect 53840 3528 53892 3534
rect 53840 3470 53892 3476
rect 53432 3420 53512 3448
rect 53380 3402 53432 3408
rect 52380 3058 52408 3402
rect 53852 3194 53880 3470
rect 53840 3188 53892 3194
rect 53840 3130 53892 3136
rect 53944 3126 53972 3590
rect 55048 3194 55076 4134
rect 55128 4072 55180 4078
rect 55128 4014 55180 4020
rect 55140 3466 55168 4014
rect 55508 3738 55536 4150
rect 55956 4004 56008 4010
rect 55956 3946 56008 3952
rect 55496 3732 55548 3738
rect 55496 3674 55548 3680
rect 55128 3460 55180 3466
rect 55128 3402 55180 3408
rect 55036 3188 55088 3194
rect 55036 3130 55088 3136
rect 53932 3120 53984 3126
rect 53932 3062 53984 3068
rect 55140 3058 55168 3402
rect 51264 3052 51316 3058
rect 51264 2994 51316 3000
rect 52368 3052 52420 3058
rect 52368 2994 52420 3000
rect 55128 3052 55180 3058
rect 55128 2994 55180 3000
rect 55508 2990 55536 3674
rect 55968 3602 55996 3946
rect 56244 3942 56272 5086
rect 56232 3936 56284 3942
rect 56232 3878 56284 3884
rect 55956 3596 56008 3602
rect 55956 3538 56008 3544
rect 55864 3460 55916 3466
rect 55864 3402 55916 3408
rect 55876 3194 55904 3402
rect 56244 3194 56272 3878
rect 55864 3188 55916 3194
rect 55864 3130 55916 3136
rect 56232 3188 56284 3194
rect 56232 3130 56284 3136
rect 54392 2984 54444 2990
rect 54392 2926 54444 2932
rect 55496 2984 55548 2990
rect 55496 2926 55548 2932
rect 54404 2650 54432 2926
rect 37372 2644 37424 2650
rect 37372 2586 37424 2592
rect 38844 2644 38896 2650
rect 38844 2586 38896 2592
rect 41328 2644 41380 2650
rect 41328 2586 41380 2592
rect 54392 2644 54444 2650
rect 54392 2586 54444 2592
rect 56336 2446 56364 10474
rect 56612 10198 56640 10678
rect 56600 10192 56652 10198
rect 56600 10134 56652 10140
rect 56980 10130 57008 13126
rect 57072 12238 57100 13824
rect 57152 13806 57204 13812
rect 57256 13530 57284 14282
rect 57348 14278 57376 16594
rect 57888 15904 57940 15910
rect 57888 15846 57940 15852
rect 57336 14272 57388 14278
rect 57336 14214 57388 14220
rect 57348 13938 57376 14214
rect 57336 13932 57388 13938
rect 57336 13874 57388 13880
rect 57244 13524 57296 13530
rect 57244 13466 57296 13472
rect 57256 13258 57284 13466
rect 57244 13252 57296 13258
rect 57244 13194 57296 13200
rect 57152 12980 57204 12986
rect 57152 12922 57204 12928
rect 57164 12434 57192 12922
rect 57348 12594 57376 13874
rect 57900 13530 57928 15846
rect 57992 15434 58020 17002
rect 58164 16448 58216 16454
rect 58164 16390 58216 16396
rect 59176 16448 59228 16454
rect 59176 16390 59228 16396
rect 57980 15428 58032 15434
rect 57980 15370 58032 15376
rect 57978 14104 58034 14113
rect 57978 14039 58034 14048
rect 57992 14006 58020 14039
rect 57980 14000 58032 14006
rect 57980 13942 58032 13948
rect 57888 13524 57940 13530
rect 57888 13466 57940 13472
rect 57704 12708 57756 12714
rect 57704 12650 57756 12656
rect 57348 12566 57652 12594
rect 57164 12406 57284 12434
rect 57060 12232 57112 12238
rect 57060 12174 57112 12180
rect 56968 10124 57020 10130
rect 56968 10066 57020 10072
rect 56784 10056 56836 10062
rect 56784 9998 56836 10004
rect 56508 9512 56560 9518
rect 56508 9454 56560 9460
rect 56520 8294 56548 9454
rect 56508 8288 56560 8294
rect 56508 8230 56560 8236
rect 56416 7200 56468 7206
rect 56416 7142 56468 7148
rect 56428 6866 56456 7142
rect 56520 6866 56548 8230
rect 56796 6934 56824 9998
rect 57152 9376 57204 9382
rect 57152 9318 57204 9324
rect 57164 7954 57192 9318
rect 57256 8634 57284 12406
rect 57348 11354 57376 12566
rect 57520 12164 57572 12170
rect 57520 12106 57572 12112
rect 57532 11830 57560 12106
rect 57520 11824 57572 11830
rect 57520 11766 57572 11772
rect 57624 11354 57652 12566
rect 57716 12481 57744 12650
rect 57702 12472 57758 12481
rect 57702 12407 57758 12416
rect 57704 12232 57756 12238
rect 57704 12174 57756 12180
rect 57900 12220 57928 13466
rect 58072 12368 58124 12374
rect 58072 12310 58124 12316
rect 57980 12232 58032 12238
rect 57900 12192 57980 12220
rect 57336 11348 57388 11354
rect 57336 11290 57388 11296
rect 57612 11348 57664 11354
rect 57612 11290 57664 11296
rect 57428 11280 57480 11286
rect 57428 11222 57480 11228
rect 57336 11144 57388 11150
rect 57334 11112 57336 11121
rect 57440 11132 57468 11222
rect 57716 11150 57744 12174
rect 57796 11756 57848 11762
rect 57796 11698 57848 11704
rect 57388 11112 57468 11132
rect 57390 11104 57468 11112
rect 57704 11144 57756 11150
rect 57704 11086 57756 11092
rect 57334 11047 57390 11056
rect 57808 10742 57836 11698
rect 57900 11558 57928 12192
rect 57980 12174 58032 12180
rect 58084 12050 58112 12310
rect 57992 12022 58112 12050
rect 57992 11558 58020 12022
rect 57888 11552 57940 11558
rect 57888 11494 57940 11500
rect 57980 11552 58032 11558
rect 57980 11494 58032 11500
rect 57992 11082 58020 11494
rect 58176 11218 58204 16390
rect 59188 16182 59216 16390
rect 59372 16182 59400 17070
rect 60740 16992 60792 16998
rect 60740 16934 60792 16940
rect 61108 16992 61160 16998
rect 61108 16934 61160 16940
rect 59542 16892 59850 16901
rect 59542 16890 59548 16892
rect 59604 16890 59628 16892
rect 59684 16890 59708 16892
rect 59764 16890 59788 16892
rect 59844 16890 59850 16892
rect 59604 16838 59606 16890
rect 59786 16838 59788 16890
rect 59542 16836 59548 16838
rect 59604 16836 59628 16838
rect 59684 16836 59708 16838
rect 59764 16836 59788 16838
rect 59844 16836 59850 16838
rect 59542 16827 59850 16836
rect 59452 16652 59504 16658
rect 59452 16594 59504 16600
rect 59176 16176 59228 16182
rect 59176 16118 59228 16124
rect 59360 16176 59412 16182
rect 59360 16118 59412 16124
rect 58624 15904 58676 15910
rect 58624 15846 58676 15852
rect 58716 15904 58768 15910
rect 58716 15846 58768 15852
rect 58256 14340 58308 14346
rect 58256 14282 58308 14288
rect 58268 14074 58296 14282
rect 58256 14068 58308 14074
rect 58256 14010 58308 14016
rect 58348 14068 58400 14074
rect 58348 14010 58400 14016
rect 58256 12640 58308 12646
rect 58360 12628 58388 14010
rect 58440 13388 58492 13394
rect 58440 13330 58492 13336
rect 58452 12714 58480 13330
rect 58440 12708 58492 12714
rect 58440 12650 58492 12656
rect 58308 12600 58388 12628
rect 58256 12582 58308 12588
rect 58360 12322 58388 12600
rect 58268 12294 58388 12322
rect 58268 11762 58296 12294
rect 58348 12232 58400 12238
rect 58348 12174 58400 12180
rect 58256 11756 58308 11762
rect 58256 11698 58308 11704
rect 58164 11212 58216 11218
rect 58164 11154 58216 11160
rect 57980 11076 58032 11082
rect 57980 11018 58032 11024
rect 58256 11076 58308 11082
rect 58256 11018 58308 11024
rect 57796 10736 57848 10742
rect 58268 10713 58296 11018
rect 57796 10678 57848 10684
rect 58254 10704 58310 10713
rect 57336 10668 57388 10674
rect 57336 10610 57388 10616
rect 57348 10266 57376 10610
rect 57428 10600 57480 10606
rect 57428 10542 57480 10548
rect 57336 10260 57388 10266
rect 57336 10202 57388 10208
rect 57440 10169 57468 10542
rect 57426 10160 57482 10169
rect 57426 10095 57482 10104
rect 57808 9926 57836 10678
rect 58254 10639 58310 10648
rect 57796 9920 57848 9926
rect 57796 9862 57848 9868
rect 58072 9580 58124 9586
rect 58124 9540 58204 9568
rect 58072 9522 58124 9528
rect 58176 9178 58204 9540
rect 57888 9172 57940 9178
rect 57888 9114 57940 9120
rect 58164 9172 58216 9178
rect 58164 9114 58216 9120
rect 57900 8974 57928 9114
rect 57888 8968 57940 8974
rect 57610 8936 57666 8945
rect 57888 8910 57940 8916
rect 57610 8871 57612 8880
rect 57664 8871 57666 8880
rect 57612 8842 57664 8848
rect 57244 8628 57296 8634
rect 57244 8570 57296 8576
rect 58176 8498 58204 9114
rect 58164 8492 58216 8498
rect 58164 8434 58216 8440
rect 57244 8288 57296 8294
rect 57244 8230 57296 8236
rect 57152 7948 57204 7954
rect 57152 7890 57204 7896
rect 57256 7410 57284 8230
rect 57704 8016 57756 8022
rect 57704 7958 57756 7964
rect 57336 7948 57388 7954
rect 57336 7890 57388 7896
rect 57348 7857 57376 7890
rect 57334 7848 57390 7857
rect 57334 7783 57390 7792
rect 57716 7546 57744 7958
rect 57704 7540 57756 7546
rect 57704 7482 57756 7488
rect 58070 7440 58126 7449
rect 57244 7404 57296 7410
rect 58070 7375 58072 7384
rect 57244 7346 57296 7352
rect 58124 7375 58126 7384
rect 58072 7346 58124 7352
rect 56784 6928 56836 6934
rect 56784 6870 56836 6876
rect 56416 6860 56468 6866
rect 56416 6802 56468 6808
rect 56508 6860 56560 6866
rect 56508 6802 56560 6808
rect 56692 5704 56744 5710
rect 56692 5646 56744 5652
rect 56600 5296 56652 5302
rect 56600 5238 56652 5244
rect 56612 4826 56640 5238
rect 56704 5216 56732 5646
rect 56796 5574 56824 6870
rect 57256 6798 57284 7346
rect 57244 6792 57296 6798
rect 56966 6760 57022 6769
rect 57244 6734 57296 6740
rect 56966 6695 56968 6704
rect 57020 6695 57022 6704
rect 56968 6666 57020 6672
rect 57888 6316 57940 6322
rect 57888 6258 57940 6264
rect 57704 6248 57756 6254
rect 57704 6190 57756 6196
rect 56968 6112 57020 6118
rect 56968 6054 57020 6060
rect 57152 6112 57204 6118
rect 57152 6054 57204 6060
rect 56980 5710 57008 6054
rect 57164 5817 57192 6054
rect 57150 5808 57206 5817
rect 57150 5743 57206 5752
rect 56968 5704 57020 5710
rect 56968 5646 57020 5652
rect 57244 5704 57296 5710
rect 57244 5646 57296 5652
rect 56784 5568 56836 5574
rect 56784 5510 56836 5516
rect 56784 5228 56836 5234
rect 56704 5188 56784 5216
rect 56784 5170 56836 5176
rect 57060 5228 57112 5234
rect 57060 5170 57112 5176
rect 56796 5137 56824 5170
rect 56782 5128 56838 5137
rect 56782 5063 56838 5072
rect 56692 5024 56744 5030
rect 56690 4992 56692 5001
rect 56744 4992 56746 5001
rect 56690 4927 56746 4936
rect 56600 4820 56652 4826
rect 56600 4762 56652 4768
rect 56416 4616 56468 4622
rect 56416 4558 56468 4564
rect 56428 4214 56456 4558
rect 56416 4208 56468 4214
rect 56416 4150 56468 4156
rect 56796 3194 56824 5063
rect 57072 4826 57100 5170
rect 57060 4820 57112 4826
rect 57060 4762 57112 4768
rect 57256 4622 57284 5646
rect 57716 5642 57744 6190
rect 57900 5642 57928 6258
rect 57704 5636 57756 5642
rect 57704 5578 57756 5584
rect 57888 5636 57940 5642
rect 57888 5578 57940 5584
rect 57716 5234 57744 5578
rect 57900 5302 57928 5578
rect 57888 5296 57940 5302
rect 57888 5238 57940 5244
rect 57336 5228 57388 5234
rect 57336 5170 57388 5176
rect 57704 5228 57756 5234
rect 57704 5170 57756 5176
rect 57348 5098 57376 5170
rect 57336 5092 57388 5098
rect 57336 5034 57388 5040
rect 57244 4616 57296 4622
rect 57336 4616 57388 4622
rect 57244 4558 57296 4564
rect 57334 4584 57336 4593
rect 57388 4584 57390 4593
rect 57334 4519 57390 4528
rect 57704 4548 57756 4554
rect 57704 4490 57756 4496
rect 57888 4548 57940 4554
rect 57888 4490 57940 4496
rect 57716 4282 57744 4490
rect 57796 4480 57848 4486
rect 57796 4422 57848 4428
rect 57704 4276 57756 4282
rect 57704 4218 57756 4224
rect 57060 4072 57112 4078
rect 57060 4014 57112 4020
rect 57072 3942 57100 4014
rect 57808 4010 57836 4422
rect 57900 4146 57928 4490
rect 58084 4146 58112 7346
rect 58176 4826 58204 8434
rect 58256 8424 58308 8430
rect 58256 8366 58308 8372
rect 58268 6458 58296 8366
rect 58360 7750 58388 12174
rect 58532 12164 58584 12170
rect 58532 12106 58584 12112
rect 58544 11762 58572 12106
rect 58636 12050 58664 15846
rect 58728 12850 58756 15846
rect 59082 15192 59138 15201
rect 59082 15127 59138 15136
rect 59096 15094 59124 15127
rect 59084 15088 59136 15094
rect 59084 15030 59136 15036
rect 58808 14816 58860 14822
rect 58808 14758 58860 14764
rect 58716 12844 58768 12850
rect 58716 12786 58768 12792
rect 58728 12238 58756 12786
rect 58716 12232 58768 12238
rect 58716 12174 58768 12180
rect 58714 12064 58770 12073
rect 58636 12022 58714 12050
rect 58714 11999 58770 12008
rect 58728 11762 58756 11999
rect 58820 11898 58848 14758
rect 59188 14634 59216 16118
rect 59464 14822 59492 16594
rect 59912 16584 59964 16590
rect 59912 16526 59964 16532
rect 59542 15804 59850 15813
rect 59542 15802 59548 15804
rect 59604 15802 59628 15804
rect 59684 15802 59708 15804
rect 59764 15802 59788 15804
rect 59844 15802 59850 15804
rect 59604 15750 59606 15802
rect 59786 15750 59788 15802
rect 59542 15748 59548 15750
rect 59604 15748 59628 15750
rect 59684 15748 59708 15750
rect 59764 15748 59788 15750
rect 59844 15748 59850 15750
rect 59542 15739 59850 15748
rect 59924 15502 59952 16526
rect 60004 16448 60056 16454
rect 60004 16390 60056 16396
rect 60096 16448 60148 16454
rect 60096 16390 60148 16396
rect 60016 16182 60044 16390
rect 60004 16176 60056 16182
rect 60004 16118 60056 16124
rect 60108 16114 60136 16390
rect 60096 16108 60148 16114
rect 60096 16050 60148 16056
rect 60752 16046 60780 16934
rect 61120 16726 61148 16934
rect 61108 16720 61160 16726
rect 61108 16662 61160 16668
rect 60832 16584 60884 16590
rect 60832 16526 60884 16532
rect 60740 16040 60792 16046
rect 60740 15982 60792 15988
rect 60844 15858 60872 16526
rect 60752 15830 60872 15858
rect 60280 15632 60332 15638
rect 60280 15574 60332 15580
rect 59912 15496 59964 15502
rect 59912 15438 59964 15444
rect 59924 15162 59952 15438
rect 60096 15360 60148 15366
rect 60096 15302 60148 15308
rect 59912 15156 59964 15162
rect 59912 15098 59964 15104
rect 59452 14816 59504 14822
rect 59452 14758 59504 14764
rect 59188 14606 59400 14634
rect 59372 14550 59400 14606
rect 59268 14544 59320 14550
rect 59268 14486 59320 14492
rect 59360 14544 59412 14550
rect 59360 14486 59412 14492
rect 58992 14408 59044 14414
rect 58992 14350 59044 14356
rect 59004 13394 59032 14350
rect 59280 14006 59308 14486
rect 59268 14000 59320 14006
rect 59174 13968 59230 13977
rect 59268 13942 59320 13948
rect 59464 13938 59492 14758
rect 59542 14716 59850 14725
rect 59542 14714 59548 14716
rect 59604 14714 59628 14716
rect 59684 14714 59708 14716
rect 59764 14714 59788 14716
rect 59844 14714 59850 14716
rect 59604 14662 59606 14714
rect 59786 14662 59788 14714
rect 59542 14660 59548 14662
rect 59604 14660 59628 14662
rect 59684 14660 59708 14662
rect 59764 14660 59788 14662
rect 59844 14660 59850 14662
rect 59542 14651 59850 14660
rect 59924 14414 59952 15098
rect 60108 15094 60136 15302
rect 60096 15088 60148 15094
rect 60096 15030 60148 15036
rect 59912 14408 59964 14414
rect 59912 14350 59964 14356
rect 60004 14272 60056 14278
rect 60004 14214 60056 14220
rect 60016 14006 60044 14214
rect 60004 14000 60056 14006
rect 60004 13942 60056 13948
rect 59174 13903 59230 13912
rect 59452 13932 59504 13938
rect 58992 13388 59044 13394
rect 58992 13330 59044 13336
rect 59188 13258 59216 13903
rect 59452 13874 59504 13880
rect 59464 13326 59492 13874
rect 60004 13796 60056 13802
rect 60004 13738 60056 13744
rect 59542 13628 59850 13637
rect 59542 13626 59548 13628
rect 59604 13626 59628 13628
rect 59684 13626 59708 13628
rect 59764 13626 59788 13628
rect 59844 13626 59850 13628
rect 59604 13574 59606 13626
rect 59786 13574 59788 13626
rect 59542 13572 59548 13574
rect 59604 13572 59628 13574
rect 59684 13572 59708 13574
rect 59764 13572 59788 13574
rect 59844 13572 59850 13574
rect 59542 13563 59850 13572
rect 59452 13320 59504 13326
rect 59452 13262 59504 13268
rect 59176 13252 59228 13258
rect 59176 13194 59228 13200
rect 59084 13184 59136 13190
rect 59084 13126 59136 13132
rect 59096 12850 59124 13126
rect 59360 12912 59412 12918
rect 59360 12854 59412 12860
rect 59084 12844 59136 12850
rect 59084 12786 59136 12792
rect 59084 12708 59136 12714
rect 59084 12650 59136 12656
rect 59096 12434 59124 12650
rect 59372 12442 59400 12854
rect 59542 12540 59850 12549
rect 59542 12538 59548 12540
rect 59604 12538 59628 12540
rect 59684 12538 59708 12540
rect 59764 12538 59788 12540
rect 59844 12538 59850 12540
rect 59604 12486 59606 12538
rect 59786 12486 59788 12538
rect 59542 12484 59548 12486
rect 59604 12484 59628 12486
rect 59684 12484 59708 12486
rect 59764 12484 59788 12486
rect 59844 12484 59850 12486
rect 59542 12475 59850 12484
rect 59360 12436 59412 12442
rect 59096 12406 59308 12434
rect 59280 12322 59308 12406
rect 59360 12378 59412 12384
rect 59910 12336 59966 12345
rect 59280 12294 59400 12322
rect 58900 12232 58952 12238
rect 58900 12174 58952 12180
rect 59174 12200 59230 12209
rect 58808 11892 58860 11898
rect 58808 11834 58860 11840
rect 58912 11762 58940 12174
rect 59174 12135 59230 12144
rect 58532 11756 58584 11762
rect 58532 11698 58584 11704
rect 58716 11756 58768 11762
rect 58716 11698 58768 11704
rect 58900 11756 58952 11762
rect 58900 11698 58952 11704
rect 58624 11552 58676 11558
rect 58624 11494 58676 11500
rect 58900 11552 58952 11558
rect 58900 11494 58952 11500
rect 58992 11552 59044 11558
rect 58992 11494 59044 11500
rect 58636 11218 58664 11494
rect 58440 11212 58492 11218
rect 58440 11154 58492 11160
rect 58624 11212 58676 11218
rect 58676 11172 58756 11200
rect 58624 11154 58676 11160
rect 58452 11082 58480 11154
rect 58440 11076 58492 11082
rect 58440 11018 58492 11024
rect 58624 9988 58676 9994
rect 58624 9930 58676 9936
rect 58636 9518 58664 9930
rect 58624 9512 58676 9518
rect 58624 9454 58676 9460
rect 58532 9104 58584 9110
rect 58532 9046 58584 9052
rect 58440 8832 58492 8838
rect 58440 8774 58492 8780
rect 58348 7744 58400 7750
rect 58348 7686 58400 7692
rect 58256 6452 58308 6458
rect 58256 6394 58308 6400
rect 58452 5710 58480 8774
rect 58544 7002 58572 9046
rect 58636 9042 58664 9454
rect 58624 9036 58676 9042
rect 58624 8978 58676 8984
rect 58624 8560 58676 8566
rect 58624 8502 58676 8508
rect 58636 7546 58664 8502
rect 58624 7540 58676 7546
rect 58624 7482 58676 7488
rect 58532 6996 58584 7002
rect 58532 6938 58584 6944
rect 58728 6497 58756 11172
rect 58912 11121 58940 11494
rect 58898 11112 58954 11121
rect 59004 11082 59032 11494
rect 59188 11286 59216 12135
rect 59372 11558 59400 12294
rect 59910 12271 59966 12280
rect 59452 12096 59504 12102
rect 59452 12038 59504 12044
rect 59360 11552 59412 11558
rect 59360 11494 59412 11500
rect 59176 11280 59228 11286
rect 59176 11222 59228 11228
rect 59084 11212 59136 11218
rect 59084 11154 59136 11160
rect 59096 11082 59124 11154
rect 58898 11047 58954 11056
rect 58992 11076 59044 11082
rect 58992 11018 59044 11024
rect 59084 11076 59136 11082
rect 59084 11018 59136 11024
rect 58808 10736 58860 10742
rect 58808 10678 58860 10684
rect 58820 9586 58848 10678
rect 59096 10470 59124 11018
rect 59464 11014 59492 12038
rect 59542 11452 59850 11461
rect 59542 11450 59548 11452
rect 59604 11450 59628 11452
rect 59684 11450 59708 11452
rect 59764 11450 59788 11452
rect 59844 11450 59850 11452
rect 59604 11398 59606 11450
rect 59786 11398 59788 11450
rect 59542 11396 59548 11398
rect 59604 11396 59628 11398
rect 59684 11396 59708 11398
rect 59764 11396 59788 11398
rect 59844 11396 59850 11398
rect 59542 11387 59850 11396
rect 59636 11348 59688 11354
rect 59636 11290 59688 11296
rect 59648 11150 59676 11290
rect 59636 11144 59688 11150
rect 59924 11121 59952 12271
rect 60016 12238 60044 13738
rect 60186 13016 60242 13025
rect 60186 12951 60242 12960
rect 60200 12617 60228 12951
rect 60186 12608 60242 12617
rect 60186 12543 60242 12552
rect 60292 12434 60320 15574
rect 60464 14544 60516 14550
rect 60464 14486 60516 14492
rect 60476 13870 60504 14486
rect 60556 14476 60608 14482
rect 60608 14436 60688 14464
rect 60556 14418 60608 14424
rect 60556 14340 60608 14346
rect 60556 14282 60608 14288
rect 60464 13864 60516 13870
rect 60464 13806 60516 13812
rect 60370 13560 60426 13569
rect 60370 13495 60426 13504
rect 60464 13524 60516 13530
rect 60384 12986 60412 13495
rect 60464 13466 60516 13472
rect 60372 12980 60424 12986
rect 60372 12922 60424 12928
rect 60476 12714 60504 13466
rect 60464 12708 60516 12714
rect 60464 12650 60516 12656
rect 60292 12406 60504 12434
rect 60004 12232 60056 12238
rect 60004 12174 60056 12180
rect 60096 11620 60148 11626
rect 60096 11562 60148 11568
rect 60004 11552 60056 11558
rect 60004 11494 60056 11500
rect 59636 11086 59688 11092
rect 59910 11112 59966 11121
rect 59452 11008 59504 11014
rect 59452 10950 59504 10956
rect 59648 10742 59676 11086
rect 59910 11047 59966 11056
rect 59636 10736 59688 10742
rect 59636 10678 59688 10684
rect 59084 10464 59136 10470
rect 59084 10406 59136 10412
rect 59542 10364 59850 10373
rect 59542 10362 59548 10364
rect 59604 10362 59628 10364
rect 59684 10362 59708 10364
rect 59764 10362 59788 10364
rect 59844 10362 59850 10364
rect 59604 10310 59606 10362
rect 59786 10310 59788 10362
rect 59542 10308 59548 10310
rect 59604 10308 59628 10310
rect 59684 10308 59708 10310
rect 59764 10308 59788 10310
rect 59844 10308 59850 10310
rect 59358 10296 59414 10305
rect 59542 10299 59850 10308
rect 59358 10231 59414 10240
rect 59372 10130 59400 10231
rect 59360 10124 59412 10130
rect 59360 10066 59412 10072
rect 58900 9988 58952 9994
rect 58900 9930 58952 9936
rect 58808 9580 58860 9586
rect 58808 9522 58860 9528
rect 58808 9376 58860 9382
rect 58808 9318 58860 9324
rect 58820 7818 58848 9318
rect 58912 8974 58940 9930
rect 59372 9761 59400 10066
rect 59358 9752 59414 9761
rect 59358 9687 59414 9696
rect 58992 9580 59044 9586
rect 58992 9522 59044 9528
rect 59004 9382 59032 9522
rect 58992 9376 59044 9382
rect 60016 9330 60044 11494
rect 60108 11393 60136 11562
rect 60372 11552 60424 11558
rect 60370 11520 60372 11529
rect 60424 11520 60426 11529
rect 60370 11455 60426 11464
rect 60094 11384 60150 11393
rect 60094 11319 60150 11328
rect 60384 10198 60412 11455
rect 60476 10198 60504 12406
rect 60568 11801 60596 14282
rect 60660 14249 60688 14436
rect 60646 14240 60702 14249
rect 60646 14175 60702 14184
rect 60752 13954 60780 15830
rect 60832 15700 60884 15706
rect 60832 15642 60884 15648
rect 60844 15094 60872 15642
rect 61120 15570 61148 16662
rect 61856 16522 61884 17070
rect 62856 17060 62908 17066
rect 62856 17002 62908 17008
rect 62028 16788 62080 16794
rect 62028 16730 62080 16736
rect 61844 16516 61896 16522
rect 61844 16458 61896 16464
rect 61856 16130 61884 16458
rect 62040 16454 62068 16730
rect 62868 16590 62896 17002
rect 62856 16584 62908 16590
rect 62856 16526 62908 16532
rect 63604 16522 63632 17070
rect 65524 16652 65576 16658
rect 65524 16594 65576 16600
rect 63592 16516 63644 16522
rect 63592 16458 63644 16464
rect 61936 16448 61988 16454
rect 61936 16390 61988 16396
rect 62028 16448 62080 16454
rect 62028 16390 62080 16396
rect 61948 16250 61976 16390
rect 61936 16244 61988 16250
rect 61936 16186 61988 16192
rect 61856 16102 61976 16130
rect 63604 16114 63632 16458
rect 64604 16448 64656 16454
rect 64604 16390 64656 16396
rect 64972 16448 65024 16454
rect 64972 16390 65024 16396
rect 61844 16040 61896 16046
rect 61844 15982 61896 15988
rect 61108 15564 61160 15570
rect 61108 15506 61160 15512
rect 61016 15496 61068 15502
rect 61068 15444 61148 15450
rect 61016 15438 61148 15444
rect 61028 15422 61148 15438
rect 60832 15088 60884 15094
rect 60832 15030 60884 15036
rect 61120 14006 61148 15422
rect 61568 15156 61620 15162
rect 61568 15098 61620 15104
rect 61476 15088 61528 15094
rect 61304 15036 61476 15042
rect 61304 15030 61528 15036
rect 61304 15026 61516 15030
rect 61580 15026 61608 15098
rect 61292 15020 61516 15026
rect 61344 15014 61516 15020
rect 61568 15020 61620 15026
rect 61292 14962 61344 14968
rect 61568 14962 61620 14968
rect 61660 14816 61712 14822
rect 61660 14758 61712 14764
rect 61672 14346 61700 14758
rect 61660 14340 61712 14346
rect 61660 14282 61712 14288
rect 61660 14068 61712 14074
rect 61660 14010 61712 14016
rect 61108 14000 61160 14006
rect 60752 13926 60872 13954
rect 61672 13977 61700 14010
rect 61108 13942 61160 13948
rect 61658 13968 61714 13977
rect 60646 13696 60702 13705
rect 60646 13631 60702 13640
rect 60660 13326 60688 13631
rect 60648 13320 60700 13326
rect 60648 13262 60700 13268
rect 60740 13184 60792 13190
rect 60740 13126 60792 13132
rect 60648 12980 60700 12986
rect 60648 12922 60700 12928
rect 60660 12646 60688 12922
rect 60752 12918 60780 13126
rect 60740 12912 60792 12918
rect 60740 12854 60792 12860
rect 60648 12640 60700 12646
rect 60648 12582 60700 12588
rect 60844 12442 60872 13926
rect 61476 13932 61528 13938
rect 61658 13903 61714 13912
rect 61476 13874 61528 13880
rect 61016 13524 61068 13530
rect 61016 13466 61068 13472
rect 61028 13274 61056 13466
rect 60936 13246 61056 13274
rect 60832 12436 60884 12442
rect 60832 12378 60884 12384
rect 60646 12336 60702 12345
rect 60646 12271 60702 12280
rect 60660 12238 60688 12271
rect 60648 12232 60700 12238
rect 60648 12174 60700 12180
rect 60648 12096 60700 12102
rect 60648 12038 60700 12044
rect 60554 11792 60610 11801
rect 60554 11727 60610 11736
rect 60660 11744 60688 12038
rect 60738 11792 60794 11801
rect 60660 11736 60738 11744
rect 60660 11727 60794 11736
rect 60568 11014 60596 11727
rect 60660 11716 60780 11727
rect 60936 11665 60964 13246
rect 61290 13152 61346 13161
rect 61290 13087 61346 13096
rect 61304 12986 61332 13087
rect 61292 12980 61344 12986
rect 61292 12922 61344 12928
rect 61016 12844 61068 12850
rect 61016 12786 61068 12792
rect 61028 12646 61056 12786
rect 61488 12764 61516 13874
rect 61568 13864 61620 13870
rect 61568 13806 61620 13812
rect 61580 12986 61608 13806
rect 61672 13326 61700 13903
rect 61660 13320 61712 13326
rect 61660 13262 61712 13268
rect 61752 13252 61804 13258
rect 61752 13194 61804 13200
rect 61568 12980 61620 12986
rect 61568 12922 61620 12928
rect 61660 12776 61712 12782
rect 61488 12736 61660 12764
rect 61660 12718 61712 12724
rect 61016 12640 61068 12646
rect 61016 12582 61068 12588
rect 61672 12238 61700 12718
rect 61764 12374 61792 13194
rect 61752 12368 61804 12374
rect 61752 12310 61804 12316
rect 61660 12232 61712 12238
rect 61660 12174 61712 12180
rect 60922 11656 60978 11665
rect 60922 11591 60978 11600
rect 60936 11218 60964 11591
rect 61672 11286 61700 12174
rect 61752 12096 61804 12102
rect 61752 12038 61804 12044
rect 61764 11286 61792 12038
rect 61660 11280 61712 11286
rect 61660 11222 61712 11228
rect 61752 11280 61804 11286
rect 61752 11222 61804 11228
rect 61856 11218 61884 15982
rect 61948 15434 61976 16102
rect 63592 16108 63644 16114
rect 63592 16050 63644 16056
rect 64616 15978 64644 16390
rect 64984 16182 65012 16390
rect 65536 16182 65564 16594
rect 65812 16522 65840 17070
rect 65904 16794 65932 17206
rect 68376 17196 68428 17202
rect 68376 17138 68428 17144
rect 67548 17060 67600 17066
rect 67548 17002 67600 17008
rect 65892 16788 65944 16794
rect 65892 16730 65944 16736
rect 67560 16590 67588 17002
rect 68192 16720 68244 16726
rect 68192 16662 68244 16668
rect 67548 16584 67600 16590
rect 67548 16526 67600 16532
rect 65800 16516 65852 16522
rect 65800 16458 65852 16464
rect 64972 16176 65024 16182
rect 64972 16118 65024 16124
rect 65524 16176 65576 16182
rect 65524 16118 65576 16124
rect 66076 16176 66128 16182
rect 66076 16118 66128 16124
rect 64604 15972 64656 15978
rect 64604 15914 64656 15920
rect 62212 15904 62264 15910
rect 62212 15846 62264 15852
rect 62948 15904 63000 15910
rect 62948 15846 63000 15852
rect 61936 15428 61988 15434
rect 61936 15370 61988 15376
rect 61948 15094 61976 15370
rect 61936 15088 61988 15094
rect 61936 15030 61988 15036
rect 61948 12646 61976 15030
rect 62224 14074 62252 15846
rect 62304 15156 62356 15162
rect 62304 15098 62356 15104
rect 62316 14890 62344 15098
rect 62304 14884 62356 14890
rect 62304 14826 62356 14832
rect 62960 14414 62988 15846
rect 64696 15564 64748 15570
rect 64696 15506 64748 15512
rect 64708 15473 64736 15506
rect 64694 15464 64750 15473
rect 64984 15434 65012 16118
rect 66088 15910 66116 16118
rect 66168 16108 66220 16114
rect 66168 16050 66220 16056
rect 65892 15904 65944 15910
rect 65892 15846 65944 15852
rect 66076 15904 66128 15910
rect 66076 15846 66128 15852
rect 65904 15502 65932 15846
rect 65984 15700 66036 15706
rect 65984 15642 66036 15648
rect 65996 15502 66024 15642
rect 65892 15496 65944 15502
rect 65892 15438 65944 15444
rect 65984 15496 66036 15502
rect 65984 15438 66036 15444
rect 64694 15399 64750 15408
rect 64972 15428 65024 15434
rect 64972 15370 65024 15376
rect 63592 15360 63644 15366
rect 63592 15302 63644 15308
rect 63132 15020 63184 15026
rect 63132 14962 63184 14968
rect 63040 14544 63092 14550
rect 63040 14486 63092 14492
rect 62948 14408 63000 14414
rect 62948 14350 63000 14356
rect 62212 14068 62264 14074
rect 62212 14010 62264 14016
rect 62120 13456 62172 13462
rect 62120 13398 62172 13404
rect 62026 13016 62082 13025
rect 62132 12986 62160 13398
rect 62960 13394 62988 14350
rect 62488 13388 62540 13394
rect 62488 13330 62540 13336
rect 62948 13388 63000 13394
rect 62948 13330 63000 13336
rect 62026 12951 62082 12960
rect 62120 12980 62172 12986
rect 62040 12850 62068 12951
rect 62120 12922 62172 12928
rect 62028 12844 62080 12850
rect 62028 12786 62080 12792
rect 61936 12640 61988 12646
rect 61936 12582 61988 12588
rect 62212 12640 62264 12646
rect 62212 12582 62264 12588
rect 62120 12300 62172 12306
rect 62120 12242 62172 12248
rect 61934 12200 61990 12209
rect 61934 12135 61990 12144
rect 61948 12102 61976 12135
rect 61936 12096 61988 12102
rect 61936 12038 61988 12044
rect 62132 11830 62160 12242
rect 62120 11824 62172 11830
rect 62120 11766 62172 11772
rect 60740 11212 60792 11218
rect 60740 11154 60792 11160
rect 60924 11212 60976 11218
rect 60924 11154 60976 11160
rect 61844 11212 61896 11218
rect 61844 11154 61896 11160
rect 60556 11008 60608 11014
rect 60556 10950 60608 10956
rect 60752 10266 60780 11154
rect 61476 11144 61528 11150
rect 61476 11086 61528 11092
rect 61488 11014 61516 11086
rect 62120 11076 62172 11082
rect 62120 11018 62172 11024
rect 61476 11008 61528 11014
rect 61476 10950 61528 10956
rect 61660 10736 61712 10742
rect 61660 10678 61712 10684
rect 61568 10600 61620 10606
rect 61568 10542 61620 10548
rect 60740 10260 60792 10266
rect 60740 10202 60792 10208
rect 60372 10192 60424 10198
rect 60372 10134 60424 10140
rect 60464 10192 60516 10198
rect 60464 10134 60516 10140
rect 60476 10010 60504 10134
rect 60384 9982 60504 10010
rect 61108 10056 61160 10062
rect 61580 10033 61608 10542
rect 61108 9998 61160 10004
rect 61566 10024 61622 10033
rect 60384 9926 60412 9982
rect 60372 9920 60424 9926
rect 60372 9862 60424 9868
rect 60464 9920 60516 9926
rect 60464 9862 60516 9868
rect 60370 9752 60426 9761
rect 60370 9687 60426 9696
rect 58992 9318 59044 9324
rect 59004 9178 59032 9318
rect 59924 9302 60044 9330
rect 59542 9276 59850 9285
rect 59542 9274 59548 9276
rect 59604 9274 59628 9276
rect 59684 9274 59708 9276
rect 59764 9274 59788 9276
rect 59844 9274 59850 9276
rect 59604 9222 59606 9274
rect 59786 9222 59788 9274
rect 59542 9220 59548 9222
rect 59604 9220 59628 9222
rect 59684 9220 59708 9222
rect 59764 9220 59788 9222
rect 59844 9220 59850 9222
rect 59542 9211 59850 9220
rect 58992 9172 59044 9178
rect 58992 9114 59044 9120
rect 59636 9104 59688 9110
rect 59636 9046 59688 9052
rect 58900 8968 58952 8974
rect 58900 8910 58952 8916
rect 58912 8090 58940 8910
rect 59648 8906 59676 9046
rect 59924 9042 59952 9302
rect 60002 9208 60058 9217
rect 60002 9143 60058 9152
rect 59912 9036 59964 9042
rect 59912 8978 59964 8984
rect 60016 8945 60044 9143
rect 60096 9104 60148 9110
rect 60096 9046 60148 9052
rect 60002 8936 60058 8945
rect 59636 8900 59688 8906
rect 60002 8871 60058 8880
rect 59636 8842 59688 8848
rect 59360 8832 59412 8838
rect 59360 8774 59412 8780
rect 59268 8628 59320 8634
rect 59268 8570 59320 8576
rect 59280 8430 59308 8570
rect 59372 8498 59400 8774
rect 59360 8492 59412 8498
rect 59360 8434 59412 8440
rect 59084 8424 59136 8430
rect 59084 8366 59136 8372
rect 59268 8424 59320 8430
rect 59268 8366 59320 8372
rect 59820 8424 59872 8430
rect 59872 8384 59952 8412
rect 59820 8366 59872 8372
rect 58900 8084 58952 8090
rect 58900 8026 58952 8032
rect 58808 7812 58860 7818
rect 58808 7754 58860 7760
rect 58714 6488 58770 6497
rect 58714 6423 58770 6432
rect 58992 6452 59044 6458
rect 58728 6390 58756 6423
rect 58992 6394 59044 6400
rect 58716 6384 58768 6390
rect 58716 6326 58768 6332
rect 58900 6316 58952 6322
rect 58900 6258 58952 6264
rect 58912 5846 58940 6258
rect 58900 5840 58952 5846
rect 58806 5808 58862 5817
rect 58900 5782 58952 5788
rect 58806 5743 58808 5752
rect 58860 5743 58862 5752
rect 58808 5714 58860 5720
rect 58440 5704 58492 5710
rect 58440 5646 58492 5652
rect 58806 5400 58862 5409
rect 58806 5335 58862 5344
rect 58348 5228 58400 5234
rect 58348 5170 58400 5176
rect 58164 4820 58216 4826
rect 58164 4762 58216 4768
rect 58360 4690 58388 5170
rect 58820 5098 58848 5335
rect 59004 5098 59032 6394
rect 58808 5092 58860 5098
rect 58808 5034 58860 5040
rect 58992 5092 59044 5098
rect 58992 5034 59044 5040
rect 59096 5030 59124 8366
rect 59360 8356 59412 8362
rect 59360 8298 59412 8304
rect 59176 8288 59228 8294
rect 59176 8230 59228 8236
rect 59188 7954 59216 8230
rect 59176 7948 59228 7954
rect 59176 7890 59228 7896
rect 59176 7744 59228 7750
rect 59176 7686 59228 7692
rect 59188 6390 59216 7686
rect 59372 7478 59400 8298
rect 59542 8188 59850 8197
rect 59542 8186 59548 8188
rect 59604 8186 59628 8188
rect 59684 8186 59708 8188
rect 59764 8186 59788 8188
rect 59844 8186 59850 8188
rect 59604 8134 59606 8186
rect 59786 8134 59788 8186
rect 59542 8132 59548 8134
rect 59604 8132 59628 8134
rect 59684 8132 59708 8134
rect 59764 8132 59788 8134
rect 59844 8132 59850 8134
rect 59542 8123 59850 8132
rect 59360 7472 59412 7478
rect 59360 7414 59412 7420
rect 59360 7268 59412 7274
rect 59360 7210 59412 7216
rect 59176 6384 59228 6390
rect 59176 6326 59228 6332
rect 59188 5574 59216 6326
rect 59372 6322 59400 7210
rect 59542 7100 59850 7109
rect 59542 7098 59548 7100
rect 59604 7098 59628 7100
rect 59684 7098 59708 7100
rect 59764 7098 59788 7100
rect 59844 7098 59850 7100
rect 59604 7046 59606 7098
rect 59786 7046 59788 7098
rect 59542 7044 59548 7046
rect 59604 7044 59628 7046
rect 59684 7044 59708 7046
rect 59764 7044 59788 7046
rect 59844 7044 59850 7046
rect 59542 7035 59850 7044
rect 59924 6882 59952 8384
rect 60016 7834 60044 8871
rect 60108 8566 60136 9046
rect 60096 8560 60148 8566
rect 60096 8502 60148 8508
rect 60096 8424 60148 8430
rect 60096 8366 60148 8372
rect 60108 8022 60136 8366
rect 60188 8288 60240 8294
rect 60188 8230 60240 8236
rect 60096 8016 60148 8022
rect 60096 7958 60148 7964
rect 60200 7886 60228 8230
rect 60188 7880 60240 7886
rect 60016 7806 60136 7834
rect 60188 7822 60240 7828
rect 59924 6854 60044 6882
rect 60016 6798 60044 6854
rect 59452 6792 59504 6798
rect 59452 6734 59504 6740
rect 59912 6792 59964 6798
rect 59912 6734 59964 6740
rect 60004 6792 60056 6798
rect 60004 6734 60056 6740
rect 59360 6316 59412 6322
rect 59360 6258 59412 6264
rect 59268 6248 59320 6254
rect 59268 6190 59320 6196
rect 59176 5568 59228 5574
rect 59176 5510 59228 5516
rect 59084 5024 59136 5030
rect 59084 4966 59136 4972
rect 58348 4684 58400 4690
rect 58348 4626 58400 4632
rect 58532 4684 58584 4690
rect 58532 4626 58584 4632
rect 57888 4140 57940 4146
rect 57888 4082 57940 4088
rect 58072 4140 58124 4146
rect 58072 4082 58124 4088
rect 57796 4004 57848 4010
rect 57796 3946 57848 3952
rect 57060 3936 57112 3942
rect 57060 3878 57112 3884
rect 56784 3188 56836 3194
rect 56784 3130 56836 3136
rect 57072 2922 57100 3878
rect 58544 3738 58572 4626
rect 59096 4622 59124 4966
rect 58716 4616 58768 4622
rect 58716 4558 58768 4564
rect 59084 4616 59136 4622
rect 59084 4558 59136 4564
rect 58728 4078 58756 4558
rect 58716 4072 58768 4078
rect 58716 4014 58768 4020
rect 59280 3738 59308 6190
rect 59464 5914 59492 6734
rect 59544 6656 59596 6662
rect 59544 6598 59596 6604
rect 59556 6458 59584 6598
rect 59544 6452 59596 6458
rect 59544 6394 59596 6400
rect 59542 6012 59850 6021
rect 59542 6010 59548 6012
rect 59604 6010 59628 6012
rect 59684 6010 59708 6012
rect 59764 6010 59788 6012
rect 59844 6010 59850 6012
rect 59604 5958 59606 6010
rect 59786 5958 59788 6010
rect 59542 5956 59548 5958
rect 59604 5956 59628 5958
rect 59684 5956 59708 5958
rect 59764 5956 59788 5958
rect 59844 5956 59850 5958
rect 59542 5947 59850 5956
rect 59452 5908 59504 5914
rect 59452 5850 59504 5856
rect 59464 5710 59492 5850
rect 59452 5704 59504 5710
rect 59452 5646 59504 5652
rect 59360 5636 59412 5642
rect 59360 5578 59412 5584
rect 59372 3942 59400 5578
rect 59820 5568 59872 5574
rect 59820 5510 59872 5516
rect 59452 5160 59504 5166
rect 59452 5102 59504 5108
rect 59464 4282 59492 5102
rect 59832 5030 59860 5510
rect 59820 5024 59872 5030
rect 59820 4966 59872 4972
rect 59542 4924 59850 4933
rect 59542 4922 59548 4924
rect 59604 4922 59628 4924
rect 59684 4922 59708 4924
rect 59764 4922 59788 4924
rect 59844 4922 59850 4924
rect 59604 4870 59606 4922
rect 59786 4870 59788 4922
rect 59542 4868 59548 4870
rect 59604 4868 59628 4870
rect 59684 4868 59708 4870
rect 59764 4868 59788 4870
rect 59844 4868 59850 4870
rect 59542 4859 59850 4868
rect 59924 4690 59952 6734
rect 60004 6656 60056 6662
rect 60004 6598 60056 6604
rect 60016 6254 60044 6598
rect 60004 6248 60056 6254
rect 60004 6190 60056 6196
rect 60108 5914 60136 7806
rect 60280 6792 60332 6798
rect 60280 6734 60332 6740
rect 60096 5908 60148 5914
rect 60096 5850 60148 5856
rect 60292 5846 60320 6734
rect 60280 5840 60332 5846
rect 60280 5782 60332 5788
rect 60292 5642 60320 5782
rect 60280 5636 60332 5642
rect 60280 5578 60332 5584
rect 60384 5574 60412 9687
rect 60476 7342 60504 9862
rect 61120 9654 61148 9998
rect 61566 9959 61622 9968
rect 61108 9648 61160 9654
rect 61108 9590 61160 9596
rect 60648 9512 60700 9518
rect 60648 9454 60700 9460
rect 60660 9042 60688 9454
rect 61016 9444 61068 9450
rect 61016 9386 61068 9392
rect 60648 9036 60700 9042
rect 60648 8978 60700 8984
rect 60924 8968 60976 8974
rect 60924 8910 60976 8916
rect 60556 8832 60608 8838
rect 60556 8774 60608 8780
rect 60568 7546 60596 8774
rect 60936 7954 60964 8910
rect 61028 8673 61056 9386
rect 61014 8664 61070 8673
rect 61014 8599 61070 8608
rect 61120 8090 61148 9590
rect 61292 9512 61344 9518
rect 61292 9454 61344 9460
rect 61304 9110 61332 9454
rect 61292 9104 61344 9110
rect 61292 9046 61344 9052
rect 61292 8900 61344 8906
rect 61292 8842 61344 8848
rect 61016 8084 61068 8090
rect 61016 8026 61068 8032
rect 61108 8084 61160 8090
rect 61108 8026 61160 8032
rect 61028 7954 61056 8026
rect 60924 7948 60976 7954
rect 60924 7890 60976 7896
rect 61016 7948 61068 7954
rect 61016 7890 61068 7896
rect 60648 7880 60700 7886
rect 60648 7822 60700 7828
rect 60660 7585 60688 7822
rect 60646 7576 60702 7585
rect 60556 7540 60608 7546
rect 60646 7511 60702 7520
rect 60832 7540 60884 7546
rect 60556 7482 60608 7488
rect 60832 7482 60884 7488
rect 60464 7336 60516 7342
rect 60464 7278 60516 7284
rect 60372 5568 60424 5574
rect 60372 5510 60424 5516
rect 60476 5166 60504 7278
rect 60648 6860 60700 6866
rect 60648 6802 60700 6808
rect 60660 6458 60688 6802
rect 60844 6798 60872 7482
rect 60924 7268 60976 7274
rect 60924 7210 60976 7216
rect 61108 7268 61160 7274
rect 61108 7210 61160 7216
rect 60936 6866 60964 7210
rect 61120 7002 61148 7210
rect 61108 6996 61160 7002
rect 61108 6938 61160 6944
rect 60924 6860 60976 6866
rect 61120 6848 61148 6938
rect 61120 6820 61240 6848
rect 60924 6802 60976 6808
rect 60832 6792 60884 6798
rect 60832 6734 60884 6740
rect 61016 6792 61068 6798
rect 61016 6734 61068 6740
rect 60648 6452 60700 6458
rect 60648 6394 60700 6400
rect 61028 6186 61056 6734
rect 61108 6724 61160 6730
rect 61108 6666 61160 6672
rect 61120 6186 61148 6666
rect 61016 6180 61068 6186
rect 61016 6122 61068 6128
rect 61108 6180 61160 6186
rect 61108 6122 61160 6128
rect 60738 5808 60794 5817
rect 60738 5743 60740 5752
rect 60792 5743 60794 5752
rect 60740 5714 60792 5720
rect 60832 5704 60884 5710
rect 60832 5646 60884 5652
rect 60464 5160 60516 5166
rect 60464 5102 60516 5108
rect 60844 5030 60872 5646
rect 60832 5024 60884 5030
rect 60832 4966 60884 4972
rect 61212 4758 61240 6820
rect 61304 4826 61332 8842
rect 61568 7540 61620 7546
rect 61568 7482 61620 7488
rect 61580 7342 61608 7482
rect 61568 7336 61620 7342
rect 61568 7278 61620 7284
rect 61672 6798 61700 10678
rect 62132 10606 62160 11018
rect 62120 10600 62172 10606
rect 62120 10542 62172 10548
rect 61936 10532 61988 10538
rect 61936 10474 61988 10480
rect 61948 9926 61976 10474
rect 61936 9920 61988 9926
rect 61936 9862 61988 9868
rect 62120 9512 62172 9518
rect 62120 9454 62172 9460
rect 61752 9376 61804 9382
rect 61752 9318 61804 9324
rect 61936 9376 61988 9382
rect 61936 9318 61988 9324
rect 61764 9110 61792 9318
rect 61752 9104 61804 9110
rect 61752 9046 61804 9052
rect 61948 7818 61976 9318
rect 62132 9042 62160 9454
rect 62120 9036 62172 9042
rect 62120 8978 62172 8984
rect 62224 8498 62252 12582
rect 62304 11892 62356 11898
rect 62304 11834 62356 11840
rect 62316 9042 62344 11834
rect 62500 11354 62528 13330
rect 62580 12368 62632 12374
rect 63052 12345 63080 14486
rect 62580 12310 62632 12316
rect 63038 12336 63094 12345
rect 62592 11558 62620 12310
rect 63038 12271 63094 12280
rect 63144 11762 63172 14962
rect 63224 14272 63276 14278
rect 63224 14214 63276 14220
rect 63236 14113 63264 14214
rect 63222 14104 63278 14113
rect 63222 14039 63278 14048
rect 63236 12850 63264 14039
rect 63500 13728 63552 13734
rect 63500 13670 63552 13676
rect 63512 13258 63540 13670
rect 63500 13252 63552 13258
rect 63500 13194 63552 13200
rect 63316 13184 63368 13190
rect 63316 13126 63368 13132
rect 63408 13184 63460 13190
rect 63408 13126 63460 13132
rect 63224 12844 63276 12850
rect 63224 12786 63276 12792
rect 63328 11898 63356 13126
rect 63316 11892 63368 11898
rect 63316 11834 63368 11840
rect 63224 11824 63276 11830
rect 63420 11778 63448 13126
rect 63276 11772 63448 11778
rect 63224 11766 63448 11772
rect 63132 11756 63184 11762
rect 63236 11750 63448 11766
rect 63132 11698 63184 11704
rect 63604 11694 63632 15302
rect 66180 15162 66208 16050
rect 66352 16040 66404 16046
rect 66352 15982 66404 15988
rect 66536 16040 66588 16046
rect 66536 15982 66588 15988
rect 66168 15156 66220 15162
rect 66168 15098 66220 15104
rect 65432 15088 65484 15094
rect 65432 15030 65484 15036
rect 64880 14952 64932 14958
rect 64880 14894 64932 14900
rect 64236 14816 64288 14822
rect 64236 14758 64288 14764
rect 64248 14278 64276 14758
rect 64892 14618 64920 14894
rect 64880 14612 64932 14618
rect 64880 14554 64932 14560
rect 65444 14414 65472 15030
rect 65892 14952 65944 14958
rect 65892 14894 65944 14900
rect 65432 14408 65484 14414
rect 65432 14350 65484 14356
rect 65904 14278 65932 14894
rect 65984 14408 66036 14414
rect 65984 14350 66036 14356
rect 66076 14408 66128 14414
rect 66076 14350 66128 14356
rect 65996 14278 66024 14350
rect 63684 14272 63736 14278
rect 63684 14214 63736 14220
rect 64236 14272 64288 14278
rect 64236 14214 64288 14220
rect 65156 14272 65208 14278
rect 65156 14214 65208 14220
rect 65892 14272 65944 14278
rect 65892 14214 65944 14220
rect 65984 14272 66036 14278
rect 66088 14249 66116 14350
rect 65984 14214 66036 14220
rect 66074 14240 66130 14249
rect 63696 12102 63724 14214
rect 63868 14000 63920 14006
rect 63868 13942 63920 13948
rect 63684 12096 63736 12102
rect 63684 12038 63736 12044
rect 63696 11898 63724 12038
rect 63684 11892 63736 11898
rect 63684 11834 63736 11840
rect 63592 11688 63644 11694
rect 63592 11630 63644 11636
rect 62580 11552 62632 11558
rect 62580 11494 62632 11500
rect 63592 11552 63644 11558
rect 63592 11494 63644 11500
rect 63604 11354 63632 11494
rect 62488 11348 62540 11354
rect 62488 11290 62540 11296
rect 63592 11348 63644 11354
rect 63592 11290 63644 11296
rect 63224 11280 63276 11286
rect 63224 11222 63276 11228
rect 62488 11212 62540 11218
rect 62488 11154 62540 11160
rect 62396 11076 62448 11082
rect 62500 11064 62528 11154
rect 62448 11036 62528 11064
rect 62396 11018 62448 11024
rect 62488 10804 62540 10810
rect 62488 10746 62540 10752
rect 62764 10804 62816 10810
rect 62764 10746 62816 10752
rect 62396 10600 62448 10606
rect 62396 10542 62448 10548
rect 62408 10130 62436 10542
rect 62500 10130 62528 10746
rect 62672 10736 62724 10742
rect 62672 10678 62724 10684
rect 62684 10266 62712 10678
rect 62672 10260 62724 10266
rect 62672 10202 62724 10208
rect 62396 10124 62448 10130
rect 62396 10066 62448 10072
rect 62488 10124 62540 10130
rect 62488 10066 62540 10072
rect 62776 10062 62804 10746
rect 63236 10674 63264 11222
rect 63224 10668 63276 10674
rect 63224 10610 63276 10616
rect 63144 10538 63632 10554
rect 63132 10532 63632 10538
rect 63184 10526 63632 10532
rect 63132 10474 63184 10480
rect 63316 10464 63368 10470
rect 63316 10406 63368 10412
rect 63328 10266 63356 10406
rect 63316 10260 63368 10266
rect 63316 10202 63368 10208
rect 63604 10146 63632 10526
rect 63880 10470 63908 13942
rect 64248 13870 64276 14214
rect 65168 14006 65196 14214
rect 66074 14175 66130 14184
rect 65156 14000 65208 14006
rect 65156 13942 65208 13948
rect 64604 13932 64656 13938
rect 64604 13874 64656 13880
rect 64236 13864 64288 13870
rect 64236 13806 64288 13812
rect 64248 13462 64276 13806
rect 64236 13456 64288 13462
rect 64236 13398 64288 13404
rect 64616 13326 64644 13874
rect 64696 13728 64748 13734
rect 64694 13696 64696 13705
rect 64748 13696 64750 13705
rect 64694 13631 64750 13640
rect 66180 13326 66208 15098
rect 66364 13818 66392 15982
rect 66548 15366 66576 15982
rect 67916 15904 67968 15910
rect 67916 15846 67968 15852
rect 68008 15904 68060 15910
rect 68008 15846 68060 15852
rect 67364 15632 67416 15638
rect 67192 15592 67364 15620
rect 66536 15360 66588 15366
rect 66536 15302 66588 15308
rect 66720 15360 66772 15366
rect 66720 15302 66772 15308
rect 66732 15094 66760 15302
rect 66720 15088 66772 15094
rect 66720 15030 66772 15036
rect 67192 15026 67220 15592
rect 67364 15574 67416 15580
rect 67640 15564 67692 15570
rect 67640 15506 67692 15512
rect 67180 15020 67232 15026
rect 67180 14962 67232 14968
rect 66444 14952 66496 14958
rect 66444 14894 66496 14900
rect 66456 13977 66484 14894
rect 66536 14408 66588 14414
rect 66536 14350 66588 14356
rect 66442 13968 66498 13977
rect 66548 13938 66576 14350
rect 66442 13903 66498 13912
rect 66536 13932 66588 13938
rect 66536 13874 66588 13880
rect 66628 13864 66680 13870
rect 66364 13812 66628 13818
rect 66364 13806 66680 13812
rect 66364 13790 66668 13806
rect 64604 13320 64656 13326
rect 64604 13262 64656 13268
rect 65984 13320 66036 13326
rect 65984 13262 66036 13268
rect 66168 13320 66220 13326
rect 66168 13262 66220 13268
rect 64420 11348 64472 11354
rect 64420 11290 64472 11296
rect 63868 10464 63920 10470
rect 63868 10406 63920 10412
rect 63408 10124 63460 10130
rect 63604 10118 63816 10146
rect 63408 10066 63460 10072
rect 62764 10056 62816 10062
rect 62764 9998 62816 10004
rect 62396 9716 62448 9722
rect 62448 9676 62528 9704
rect 62396 9658 62448 9664
rect 62500 9636 62528 9676
rect 63316 9648 63368 9654
rect 62500 9608 62712 9636
rect 62396 9580 62448 9586
rect 62396 9522 62448 9528
rect 62408 9178 62436 9522
rect 62580 9376 62632 9382
rect 62580 9318 62632 9324
rect 62396 9172 62448 9178
rect 62396 9114 62448 9120
rect 62304 9036 62356 9042
rect 62304 8978 62356 8984
rect 62592 8634 62620 9318
rect 62580 8628 62632 8634
rect 62580 8570 62632 8576
rect 62212 8492 62264 8498
rect 62212 8434 62264 8440
rect 62224 7970 62252 8434
rect 62040 7942 62252 7970
rect 61936 7812 61988 7818
rect 61936 7754 61988 7760
rect 61936 7404 61988 7410
rect 61936 7346 61988 7352
rect 61948 6798 61976 7346
rect 61660 6792 61712 6798
rect 61660 6734 61712 6740
rect 61936 6792 61988 6798
rect 61936 6734 61988 6740
rect 61660 6656 61712 6662
rect 61660 6598 61712 6604
rect 61672 6322 61700 6598
rect 61948 6322 61976 6734
rect 61660 6316 61712 6322
rect 61660 6258 61712 6264
rect 61936 6316 61988 6322
rect 61936 6258 61988 6264
rect 61292 4820 61344 4826
rect 61292 4762 61344 4768
rect 61200 4752 61252 4758
rect 61200 4694 61252 4700
rect 59912 4684 59964 4690
rect 59912 4626 59964 4632
rect 59452 4276 59504 4282
rect 59452 4218 59504 4224
rect 59360 3936 59412 3942
rect 59360 3878 59412 3884
rect 59542 3836 59850 3845
rect 59542 3834 59548 3836
rect 59604 3834 59628 3836
rect 59684 3834 59708 3836
rect 59764 3834 59788 3836
rect 59844 3834 59850 3836
rect 59604 3782 59606 3834
rect 59786 3782 59788 3834
rect 59542 3780 59548 3782
rect 59604 3780 59628 3782
rect 59684 3780 59708 3782
rect 59764 3780 59788 3782
rect 59844 3780 59850 3782
rect 59542 3771 59850 3780
rect 61212 3738 61240 4694
rect 62040 4146 62068 7942
rect 62212 7880 62264 7886
rect 62212 7822 62264 7828
rect 62120 7268 62172 7274
rect 62120 7210 62172 7216
rect 62132 6798 62160 7210
rect 62120 6792 62172 6798
rect 62120 6734 62172 6740
rect 62132 6458 62160 6734
rect 62120 6452 62172 6458
rect 62120 6394 62172 6400
rect 62120 6112 62172 6118
rect 62120 6054 62172 6060
rect 62132 5914 62160 6054
rect 62120 5908 62172 5914
rect 62120 5850 62172 5856
rect 62224 4282 62252 7822
rect 62684 7818 62712 9608
rect 63316 9590 63368 9596
rect 63040 9580 63092 9586
rect 63040 9522 63092 9528
rect 63224 9580 63276 9586
rect 63224 9522 63276 9528
rect 62672 7812 62724 7818
rect 62672 7754 62724 7760
rect 62578 7576 62634 7585
rect 62578 7511 62634 7520
rect 62488 7200 62540 7206
rect 62488 7142 62540 7148
rect 62500 6866 62528 7142
rect 62488 6860 62540 6866
rect 62488 6802 62540 6808
rect 62304 5908 62356 5914
rect 62304 5850 62356 5856
rect 62316 5302 62344 5850
rect 62396 5568 62448 5574
rect 62396 5510 62448 5516
rect 62408 5302 62436 5510
rect 62304 5296 62356 5302
rect 62304 5238 62356 5244
rect 62396 5296 62448 5302
rect 62396 5238 62448 5244
rect 62212 4276 62264 4282
rect 62212 4218 62264 4224
rect 62028 4140 62080 4146
rect 62028 4082 62080 4088
rect 61292 4072 61344 4078
rect 61292 4014 61344 4020
rect 58532 3732 58584 3738
rect 58532 3674 58584 3680
rect 59268 3732 59320 3738
rect 59268 3674 59320 3680
rect 61200 3732 61252 3738
rect 61200 3674 61252 3680
rect 57336 3528 57388 3534
rect 57336 3470 57388 3476
rect 57348 3194 57376 3470
rect 57428 3392 57480 3398
rect 57428 3334 57480 3340
rect 57440 3194 57468 3334
rect 57336 3188 57388 3194
rect 57336 3130 57388 3136
rect 57428 3188 57480 3194
rect 57428 3130 57480 3136
rect 61304 3126 61332 4014
rect 62040 4010 62068 4082
rect 62028 4004 62080 4010
rect 62028 3946 62080 3952
rect 62224 3534 62252 4218
rect 62316 4214 62344 5238
rect 62304 4208 62356 4214
rect 62304 4150 62356 4156
rect 62212 3528 62264 3534
rect 62212 3470 62264 3476
rect 62316 3466 62344 4150
rect 62592 4146 62620 7511
rect 62684 7410 62712 7754
rect 63052 7546 63080 9522
rect 63130 9480 63186 9489
rect 63130 9415 63132 9424
rect 63184 9415 63186 9424
rect 63132 9386 63184 9392
rect 63236 8838 63264 9522
rect 63224 8832 63276 8838
rect 63224 8774 63276 8780
rect 63040 7540 63092 7546
rect 63040 7482 63092 7488
rect 62672 7404 62724 7410
rect 62672 7346 62724 7352
rect 62580 4140 62632 4146
rect 62580 4082 62632 4088
rect 62684 3942 62712 7346
rect 63236 6866 63264 8774
rect 63328 8294 63356 9590
rect 63420 8820 63448 10066
rect 63684 10056 63736 10062
rect 63512 10016 63684 10044
rect 63512 9926 63540 10016
rect 63684 9998 63736 10004
rect 63500 9920 63552 9926
rect 63500 9862 63552 9868
rect 63512 9042 63540 9862
rect 63788 9382 63816 10118
rect 64328 9648 64380 9654
rect 64328 9590 64380 9596
rect 64144 9512 64196 9518
rect 64144 9454 64196 9460
rect 63776 9376 63828 9382
rect 63776 9318 63828 9324
rect 63500 9036 63552 9042
rect 63500 8978 63552 8984
rect 63788 8974 63816 9318
rect 63776 8968 63828 8974
rect 63776 8910 63828 8916
rect 63420 8792 63724 8820
rect 63498 8664 63554 8673
rect 63498 8599 63554 8608
rect 63408 8356 63460 8362
rect 63408 8298 63460 8304
rect 63316 8288 63368 8294
rect 63316 8230 63368 8236
rect 63328 7449 63356 8230
rect 63314 7440 63370 7449
rect 63314 7375 63370 7384
rect 62948 6860 63000 6866
rect 62948 6802 63000 6808
rect 63224 6860 63276 6866
rect 63224 6802 63276 6808
rect 62960 4622 62988 6802
rect 63328 6118 63356 7375
rect 63316 6112 63368 6118
rect 63316 6054 63368 6060
rect 63328 5302 63356 6054
rect 63420 5914 63448 8298
rect 63512 7478 63540 8599
rect 63696 8498 63724 8792
rect 63774 8528 63830 8537
rect 63684 8492 63736 8498
rect 63774 8463 63830 8472
rect 63684 8434 63736 8440
rect 63696 8401 63724 8434
rect 63788 8430 63816 8463
rect 63776 8424 63828 8430
rect 63682 8392 63738 8401
rect 63776 8366 63828 8372
rect 64050 8392 64106 8401
rect 63682 8327 63738 8336
rect 64050 8327 64106 8336
rect 63500 7472 63552 7478
rect 63500 7414 63552 7420
rect 63868 7404 63920 7410
rect 63868 7346 63920 7352
rect 63500 6792 63552 6798
rect 63500 6734 63552 6740
rect 63512 6118 63540 6734
rect 63592 6316 63644 6322
rect 63592 6258 63644 6264
rect 63776 6316 63828 6322
rect 63776 6258 63828 6264
rect 63500 6112 63552 6118
rect 63500 6054 63552 6060
rect 63408 5908 63460 5914
rect 63408 5850 63460 5856
rect 63420 5642 63448 5850
rect 63512 5778 63540 6054
rect 63604 5846 63632 6258
rect 63592 5840 63644 5846
rect 63592 5782 63644 5788
rect 63500 5772 63552 5778
rect 63500 5714 63552 5720
rect 63408 5636 63460 5642
rect 63408 5578 63460 5584
rect 63316 5296 63368 5302
rect 63316 5238 63368 5244
rect 63512 5234 63540 5714
rect 63684 5704 63736 5710
rect 63684 5646 63736 5652
rect 63500 5228 63552 5234
rect 63500 5170 63552 5176
rect 63512 4826 63540 5170
rect 63696 5030 63724 5646
rect 63684 5024 63736 5030
rect 63684 4966 63736 4972
rect 63590 4856 63646 4865
rect 63500 4820 63552 4826
rect 63696 4826 63724 4966
rect 63590 4791 63646 4800
rect 63684 4820 63736 4826
rect 63500 4762 63552 4768
rect 62948 4616 63000 4622
rect 62948 4558 63000 4564
rect 62960 4146 62988 4558
rect 63512 4282 63540 4762
rect 63604 4690 63632 4791
rect 63684 4762 63736 4768
rect 63592 4684 63644 4690
rect 63592 4626 63644 4632
rect 63500 4276 63552 4282
rect 63500 4218 63552 4224
rect 62948 4140 63000 4146
rect 62948 4082 63000 4088
rect 63788 4010 63816 6258
rect 63880 5166 63908 7346
rect 63868 5160 63920 5166
rect 63868 5102 63920 5108
rect 63880 4622 63908 5102
rect 64064 4690 64092 8327
rect 64156 8294 64184 9454
rect 64340 8974 64368 9590
rect 64432 9518 64460 11290
rect 64616 11150 64644 13262
rect 64696 13184 64748 13190
rect 64696 13126 64748 13132
rect 65892 13184 65944 13190
rect 65892 13126 65944 13132
rect 64708 12306 64736 13126
rect 65904 12918 65932 13126
rect 65892 12912 65944 12918
rect 65892 12854 65944 12860
rect 64696 12300 64748 12306
rect 64696 12242 64748 12248
rect 65996 12238 66024 13262
rect 66180 12850 66208 13262
rect 66168 12844 66220 12850
rect 66168 12786 66220 12792
rect 65984 12232 66036 12238
rect 64786 12200 64842 12209
rect 65984 12174 66036 12180
rect 64786 12135 64842 12144
rect 64800 12102 64828 12135
rect 64788 12096 64840 12102
rect 64788 12038 64840 12044
rect 65892 12096 65944 12102
rect 65892 12038 65944 12044
rect 64800 11694 64828 12038
rect 65062 11928 65118 11937
rect 65062 11863 65118 11872
rect 65076 11694 65104 11863
rect 65904 11830 65932 12038
rect 65892 11824 65944 11830
rect 65892 11766 65944 11772
rect 66076 11824 66128 11830
rect 66076 11766 66128 11772
rect 64788 11688 64840 11694
rect 64788 11630 64840 11636
rect 65064 11688 65116 11694
rect 65064 11630 65116 11636
rect 64972 11620 65024 11626
rect 64972 11562 65024 11568
rect 65892 11620 65944 11626
rect 65892 11562 65944 11568
rect 64984 11354 65012 11562
rect 64972 11348 65024 11354
rect 64972 11290 65024 11296
rect 64604 11144 64656 11150
rect 64604 11086 64656 11092
rect 65432 11144 65484 11150
rect 65432 11086 65484 11092
rect 65444 10742 65472 11086
rect 65432 10736 65484 10742
rect 65432 10678 65484 10684
rect 65432 10192 65484 10198
rect 65432 10134 65484 10140
rect 64696 9988 64748 9994
rect 64696 9930 64748 9936
rect 64708 9654 64736 9930
rect 65444 9926 65472 10134
rect 65432 9920 65484 9926
rect 65432 9862 65484 9868
rect 65444 9722 65472 9862
rect 65432 9716 65484 9722
rect 65432 9658 65484 9664
rect 64696 9648 64748 9654
rect 64696 9590 64748 9596
rect 64420 9512 64472 9518
rect 64420 9454 64472 9460
rect 65800 9444 65852 9450
rect 65800 9386 65852 9392
rect 64236 8968 64288 8974
rect 64234 8936 64236 8945
rect 64328 8968 64380 8974
rect 64288 8936 64290 8945
rect 64328 8910 64380 8916
rect 64234 8871 64290 8880
rect 65812 8809 65840 9386
rect 65798 8800 65854 8809
rect 65798 8735 65854 8744
rect 64510 8664 64566 8673
rect 64510 8599 64566 8608
rect 64524 8498 64552 8599
rect 64512 8492 64564 8498
rect 64432 8452 64512 8480
rect 64144 8288 64196 8294
rect 64144 8230 64196 8236
rect 64156 7342 64184 8230
rect 64144 7336 64196 7342
rect 64144 7278 64196 7284
rect 64432 5098 64460 8452
rect 64512 8434 64564 8440
rect 64788 8424 64840 8430
rect 64788 8366 64840 8372
rect 64800 7750 64828 8366
rect 65156 7880 65208 7886
rect 65156 7822 65208 7828
rect 64788 7744 64840 7750
rect 64788 7686 64840 7692
rect 64512 7404 64564 7410
rect 64512 7346 64564 7352
rect 64696 7404 64748 7410
rect 64696 7346 64748 7352
rect 64524 6322 64552 7346
rect 64708 6322 64736 7346
rect 64512 6316 64564 6322
rect 64512 6258 64564 6264
rect 64696 6316 64748 6322
rect 64696 6258 64748 6264
rect 64524 5574 64552 6258
rect 64604 6180 64656 6186
rect 64604 6122 64656 6128
rect 64616 5778 64644 6122
rect 64708 5846 64736 6258
rect 64696 5840 64748 5846
rect 64696 5782 64748 5788
rect 64604 5772 64656 5778
rect 64604 5714 64656 5720
rect 64512 5568 64564 5574
rect 64512 5510 64564 5516
rect 64420 5092 64472 5098
rect 64420 5034 64472 5040
rect 64432 4690 64460 5034
rect 64052 4684 64104 4690
rect 64052 4626 64104 4632
rect 64420 4684 64472 4690
rect 64420 4626 64472 4632
rect 63868 4616 63920 4622
rect 63868 4558 63920 4564
rect 63776 4004 63828 4010
rect 63776 3946 63828 3952
rect 62672 3936 62724 3942
rect 62672 3878 62724 3884
rect 64616 3738 64644 5714
rect 64708 5302 64736 5782
rect 64696 5296 64748 5302
rect 64696 5238 64748 5244
rect 64708 4758 64736 5238
rect 64696 4752 64748 4758
rect 64696 4694 64748 4700
rect 64604 3732 64656 3738
rect 64604 3674 64656 3680
rect 64328 3596 64380 3602
rect 64328 3538 64380 3544
rect 62304 3460 62356 3466
rect 62304 3402 62356 3408
rect 62316 3126 62344 3402
rect 61292 3120 61344 3126
rect 61292 3062 61344 3068
rect 62304 3120 62356 3126
rect 62304 3062 62356 3068
rect 57060 2916 57112 2922
rect 57060 2858 57112 2864
rect 59542 2748 59850 2757
rect 59542 2746 59548 2748
rect 59604 2746 59628 2748
rect 59684 2746 59708 2748
rect 59764 2746 59788 2748
rect 59844 2746 59850 2748
rect 59604 2694 59606 2746
rect 59786 2694 59788 2746
rect 59542 2692 59548 2694
rect 59604 2692 59628 2694
rect 59684 2692 59708 2694
rect 59764 2692 59788 2694
rect 59844 2692 59850 2694
rect 59542 2683 59850 2692
rect 64340 2650 64368 3538
rect 64616 3534 64644 3674
rect 64708 3670 64736 4694
rect 64800 4078 64828 7686
rect 65168 7206 65196 7822
rect 65616 7404 65668 7410
rect 65616 7346 65668 7352
rect 65340 7336 65392 7342
rect 65340 7278 65392 7284
rect 65156 7200 65208 7206
rect 65156 7142 65208 7148
rect 65168 7002 65196 7142
rect 65156 6996 65208 7002
rect 65156 6938 65208 6944
rect 65156 6860 65208 6866
rect 65156 6802 65208 6808
rect 64880 6792 64932 6798
rect 64880 6734 64932 6740
rect 64892 5642 64920 6734
rect 65168 6322 65196 6802
rect 65248 6656 65300 6662
rect 65248 6598 65300 6604
rect 65156 6316 65208 6322
rect 65156 6258 65208 6264
rect 65260 6118 65288 6598
rect 65352 6322 65380 7278
rect 65432 6860 65484 6866
rect 65432 6802 65484 6808
rect 65444 6730 65472 6802
rect 65432 6724 65484 6730
rect 65432 6666 65484 6672
rect 65628 6458 65656 7346
rect 65616 6452 65668 6458
rect 65616 6394 65668 6400
rect 65708 6452 65760 6458
rect 65708 6394 65760 6400
rect 65340 6316 65392 6322
rect 65340 6258 65392 6264
rect 65248 6112 65300 6118
rect 65248 6054 65300 6060
rect 64880 5636 64932 5642
rect 64880 5578 64932 5584
rect 65352 5234 65380 6258
rect 65720 5846 65748 6394
rect 65904 6118 65932 11562
rect 65984 11144 66036 11150
rect 65984 11086 66036 11092
rect 65996 9761 66024 11086
rect 66088 10538 66116 11766
rect 66168 11688 66220 11694
rect 66168 11630 66220 11636
rect 66076 10532 66128 10538
rect 66076 10474 66128 10480
rect 65982 9752 66038 9761
rect 65982 9687 66038 9696
rect 66180 9042 66208 11630
rect 66168 9036 66220 9042
rect 66168 8978 66220 8984
rect 66260 9036 66312 9042
rect 66260 8978 66312 8984
rect 66076 8288 66128 8294
rect 66076 8230 66128 8236
rect 66088 7954 66116 8230
rect 66272 8022 66300 8978
rect 66260 8016 66312 8022
rect 66260 7958 66312 7964
rect 66364 7954 66392 13790
rect 66536 13728 66588 13734
rect 66536 13670 66588 13676
rect 66548 12986 66576 13670
rect 66718 13560 66774 13569
rect 66718 13495 66774 13504
rect 66628 13252 66680 13258
rect 66628 13194 66680 13200
rect 66640 12986 66668 13194
rect 66536 12980 66588 12986
rect 66536 12922 66588 12928
rect 66628 12980 66680 12986
rect 66628 12922 66680 12928
rect 66732 12918 66760 13495
rect 67088 13184 67140 13190
rect 67088 13126 67140 13132
rect 66720 12912 66772 12918
rect 66720 12854 66772 12860
rect 66904 12844 66956 12850
rect 66904 12786 66956 12792
rect 66628 12232 66680 12238
rect 66628 12174 66680 12180
rect 66536 12164 66588 12170
rect 66536 12106 66588 12112
rect 66442 11384 66498 11393
rect 66548 11354 66576 12106
rect 66442 11319 66498 11328
rect 66536 11348 66588 11354
rect 66456 11286 66484 11319
rect 66536 11290 66588 11296
rect 66444 11280 66496 11286
rect 66444 11222 66496 11228
rect 66640 11218 66668 12174
rect 66916 11626 66944 12786
rect 67100 12782 67128 13126
rect 67192 13025 67220 14962
rect 67652 14482 67680 15506
rect 67928 15502 67956 15846
rect 67916 15496 67968 15502
rect 67916 15438 67968 15444
rect 67824 15428 67876 15434
rect 67824 15370 67876 15376
rect 67732 14816 67784 14822
rect 67732 14758 67784 14764
rect 67640 14476 67692 14482
rect 67640 14418 67692 14424
rect 67744 14414 67772 14758
rect 67272 14408 67324 14414
rect 67272 14350 67324 14356
rect 67732 14408 67784 14414
rect 67732 14350 67784 14356
rect 67178 13016 67234 13025
rect 67178 12951 67234 12960
rect 67088 12776 67140 12782
rect 67088 12718 67140 12724
rect 67100 12442 67128 12718
rect 67088 12436 67140 12442
rect 67088 12378 67140 12384
rect 67086 12064 67142 12073
rect 67086 11999 67142 12008
rect 67100 11626 67128 11999
rect 66904 11620 66956 11626
rect 66904 11562 66956 11568
rect 67088 11620 67140 11626
rect 67088 11562 67140 11568
rect 66628 11212 66680 11218
rect 66628 11154 66680 11160
rect 67088 11076 67140 11082
rect 67088 11018 67140 11024
rect 66628 9988 66680 9994
rect 66628 9930 66680 9936
rect 66444 9580 66496 9586
rect 66444 9522 66496 9528
rect 66076 7948 66128 7954
rect 66076 7890 66128 7896
rect 66352 7948 66404 7954
rect 66352 7890 66404 7896
rect 66456 7834 66484 9522
rect 66536 8900 66588 8906
rect 66536 8842 66588 8848
rect 66548 8294 66576 8842
rect 66640 8838 66668 9930
rect 66720 9376 66772 9382
rect 66720 9318 66772 9324
rect 66732 9110 66760 9318
rect 66720 9104 66772 9110
rect 67100 9081 67128 11018
rect 66720 9046 66772 9052
rect 67086 9072 67142 9081
rect 67086 9007 67142 9016
rect 66996 8900 67048 8906
rect 66996 8842 67048 8848
rect 66628 8832 66680 8838
rect 66628 8774 66680 8780
rect 66812 8560 66864 8566
rect 66812 8502 66864 8508
rect 66548 8266 66760 8294
rect 66732 7857 66760 8266
rect 66364 7806 66484 7834
rect 66718 7848 66774 7857
rect 66364 7410 66392 7806
rect 66718 7783 66774 7792
rect 66626 7440 66682 7449
rect 66352 7404 66404 7410
rect 66732 7410 66760 7783
rect 66626 7375 66682 7384
rect 66720 7404 66772 7410
rect 66352 7346 66404 7352
rect 66640 7206 66668 7375
rect 66720 7346 66772 7352
rect 66628 7200 66680 7206
rect 66628 7142 66680 7148
rect 66824 6798 66852 8502
rect 67008 8294 67036 8842
rect 66996 8288 67048 8294
rect 66996 8230 67048 8236
rect 67088 7268 67140 7274
rect 67088 7210 67140 7216
rect 67100 7177 67128 7210
rect 67086 7168 67142 7177
rect 67086 7103 67142 7112
rect 67192 7041 67220 12951
rect 67284 11694 67312 14350
rect 67454 14104 67510 14113
rect 67454 14039 67456 14048
rect 67508 14039 67510 14048
rect 67456 14010 67508 14016
rect 67364 11756 67416 11762
rect 67364 11698 67416 11704
rect 67272 11688 67324 11694
rect 67272 11630 67324 11636
rect 67284 11558 67312 11630
rect 67272 11552 67324 11558
rect 67272 11494 67324 11500
rect 67272 11348 67324 11354
rect 67272 11290 67324 11296
rect 67284 9178 67312 11290
rect 67376 10606 67404 11698
rect 67468 11354 67496 14010
rect 67744 14006 67772 14350
rect 67732 14000 67784 14006
rect 67732 13942 67784 13948
rect 67836 12850 67864 15370
rect 68020 15348 68048 15846
rect 67928 15320 68048 15348
rect 67928 13161 67956 15320
rect 68204 14414 68232 16662
rect 68388 15162 68416 17138
rect 68744 16516 68796 16522
rect 68744 16458 68796 16464
rect 68756 15366 68784 16458
rect 69020 15904 69072 15910
rect 69020 15846 69072 15852
rect 68744 15360 68796 15366
rect 68744 15302 68796 15308
rect 68376 15156 68428 15162
rect 68376 15098 68428 15104
rect 68468 14816 68520 14822
rect 68468 14758 68520 14764
rect 68480 14521 68508 14758
rect 68466 14512 68522 14521
rect 68466 14447 68522 14456
rect 68560 14476 68612 14482
rect 68560 14418 68612 14424
rect 68192 14408 68244 14414
rect 68190 14376 68192 14385
rect 68244 14376 68246 14385
rect 68190 14311 68246 14320
rect 68468 14340 68520 14346
rect 68468 14282 68520 14288
rect 68008 13728 68060 13734
rect 68480 13705 68508 14282
rect 68008 13670 68060 13676
rect 68466 13696 68522 13705
rect 67914 13152 67970 13161
rect 67914 13087 67970 13096
rect 67928 12850 67956 13087
rect 67824 12844 67876 12850
rect 67824 12786 67876 12792
rect 67916 12844 67968 12850
rect 67916 12786 67968 12792
rect 67640 12436 67692 12442
rect 68020 12434 68048 13670
rect 68466 13631 68522 13640
rect 68282 13560 68338 13569
rect 68282 13495 68338 13504
rect 68296 12782 68324 13495
rect 68468 12844 68520 12850
rect 68468 12786 68520 12792
rect 68284 12776 68336 12782
rect 68284 12718 68336 12724
rect 68376 12708 68428 12714
rect 68376 12650 68428 12656
rect 67640 12378 67692 12384
rect 67928 12406 68048 12434
rect 67548 12300 67600 12306
rect 67548 12242 67600 12248
rect 67560 12209 67588 12242
rect 67546 12200 67602 12209
rect 67546 12135 67602 12144
rect 67652 12102 67680 12378
rect 67640 12096 67692 12102
rect 67640 12038 67692 12044
rect 67732 12096 67784 12102
rect 67732 12038 67784 12044
rect 67744 11830 67772 12038
rect 67732 11824 67784 11830
rect 67732 11766 67784 11772
rect 67824 11756 67876 11762
rect 67824 11698 67876 11704
rect 67456 11348 67508 11354
rect 67456 11290 67508 11296
rect 67456 11008 67508 11014
rect 67456 10950 67508 10956
rect 67364 10600 67416 10606
rect 67364 10542 67416 10548
rect 67376 10062 67404 10542
rect 67468 10266 67496 10950
rect 67732 10668 67784 10674
rect 67732 10610 67784 10616
rect 67640 10464 67692 10470
rect 67640 10406 67692 10412
rect 67456 10260 67508 10266
rect 67456 10202 67508 10208
rect 67364 10056 67416 10062
rect 67364 9998 67416 10004
rect 67652 9654 67680 10406
rect 67640 9648 67692 9654
rect 67640 9590 67692 9596
rect 67454 9480 67510 9489
rect 67454 9415 67510 9424
rect 67638 9480 67694 9489
rect 67638 9415 67694 9424
rect 67364 9376 67416 9382
rect 67364 9318 67416 9324
rect 67272 9172 67324 9178
rect 67272 9114 67324 9120
rect 67272 7948 67324 7954
rect 67272 7890 67324 7896
rect 67284 7206 67312 7890
rect 67376 7342 67404 9318
rect 67468 9024 67496 9415
rect 67652 9024 67680 9415
rect 67468 8996 67680 9024
rect 67548 8832 67600 8838
rect 67548 8774 67600 8780
rect 67640 8832 67692 8838
rect 67640 8774 67692 8780
rect 67560 8566 67588 8774
rect 67548 8560 67600 8566
rect 67548 8502 67600 8508
rect 67548 8424 67600 8430
rect 67548 8366 67600 8372
rect 67456 8288 67508 8294
rect 67456 8230 67508 8236
rect 67468 7410 67496 8230
rect 67560 7698 67588 8366
rect 67652 7818 67680 8774
rect 67640 7812 67692 7818
rect 67640 7754 67692 7760
rect 67744 7750 67772 10610
rect 67836 10470 67864 11698
rect 67824 10464 67876 10470
rect 67824 10406 67876 10412
rect 67836 10198 67864 10406
rect 67824 10192 67876 10198
rect 67824 10134 67876 10140
rect 67928 9897 67956 12406
rect 68388 11830 68416 12650
rect 68376 11824 68428 11830
rect 68376 11766 68428 11772
rect 68008 11756 68060 11762
rect 68008 11698 68060 11704
rect 67914 9888 67970 9897
rect 67914 9823 67970 9832
rect 67916 9648 67968 9654
rect 67916 9590 67968 9596
rect 67824 9580 67876 9586
rect 67824 9522 67876 9528
rect 67836 9353 67864 9522
rect 67822 9344 67878 9353
rect 67822 9279 67878 9288
rect 67928 7750 67956 9590
rect 68020 9489 68048 11698
rect 68282 10840 68338 10849
rect 68282 10775 68338 10784
rect 68296 10674 68324 10775
rect 68284 10668 68336 10674
rect 68284 10610 68336 10616
rect 68376 10600 68428 10606
rect 68376 10542 68428 10548
rect 68388 10062 68416 10542
rect 68480 10441 68508 12786
rect 68572 11150 68600 14418
rect 68756 14090 68784 15302
rect 69032 15026 69060 15846
rect 69020 15020 69072 15026
rect 69020 14962 69072 14968
rect 69296 14272 69348 14278
rect 69296 14214 69348 14220
rect 68756 14062 68876 14090
rect 68652 13796 68704 13802
rect 68652 13738 68704 13744
rect 68664 12714 68692 13738
rect 68848 12968 68876 14062
rect 69020 13524 69072 13530
rect 69020 13466 69072 13472
rect 68756 12940 68876 12968
rect 68652 12708 68704 12714
rect 68652 12650 68704 12656
rect 68756 12170 68784 12940
rect 69032 12918 69060 13466
rect 69020 12912 69072 12918
rect 69020 12854 69072 12860
rect 68836 12844 68888 12850
rect 68836 12786 68888 12792
rect 68744 12164 68796 12170
rect 68744 12106 68796 12112
rect 68560 11144 68612 11150
rect 68560 11086 68612 11092
rect 68744 10736 68796 10742
rect 68744 10678 68796 10684
rect 68756 10606 68784 10678
rect 68652 10600 68704 10606
rect 68652 10542 68704 10548
rect 68744 10600 68796 10606
rect 68744 10542 68796 10548
rect 68466 10432 68522 10441
rect 68466 10367 68522 10376
rect 68664 10266 68692 10542
rect 68652 10260 68704 10266
rect 68652 10202 68704 10208
rect 68376 10056 68428 10062
rect 68376 9998 68428 10004
rect 68468 9988 68520 9994
rect 68468 9930 68520 9936
rect 68006 9480 68062 9489
rect 68006 9415 68062 9424
rect 68480 9042 68508 9930
rect 68848 9926 68876 12786
rect 69308 12782 69336 14214
rect 69296 12776 69348 12782
rect 69296 12718 69348 12724
rect 69570 12472 69626 12481
rect 69570 12407 69626 12416
rect 69676 12434 69704 17478
rect 71260 17436 71568 17445
rect 71260 17434 71266 17436
rect 71322 17434 71346 17436
rect 71402 17434 71426 17436
rect 71482 17434 71506 17436
rect 71562 17434 71568 17436
rect 71322 17382 71324 17434
rect 71504 17382 71506 17434
rect 71260 17380 71266 17382
rect 71322 17380 71346 17382
rect 71402 17380 71426 17382
rect 71482 17380 71506 17382
rect 71562 17380 71568 17382
rect 71260 17371 71568 17380
rect 75656 17338 75684 19200
rect 75644 17332 75696 17338
rect 75644 17274 75696 17280
rect 76104 17196 76156 17202
rect 76104 17138 76156 17144
rect 71964 16448 72016 16454
rect 71964 16390 72016 16396
rect 71260 16348 71568 16357
rect 71260 16346 71266 16348
rect 71322 16346 71346 16348
rect 71402 16346 71426 16348
rect 71482 16346 71506 16348
rect 71562 16346 71568 16348
rect 71322 16294 71324 16346
rect 71504 16294 71506 16346
rect 71260 16292 71266 16294
rect 71322 16292 71346 16294
rect 71402 16292 71426 16294
rect 71482 16292 71506 16294
rect 71562 16292 71568 16294
rect 71260 16283 71568 16292
rect 71976 16250 72004 16390
rect 71964 16244 72016 16250
rect 71964 16186 72016 16192
rect 72148 16244 72200 16250
rect 72148 16186 72200 16192
rect 72056 16176 72108 16182
rect 72056 16118 72108 16124
rect 71136 16108 71188 16114
rect 71136 16050 71188 16056
rect 69756 15904 69808 15910
rect 69756 15846 69808 15852
rect 71044 15904 71096 15910
rect 71044 15846 71096 15852
rect 69768 14958 69796 15846
rect 70492 15632 70544 15638
rect 70492 15574 70544 15580
rect 70308 15564 70360 15570
rect 70308 15506 70360 15512
rect 69848 15360 69900 15366
rect 69848 15302 69900 15308
rect 69756 14952 69808 14958
rect 69756 14894 69808 14900
rect 69768 13433 69796 14894
rect 69754 13424 69810 13433
rect 69754 13359 69810 13368
rect 69860 13326 69888 15302
rect 69940 14272 69992 14278
rect 69940 14214 69992 14220
rect 69848 13320 69900 13326
rect 69848 13262 69900 13268
rect 69204 12368 69256 12374
rect 69204 12310 69256 12316
rect 69216 11150 69244 12310
rect 69478 12200 69534 12209
rect 69478 12135 69534 12144
rect 69492 11558 69520 12135
rect 69480 11552 69532 11558
rect 69480 11494 69532 11500
rect 69204 11144 69256 11150
rect 69204 11086 69256 11092
rect 69480 11144 69532 11150
rect 69480 11086 69532 11092
rect 68836 9920 68888 9926
rect 68836 9862 68888 9868
rect 68836 9512 68888 9518
rect 68836 9454 68888 9460
rect 68192 9036 68244 9042
rect 68192 8978 68244 8984
rect 68468 9036 68520 9042
rect 68468 8978 68520 8984
rect 68204 8906 68232 8978
rect 68192 8900 68244 8906
rect 68192 8842 68244 8848
rect 68192 8424 68244 8430
rect 68192 8366 68244 8372
rect 68560 8424 68612 8430
rect 68560 8366 68612 8372
rect 67732 7744 67784 7750
rect 67560 7670 67680 7698
rect 67916 7744 67968 7750
rect 67732 7686 67784 7692
rect 67836 7704 67916 7732
rect 67652 7546 67680 7670
rect 67548 7540 67600 7546
rect 67548 7482 67600 7488
rect 67640 7540 67692 7546
rect 67640 7482 67692 7488
rect 67560 7426 67588 7482
rect 67836 7426 67864 7704
rect 67916 7686 67968 7692
rect 68008 7540 68060 7546
rect 68008 7482 68060 7488
rect 68020 7449 68048 7482
rect 67456 7404 67508 7410
rect 67560 7398 67864 7426
rect 68006 7440 68062 7449
rect 68006 7375 68062 7384
rect 68100 7404 68152 7410
rect 67456 7346 67508 7352
rect 68100 7346 68152 7352
rect 67364 7336 67416 7342
rect 67364 7278 67416 7284
rect 67272 7200 67324 7206
rect 67272 7142 67324 7148
rect 67178 7032 67234 7041
rect 67178 6967 67234 6976
rect 67824 6996 67876 7002
rect 66812 6792 66864 6798
rect 66812 6734 66864 6740
rect 66076 6724 66128 6730
rect 66076 6666 66128 6672
rect 66088 6322 66116 6666
rect 66626 6488 66682 6497
rect 66626 6423 66682 6432
rect 66076 6316 66128 6322
rect 66076 6258 66128 6264
rect 66168 6248 66220 6254
rect 66168 6190 66220 6196
rect 65892 6112 65944 6118
rect 65892 6054 65944 6060
rect 66076 6112 66128 6118
rect 66076 6054 66128 6060
rect 65708 5840 65760 5846
rect 65708 5782 65760 5788
rect 65904 5302 65932 6054
rect 66088 5778 66116 6054
rect 66180 5778 66208 6190
rect 66640 6186 66668 6423
rect 66628 6180 66680 6186
rect 66628 6122 66680 6128
rect 66076 5772 66128 5778
rect 66076 5714 66128 5720
rect 66168 5772 66220 5778
rect 66168 5714 66220 5720
rect 65892 5296 65944 5302
rect 65892 5238 65944 5244
rect 65340 5228 65392 5234
rect 65340 5170 65392 5176
rect 65352 4758 65380 5170
rect 65340 4752 65392 4758
rect 65340 4694 65392 4700
rect 66824 4554 66852 6734
rect 66812 4548 66864 4554
rect 66812 4490 66864 4496
rect 64788 4072 64840 4078
rect 64788 4014 64840 4020
rect 64880 4004 64932 4010
rect 64880 3946 64932 3952
rect 64892 3890 64920 3946
rect 64800 3862 64920 3890
rect 64696 3664 64748 3670
rect 64696 3606 64748 3612
rect 64604 3528 64656 3534
rect 64604 3470 64656 3476
rect 64800 3194 64828 3862
rect 67192 3738 67220 6967
rect 67824 6938 67876 6944
rect 67836 6905 67864 6938
rect 67822 6896 67878 6905
rect 67822 6831 67878 6840
rect 67640 6656 67692 6662
rect 67640 6598 67692 6604
rect 67652 6458 67680 6598
rect 67640 6452 67692 6458
rect 67640 6394 67692 6400
rect 67456 6384 67508 6390
rect 67456 6326 67508 6332
rect 67732 6384 67784 6390
rect 67732 6326 67784 6332
rect 67364 5908 67416 5914
rect 67364 5850 67416 5856
rect 67376 4690 67404 5850
rect 67468 5642 67496 6326
rect 67548 6316 67600 6322
rect 67548 6258 67600 6264
rect 67560 5846 67588 6258
rect 67548 5840 67600 5846
rect 67548 5782 67600 5788
rect 67744 5710 67772 6326
rect 68112 6118 68140 7346
rect 68204 6798 68232 8366
rect 68284 7200 68336 7206
rect 68284 7142 68336 7148
rect 68468 7200 68520 7206
rect 68468 7142 68520 7148
rect 68296 6934 68324 7142
rect 68480 7002 68508 7142
rect 68468 6996 68520 7002
rect 68468 6938 68520 6944
rect 68284 6928 68336 6934
rect 68284 6870 68336 6876
rect 68192 6792 68244 6798
rect 68192 6734 68244 6740
rect 68100 6112 68152 6118
rect 68100 6054 68152 6060
rect 68112 5914 68140 6054
rect 68100 5908 68152 5914
rect 68100 5850 68152 5856
rect 67732 5704 67784 5710
rect 67732 5646 67784 5652
rect 67456 5636 67508 5642
rect 67456 5578 67508 5584
rect 67640 5568 67692 5574
rect 67640 5510 67692 5516
rect 67652 4690 67680 5510
rect 67744 5302 67772 5646
rect 68204 5574 68232 6734
rect 68572 6458 68600 8366
rect 68848 7585 68876 9454
rect 69112 8288 69164 8294
rect 69112 8230 69164 8236
rect 69124 8022 69152 8230
rect 69112 8016 69164 8022
rect 69112 7958 69164 7964
rect 68834 7576 68890 7585
rect 68834 7511 68890 7520
rect 68652 7336 68704 7342
rect 68652 7278 68704 7284
rect 68836 7336 68888 7342
rect 69492 7313 69520 11086
rect 69584 10305 69612 12407
rect 69676 12406 69796 12434
rect 69768 11665 69796 12406
rect 69860 11898 69888 13262
rect 69952 12442 69980 14214
rect 70320 13326 70348 15506
rect 70308 13320 70360 13326
rect 70308 13262 70360 13268
rect 70504 12850 70532 15574
rect 70860 15496 70912 15502
rect 70860 15438 70912 15444
rect 70872 15366 70900 15438
rect 70860 15360 70912 15366
rect 70860 15302 70912 15308
rect 70872 14260 70900 15302
rect 70952 15156 71004 15162
rect 70952 15098 71004 15104
rect 70964 14414 70992 15098
rect 71056 15094 71084 15846
rect 71148 15570 71176 16050
rect 72068 15570 72096 16118
rect 71136 15564 71188 15570
rect 71136 15506 71188 15512
rect 72056 15564 72108 15570
rect 72056 15506 72108 15512
rect 71596 15360 71648 15366
rect 71596 15302 71648 15308
rect 71260 15260 71568 15269
rect 71260 15258 71266 15260
rect 71322 15258 71346 15260
rect 71402 15258 71426 15260
rect 71482 15258 71506 15260
rect 71562 15258 71568 15260
rect 71322 15206 71324 15258
rect 71504 15206 71506 15258
rect 71260 15204 71266 15206
rect 71322 15204 71346 15206
rect 71402 15204 71426 15206
rect 71482 15204 71506 15206
rect 71562 15204 71568 15206
rect 71260 15195 71568 15204
rect 71044 15088 71096 15094
rect 71044 15030 71096 15036
rect 71504 15020 71556 15026
rect 71504 14962 71556 14968
rect 71044 14952 71096 14958
rect 71044 14894 71096 14900
rect 71056 14482 71084 14894
rect 71516 14550 71544 14962
rect 71504 14544 71556 14550
rect 71504 14486 71556 14492
rect 71044 14476 71096 14482
rect 71044 14418 71096 14424
rect 70952 14408 71004 14414
rect 70952 14350 71004 14356
rect 71044 14340 71096 14346
rect 71044 14282 71096 14288
rect 70872 14232 70992 14260
rect 70674 13968 70730 13977
rect 70674 13903 70730 13912
rect 70688 13802 70716 13903
rect 70676 13796 70728 13802
rect 70676 13738 70728 13744
rect 70768 13796 70820 13802
rect 70768 13738 70820 13744
rect 70780 12918 70808 13738
rect 70860 13728 70912 13734
rect 70860 13670 70912 13676
rect 70872 13530 70900 13670
rect 70860 13524 70912 13530
rect 70860 13466 70912 13472
rect 70768 12912 70820 12918
rect 70768 12854 70820 12860
rect 70492 12844 70544 12850
rect 70492 12786 70544 12792
rect 70964 12646 70992 14232
rect 71056 13530 71084 14282
rect 71260 14172 71568 14181
rect 71260 14170 71266 14172
rect 71322 14170 71346 14172
rect 71402 14170 71426 14172
rect 71482 14170 71506 14172
rect 71562 14170 71568 14172
rect 71322 14118 71324 14170
rect 71504 14118 71506 14170
rect 71260 14116 71266 14118
rect 71322 14116 71346 14118
rect 71402 14116 71426 14118
rect 71482 14116 71506 14118
rect 71562 14116 71568 14118
rect 71260 14107 71568 14116
rect 71608 14006 71636 15302
rect 72068 15026 72096 15506
rect 72160 15502 72188 16186
rect 74264 15904 74316 15910
rect 74264 15846 74316 15852
rect 73252 15700 73304 15706
rect 73252 15642 73304 15648
rect 72424 15632 72476 15638
rect 72608 15632 72660 15638
rect 72476 15580 72608 15586
rect 72424 15574 72660 15580
rect 72436 15558 72648 15574
rect 72148 15496 72200 15502
rect 72148 15438 72200 15444
rect 72056 15020 72108 15026
rect 72056 14962 72108 14968
rect 72160 14890 72188 15438
rect 73264 14958 73292 15642
rect 74172 15496 74224 15502
rect 74172 15438 74224 15444
rect 74184 15162 74212 15438
rect 74172 15156 74224 15162
rect 74172 15098 74224 15104
rect 74276 15026 74304 15846
rect 74632 15632 74684 15638
rect 74632 15574 74684 15580
rect 74540 15156 74592 15162
rect 74540 15098 74592 15104
rect 74264 15020 74316 15026
rect 74264 14962 74316 14968
rect 73252 14952 73304 14958
rect 73252 14894 73304 14900
rect 72148 14884 72200 14890
rect 72148 14826 72200 14832
rect 73528 14408 73580 14414
rect 73528 14350 73580 14356
rect 71872 14340 71924 14346
rect 71872 14282 71924 14288
rect 71596 14000 71648 14006
rect 71596 13942 71648 13948
rect 71884 13530 71912 14282
rect 72056 14272 72108 14278
rect 72056 14214 72108 14220
rect 72332 14272 72384 14278
rect 72332 14214 72384 14220
rect 71044 13524 71096 13530
rect 71044 13466 71096 13472
rect 71872 13524 71924 13530
rect 71872 13466 71924 13472
rect 71134 13424 71190 13433
rect 71134 13359 71190 13368
rect 70124 12640 70176 12646
rect 70124 12582 70176 12588
rect 70952 12640 71004 12646
rect 71148 12617 71176 13359
rect 71780 13252 71832 13258
rect 71780 13194 71832 13200
rect 71688 13184 71740 13190
rect 71688 13126 71740 13132
rect 71260 13084 71568 13093
rect 71260 13082 71266 13084
rect 71322 13082 71346 13084
rect 71402 13082 71426 13084
rect 71482 13082 71506 13084
rect 71562 13082 71568 13084
rect 71322 13030 71324 13082
rect 71504 13030 71506 13082
rect 71260 13028 71266 13030
rect 71322 13028 71346 13030
rect 71402 13028 71426 13030
rect 71482 13028 71506 13030
rect 71562 13028 71568 13030
rect 71260 13019 71568 13028
rect 71700 13025 71728 13126
rect 71686 13016 71742 13025
rect 71686 12951 71742 12960
rect 71228 12640 71280 12646
rect 70952 12582 71004 12588
rect 71134 12608 71190 12617
rect 69940 12436 69992 12442
rect 69940 12378 69992 12384
rect 69848 11892 69900 11898
rect 69848 11834 69900 11840
rect 69952 11830 69980 12378
rect 69940 11824 69992 11830
rect 69940 11766 69992 11772
rect 69754 11656 69810 11665
rect 69754 11591 69810 11600
rect 69664 11552 69716 11558
rect 69664 11494 69716 11500
rect 69676 10810 69704 11494
rect 69768 11218 69796 11591
rect 69756 11212 69808 11218
rect 69756 11154 69808 11160
rect 69664 10804 69716 10810
rect 69664 10746 69716 10752
rect 69664 10532 69716 10538
rect 69664 10474 69716 10480
rect 69570 10296 69626 10305
rect 69570 10231 69626 10240
rect 69676 10130 69704 10474
rect 70136 10130 70164 12582
rect 70768 12164 70820 12170
rect 70768 12106 70820 12112
rect 70308 12096 70360 12102
rect 70308 12038 70360 12044
rect 70320 10742 70348 12038
rect 70676 11688 70728 11694
rect 70676 11630 70728 11636
rect 70688 11150 70716 11630
rect 70676 11144 70728 11150
rect 70676 11086 70728 11092
rect 70582 10840 70638 10849
rect 70582 10775 70638 10784
rect 70308 10736 70360 10742
rect 70308 10678 70360 10684
rect 70596 10724 70624 10775
rect 70676 10736 70728 10742
rect 70596 10696 70676 10724
rect 70400 10600 70452 10606
rect 70400 10542 70452 10548
rect 69664 10124 69716 10130
rect 69664 10066 69716 10072
rect 70124 10124 70176 10130
rect 70124 10066 70176 10072
rect 70306 9752 70362 9761
rect 70412 9722 70440 10542
rect 70492 10464 70544 10470
rect 70492 10406 70544 10412
rect 70306 9687 70362 9696
rect 70400 9716 70452 9722
rect 70214 9480 70270 9489
rect 70214 9415 70270 9424
rect 70228 9178 70256 9415
rect 70320 9178 70348 9687
rect 70400 9658 70452 9664
rect 70504 9654 70532 10406
rect 70492 9648 70544 9654
rect 70492 9590 70544 9596
rect 70400 9580 70452 9586
rect 70400 9522 70452 9528
rect 70412 9382 70440 9522
rect 70400 9376 70452 9382
rect 70400 9318 70452 9324
rect 70216 9172 70268 9178
rect 70216 9114 70268 9120
rect 70308 9172 70360 9178
rect 70308 9114 70360 9120
rect 69940 8968 69992 8974
rect 69940 8910 69992 8916
rect 69952 8838 69980 8910
rect 69940 8832 69992 8838
rect 69940 8774 69992 8780
rect 69756 8560 69808 8566
rect 69756 8502 69808 8508
rect 69768 7886 69796 8502
rect 70596 7886 70624 10696
rect 70676 10678 70728 10684
rect 70780 10554 70808 12106
rect 70964 11370 70992 12582
rect 71228 12582 71280 12588
rect 71318 12608 71374 12617
rect 71134 12543 71190 12552
rect 71042 12472 71098 12481
rect 71042 12407 71098 12416
rect 71056 12306 71084 12407
rect 71240 12374 71268 12582
rect 71318 12543 71374 12552
rect 71228 12368 71280 12374
rect 71228 12310 71280 12316
rect 71044 12300 71096 12306
rect 71044 12242 71096 12248
rect 71332 12102 71360 12543
rect 71504 12232 71556 12238
rect 71556 12180 71636 12186
rect 71504 12174 71636 12180
rect 71516 12158 71636 12174
rect 71136 12096 71188 12102
rect 71136 12038 71188 12044
rect 71320 12096 71372 12102
rect 71320 12038 71372 12044
rect 71148 11762 71176 12038
rect 71260 11996 71568 12005
rect 71260 11994 71266 11996
rect 71322 11994 71346 11996
rect 71402 11994 71426 11996
rect 71482 11994 71506 11996
rect 71562 11994 71568 11996
rect 71322 11942 71324 11994
rect 71504 11942 71506 11994
rect 71260 11940 71266 11942
rect 71322 11940 71346 11942
rect 71402 11940 71426 11942
rect 71482 11940 71506 11942
rect 71562 11940 71568 11942
rect 71260 11931 71568 11940
rect 71136 11756 71188 11762
rect 71136 11698 71188 11704
rect 71608 11558 71636 12158
rect 71792 11898 71820 13194
rect 71962 13152 72018 13161
rect 71962 13087 72018 13096
rect 71976 12782 72004 13087
rect 72068 12918 72096 14214
rect 72056 12912 72108 12918
rect 72056 12854 72108 12860
rect 71964 12776 72016 12782
rect 71964 12718 72016 12724
rect 72240 12300 72292 12306
rect 72240 12242 72292 12248
rect 71780 11892 71832 11898
rect 71780 11834 71832 11840
rect 72252 11762 72280 12242
rect 72056 11756 72108 11762
rect 72056 11698 72108 11704
rect 72240 11756 72292 11762
rect 72240 11698 72292 11704
rect 71596 11552 71648 11558
rect 71596 11494 71648 11500
rect 71134 11384 71190 11393
rect 70964 11342 71134 11370
rect 71134 11319 71190 11328
rect 71148 11150 71176 11319
rect 71136 11144 71188 11150
rect 71136 11086 71188 11092
rect 71872 11076 71924 11082
rect 71872 11018 71924 11024
rect 71044 11008 71096 11014
rect 71136 11008 71188 11014
rect 71044 10950 71096 10956
rect 71134 10976 71136 10985
rect 71188 10976 71190 10985
rect 71056 10810 71084 10950
rect 71134 10911 71190 10920
rect 71260 10908 71568 10917
rect 71260 10906 71266 10908
rect 71322 10906 71346 10908
rect 71402 10906 71426 10908
rect 71482 10906 71506 10908
rect 71562 10906 71568 10908
rect 71322 10854 71324 10906
rect 71504 10854 71506 10906
rect 71260 10852 71266 10854
rect 71322 10852 71346 10854
rect 71402 10852 71426 10854
rect 71482 10852 71506 10854
rect 71562 10852 71568 10854
rect 71260 10843 71568 10852
rect 71044 10804 71096 10810
rect 71044 10746 71096 10752
rect 71780 10668 71832 10674
rect 71780 10610 71832 10616
rect 70688 10526 70808 10554
rect 70688 10062 70716 10526
rect 70950 10432 71006 10441
rect 70950 10367 71006 10376
rect 70964 10062 70992 10367
rect 71688 10260 71740 10266
rect 71688 10202 71740 10208
rect 71700 10130 71728 10202
rect 71688 10124 71740 10130
rect 71688 10066 71740 10072
rect 70676 10056 70728 10062
rect 70676 9998 70728 10004
rect 70952 10056 71004 10062
rect 70952 9998 71004 10004
rect 69756 7880 69808 7886
rect 69570 7848 69626 7857
rect 69756 7822 69808 7828
rect 70584 7880 70636 7886
rect 70584 7822 70636 7828
rect 69570 7783 69626 7792
rect 69584 7410 69612 7783
rect 69572 7404 69624 7410
rect 69572 7346 69624 7352
rect 68836 7278 68888 7284
rect 69478 7304 69534 7313
rect 68664 6866 68692 7278
rect 68848 7177 68876 7278
rect 69478 7239 69534 7248
rect 68834 7168 68890 7177
rect 68834 7103 68890 7112
rect 69846 7168 69902 7177
rect 69846 7103 69902 7112
rect 68744 6996 68796 7002
rect 68744 6938 68796 6944
rect 68756 6905 68784 6938
rect 69204 6928 69256 6934
rect 68742 6896 68798 6905
rect 68652 6860 68704 6866
rect 69204 6870 69256 6876
rect 68742 6831 68798 6840
rect 68652 6802 68704 6808
rect 68560 6452 68612 6458
rect 68560 6394 68612 6400
rect 69216 5914 69244 6870
rect 69296 6860 69348 6866
rect 69296 6802 69348 6808
rect 69308 5914 69336 6802
rect 69204 5908 69256 5914
rect 69204 5850 69256 5856
rect 69296 5908 69348 5914
rect 69296 5850 69348 5856
rect 69216 5817 69244 5850
rect 69202 5808 69258 5817
rect 69202 5743 69258 5752
rect 68192 5568 68244 5574
rect 68192 5510 68244 5516
rect 67732 5296 67784 5302
rect 67732 5238 67784 5244
rect 67364 4684 67416 4690
rect 67364 4626 67416 4632
rect 67640 4684 67692 4690
rect 67640 4626 67692 4632
rect 67744 4554 67772 5238
rect 69308 5166 69336 5850
rect 69860 5710 69888 7103
rect 70308 6792 70360 6798
rect 70308 6734 70360 6740
rect 70320 6322 70348 6734
rect 70400 6656 70452 6662
rect 70400 6598 70452 6604
rect 70308 6316 70360 6322
rect 70308 6258 70360 6264
rect 70124 5908 70176 5914
rect 70124 5850 70176 5856
rect 70136 5710 70164 5850
rect 69848 5704 69900 5710
rect 69848 5646 69900 5652
rect 70124 5704 70176 5710
rect 70124 5646 70176 5652
rect 69296 5160 69348 5166
rect 69296 5102 69348 5108
rect 69860 5030 69888 5646
rect 70320 5302 70348 6258
rect 70412 6118 70440 6598
rect 70400 6112 70452 6118
rect 70400 6054 70452 6060
rect 70596 5914 70624 7822
rect 70688 6662 70716 9998
rect 70860 9988 70912 9994
rect 70860 9930 70912 9936
rect 70872 9042 70900 9930
rect 70860 9036 70912 9042
rect 70860 8978 70912 8984
rect 70768 8900 70820 8906
rect 70768 8842 70820 8848
rect 70780 8430 70808 8842
rect 70768 8424 70820 8430
rect 70768 8366 70820 8372
rect 70676 6656 70728 6662
rect 70676 6598 70728 6604
rect 70768 6656 70820 6662
rect 70768 6598 70820 6604
rect 70780 6322 70808 6598
rect 70768 6316 70820 6322
rect 70768 6258 70820 6264
rect 70964 5914 70992 9998
rect 71596 9920 71648 9926
rect 71596 9862 71648 9868
rect 71260 9820 71568 9829
rect 71260 9818 71266 9820
rect 71322 9818 71346 9820
rect 71402 9818 71426 9820
rect 71482 9818 71506 9820
rect 71562 9818 71568 9820
rect 71322 9766 71324 9818
rect 71504 9766 71506 9818
rect 71260 9764 71266 9766
rect 71322 9764 71346 9766
rect 71402 9764 71426 9766
rect 71482 9764 71506 9766
rect 71562 9764 71568 9766
rect 71260 9755 71568 9764
rect 71412 9512 71464 9518
rect 71134 9480 71190 9489
rect 71412 9454 71464 9460
rect 71134 9415 71190 9424
rect 71148 9382 71176 9415
rect 71044 9376 71096 9382
rect 71044 9318 71096 9324
rect 71136 9376 71188 9382
rect 71136 9318 71188 9324
rect 71056 9178 71084 9318
rect 71044 9172 71096 9178
rect 71044 9114 71096 9120
rect 71424 9042 71452 9454
rect 71608 9178 71636 9862
rect 71596 9172 71648 9178
rect 71596 9114 71648 9120
rect 71412 9036 71464 9042
rect 71412 8978 71464 8984
rect 71700 8974 71728 10066
rect 71792 8974 71820 10610
rect 71884 9217 71912 11018
rect 72068 10010 72096 11698
rect 72252 11257 72280 11698
rect 72238 11248 72294 11257
rect 72238 11183 72294 11192
rect 72344 11150 72372 14214
rect 72606 14104 72662 14113
rect 72606 14039 72662 14048
rect 72620 13938 72648 14039
rect 73540 13938 73568 14350
rect 73988 14272 74040 14278
rect 73988 14214 74040 14220
rect 73712 14000 73764 14006
rect 73712 13942 73764 13948
rect 73802 13968 73858 13977
rect 72608 13932 72660 13938
rect 72608 13874 72660 13880
rect 73528 13932 73580 13938
rect 73528 13874 73580 13880
rect 72976 13864 73028 13870
rect 72976 13806 73028 13812
rect 72516 13524 72568 13530
rect 72516 13466 72568 13472
rect 72424 12912 72476 12918
rect 72424 12854 72476 12860
rect 72436 12617 72464 12854
rect 72528 12782 72556 13466
rect 72988 13326 73016 13806
rect 73068 13728 73120 13734
rect 73068 13670 73120 13676
rect 73080 13462 73108 13670
rect 73250 13560 73306 13569
rect 73250 13495 73306 13504
rect 73068 13456 73120 13462
rect 73068 13398 73120 13404
rect 72976 13320 73028 13326
rect 72976 13262 73028 13268
rect 72516 12776 72568 12782
rect 72516 12718 72568 12724
rect 72422 12608 72478 12617
rect 72422 12543 72478 12552
rect 72606 12336 72662 12345
rect 72606 12271 72662 12280
rect 72516 12164 72568 12170
rect 72516 12106 72568 12112
rect 72528 12073 72556 12106
rect 72514 12064 72570 12073
rect 72514 11999 72570 12008
rect 72620 11898 72648 12271
rect 72698 12200 72754 12209
rect 72698 12135 72700 12144
rect 72752 12135 72754 12144
rect 72700 12106 72752 12112
rect 72608 11892 72660 11898
rect 72608 11834 72660 11840
rect 72620 11762 72648 11834
rect 72608 11756 72660 11762
rect 72608 11698 72660 11704
rect 72792 11756 72844 11762
rect 72792 11698 72844 11704
rect 72332 11144 72384 11150
rect 72332 11086 72384 11092
rect 72240 10736 72292 10742
rect 72240 10678 72292 10684
rect 72252 10266 72280 10678
rect 72240 10260 72292 10266
rect 72240 10202 72292 10208
rect 72068 9982 72188 10010
rect 72160 9382 72188 9982
rect 72148 9376 72200 9382
rect 72148 9318 72200 9324
rect 72422 9344 72478 9353
rect 72422 9279 72478 9288
rect 71870 9208 71926 9217
rect 71870 9143 71926 9152
rect 71688 8968 71740 8974
rect 71688 8910 71740 8916
rect 71780 8968 71832 8974
rect 71780 8910 71832 8916
rect 71260 8732 71568 8741
rect 71260 8730 71266 8732
rect 71322 8730 71346 8732
rect 71402 8730 71426 8732
rect 71482 8730 71506 8732
rect 71562 8730 71568 8732
rect 71322 8678 71324 8730
rect 71504 8678 71506 8730
rect 71260 8676 71266 8678
rect 71322 8676 71346 8678
rect 71402 8676 71426 8678
rect 71482 8676 71506 8678
rect 71562 8676 71568 8678
rect 71260 8667 71568 8676
rect 71872 8016 71924 8022
rect 71502 7984 71558 7993
rect 71924 7964 72004 7970
rect 71872 7958 72004 7964
rect 71884 7942 72004 7958
rect 71502 7919 71558 7928
rect 71516 7886 71544 7919
rect 71504 7880 71556 7886
rect 71504 7822 71556 7828
rect 71872 7880 71924 7886
rect 71872 7822 71924 7828
rect 71260 7644 71568 7653
rect 71260 7642 71266 7644
rect 71322 7642 71346 7644
rect 71402 7642 71426 7644
rect 71482 7642 71506 7644
rect 71562 7642 71568 7644
rect 71322 7590 71324 7642
rect 71504 7590 71506 7642
rect 71260 7588 71266 7590
rect 71322 7588 71346 7590
rect 71402 7588 71426 7590
rect 71482 7588 71506 7590
rect 71562 7588 71568 7590
rect 71260 7579 71568 7588
rect 71884 7188 71912 7822
rect 71976 7732 72004 7942
rect 72436 7886 72464 9279
rect 72516 8832 72568 8838
rect 72516 8774 72568 8780
rect 72528 8430 72556 8774
rect 72516 8424 72568 8430
rect 72516 8366 72568 8372
rect 72424 7880 72476 7886
rect 72424 7822 72476 7828
rect 72424 7744 72476 7750
rect 71976 7704 72424 7732
rect 71976 7478 72004 7704
rect 72424 7686 72476 7692
rect 71964 7472 72016 7478
rect 71964 7414 72016 7420
rect 72424 7472 72476 7478
rect 72424 7414 72476 7420
rect 71976 7290 72004 7414
rect 71976 7262 72096 7290
rect 71964 7200 72016 7206
rect 71884 7177 71964 7188
rect 71870 7168 71964 7177
rect 71926 7160 71964 7168
rect 71964 7142 72016 7148
rect 71870 7103 71926 7112
rect 71870 6896 71926 6905
rect 71870 6831 71926 6840
rect 71136 6792 71188 6798
rect 71136 6734 71188 6740
rect 70584 5908 70636 5914
rect 70584 5850 70636 5856
rect 70952 5908 71004 5914
rect 70952 5850 71004 5856
rect 70308 5296 70360 5302
rect 70308 5238 70360 5244
rect 69848 5024 69900 5030
rect 69848 4966 69900 4972
rect 67732 4548 67784 4554
rect 67732 4490 67784 4496
rect 67744 3942 67772 4490
rect 71148 4162 71176 6734
rect 71884 6730 71912 6831
rect 72068 6730 72096 7262
rect 71872 6724 71924 6730
rect 71872 6666 71924 6672
rect 72056 6724 72108 6730
rect 72056 6666 72108 6672
rect 72068 6610 72096 6666
rect 72436 6662 72464 7414
rect 72620 7313 72648 11698
rect 72700 11552 72752 11558
rect 72700 11494 72752 11500
rect 72712 11354 72740 11494
rect 72700 11348 72752 11354
rect 72700 11290 72752 11296
rect 72804 11218 72832 11698
rect 72884 11552 72936 11558
rect 72884 11494 72936 11500
rect 72792 11212 72844 11218
rect 72792 11154 72844 11160
rect 72896 10169 72924 11494
rect 73080 11150 73108 13398
rect 73264 13190 73292 13495
rect 73252 13184 73304 13190
rect 73252 13126 73304 13132
rect 73540 12850 73568 13874
rect 73724 13802 73752 13942
rect 73802 13903 73804 13912
rect 73856 13903 73858 13912
rect 73804 13874 73856 13880
rect 73896 13864 73948 13870
rect 73896 13806 73948 13812
rect 73712 13796 73764 13802
rect 73712 13738 73764 13744
rect 73528 12844 73580 12850
rect 73528 12786 73580 12792
rect 73540 12730 73568 12786
rect 73540 12702 73660 12730
rect 73908 12714 73936 13806
rect 74000 13394 74028 14214
rect 74276 13802 74304 14962
rect 74552 14822 74580 15098
rect 74644 14822 74672 15574
rect 75828 15020 75880 15026
rect 75828 14962 75880 14968
rect 75274 14920 75330 14929
rect 75274 14855 75276 14864
rect 75328 14855 75330 14864
rect 75276 14826 75328 14832
rect 74540 14816 74592 14822
rect 74540 14758 74592 14764
rect 74632 14816 74684 14822
rect 74632 14758 74684 14764
rect 74356 13932 74408 13938
rect 74356 13874 74408 13880
rect 74264 13796 74316 13802
rect 74264 13738 74316 13744
rect 73988 13388 74040 13394
rect 73988 13330 74040 13336
rect 73528 12640 73580 12646
rect 73528 12582 73580 12588
rect 73540 12306 73568 12582
rect 73528 12300 73580 12306
rect 73528 12242 73580 12248
rect 73632 12186 73660 12702
rect 73896 12708 73948 12714
rect 73896 12650 73948 12656
rect 73988 12640 74040 12646
rect 73988 12582 74040 12588
rect 73540 12158 73660 12186
rect 73896 12164 73948 12170
rect 73540 11762 73568 12158
rect 73896 12106 73948 12112
rect 73618 12064 73674 12073
rect 73618 11999 73674 12008
rect 73632 11898 73660 11999
rect 73620 11892 73672 11898
rect 73620 11834 73672 11840
rect 73528 11756 73580 11762
rect 73528 11698 73580 11704
rect 73068 11144 73120 11150
rect 73068 11086 73120 11092
rect 73540 10742 73568 11698
rect 73804 11280 73856 11286
rect 73908 11268 73936 12106
rect 74000 11830 74028 12582
rect 73988 11824 74040 11830
rect 73988 11766 74040 11772
rect 74172 11824 74224 11830
rect 74172 11766 74224 11772
rect 74080 11688 74132 11694
rect 74080 11630 74132 11636
rect 73988 11552 74040 11558
rect 73988 11494 74040 11500
rect 73856 11240 73936 11268
rect 73804 11222 73856 11228
rect 74000 11150 74028 11494
rect 74092 11354 74120 11630
rect 74080 11348 74132 11354
rect 74080 11290 74132 11296
rect 74184 11286 74212 11766
rect 74172 11280 74224 11286
rect 74172 11222 74224 11228
rect 73620 11144 73672 11150
rect 73620 11086 73672 11092
rect 73988 11144 74040 11150
rect 73988 11086 74040 11092
rect 73528 10736 73580 10742
rect 73528 10678 73580 10684
rect 73632 10554 73660 11086
rect 74080 10668 74132 10674
rect 74184 10656 74212 11222
rect 74276 11132 74304 13738
rect 74368 11286 74396 13874
rect 74644 12345 74672 14758
rect 74816 14408 74868 14414
rect 74816 14350 74868 14356
rect 74828 14074 74856 14350
rect 75092 14272 75144 14278
rect 75092 14214 75144 14220
rect 75184 14272 75236 14278
rect 75184 14214 75236 14220
rect 74816 14068 74868 14074
rect 74816 14010 74868 14016
rect 74630 12336 74686 12345
rect 74828 12306 74856 14010
rect 75000 12640 75052 12646
rect 75000 12582 75052 12588
rect 75012 12442 75040 12582
rect 75000 12436 75052 12442
rect 75000 12378 75052 12384
rect 74630 12271 74686 12280
rect 74816 12300 74868 12306
rect 74816 12242 74868 12248
rect 75012 12186 75040 12378
rect 74552 12170 75040 12186
rect 74540 12164 75040 12170
rect 74592 12158 75040 12164
rect 74540 12106 74592 12112
rect 74448 11348 74500 11354
rect 74448 11290 74500 11296
rect 74356 11280 74408 11286
rect 74356 11222 74408 11228
rect 74356 11144 74408 11150
rect 74276 11104 74356 11132
rect 74356 11086 74408 11092
rect 74132 10628 74212 10656
rect 74080 10610 74132 10616
rect 73540 10538 73660 10554
rect 73528 10532 73660 10538
rect 73580 10526 73660 10532
rect 73528 10474 73580 10480
rect 72976 10464 73028 10470
rect 72976 10406 73028 10412
rect 72882 10160 72938 10169
rect 72882 10095 72938 10104
rect 72988 10062 73016 10406
rect 72976 10056 73028 10062
rect 72976 9998 73028 10004
rect 73160 10056 73212 10062
rect 73160 9998 73212 10004
rect 73172 9722 73200 9998
rect 73436 9988 73488 9994
rect 73436 9930 73488 9936
rect 73160 9716 73212 9722
rect 73160 9658 73212 9664
rect 73448 9654 73476 9930
rect 73632 9722 73660 10526
rect 73620 9716 73672 9722
rect 74092 9674 74120 10610
rect 74460 10606 74488 11290
rect 74448 10600 74500 10606
rect 74448 10542 74500 10548
rect 74172 10464 74224 10470
rect 74172 10406 74224 10412
rect 74184 10266 74212 10406
rect 74172 10260 74224 10266
rect 74172 10202 74224 10208
rect 73620 9658 73672 9664
rect 73436 9648 73488 9654
rect 73436 9590 73488 9596
rect 74000 9646 74120 9674
rect 74184 9654 74212 10202
rect 74172 9648 74224 9654
rect 72700 9580 72752 9586
rect 72700 9522 72752 9528
rect 73620 9580 73672 9586
rect 73620 9522 73672 9528
rect 72712 9042 72740 9522
rect 72700 9036 72752 9042
rect 72700 8978 72752 8984
rect 73068 8900 73120 8906
rect 73068 8842 73120 8848
rect 73080 8430 73108 8842
rect 73632 8498 73660 9522
rect 74000 9489 74028 9646
rect 74172 9590 74224 9596
rect 73986 9480 74042 9489
rect 73986 9415 74042 9424
rect 73804 8968 73856 8974
rect 73804 8910 73856 8916
rect 74000 8922 74028 9415
rect 74080 9376 74132 9382
rect 74080 9318 74132 9324
rect 74092 9042 74120 9318
rect 74552 9042 74580 12106
rect 75104 12102 75132 14214
rect 75196 13938 75224 14214
rect 75184 13932 75236 13938
rect 75184 13874 75236 13880
rect 75288 12850 75316 14826
rect 75840 14618 75868 14962
rect 75920 14816 75972 14822
rect 75920 14758 75972 14764
rect 75828 14612 75880 14618
rect 75828 14554 75880 14560
rect 75932 14278 75960 14758
rect 75920 14272 75972 14278
rect 75920 14214 75972 14220
rect 75734 13696 75790 13705
rect 75734 13631 75790 13640
rect 75748 12918 75776 13631
rect 76116 13530 76144 17138
rect 83372 17128 83424 17134
rect 83372 17070 83424 17076
rect 82979 16892 83287 16901
rect 82979 16890 82985 16892
rect 83041 16890 83065 16892
rect 83121 16890 83145 16892
rect 83201 16890 83225 16892
rect 83281 16890 83287 16892
rect 83041 16838 83043 16890
rect 83223 16838 83225 16890
rect 82979 16836 82985 16838
rect 83041 16836 83065 16838
rect 83121 16836 83145 16838
rect 83201 16836 83225 16838
rect 83281 16836 83287 16838
rect 82979 16827 83287 16836
rect 83384 16726 83412 17070
rect 83372 16720 83424 16726
rect 83372 16662 83424 16668
rect 77300 16652 77352 16658
rect 77300 16594 77352 16600
rect 77208 16040 77260 16046
rect 77208 15982 77260 15988
rect 76748 15972 76800 15978
rect 76748 15914 76800 15920
rect 77116 15972 77168 15978
rect 77116 15914 77168 15920
rect 76564 15904 76616 15910
rect 76564 15846 76616 15852
rect 76472 15360 76524 15366
rect 76472 15302 76524 15308
rect 76484 15094 76512 15302
rect 76472 15088 76524 15094
rect 76472 15030 76524 15036
rect 76196 14272 76248 14278
rect 76196 14214 76248 14220
rect 76104 13524 76156 13530
rect 76104 13466 76156 13472
rect 75736 12912 75788 12918
rect 75736 12854 75788 12860
rect 75276 12844 75328 12850
rect 75276 12786 75328 12792
rect 75828 12708 75880 12714
rect 75828 12650 75880 12656
rect 75184 12640 75236 12646
rect 75184 12582 75236 12588
rect 75196 12481 75224 12582
rect 75182 12472 75238 12481
rect 75182 12407 75238 12416
rect 75368 12300 75420 12306
rect 75368 12242 75420 12248
rect 75644 12300 75696 12306
rect 75644 12242 75696 12248
rect 75092 12096 75144 12102
rect 75092 12038 75144 12044
rect 75380 11898 75408 12242
rect 75552 12164 75604 12170
rect 75552 12106 75604 12112
rect 75368 11892 75420 11898
rect 75368 11834 75420 11840
rect 75564 11762 75592 12106
rect 75656 12102 75684 12242
rect 75644 12096 75696 12102
rect 75644 12038 75696 12044
rect 75368 11756 75420 11762
rect 75552 11756 75604 11762
rect 75368 11698 75420 11704
rect 75472 11716 75552 11744
rect 74724 11688 74776 11694
rect 74722 11656 74724 11665
rect 74776 11656 74778 11665
rect 74722 11591 74778 11600
rect 75276 11348 75328 11354
rect 75276 11290 75328 11296
rect 75182 11248 75238 11257
rect 75182 11183 75238 11192
rect 75196 11082 75224 11183
rect 75288 11150 75316 11290
rect 75380 11218 75408 11698
rect 75472 11393 75500 11716
rect 75552 11698 75604 11704
rect 75458 11384 75514 11393
rect 75458 11319 75514 11328
rect 75368 11212 75420 11218
rect 75368 11154 75420 11160
rect 75276 11144 75328 11150
rect 75276 11086 75328 11092
rect 75656 11082 75684 12038
rect 75736 11824 75788 11830
rect 75736 11766 75788 11772
rect 75748 11218 75776 11766
rect 75840 11694 75868 12650
rect 75920 12164 75972 12170
rect 75920 12106 75972 12112
rect 75932 11762 75960 12106
rect 76208 12102 76236 14214
rect 76576 13326 76604 15846
rect 76564 13320 76616 13326
rect 76564 13262 76616 13268
rect 76380 12232 76432 12238
rect 76378 12200 76380 12209
rect 76432 12200 76434 12209
rect 76378 12135 76434 12144
rect 76196 12096 76248 12102
rect 76196 12038 76248 12044
rect 76194 11928 76250 11937
rect 76194 11863 76250 11872
rect 75920 11756 75972 11762
rect 75920 11698 75972 11704
rect 75828 11688 75880 11694
rect 75828 11630 75880 11636
rect 75736 11212 75788 11218
rect 75736 11154 75788 11160
rect 75184 11076 75236 11082
rect 75184 11018 75236 11024
rect 75644 11076 75696 11082
rect 75644 11018 75696 11024
rect 75932 10266 75960 11698
rect 76208 11694 76236 11863
rect 76196 11688 76248 11694
rect 76196 11630 76248 11636
rect 76208 11558 76236 11630
rect 76196 11552 76248 11558
rect 76196 11494 76248 11500
rect 76104 11144 76156 11150
rect 76208 11132 76236 11494
rect 76156 11104 76236 11132
rect 76104 11086 76156 11092
rect 76012 10736 76064 10742
rect 76012 10678 76064 10684
rect 75920 10260 75972 10266
rect 75920 10202 75972 10208
rect 75920 10056 75972 10062
rect 75920 9998 75972 10004
rect 75276 9988 75328 9994
rect 75276 9930 75328 9936
rect 74816 9920 74868 9926
rect 74816 9862 74868 9868
rect 74828 9586 74856 9862
rect 75288 9654 75316 9930
rect 75932 9722 75960 9998
rect 75920 9716 75972 9722
rect 75920 9658 75972 9664
rect 76024 9654 76052 10678
rect 76102 10296 76158 10305
rect 76102 10231 76158 10240
rect 76116 10062 76144 10231
rect 76104 10056 76156 10062
rect 76104 9998 76156 10004
rect 75276 9648 75328 9654
rect 75276 9590 75328 9596
rect 76012 9648 76064 9654
rect 76012 9590 76064 9596
rect 74816 9580 74868 9586
rect 74816 9522 74868 9528
rect 75460 9580 75512 9586
rect 75460 9522 75512 9528
rect 74828 9178 74856 9522
rect 75472 9489 75500 9522
rect 75458 9480 75514 9489
rect 75458 9415 75514 9424
rect 75920 9444 75972 9450
rect 75920 9386 75972 9392
rect 74816 9172 74868 9178
rect 74816 9114 74868 9120
rect 74080 9036 74132 9042
rect 74080 8978 74132 8984
rect 74540 9036 74592 9042
rect 74540 8978 74592 8984
rect 75276 9036 75328 9042
rect 75276 8978 75328 8984
rect 73816 8634 73844 8910
rect 74000 8894 74120 8922
rect 73804 8628 73856 8634
rect 73804 8570 73856 8576
rect 73620 8492 73672 8498
rect 73620 8434 73672 8440
rect 72792 8424 72844 8430
rect 72792 8366 72844 8372
rect 72976 8424 73028 8430
rect 72976 8366 73028 8372
rect 73068 8424 73120 8430
rect 73068 8366 73120 8372
rect 72606 7304 72662 7313
rect 72606 7239 72662 7248
rect 72804 6769 72832 8366
rect 72988 8022 73016 8366
rect 72976 8016 73028 8022
rect 72976 7958 73028 7964
rect 72988 7002 73016 7958
rect 72976 6996 73028 7002
rect 72976 6938 73028 6944
rect 72790 6760 72846 6769
rect 73080 6746 73108 8366
rect 73160 8356 73212 8362
rect 73160 8298 73212 8304
rect 73172 8090 73200 8298
rect 73632 8294 73660 8434
rect 73620 8288 73672 8294
rect 73620 8230 73672 8236
rect 73160 8084 73212 8090
rect 73160 8026 73212 8032
rect 73172 7886 73200 8026
rect 73160 7880 73212 7886
rect 73212 7840 73292 7868
rect 73160 7822 73212 7828
rect 73080 6730 73200 6746
rect 73080 6724 73212 6730
rect 73080 6718 73160 6724
rect 72790 6695 72846 6704
rect 73160 6666 73212 6672
rect 71884 6582 72096 6610
rect 72424 6656 72476 6662
rect 73264 6610 73292 7840
rect 73528 7336 73580 7342
rect 73526 7304 73528 7313
rect 73580 7304 73582 7313
rect 73526 7239 73582 7248
rect 72424 6598 72476 6604
rect 73172 6582 73292 6610
rect 71260 6556 71568 6565
rect 71260 6554 71266 6556
rect 71322 6554 71346 6556
rect 71402 6554 71426 6556
rect 71482 6554 71506 6556
rect 71562 6554 71568 6556
rect 71322 6502 71324 6554
rect 71504 6502 71506 6554
rect 71260 6500 71266 6502
rect 71322 6500 71346 6502
rect 71402 6500 71426 6502
rect 71482 6500 71506 6502
rect 71562 6500 71568 6502
rect 71260 6491 71568 6500
rect 71504 6452 71556 6458
rect 71504 6394 71556 6400
rect 71412 6316 71464 6322
rect 71412 6258 71464 6264
rect 71424 5914 71452 6258
rect 71516 6254 71544 6394
rect 71688 6316 71740 6322
rect 71688 6258 71740 6264
rect 71504 6248 71556 6254
rect 71504 6190 71556 6196
rect 71412 5908 71464 5914
rect 71412 5850 71464 5856
rect 71424 5710 71452 5850
rect 71412 5704 71464 5710
rect 71412 5646 71464 5652
rect 71260 5468 71568 5477
rect 71260 5466 71266 5468
rect 71322 5466 71346 5468
rect 71402 5466 71426 5468
rect 71482 5466 71506 5468
rect 71562 5466 71568 5468
rect 71322 5414 71324 5466
rect 71504 5414 71506 5466
rect 71260 5412 71266 5414
rect 71322 5412 71346 5414
rect 71402 5412 71426 5414
rect 71482 5412 71506 5414
rect 71562 5412 71568 5414
rect 71260 5403 71568 5412
rect 71700 4826 71728 6258
rect 71780 5704 71832 5710
rect 71780 5646 71832 5652
rect 71792 5545 71820 5646
rect 71778 5536 71834 5545
rect 71778 5471 71834 5480
rect 71792 5234 71820 5471
rect 71884 5302 71912 6582
rect 71962 6488 72018 6497
rect 71962 6423 72018 6432
rect 72056 6452 72108 6458
rect 71976 5778 72004 6423
rect 72056 6394 72108 6400
rect 71964 5772 72016 5778
rect 71964 5714 72016 5720
rect 72068 5302 72096 6394
rect 72148 6112 72200 6118
rect 72148 6054 72200 6060
rect 71872 5296 71924 5302
rect 71872 5238 71924 5244
rect 72056 5296 72108 5302
rect 72056 5238 72108 5244
rect 71780 5228 71832 5234
rect 71780 5170 71832 5176
rect 71792 5098 71820 5170
rect 71780 5092 71832 5098
rect 71780 5034 71832 5040
rect 71688 4820 71740 4826
rect 71688 4762 71740 4768
rect 71596 4480 71648 4486
rect 71596 4422 71648 4428
rect 71260 4380 71568 4389
rect 71260 4378 71266 4380
rect 71322 4378 71346 4380
rect 71402 4378 71426 4380
rect 71482 4378 71506 4380
rect 71562 4378 71568 4380
rect 71322 4326 71324 4378
rect 71504 4326 71506 4378
rect 71260 4324 71266 4326
rect 71322 4324 71346 4326
rect 71402 4324 71426 4326
rect 71482 4324 71506 4326
rect 71562 4324 71568 4326
rect 71260 4315 71568 4324
rect 71608 4214 71636 4422
rect 71884 4282 71912 5238
rect 72160 5166 72188 6054
rect 73172 5778 73200 6582
rect 73528 6316 73580 6322
rect 73528 6258 73580 6264
rect 73540 6118 73568 6258
rect 73528 6112 73580 6118
rect 73528 6054 73580 6060
rect 73988 6112 74040 6118
rect 73988 6054 74040 6060
rect 73160 5772 73212 5778
rect 73160 5714 73212 5720
rect 73252 5772 73304 5778
rect 73252 5714 73304 5720
rect 72148 5160 72200 5166
rect 72148 5102 72200 5108
rect 73264 4826 73292 5714
rect 73344 5704 73396 5710
rect 73344 5646 73396 5652
rect 73252 4820 73304 4826
rect 73252 4762 73304 4768
rect 72056 4684 72108 4690
rect 72056 4626 72108 4632
rect 71872 4276 71924 4282
rect 71872 4218 71924 4224
rect 71596 4208 71648 4214
rect 71148 4146 71268 4162
rect 71596 4150 71648 4156
rect 71148 4140 71280 4146
rect 71148 4134 71228 4140
rect 71228 4082 71280 4088
rect 68652 4072 68704 4078
rect 68652 4014 68704 4020
rect 67732 3936 67784 3942
rect 67732 3878 67784 3884
rect 68664 3738 68692 4014
rect 67180 3732 67232 3738
rect 67180 3674 67232 3680
rect 68652 3732 68704 3738
rect 68652 3674 68704 3680
rect 65892 3460 65944 3466
rect 65892 3402 65944 3408
rect 64788 3188 64840 3194
rect 64788 3130 64840 3136
rect 64972 2984 65024 2990
rect 64972 2926 65024 2932
rect 64984 2650 65012 2926
rect 64328 2644 64380 2650
rect 64328 2586 64380 2592
rect 64972 2644 65024 2650
rect 64972 2586 65024 2592
rect 65904 2582 65932 3402
rect 71240 3398 71268 4082
rect 72068 3670 72096 4626
rect 73252 4616 73304 4622
rect 73356 4604 73384 5646
rect 74000 5234 74028 6054
rect 74092 5953 74120 8894
rect 74356 8900 74408 8906
rect 74356 8842 74408 8848
rect 74368 8498 74396 8842
rect 74356 8492 74408 8498
rect 74356 8434 74408 8440
rect 74356 8288 74408 8294
rect 74356 8230 74408 8236
rect 74368 7546 74396 8230
rect 74552 7993 74580 8978
rect 75184 8968 75236 8974
rect 75184 8910 75236 8916
rect 75196 8634 75224 8910
rect 75184 8628 75236 8634
rect 75184 8570 75236 8576
rect 75288 8498 75316 8978
rect 75552 8832 75604 8838
rect 75552 8774 75604 8780
rect 75736 8832 75788 8838
rect 75736 8774 75788 8780
rect 75564 8566 75592 8774
rect 75552 8560 75604 8566
rect 75552 8502 75604 8508
rect 75748 8498 75776 8774
rect 75276 8492 75328 8498
rect 75276 8434 75328 8440
rect 75736 8492 75788 8498
rect 75736 8434 75788 8440
rect 74724 8424 74776 8430
rect 74724 8366 74776 8372
rect 74816 8424 74868 8430
rect 74816 8366 74868 8372
rect 74538 7984 74594 7993
rect 74736 7954 74764 8366
rect 74538 7919 74594 7928
rect 74724 7948 74776 7954
rect 74724 7890 74776 7896
rect 74632 7744 74684 7750
rect 74632 7686 74684 7692
rect 74356 7540 74408 7546
rect 74356 7482 74408 7488
rect 74644 7342 74672 7686
rect 74828 7546 74856 8366
rect 74908 7880 74960 7886
rect 74908 7822 74960 7828
rect 74816 7540 74868 7546
rect 74816 7482 74868 7488
rect 74632 7336 74684 7342
rect 74632 7278 74684 7284
rect 74540 7268 74592 7274
rect 74540 7210 74592 7216
rect 74356 6860 74408 6866
rect 74356 6802 74408 6808
rect 74368 6322 74396 6802
rect 74552 6798 74580 7210
rect 74540 6792 74592 6798
rect 74540 6734 74592 6740
rect 74632 6656 74684 6662
rect 74632 6598 74684 6604
rect 74644 6390 74672 6598
rect 74632 6384 74684 6390
rect 74632 6326 74684 6332
rect 74356 6316 74408 6322
rect 74356 6258 74408 6264
rect 74078 5944 74134 5953
rect 74368 5914 74396 6258
rect 74078 5879 74134 5888
rect 74356 5908 74408 5914
rect 74092 5574 74120 5879
rect 74356 5850 74408 5856
rect 74080 5568 74132 5574
rect 74080 5510 74132 5516
rect 73804 5228 73856 5234
rect 73804 5170 73856 5176
rect 73988 5228 74040 5234
rect 73988 5170 74040 5176
rect 73528 5092 73580 5098
rect 73528 5034 73580 5040
rect 73540 4622 73568 5034
rect 73620 4820 73672 4826
rect 73620 4762 73672 4768
rect 73304 4576 73384 4604
rect 73436 4616 73488 4622
rect 73252 4558 73304 4564
rect 73436 4558 73488 4564
rect 73528 4616 73580 4622
rect 73528 4558 73580 4564
rect 73448 4214 73476 4558
rect 73540 4486 73568 4558
rect 73528 4480 73580 4486
rect 73528 4422 73580 4428
rect 73436 4208 73488 4214
rect 73436 4150 73488 4156
rect 73540 4078 73568 4422
rect 73528 4072 73580 4078
rect 73528 4014 73580 4020
rect 73632 4026 73660 4762
rect 73816 4758 73844 5170
rect 73804 4752 73856 4758
rect 73804 4694 73856 4700
rect 73712 4548 73764 4554
rect 73712 4490 73764 4496
rect 73724 4146 73752 4490
rect 73712 4140 73764 4146
rect 73712 4082 73764 4088
rect 73632 4010 73752 4026
rect 73632 4004 73764 4010
rect 73632 3998 73712 4004
rect 73712 3946 73764 3952
rect 73620 3936 73672 3942
rect 73620 3878 73672 3884
rect 73632 3670 73660 3878
rect 72056 3664 72108 3670
rect 72056 3606 72108 3612
rect 73620 3664 73672 3670
rect 73620 3606 73672 3612
rect 73724 3466 73752 3946
rect 73816 3534 73844 4694
rect 74000 4282 74028 5170
rect 74264 5024 74316 5030
rect 74264 4966 74316 4972
rect 74276 4690 74304 4966
rect 74264 4684 74316 4690
rect 74264 4626 74316 4632
rect 74172 4548 74224 4554
rect 74172 4490 74224 4496
rect 73988 4276 74040 4282
rect 73988 4218 74040 4224
rect 73804 3528 73856 3534
rect 73804 3470 73856 3476
rect 73712 3460 73764 3466
rect 73712 3402 73764 3408
rect 74000 3398 74028 4218
rect 74184 4214 74212 4490
rect 74172 4208 74224 4214
rect 74172 4150 74224 4156
rect 74368 4078 74396 5850
rect 74448 5228 74500 5234
rect 74448 5170 74500 5176
rect 74460 4758 74488 5170
rect 74448 4752 74500 4758
rect 74448 4694 74500 4700
rect 74632 4684 74684 4690
rect 74632 4626 74684 4632
rect 74356 4072 74408 4078
rect 74356 4014 74408 4020
rect 74448 4072 74500 4078
rect 74448 4014 74500 4020
rect 74460 3602 74488 4014
rect 74448 3596 74500 3602
rect 74448 3538 74500 3544
rect 68376 3392 68428 3398
rect 68376 3334 68428 3340
rect 71228 3392 71280 3398
rect 71228 3334 71280 3340
rect 72884 3392 72936 3398
rect 72884 3334 72936 3340
rect 73988 3392 74040 3398
rect 73988 3334 74040 3340
rect 65892 2576 65944 2582
rect 65892 2518 65944 2524
rect 68388 2446 68416 3334
rect 71260 3292 71568 3301
rect 71260 3290 71266 3292
rect 71322 3290 71346 3292
rect 71402 3290 71426 3292
rect 71482 3290 71506 3292
rect 71562 3290 71568 3292
rect 71322 3238 71324 3290
rect 71504 3238 71506 3290
rect 71260 3236 71266 3238
rect 71322 3236 71346 3238
rect 71402 3236 71426 3238
rect 71482 3236 71506 3238
rect 71562 3236 71568 3238
rect 71260 3227 71568 3236
rect 72896 3126 72924 3334
rect 74644 3126 74672 4626
rect 72884 3120 72936 3126
rect 72884 3062 72936 3068
rect 74632 3120 74684 3126
rect 74632 3062 74684 3068
rect 74828 2446 74856 7482
rect 74920 5914 74948 7822
rect 75932 7041 75960 9386
rect 76196 9036 76248 9042
rect 76196 8978 76248 8984
rect 76104 8424 76156 8430
rect 76104 8366 76156 8372
rect 76116 7546 76144 8366
rect 76104 7540 76156 7546
rect 76104 7482 76156 7488
rect 76012 7404 76064 7410
rect 76012 7346 76064 7352
rect 75918 7032 75974 7041
rect 75918 6967 75974 6976
rect 75184 6792 75236 6798
rect 75184 6734 75236 6740
rect 75460 6792 75512 6798
rect 75460 6734 75512 6740
rect 74998 6624 75054 6633
rect 74998 6559 75054 6568
rect 75012 6322 75040 6559
rect 75000 6316 75052 6322
rect 75000 6258 75052 6264
rect 74908 5908 74960 5914
rect 74908 5850 74960 5856
rect 74920 5710 74948 5850
rect 75012 5846 75040 6258
rect 75000 5840 75052 5846
rect 75000 5782 75052 5788
rect 74908 5704 74960 5710
rect 74908 5646 74960 5652
rect 75196 5642 75224 6734
rect 75472 6458 75500 6734
rect 75644 6724 75696 6730
rect 75644 6666 75696 6672
rect 75368 6452 75420 6458
rect 75368 6394 75420 6400
rect 75460 6452 75512 6458
rect 75460 6394 75512 6400
rect 75276 5704 75328 5710
rect 75276 5646 75328 5652
rect 75184 5636 75236 5642
rect 75184 5578 75236 5584
rect 75196 4078 75224 5578
rect 75288 5574 75316 5646
rect 75276 5568 75328 5574
rect 75274 5536 75276 5545
rect 75328 5536 75330 5545
rect 75274 5471 75330 5480
rect 75288 5234 75316 5471
rect 75276 5228 75328 5234
rect 75276 5170 75328 5176
rect 75380 5080 75408 6394
rect 75460 6248 75512 6254
rect 75656 6236 75684 6666
rect 76024 6390 76052 7346
rect 76012 6384 76064 6390
rect 76012 6326 76064 6332
rect 75512 6208 75684 6236
rect 75460 6190 75512 6196
rect 75472 6118 75500 6149
rect 75460 6112 75512 6118
rect 75458 6080 75460 6089
rect 75512 6080 75514 6089
rect 75458 6015 75514 6024
rect 75472 5642 75500 6015
rect 76024 5846 76052 6326
rect 76012 5840 76064 5846
rect 76012 5782 76064 5788
rect 75552 5704 75604 5710
rect 75552 5646 75604 5652
rect 75460 5636 75512 5642
rect 75460 5578 75512 5584
rect 75564 5273 75592 5646
rect 75828 5636 75880 5642
rect 75828 5578 75880 5584
rect 75920 5636 75972 5642
rect 75920 5578 75972 5584
rect 75550 5264 75606 5273
rect 75840 5234 75868 5578
rect 75550 5199 75606 5208
rect 75828 5228 75880 5234
rect 75828 5170 75880 5176
rect 75460 5092 75512 5098
rect 75380 5052 75460 5080
rect 75460 5034 75512 5040
rect 75840 5030 75868 5170
rect 75932 5166 75960 5578
rect 75920 5160 75972 5166
rect 75920 5102 75972 5108
rect 75828 5024 75880 5030
rect 75828 4966 75880 4972
rect 75840 4264 75868 4966
rect 76208 4826 76236 8978
rect 76576 8974 76604 13262
rect 76760 12434 76788 15914
rect 77128 14618 77156 15914
rect 77116 14612 77168 14618
rect 77116 14554 77168 14560
rect 76932 14340 76984 14346
rect 76932 14282 76984 14288
rect 76944 13938 76972 14282
rect 76932 13932 76984 13938
rect 76932 13874 76984 13880
rect 77220 13734 77248 15982
rect 77312 15094 77340 16594
rect 77852 16244 77904 16250
rect 77852 16186 77904 16192
rect 77484 15904 77536 15910
rect 77484 15846 77536 15852
rect 77392 15360 77444 15366
rect 77392 15302 77444 15308
rect 77300 15088 77352 15094
rect 77300 15030 77352 15036
rect 76840 13728 76892 13734
rect 76840 13670 76892 13676
rect 77208 13728 77260 13734
rect 77208 13670 77260 13676
rect 76852 13258 76880 13670
rect 77022 13424 77078 13433
rect 77022 13359 77078 13368
rect 77036 13326 77064 13359
rect 77024 13320 77076 13326
rect 77024 13262 77076 13268
rect 76840 13252 76892 13258
rect 76840 13194 76892 13200
rect 76932 13252 76984 13258
rect 76932 13194 76984 13200
rect 76944 12986 76972 13194
rect 77022 13152 77078 13161
rect 77022 13087 77078 13096
rect 77036 12986 77064 13087
rect 77114 13016 77170 13025
rect 76932 12980 76984 12986
rect 76932 12922 76984 12928
rect 77024 12980 77076 12986
rect 77114 12951 77170 12960
rect 77024 12922 77076 12928
rect 77128 12850 77156 12951
rect 77220 12918 77248 13670
rect 77208 12912 77260 12918
rect 77208 12854 77260 12860
rect 77116 12844 77168 12850
rect 77116 12786 77168 12792
rect 77220 12434 77248 12854
rect 76760 12406 76880 12434
rect 76656 12232 76708 12238
rect 76656 12174 76708 12180
rect 76668 11354 76696 12174
rect 76748 11756 76800 11762
rect 76748 11698 76800 11704
rect 76656 11348 76708 11354
rect 76656 11290 76708 11296
rect 76760 10674 76788 11698
rect 76852 11218 76880 12406
rect 77036 12406 77248 12434
rect 77036 12238 77064 12406
rect 77116 12300 77168 12306
rect 77116 12242 77168 12248
rect 77024 12232 77076 12238
rect 77024 12174 77076 12180
rect 77128 11898 77156 12242
rect 77116 11892 77168 11898
rect 77116 11834 77168 11840
rect 77116 11756 77168 11762
rect 77116 11698 77168 11704
rect 76932 11620 76984 11626
rect 76932 11562 76984 11568
rect 76944 11354 76972 11562
rect 77128 11354 77156 11698
rect 77208 11552 77260 11558
rect 77208 11494 77260 11500
rect 76932 11348 76984 11354
rect 76932 11290 76984 11296
rect 77116 11348 77168 11354
rect 77116 11290 77168 11296
rect 77220 11257 77248 11494
rect 77206 11248 77262 11257
rect 76840 11212 76892 11218
rect 77206 11183 77262 11192
rect 76840 11154 76892 11160
rect 76748 10668 76800 10674
rect 76748 10610 76800 10616
rect 76852 9722 76880 11154
rect 77220 11150 77248 11183
rect 77208 11144 77260 11150
rect 77208 11086 77260 11092
rect 77116 11008 77168 11014
rect 77116 10950 77168 10956
rect 77128 10674 77156 10950
rect 77116 10668 77168 10674
rect 77116 10610 77168 10616
rect 76932 10464 76984 10470
rect 76932 10406 76984 10412
rect 76944 9722 76972 10406
rect 77128 10266 77156 10610
rect 77116 10260 77168 10266
rect 77116 10202 77168 10208
rect 76840 9716 76892 9722
rect 76840 9658 76892 9664
rect 76932 9716 76984 9722
rect 76932 9658 76984 9664
rect 76656 9104 76708 9110
rect 76656 9046 76708 9052
rect 76564 8968 76616 8974
rect 76564 8910 76616 8916
rect 76472 8560 76524 8566
rect 76472 8502 76524 8508
rect 76380 8424 76432 8430
rect 76380 8366 76432 8372
rect 76288 7948 76340 7954
rect 76288 7890 76340 7896
rect 76300 7410 76328 7890
rect 76392 7478 76420 8366
rect 76484 8090 76512 8502
rect 76472 8084 76524 8090
rect 76472 8026 76524 8032
rect 76484 7818 76512 8026
rect 76472 7812 76524 7818
rect 76472 7754 76524 7760
rect 76380 7472 76432 7478
rect 76380 7414 76432 7420
rect 76288 7404 76340 7410
rect 76288 7346 76340 7352
rect 76300 6633 76328 7346
rect 76576 7290 76604 8910
rect 76668 7546 76696 9046
rect 76656 7540 76708 7546
rect 76656 7482 76708 7488
rect 76392 7262 76604 7290
rect 76286 6624 76342 6633
rect 76286 6559 76342 6568
rect 76392 6458 76420 7262
rect 76472 7200 76524 7206
rect 76472 7142 76524 7148
rect 76484 6662 76512 7142
rect 76748 6724 76800 6730
rect 76748 6666 76800 6672
rect 76472 6656 76524 6662
rect 76564 6656 76616 6662
rect 76472 6598 76524 6604
rect 76562 6624 76564 6633
rect 76616 6624 76618 6633
rect 76380 6452 76432 6458
rect 76380 6394 76432 6400
rect 76286 5944 76342 5953
rect 76286 5879 76288 5888
rect 76340 5879 76342 5888
rect 76288 5850 76340 5856
rect 76288 5568 76340 5574
rect 76288 5510 76340 5516
rect 76300 5234 76328 5510
rect 76288 5228 76340 5234
rect 76288 5170 76340 5176
rect 76196 4820 76248 4826
rect 76196 4762 76248 4768
rect 75920 4276 75972 4282
rect 75840 4236 75920 4264
rect 75920 4218 75972 4224
rect 75184 4072 75236 4078
rect 75184 4014 75236 4020
rect 75932 3670 75960 4218
rect 76208 4010 76236 4762
rect 76392 4690 76420 6394
rect 76484 6236 76512 6598
rect 76618 6582 76696 6610
rect 76562 6559 76618 6568
rect 76564 6248 76616 6254
rect 76484 6208 76564 6236
rect 76564 6190 76616 6196
rect 76668 6118 76696 6582
rect 76656 6112 76708 6118
rect 76760 6089 76788 6666
rect 76852 6662 76880 9658
rect 76932 9512 76984 9518
rect 76932 9454 76984 9460
rect 76944 8974 76972 9454
rect 76932 8968 76984 8974
rect 76932 8910 76984 8916
rect 77312 6914 77340 15030
rect 77404 14550 77432 15302
rect 77392 14544 77444 14550
rect 77392 14486 77444 14492
rect 77496 13433 77524 15846
rect 77864 15473 77892 16186
rect 78864 16108 78916 16114
rect 78864 16050 78916 16056
rect 78772 15904 78824 15910
rect 78772 15846 78824 15852
rect 77850 15464 77906 15473
rect 78784 15434 78812 15846
rect 77850 15399 77906 15408
rect 78772 15428 78824 15434
rect 77864 15094 77892 15399
rect 78772 15370 78824 15376
rect 77852 15088 77904 15094
rect 78680 15088 78732 15094
rect 77852 15030 77904 15036
rect 78678 15056 78680 15065
rect 78732 15056 78734 15065
rect 78876 15026 78904 16050
rect 82174 16008 82230 16017
rect 80704 15972 80756 15978
rect 82174 15943 82230 15952
rect 80704 15914 80756 15920
rect 80612 15904 80664 15910
rect 80612 15846 80664 15852
rect 80244 15564 80296 15570
rect 80244 15506 80296 15512
rect 80152 15360 80204 15366
rect 80152 15302 80204 15308
rect 80164 15094 80192 15302
rect 80152 15088 80204 15094
rect 80152 15030 80204 15036
rect 78678 14991 78734 15000
rect 78864 15020 78916 15026
rect 78220 14816 78272 14822
rect 78220 14758 78272 14764
rect 77668 14612 77720 14618
rect 77720 14572 77800 14600
rect 77668 14554 77720 14560
rect 77482 13424 77538 13433
rect 77482 13359 77538 13368
rect 77574 12336 77630 12345
rect 77574 12271 77576 12280
rect 77628 12271 77630 12280
rect 77576 12242 77628 12248
rect 77484 12232 77536 12238
rect 77484 12174 77536 12180
rect 77496 11762 77524 12174
rect 77484 11756 77536 11762
rect 77484 11698 77536 11704
rect 77484 11348 77536 11354
rect 77484 11290 77536 11296
rect 77496 11082 77524 11290
rect 77484 11076 77536 11082
rect 77484 11018 77536 11024
rect 77588 10470 77616 12242
rect 77772 11286 77800 14572
rect 78232 14346 78260 14758
rect 78496 14612 78548 14618
rect 78496 14554 78548 14560
rect 78220 14340 78272 14346
rect 78220 14282 78272 14288
rect 78404 14340 78456 14346
rect 78404 14282 78456 14288
rect 78416 14074 78444 14282
rect 78404 14068 78456 14074
rect 78404 14010 78456 14016
rect 78220 13932 78272 13938
rect 78220 13874 78272 13880
rect 78128 13864 78180 13870
rect 78128 13806 78180 13812
rect 77944 12368 77996 12374
rect 77944 12310 77996 12316
rect 77956 12102 77984 12310
rect 77852 12096 77904 12102
rect 77852 12038 77904 12044
rect 77944 12096 77996 12102
rect 77944 12038 77996 12044
rect 77760 11280 77812 11286
rect 77760 11222 77812 11228
rect 77864 11218 77892 12038
rect 77942 11928 77998 11937
rect 77942 11863 77998 11872
rect 77956 11762 77984 11863
rect 77944 11756 77996 11762
rect 77944 11698 77996 11704
rect 77852 11212 77904 11218
rect 77852 11154 77904 11160
rect 77760 11144 77812 11150
rect 77680 11104 77760 11132
rect 77576 10464 77628 10470
rect 77680 10441 77708 11104
rect 77760 11086 77812 11092
rect 77956 10538 77984 11698
rect 78140 11354 78168 13806
rect 78232 12782 78260 13874
rect 78508 13546 78536 14554
rect 78588 14476 78640 14482
rect 78588 14418 78640 14424
rect 78600 14074 78628 14418
rect 78588 14068 78640 14074
rect 78588 14010 78640 14016
rect 78416 13518 78536 13546
rect 78312 13456 78364 13462
rect 78312 13398 78364 13404
rect 78220 12776 78272 12782
rect 78220 12718 78272 12724
rect 78324 12646 78352 13398
rect 78312 12640 78364 12646
rect 78312 12582 78364 12588
rect 78416 12238 78444 13518
rect 78600 13138 78628 14010
rect 78692 13938 78720 14991
rect 78864 14962 78916 14968
rect 79600 15020 79652 15026
rect 79600 14962 79652 14968
rect 79324 14816 79376 14822
rect 79324 14758 79376 14764
rect 79232 14340 79284 14346
rect 79232 14282 79284 14288
rect 78864 14272 78916 14278
rect 78864 14214 78916 14220
rect 78680 13932 78732 13938
rect 78680 13874 78732 13880
rect 78876 13682 78904 14214
rect 79048 14000 79100 14006
rect 79048 13942 79100 13948
rect 78508 13110 78628 13138
rect 78784 13654 78904 13682
rect 78508 12306 78536 13110
rect 78784 12968 78812 13654
rect 79060 13530 79088 13942
rect 78956 13524 79008 13530
rect 78956 13466 79008 13472
rect 79048 13524 79100 13530
rect 79048 13466 79100 13472
rect 78968 13326 78996 13466
rect 78956 13320 79008 13326
rect 78956 13262 79008 13268
rect 78600 12940 78812 12968
rect 78600 12646 78628 12940
rect 78680 12844 78732 12850
rect 78680 12786 78732 12792
rect 78588 12640 78640 12646
rect 78588 12582 78640 12588
rect 78692 12442 78720 12786
rect 78588 12436 78640 12442
rect 78588 12378 78640 12384
rect 78680 12436 78732 12442
rect 78680 12378 78732 12384
rect 78600 12322 78628 12378
rect 78956 12368 79008 12374
rect 78600 12316 78956 12322
rect 78600 12310 79008 12316
rect 78496 12300 78548 12306
rect 78600 12294 78996 12310
rect 79244 12306 79272 14282
rect 79232 12300 79284 12306
rect 78496 12242 78548 12248
rect 79232 12242 79284 12248
rect 78404 12232 78456 12238
rect 78404 12174 78456 12180
rect 78692 12158 78996 12186
rect 78692 12102 78720 12158
rect 78680 12096 78732 12102
rect 78680 12038 78732 12044
rect 78680 11892 78732 11898
rect 78680 11834 78732 11840
rect 78128 11348 78180 11354
rect 78128 11290 78180 11296
rect 78588 11348 78640 11354
rect 78588 11290 78640 11296
rect 78496 11280 78548 11286
rect 78600 11257 78628 11290
rect 78496 11222 78548 11228
rect 78586 11248 78642 11257
rect 78508 10674 78536 11222
rect 78586 11183 78642 11192
rect 78600 11150 78628 11183
rect 78692 11150 78720 11834
rect 78864 11620 78916 11626
rect 78864 11562 78916 11568
rect 78876 11354 78904 11562
rect 78864 11348 78916 11354
rect 78864 11290 78916 11296
rect 78968 11234 78996 12158
rect 79048 12164 79100 12170
rect 79048 12106 79100 12112
rect 79060 11937 79088 12106
rect 79046 11928 79102 11937
rect 79336 11898 79364 14758
rect 79612 14414 79640 14962
rect 79600 14408 79652 14414
rect 79600 14350 79652 14356
rect 79508 14272 79560 14278
rect 79508 14214 79560 14220
rect 79416 13320 79468 13326
rect 79416 13262 79468 13268
rect 79428 13161 79456 13262
rect 79414 13152 79470 13161
rect 79414 13087 79470 13096
rect 79520 12918 79548 14214
rect 79612 13394 79640 14350
rect 80060 14272 80112 14278
rect 80060 14214 80112 14220
rect 80072 13938 80100 14214
rect 80060 13932 80112 13938
rect 80060 13874 80112 13880
rect 79692 13728 79744 13734
rect 79744 13676 79916 13682
rect 79692 13670 79916 13676
rect 79704 13654 79916 13670
rect 79888 13546 79916 13654
rect 79692 13524 79744 13530
rect 79888 13518 80008 13546
rect 79692 13466 79744 13472
rect 79600 13388 79652 13394
rect 79600 13330 79652 13336
rect 79508 12912 79560 12918
rect 79508 12854 79560 12860
rect 79600 12368 79652 12374
rect 79600 12310 79652 12316
rect 79612 12102 79640 12310
rect 79600 12096 79652 12102
rect 79600 12038 79652 12044
rect 79046 11863 79102 11872
rect 79324 11892 79376 11898
rect 79324 11834 79376 11840
rect 79600 11824 79652 11830
rect 79600 11766 79652 11772
rect 79048 11756 79100 11762
rect 79048 11698 79100 11704
rect 79508 11756 79560 11762
rect 79508 11698 79560 11704
rect 78876 11206 78996 11234
rect 78588 11144 78640 11150
rect 78588 11086 78640 11092
rect 78680 11144 78732 11150
rect 78680 11086 78732 11092
rect 78496 10668 78548 10674
rect 78496 10610 78548 10616
rect 77944 10532 77996 10538
rect 77944 10474 77996 10480
rect 77576 10406 77628 10412
rect 77666 10432 77722 10441
rect 77666 10367 77722 10376
rect 77680 10062 77708 10367
rect 77668 10056 77720 10062
rect 77668 9998 77720 10004
rect 77392 9988 77444 9994
rect 77392 9930 77444 9936
rect 77760 9988 77812 9994
rect 77760 9930 77812 9936
rect 77404 9178 77432 9930
rect 77668 9920 77720 9926
rect 77668 9862 77720 9868
rect 77392 9172 77444 9178
rect 77392 9114 77444 9120
rect 77680 7834 77708 9862
rect 77772 9518 77800 9930
rect 78128 9920 78180 9926
rect 78128 9862 78180 9868
rect 78140 9586 78168 9862
rect 78128 9580 78180 9586
rect 78128 9522 78180 9528
rect 77760 9512 77812 9518
rect 77760 9454 77812 9460
rect 77944 9512 77996 9518
rect 77944 9454 77996 9460
rect 77956 9194 77984 9454
rect 78128 9376 78180 9382
rect 78128 9318 78180 9324
rect 77864 9166 77984 9194
rect 77864 9042 77892 9166
rect 77852 9036 77904 9042
rect 77852 8978 77904 8984
rect 77944 9036 77996 9042
rect 77944 8978 77996 8984
rect 77956 8566 77984 8978
rect 78140 8906 78168 9318
rect 78128 8900 78180 8906
rect 78128 8842 78180 8848
rect 77944 8560 77996 8566
rect 77944 8502 77996 8508
rect 78128 7948 78180 7954
rect 78128 7890 78180 7896
rect 77680 7806 77800 7834
rect 77668 7744 77720 7750
rect 77668 7686 77720 7692
rect 77680 7410 77708 7686
rect 77668 7404 77720 7410
rect 77668 7346 77720 7352
rect 77312 6886 77616 6914
rect 76932 6792 76984 6798
rect 77300 6792 77352 6798
rect 76932 6734 76984 6740
rect 77298 6760 77300 6769
rect 77352 6760 77354 6769
rect 76840 6656 76892 6662
rect 76840 6598 76892 6604
rect 76656 6054 76708 6060
rect 76746 6080 76802 6089
rect 76746 6015 76802 6024
rect 76748 5840 76800 5846
rect 76748 5782 76800 5788
rect 76472 5568 76524 5574
rect 76472 5510 76524 5516
rect 76484 4758 76512 5510
rect 76760 5302 76788 5782
rect 76944 5574 76972 6734
rect 77354 6718 77432 6746
rect 77298 6695 77354 6704
rect 77404 6458 77432 6718
rect 77392 6452 77444 6458
rect 77392 6394 77444 6400
rect 76932 5568 76984 5574
rect 76932 5510 76984 5516
rect 76748 5296 76800 5302
rect 76748 5238 76800 5244
rect 76838 5264 76894 5273
rect 76944 5234 76972 5510
rect 76838 5199 76840 5208
rect 76892 5199 76894 5208
rect 76932 5228 76984 5234
rect 76840 5170 76892 5176
rect 76932 5170 76984 5176
rect 77484 4820 77536 4826
rect 77484 4762 77536 4768
rect 76472 4752 76524 4758
rect 76472 4694 76524 4700
rect 76380 4684 76432 4690
rect 76380 4626 76432 4632
rect 76196 4004 76248 4010
rect 76196 3946 76248 3952
rect 76392 3942 76420 4626
rect 76932 4616 76984 4622
rect 76932 4558 76984 4564
rect 76944 4214 76972 4558
rect 77392 4480 77444 4486
rect 77312 4428 77392 4434
rect 77312 4422 77444 4428
rect 77312 4406 77432 4422
rect 77312 4282 77340 4406
rect 77496 4282 77524 4762
rect 77300 4276 77352 4282
rect 77300 4218 77352 4224
rect 77484 4276 77536 4282
rect 77484 4218 77536 4224
rect 76932 4208 76984 4214
rect 77588 4185 77616 6886
rect 77772 6798 77800 7806
rect 78140 7546 78168 7890
rect 78128 7540 78180 7546
rect 78128 7482 78180 7488
rect 77944 7404 77996 7410
rect 77944 7346 77996 7352
rect 77956 7002 77984 7346
rect 77944 6996 77996 7002
rect 77944 6938 77996 6944
rect 78036 6928 78088 6934
rect 78036 6870 78088 6876
rect 77760 6792 77812 6798
rect 77760 6734 77812 6740
rect 77852 6112 77904 6118
rect 77852 6054 77904 6060
rect 77864 5953 77892 6054
rect 77850 5944 77906 5953
rect 77850 5879 77852 5888
rect 77904 5879 77906 5888
rect 77852 5850 77904 5856
rect 77864 5819 77892 5850
rect 77668 5568 77720 5574
rect 77668 5510 77720 5516
rect 77680 5234 77708 5510
rect 77668 5228 77720 5234
rect 77668 5170 77720 5176
rect 78048 5166 78076 6870
rect 78508 6730 78536 10610
rect 78692 10198 78720 11086
rect 78876 11082 78904 11206
rect 78864 11076 78916 11082
rect 78864 11018 78916 11024
rect 78876 10674 78904 11018
rect 78864 10668 78916 10674
rect 78864 10610 78916 10616
rect 78772 10532 78824 10538
rect 78772 10474 78824 10480
rect 78680 10192 78732 10198
rect 78680 10134 78732 10140
rect 78680 8424 78732 8430
rect 78680 8366 78732 8372
rect 78692 7886 78720 8366
rect 78680 7880 78732 7886
rect 78680 7822 78732 7828
rect 78588 7812 78640 7818
rect 78588 7754 78640 7760
rect 78496 6724 78548 6730
rect 78496 6666 78548 6672
rect 78600 6186 78628 7754
rect 78680 7540 78732 7546
rect 78680 7482 78732 7488
rect 78692 7410 78720 7482
rect 78680 7404 78732 7410
rect 78680 7346 78732 7352
rect 78784 6390 78812 10474
rect 78876 9382 78904 10610
rect 79060 9926 79088 11698
rect 79520 10810 79548 11698
rect 79612 11150 79640 11766
rect 79600 11144 79652 11150
rect 79600 11086 79652 11092
rect 79508 10804 79560 10810
rect 79508 10746 79560 10752
rect 79612 10606 79640 11086
rect 79704 11082 79732 13466
rect 79980 13462 80008 13518
rect 79968 13456 80020 13462
rect 79968 13398 80020 13404
rect 80256 13376 80284 15506
rect 80624 15162 80652 15846
rect 80612 15156 80664 15162
rect 80612 15098 80664 15104
rect 80624 15026 80652 15098
rect 80612 15020 80664 15026
rect 80612 14962 80664 14968
rect 80336 14816 80388 14822
rect 80336 14758 80388 14764
rect 80348 14482 80376 14758
rect 80624 14482 80652 14962
rect 80716 14958 80744 15914
rect 81256 15496 81308 15502
rect 81256 15438 81308 15444
rect 80704 14952 80756 14958
rect 80704 14894 80756 14900
rect 80336 14476 80388 14482
rect 80336 14418 80388 14424
rect 80612 14476 80664 14482
rect 80612 14418 80664 14424
rect 80612 14272 80664 14278
rect 80612 14214 80664 14220
rect 80520 13728 80572 13734
rect 80520 13670 80572 13676
rect 80336 13388 80388 13394
rect 80256 13348 80336 13376
rect 80336 13330 80388 13336
rect 79876 13184 79928 13190
rect 79876 13126 79928 13132
rect 79968 13184 80020 13190
rect 79968 13126 80020 13132
rect 79888 12986 79916 13126
rect 79876 12980 79928 12986
rect 79876 12922 79928 12928
rect 79980 12442 80008 13126
rect 80152 12640 80204 12646
rect 80152 12582 80204 12588
rect 79968 12436 80020 12442
rect 79968 12378 80020 12384
rect 79876 12368 79928 12374
rect 79876 12310 79928 12316
rect 79784 12300 79836 12306
rect 79784 12242 79836 12248
rect 79796 12170 79824 12242
rect 79888 12238 79916 12310
rect 79876 12232 79928 12238
rect 79876 12174 79928 12180
rect 79784 12164 79836 12170
rect 79784 12106 79836 12112
rect 79980 11354 80008 12378
rect 80164 11830 80192 12582
rect 80244 12436 80296 12442
rect 80244 12378 80296 12384
rect 80152 11824 80204 11830
rect 80152 11766 80204 11772
rect 80256 11694 80284 12378
rect 80348 12306 80376 13330
rect 80532 12850 80560 13670
rect 80624 13190 80652 14214
rect 80716 13841 80744 14894
rect 80702 13832 80758 13841
rect 80702 13767 80758 13776
rect 80796 13796 80848 13802
rect 80796 13738 80848 13744
rect 80612 13184 80664 13190
rect 80612 13126 80664 13132
rect 80520 12844 80572 12850
rect 80520 12786 80572 12792
rect 80336 12300 80388 12306
rect 80336 12242 80388 12248
rect 80624 11898 80652 13126
rect 80808 12442 80836 13738
rect 81072 13728 81124 13734
rect 81072 13670 81124 13676
rect 80796 12436 80848 12442
rect 80796 12378 80848 12384
rect 81084 12374 81112 13670
rect 81164 13456 81216 13462
rect 81164 13398 81216 13404
rect 81176 13190 81204 13398
rect 81164 13184 81216 13190
rect 81164 13126 81216 13132
rect 81268 12374 81296 15438
rect 81624 15360 81676 15366
rect 81624 15302 81676 15308
rect 81348 14272 81400 14278
rect 81348 14214 81400 14220
rect 81360 14074 81388 14214
rect 81348 14068 81400 14074
rect 81348 14010 81400 14016
rect 81348 13932 81400 13938
rect 81348 13874 81400 13880
rect 81072 12368 81124 12374
rect 81072 12310 81124 12316
rect 81256 12368 81308 12374
rect 81256 12310 81308 12316
rect 81164 12164 81216 12170
rect 81164 12106 81216 12112
rect 80612 11892 80664 11898
rect 80612 11834 80664 11840
rect 80704 11756 80756 11762
rect 80704 11698 80756 11704
rect 80244 11688 80296 11694
rect 80244 11630 80296 11636
rect 79968 11348 80020 11354
rect 79968 11290 80020 11296
rect 80716 11286 80744 11698
rect 80704 11280 80756 11286
rect 80704 11222 80756 11228
rect 81176 11218 81204 12106
rect 81256 11824 81308 11830
rect 81360 11812 81388 13874
rect 81532 12640 81584 12646
rect 81532 12582 81584 12588
rect 81308 11784 81388 11812
rect 81438 11792 81494 11801
rect 81256 11766 81308 11772
rect 80152 11212 80204 11218
rect 80152 11154 80204 11160
rect 81164 11212 81216 11218
rect 81164 11154 81216 11160
rect 79692 11076 79744 11082
rect 79692 11018 79744 11024
rect 79600 10600 79652 10606
rect 79600 10542 79652 10548
rect 79966 10160 80022 10169
rect 79784 10124 79836 10130
rect 79966 10095 80022 10104
rect 79784 10066 79836 10072
rect 79140 10056 79192 10062
rect 79140 9998 79192 10004
rect 79048 9920 79100 9926
rect 79048 9862 79100 9868
rect 78956 9648 79008 9654
rect 78956 9590 79008 9596
rect 78864 9376 78916 9382
rect 78864 9318 78916 9324
rect 78862 8936 78918 8945
rect 78862 8871 78918 8880
rect 78968 8922 78996 9590
rect 79152 9586 79180 9998
rect 79416 9920 79468 9926
rect 79416 9862 79468 9868
rect 79232 9648 79284 9654
rect 79232 9590 79284 9596
rect 79140 9580 79192 9586
rect 79140 9522 79192 9528
rect 79152 9178 79180 9522
rect 79244 9450 79272 9590
rect 79232 9444 79284 9450
rect 79232 9386 79284 9392
rect 79140 9172 79192 9178
rect 79140 9114 79192 9120
rect 79140 8968 79192 8974
rect 78968 8916 79140 8922
rect 78968 8910 79192 8916
rect 78968 8894 79180 8910
rect 78876 8566 78904 8871
rect 78864 8560 78916 8566
rect 78864 8502 78916 8508
rect 78864 8424 78916 8430
rect 78864 8366 78916 8372
rect 78876 8022 78904 8366
rect 78864 8016 78916 8022
rect 78864 7958 78916 7964
rect 78864 7404 78916 7410
rect 78864 7346 78916 7352
rect 78876 6866 78904 7346
rect 78864 6860 78916 6866
rect 78864 6802 78916 6808
rect 78968 6798 78996 8894
rect 79048 8084 79100 8090
rect 79048 8026 79100 8032
rect 78956 6792 79008 6798
rect 78956 6734 79008 6740
rect 78772 6384 78824 6390
rect 78772 6326 78824 6332
rect 78588 6180 78640 6186
rect 78588 6122 78640 6128
rect 79060 5710 79088 8026
rect 79244 6390 79272 9386
rect 79428 9178 79456 9862
rect 79600 9376 79652 9382
rect 79600 9318 79652 9324
rect 79416 9172 79468 9178
rect 79416 9114 79468 9120
rect 79232 6384 79284 6390
rect 79232 6326 79284 6332
rect 79048 5704 79100 5710
rect 79048 5646 79100 5652
rect 78772 5636 78824 5642
rect 78772 5578 78824 5584
rect 78036 5160 78088 5166
rect 78036 5102 78088 5108
rect 78048 4758 78076 5102
rect 78036 4752 78088 4758
rect 78036 4694 78088 4700
rect 76932 4150 76984 4156
rect 77574 4176 77630 4185
rect 77574 4111 77630 4120
rect 78048 4078 78076 4694
rect 78784 4554 78812 5578
rect 78404 4548 78456 4554
rect 78404 4490 78456 4496
rect 78772 4548 78824 4554
rect 78772 4490 78824 4496
rect 78416 4214 78444 4490
rect 78680 4480 78732 4486
rect 78680 4422 78732 4428
rect 78404 4208 78456 4214
rect 78404 4150 78456 4156
rect 78036 4072 78088 4078
rect 78036 4014 78088 4020
rect 78588 4072 78640 4078
rect 78588 4014 78640 4020
rect 76380 3936 76432 3942
rect 76380 3878 76432 3884
rect 75920 3664 75972 3670
rect 75920 3606 75972 3612
rect 76288 3664 76340 3670
rect 76288 3606 76340 3612
rect 76300 3126 76328 3606
rect 76392 3534 76420 3878
rect 76380 3528 76432 3534
rect 76380 3470 76432 3476
rect 77852 3392 77904 3398
rect 77852 3334 77904 3340
rect 76288 3120 76340 3126
rect 76288 3062 76340 3068
rect 77864 3058 77892 3334
rect 78048 3126 78076 4014
rect 78600 3194 78628 4014
rect 78588 3188 78640 3194
rect 78588 3130 78640 3136
rect 78036 3120 78088 3126
rect 78036 3062 78088 3068
rect 77852 3052 77904 3058
rect 77852 2994 77904 3000
rect 78692 2990 78720 4422
rect 78784 3602 78812 4490
rect 78772 3596 78824 3602
rect 78772 3538 78824 3544
rect 78680 2984 78732 2990
rect 78680 2926 78732 2932
rect 78680 2848 78732 2854
rect 78680 2790 78732 2796
rect 78692 2666 78720 2790
rect 78600 2650 78720 2666
rect 78784 2650 78812 3538
rect 79060 3466 79088 5646
rect 79612 4842 79640 9318
rect 79796 8537 79824 10066
rect 79980 10062 80008 10095
rect 79968 10056 80020 10062
rect 79968 9998 80020 10004
rect 79980 9674 80008 9998
rect 79888 9646 80008 9674
rect 79782 8528 79838 8537
rect 79782 8463 79838 8472
rect 79888 8401 79916 9646
rect 79874 8392 79930 8401
rect 79874 8327 79930 8336
rect 79876 7880 79928 7886
rect 79876 7822 79928 7828
rect 80060 7880 80112 7886
rect 80060 7822 80112 7828
rect 79888 7206 79916 7822
rect 80072 7206 80100 7822
rect 79876 7200 79928 7206
rect 79876 7142 79928 7148
rect 80060 7200 80112 7206
rect 80060 7142 80112 7148
rect 79784 6792 79836 6798
rect 79784 6734 79836 6740
rect 79692 6384 79744 6390
rect 79692 6326 79744 6332
rect 79704 5710 79732 6326
rect 79692 5704 79744 5710
rect 79692 5646 79744 5652
rect 79796 5658 79824 6734
rect 79888 6662 79916 7142
rect 79968 6996 80020 7002
rect 79968 6938 80020 6944
rect 79876 6656 79928 6662
rect 79980 6633 80008 6938
rect 79876 6598 79928 6604
rect 79966 6624 80022 6633
rect 79966 6559 80022 6568
rect 79796 5630 80008 5658
rect 79980 5574 80008 5630
rect 79876 5568 79928 5574
rect 79876 5510 79928 5516
rect 79968 5568 80020 5574
rect 80060 5568 80112 5574
rect 79968 5510 80020 5516
rect 80058 5536 80060 5545
rect 80112 5536 80114 5545
rect 79612 4814 79732 4842
rect 79888 4826 79916 5510
rect 80058 5471 80114 5480
rect 80060 5364 80112 5370
rect 80060 5306 80112 5312
rect 79704 4554 79732 4814
rect 79876 4820 79928 4826
rect 79876 4762 79928 4768
rect 79692 4548 79744 4554
rect 79692 4490 79744 4496
rect 79888 3466 79916 4762
rect 79968 4684 80020 4690
rect 79968 4626 80020 4632
rect 79980 4282 80008 4626
rect 80072 4570 80100 5306
rect 80164 5030 80192 11154
rect 80428 11008 80480 11014
rect 80428 10950 80480 10956
rect 80440 10810 80468 10950
rect 80428 10804 80480 10810
rect 80428 10746 80480 10752
rect 80796 10124 80848 10130
rect 80796 10066 80848 10072
rect 80244 9920 80296 9926
rect 80244 9862 80296 9868
rect 80256 8498 80284 9862
rect 80704 9512 80756 9518
rect 80704 9454 80756 9460
rect 80612 9444 80664 9450
rect 80612 9386 80664 9392
rect 80624 9110 80652 9386
rect 80612 9104 80664 9110
rect 80612 9046 80664 9052
rect 80520 8968 80572 8974
rect 80518 8936 80520 8945
rect 80572 8936 80574 8945
rect 80518 8871 80574 8880
rect 80532 8634 80560 8871
rect 80520 8628 80572 8634
rect 80520 8570 80572 8576
rect 80244 8492 80296 8498
rect 80244 8434 80296 8440
rect 80520 7880 80572 7886
rect 80520 7822 80572 7828
rect 80428 7744 80480 7750
rect 80428 7686 80480 7692
rect 80336 7404 80388 7410
rect 80336 7346 80388 7352
rect 80348 7002 80376 7346
rect 80336 6996 80388 7002
rect 80336 6938 80388 6944
rect 80440 6866 80468 7686
rect 80532 6934 80560 7822
rect 80716 7478 80744 9454
rect 80808 8537 80836 10066
rect 81268 8974 81296 11766
rect 81438 11727 81494 11736
rect 81452 11218 81480 11727
rect 81440 11212 81492 11218
rect 81440 11154 81492 11160
rect 81348 10736 81400 10742
rect 81348 10678 81400 10684
rect 81360 10266 81388 10678
rect 81348 10260 81400 10266
rect 81348 10202 81400 10208
rect 81544 9625 81572 12582
rect 81636 11665 81664 15302
rect 82188 15162 82216 15943
rect 82979 15804 83287 15813
rect 82979 15802 82985 15804
rect 83041 15802 83065 15804
rect 83121 15802 83145 15804
rect 83201 15802 83225 15804
rect 83281 15802 83287 15804
rect 83041 15750 83043 15802
rect 83223 15750 83225 15802
rect 82979 15748 82985 15750
rect 83041 15748 83065 15750
rect 83121 15748 83145 15750
rect 83201 15748 83225 15750
rect 83281 15748 83287 15750
rect 82979 15739 83287 15748
rect 82820 15496 82872 15502
rect 82820 15438 82872 15444
rect 82176 15156 82228 15162
rect 82176 15098 82228 15104
rect 82544 15020 82596 15026
rect 82544 14962 82596 14968
rect 81716 14816 81768 14822
rect 81716 14758 81768 14764
rect 81728 12306 81756 14758
rect 81808 14408 81860 14414
rect 81808 14350 81860 14356
rect 81716 12300 81768 12306
rect 81716 12242 81768 12248
rect 81622 11656 81678 11665
rect 81622 11591 81678 11600
rect 81728 10130 81756 12242
rect 81820 12238 81848 14350
rect 82556 14346 82584 14962
rect 82832 14958 82860 15438
rect 83004 15428 83056 15434
rect 83004 15370 83056 15376
rect 83016 14958 83044 15370
rect 82820 14952 82872 14958
rect 82820 14894 82872 14900
rect 83004 14952 83056 14958
rect 83004 14894 83056 14900
rect 82979 14716 83287 14725
rect 82979 14714 82985 14716
rect 83041 14714 83065 14716
rect 83121 14714 83145 14716
rect 83201 14714 83225 14716
rect 83281 14714 83287 14716
rect 83041 14662 83043 14714
rect 83223 14662 83225 14714
rect 82979 14660 82985 14662
rect 83041 14660 83065 14662
rect 83121 14660 83145 14662
rect 83201 14660 83225 14662
rect 83281 14660 83287 14662
rect 82979 14651 83287 14660
rect 82544 14340 82596 14346
rect 82544 14282 82596 14288
rect 82979 13628 83287 13637
rect 82979 13626 82985 13628
rect 83041 13626 83065 13628
rect 83121 13626 83145 13628
rect 83201 13626 83225 13628
rect 83281 13626 83287 13628
rect 83041 13574 83043 13626
rect 83223 13574 83225 13626
rect 82979 13572 82985 13574
rect 83041 13572 83065 13574
rect 83121 13572 83145 13574
rect 83201 13572 83225 13574
rect 83281 13572 83287 13574
rect 82979 13563 83287 13572
rect 83188 13252 83240 13258
rect 83188 13194 83240 13200
rect 82266 13152 82322 13161
rect 82266 13087 82322 13096
rect 82280 12850 82308 13087
rect 83200 12986 83228 13194
rect 83188 12980 83240 12986
rect 83188 12922 83240 12928
rect 82268 12844 82320 12850
rect 82268 12786 82320 12792
rect 82979 12540 83287 12549
rect 82979 12538 82985 12540
rect 83041 12538 83065 12540
rect 83121 12538 83145 12540
rect 83201 12538 83225 12540
rect 83281 12538 83287 12540
rect 83041 12486 83043 12538
rect 83223 12486 83225 12538
rect 82979 12484 82985 12486
rect 83041 12484 83065 12486
rect 83121 12484 83145 12486
rect 83201 12484 83225 12486
rect 83281 12484 83287 12486
rect 82979 12475 83287 12484
rect 83384 12434 83412 16662
rect 83568 16590 83596 19200
rect 84016 17264 84068 17270
rect 84016 17206 84068 17212
rect 83740 17060 83792 17066
rect 83740 17002 83792 17008
rect 83752 16794 83780 17002
rect 83740 16788 83792 16794
rect 83740 16730 83792 16736
rect 83556 16584 83608 16590
rect 83556 16526 83608 16532
rect 83464 15904 83516 15910
rect 83464 15846 83516 15852
rect 83924 15904 83976 15910
rect 83924 15846 83976 15852
rect 83476 14414 83504 15846
rect 83740 15360 83792 15366
rect 83740 15302 83792 15308
rect 83464 14408 83516 14414
rect 83464 14350 83516 14356
rect 83476 14074 83504 14350
rect 83464 14068 83516 14074
rect 83464 14010 83516 14016
rect 83556 13864 83608 13870
rect 83556 13806 83608 13812
rect 83384 12406 83504 12434
rect 81808 12232 81860 12238
rect 81808 12174 81860 12180
rect 81820 10169 81848 12174
rect 82360 12096 82412 12102
rect 82360 12038 82412 12044
rect 82372 11830 82400 12038
rect 82360 11824 82412 11830
rect 82360 11766 82412 11772
rect 83004 11688 83056 11694
rect 82542 11656 82598 11665
rect 83004 11630 83056 11636
rect 82542 11591 82598 11600
rect 82556 11150 82584 11591
rect 83016 11558 83044 11630
rect 83004 11552 83056 11558
rect 83004 11494 83056 11500
rect 82979 11452 83287 11461
rect 82979 11450 82985 11452
rect 83041 11450 83065 11452
rect 83121 11450 83145 11452
rect 83201 11450 83225 11452
rect 83281 11450 83287 11452
rect 83041 11398 83043 11450
rect 83223 11398 83225 11450
rect 82979 11396 82985 11398
rect 83041 11396 83065 11398
rect 83121 11396 83145 11398
rect 83201 11396 83225 11398
rect 83281 11396 83287 11398
rect 82979 11387 83287 11396
rect 82544 11144 82596 11150
rect 82544 11086 82596 11092
rect 82176 11076 82228 11082
rect 82228 11036 82308 11064
rect 82176 11018 82228 11024
rect 82280 10810 82308 11036
rect 82268 10804 82320 10810
rect 82268 10746 82320 10752
rect 82280 10674 82308 10746
rect 82268 10668 82320 10674
rect 82268 10610 82320 10616
rect 83372 10668 83424 10674
rect 83372 10610 83424 10616
rect 82360 10464 82412 10470
rect 82360 10406 82412 10412
rect 81806 10160 81862 10169
rect 81716 10124 81768 10130
rect 81806 10095 81862 10104
rect 81716 10066 81768 10072
rect 82372 10062 82400 10406
rect 82979 10364 83287 10373
rect 82979 10362 82985 10364
rect 83041 10362 83065 10364
rect 83121 10362 83145 10364
rect 83201 10362 83225 10364
rect 83281 10362 83287 10364
rect 83041 10310 83043 10362
rect 83223 10310 83225 10362
rect 82979 10308 82985 10310
rect 83041 10308 83065 10310
rect 83121 10308 83145 10310
rect 83201 10308 83225 10310
rect 83281 10308 83287 10310
rect 82979 10299 83287 10308
rect 83384 10130 83412 10610
rect 83372 10124 83424 10130
rect 83372 10066 83424 10072
rect 82360 10056 82412 10062
rect 82360 9998 82412 10004
rect 81530 9616 81586 9625
rect 83384 9586 83412 10066
rect 83476 9674 83504 12406
rect 83568 11694 83596 13806
rect 83648 12164 83700 12170
rect 83648 12106 83700 12112
rect 83556 11688 83608 11694
rect 83556 11630 83608 11636
rect 83568 10674 83596 11630
rect 83556 10668 83608 10674
rect 83556 10610 83608 10616
rect 83476 9646 83596 9674
rect 81530 9551 81586 9560
rect 82820 9580 82872 9586
rect 82820 9522 82872 9528
rect 83372 9580 83424 9586
rect 83372 9522 83424 9528
rect 82728 9512 82780 9518
rect 82728 9454 82780 9460
rect 81440 9444 81492 9450
rect 81440 9386 81492 9392
rect 81256 8968 81308 8974
rect 81256 8910 81308 8916
rect 80794 8528 80850 8537
rect 80794 8463 80850 8472
rect 80704 7472 80756 7478
rect 80704 7414 80756 7420
rect 80520 6928 80572 6934
rect 80520 6870 80572 6876
rect 80428 6860 80480 6866
rect 80428 6802 80480 6808
rect 80336 6792 80388 6798
rect 80334 6760 80336 6769
rect 80388 6760 80390 6769
rect 80334 6695 80390 6704
rect 80334 6624 80390 6633
rect 80334 6559 80390 6568
rect 80244 6248 80296 6254
rect 80244 6190 80296 6196
rect 80256 5166 80284 6190
rect 80348 5642 80376 6559
rect 80336 5636 80388 5642
rect 80336 5578 80388 5584
rect 80244 5160 80296 5166
rect 80244 5102 80296 5108
rect 80152 5024 80204 5030
rect 80152 4966 80204 4972
rect 80072 4542 80284 4570
rect 80256 4282 80284 4542
rect 79968 4276 80020 4282
rect 79968 4218 80020 4224
rect 80244 4276 80296 4282
rect 80244 4218 80296 4224
rect 79980 4078 80008 4218
rect 80532 4146 80560 6870
rect 80704 6384 80756 6390
rect 80624 6344 80704 6372
rect 80624 5302 80652 6344
rect 80704 6326 80756 6332
rect 80808 5846 80836 8463
rect 81268 8362 81296 8910
rect 81256 8356 81308 8362
rect 81256 8298 81308 8304
rect 81268 6254 81296 8298
rect 81452 8106 81480 9386
rect 81532 8900 81584 8906
rect 81532 8842 81584 8848
rect 81544 8634 81572 8842
rect 81532 8628 81584 8634
rect 81532 8570 81584 8576
rect 82636 8628 82688 8634
rect 82636 8570 82688 8576
rect 82648 8498 82676 8570
rect 82636 8492 82688 8498
rect 82636 8434 82688 8440
rect 81716 8424 81768 8430
rect 81716 8366 81768 8372
rect 81452 8078 81572 8106
rect 81440 7948 81492 7954
rect 81440 7890 81492 7896
rect 81348 7472 81400 7478
rect 81348 7414 81400 7420
rect 81256 6248 81308 6254
rect 81256 6190 81308 6196
rect 80980 5908 81032 5914
rect 80980 5850 81032 5856
rect 80796 5840 80848 5846
rect 80796 5782 80848 5788
rect 80704 5772 80756 5778
rect 80704 5714 80756 5720
rect 80612 5296 80664 5302
rect 80612 5238 80664 5244
rect 80624 4214 80652 5238
rect 80716 4622 80744 5714
rect 80992 5166 81020 5850
rect 81268 5817 81296 6190
rect 81254 5808 81310 5817
rect 81254 5743 81310 5752
rect 81360 5710 81388 7414
rect 81348 5704 81400 5710
rect 81452 5681 81480 7890
rect 81544 6118 81572 8078
rect 81728 8022 81756 8366
rect 81716 8016 81768 8022
rect 81716 7958 81768 7964
rect 81728 7342 81756 7958
rect 82648 7886 82676 8434
rect 82740 8294 82768 9454
rect 82832 8838 82860 9522
rect 82979 9276 83287 9285
rect 82979 9274 82985 9276
rect 83041 9274 83065 9276
rect 83121 9274 83145 9276
rect 83201 9274 83225 9276
rect 83281 9274 83287 9276
rect 83041 9222 83043 9274
rect 83223 9222 83225 9274
rect 82979 9220 82985 9222
rect 83041 9220 83065 9222
rect 83121 9220 83145 9222
rect 83201 9220 83225 9222
rect 83281 9220 83287 9222
rect 82979 9211 83287 9220
rect 82820 8832 82872 8838
rect 82820 8774 82872 8780
rect 83464 8832 83516 8838
rect 83464 8774 83516 8780
rect 82728 8288 82780 8294
rect 82728 8230 82780 8236
rect 82636 7880 82688 7886
rect 82636 7822 82688 7828
rect 82176 7812 82228 7818
rect 82176 7754 82228 7760
rect 81624 7336 81676 7342
rect 81624 7278 81676 7284
rect 81716 7336 81768 7342
rect 81716 7278 81768 7284
rect 81636 6798 81664 7278
rect 82188 6798 82216 7754
rect 82636 7540 82688 7546
rect 82636 7482 82688 7488
rect 82648 7002 82676 7482
rect 82636 6996 82688 7002
rect 82636 6938 82688 6944
rect 82544 6860 82596 6866
rect 82544 6802 82596 6808
rect 81624 6792 81676 6798
rect 82176 6792 82228 6798
rect 81624 6734 81676 6740
rect 81714 6760 81770 6769
rect 82176 6734 82228 6740
rect 81714 6695 81716 6704
rect 81768 6695 81770 6704
rect 81716 6666 81768 6672
rect 81624 6248 81676 6254
rect 81624 6190 81676 6196
rect 81992 6248 82044 6254
rect 81992 6190 82044 6196
rect 81532 6112 81584 6118
rect 81532 6054 81584 6060
rect 81544 5778 81572 6054
rect 81636 5778 81664 6190
rect 81532 5772 81584 5778
rect 81532 5714 81584 5720
rect 81624 5772 81676 5778
rect 81624 5714 81676 5720
rect 81348 5646 81400 5652
rect 81438 5672 81494 5681
rect 81438 5607 81494 5616
rect 81440 5568 81492 5574
rect 81440 5510 81492 5516
rect 81452 5166 81480 5510
rect 80980 5160 81032 5166
rect 80980 5102 81032 5108
rect 81440 5160 81492 5166
rect 81440 5102 81492 5108
rect 81440 5024 81492 5030
rect 81440 4966 81492 4972
rect 80704 4616 80756 4622
rect 80704 4558 80756 4564
rect 80612 4208 80664 4214
rect 80612 4150 80664 4156
rect 80520 4140 80572 4146
rect 80520 4082 80572 4088
rect 79968 4072 80020 4078
rect 79968 4014 80020 4020
rect 80704 4072 80756 4078
rect 80704 4014 80756 4020
rect 80716 3670 80744 4014
rect 80704 3664 80756 3670
rect 80704 3606 80756 3612
rect 79048 3460 79100 3466
rect 79048 3402 79100 3408
rect 79232 3460 79284 3466
rect 79232 3402 79284 3408
rect 79876 3460 79928 3466
rect 79876 3402 79928 3408
rect 79244 3194 79272 3402
rect 79232 3188 79284 3194
rect 79232 3130 79284 3136
rect 79888 3058 79916 3402
rect 80716 3398 80744 3606
rect 80704 3392 80756 3398
rect 80704 3334 80756 3340
rect 81452 3194 81480 4966
rect 81544 4622 81572 5714
rect 82004 5710 82032 6190
rect 81992 5704 82044 5710
rect 81992 5646 82044 5652
rect 81624 5568 81676 5574
rect 81622 5536 81624 5545
rect 81676 5536 81678 5545
rect 81622 5471 81678 5480
rect 82004 5370 82032 5646
rect 81992 5364 82044 5370
rect 81992 5306 82044 5312
rect 81532 4616 81584 4622
rect 81532 4558 81584 4564
rect 81544 3194 81572 4558
rect 81716 4548 81768 4554
rect 81716 4490 81768 4496
rect 81728 3534 81756 4490
rect 82004 4146 82032 5306
rect 82188 5030 82216 6734
rect 82556 6662 82584 6802
rect 82544 6656 82596 6662
rect 82544 6598 82596 6604
rect 82740 6066 82768 8230
rect 82832 7886 82860 8774
rect 83372 8492 83424 8498
rect 83372 8434 83424 8440
rect 82979 8188 83287 8197
rect 82979 8186 82985 8188
rect 83041 8186 83065 8188
rect 83121 8186 83145 8188
rect 83201 8186 83225 8188
rect 83281 8186 83287 8188
rect 83041 8134 83043 8186
rect 83223 8134 83225 8186
rect 82979 8132 82985 8134
rect 83041 8132 83065 8134
rect 83121 8132 83145 8134
rect 83201 8132 83225 8134
rect 83281 8132 83287 8134
rect 82979 8123 83287 8132
rect 82820 7880 82872 7886
rect 82820 7822 82872 7828
rect 83280 7540 83332 7546
rect 83280 7482 83332 7488
rect 83292 7410 83320 7482
rect 83280 7404 83332 7410
rect 83280 7346 83332 7352
rect 82820 7200 82872 7206
rect 82820 7142 82872 7148
rect 82832 6254 82860 7142
rect 82979 7100 83287 7109
rect 82979 7098 82985 7100
rect 83041 7098 83065 7100
rect 83121 7098 83145 7100
rect 83201 7098 83225 7100
rect 83281 7098 83287 7100
rect 83041 7046 83043 7098
rect 83223 7046 83225 7098
rect 82979 7044 82985 7046
rect 83041 7044 83065 7046
rect 83121 7044 83145 7046
rect 83201 7044 83225 7046
rect 83281 7044 83287 7046
rect 82979 7035 83287 7044
rect 83188 6452 83240 6458
rect 83188 6394 83240 6400
rect 82820 6248 82872 6254
rect 82820 6190 82872 6196
rect 83200 6202 83228 6394
rect 83384 6322 83412 8434
rect 83372 6316 83424 6322
rect 83372 6258 83424 6264
rect 83476 6202 83504 8774
rect 83568 8566 83596 9646
rect 83556 8560 83608 8566
rect 83556 8502 83608 8508
rect 83568 7585 83596 8502
rect 83660 8498 83688 12106
rect 83752 11801 83780 15302
rect 83936 15094 83964 15846
rect 83924 15088 83976 15094
rect 83924 15030 83976 15036
rect 83832 12708 83884 12714
rect 83832 12650 83884 12656
rect 83738 11792 83794 11801
rect 83738 11727 83740 11736
rect 83792 11727 83794 11736
rect 83740 11698 83792 11704
rect 83844 11694 83872 12650
rect 83832 11688 83884 11694
rect 83832 11630 83884 11636
rect 83740 11212 83792 11218
rect 83740 11154 83792 11160
rect 83648 8492 83700 8498
rect 83648 8434 83700 8440
rect 83648 7880 83700 7886
rect 83648 7822 83700 7828
rect 83554 7576 83610 7585
rect 83554 7511 83610 7520
rect 83660 7002 83688 7822
rect 83648 6996 83700 7002
rect 83648 6938 83700 6944
rect 83752 6322 83780 11154
rect 83830 10024 83886 10033
rect 83830 9959 83832 9968
rect 83884 9959 83886 9968
rect 83832 9930 83884 9936
rect 83832 9512 83884 9518
rect 83832 9454 83884 9460
rect 83844 7954 83872 9454
rect 83832 7948 83884 7954
rect 83832 7890 83884 7896
rect 83832 6724 83884 6730
rect 83832 6666 83884 6672
rect 83740 6316 83792 6322
rect 83740 6258 83792 6264
rect 83200 6174 83504 6202
rect 83464 6112 83516 6118
rect 82740 6038 82860 6066
rect 83464 6054 83516 6060
rect 82726 5944 82782 5953
rect 82832 5914 82860 6038
rect 82979 6012 83287 6021
rect 82979 6010 82985 6012
rect 83041 6010 83065 6012
rect 83121 6010 83145 6012
rect 83201 6010 83225 6012
rect 83281 6010 83287 6012
rect 83041 5958 83043 6010
rect 83223 5958 83225 6010
rect 82979 5956 82985 5958
rect 83041 5956 83065 5958
rect 83121 5956 83145 5958
rect 83201 5956 83225 5958
rect 83281 5956 83287 5958
rect 82979 5947 83287 5956
rect 83476 5914 83504 6054
rect 82726 5879 82782 5888
rect 82820 5908 82872 5914
rect 82740 5846 82768 5879
rect 82820 5850 82872 5856
rect 83464 5908 83516 5914
rect 83464 5850 83516 5856
rect 82728 5840 82780 5846
rect 82728 5782 82780 5788
rect 82176 5024 82228 5030
rect 82176 4966 82228 4972
rect 83372 5024 83424 5030
rect 83372 4966 83424 4972
rect 82979 4924 83287 4933
rect 82979 4922 82985 4924
rect 83041 4922 83065 4924
rect 83121 4922 83145 4924
rect 83201 4922 83225 4924
rect 83281 4922 83287 4924
rect 83041 4870 83043 4922
rect 83223 4870 83225 4922
rect 82979 4868 82985 4870
rect 83041 4868 83065 4870
rect 83121 4868 83145 4870
rect 83201 4868 83225 4870
rect 83281 4868 83287 4870
rect 82979 4859 83287 4868
rect 82452 4820 82504 4826
rect 82452 4762 82504 4768
rect 82464 4486 82492 4762
rect 83384 4622 83412 4966
rect 83752 4706 83780 6258
rect 83844 6118 83872 6666
rect 83832 6112 83884 6118
rect 83832 6054 83884 6060
rect 83936 4729 83964 15030
rect 84028 12374 84056 17206
rect 91480 17202 91508 19200
rect 94697 17436 95005 17445
rect 94697 17434 94703 17436
rect 94759 17434 94783 17436
rect 94839 17434 94863 17436
rect 94919 17434 94943 17436
rect 94999 17434 95005 17436
rect 94759 17382 94761 17434
rect 94941 17382 94943 17434
rect 94697 17380 94703 17382
rect 94759 17380 94783 17382
rect 94839 17380 94863 17382
rect 94919 17380 94943 17382
rect 94999 17380 95005 17382
rect 94697 17371 95005 17380
rect 91468 17196 91520 17202
rect 91468 17138 91520 17144
rect 94226 16824 94282 16833
rect 94226 16759 94228 16768
rect 94280 16759 94282 16768
rect 94228 16730 94280 16736
rect 87880 16720 87932 16726
rect 87880 16662 87932 16668
rect 86314 16144 86370 16153
rect 86314 16079 86370 16088
rect 84108 15360 84160 15366
rect 84108 15302 84160 15308
rect 84120 14482 84148 15302
rect 84936 15156 84988 15162
rect 84936 15098 84988 15104
rect 84108 14476 84160 14482
rect 84108 14418 84160 14424
rect 84120 13938 84148 14418
rect 84948 14414 84976 15098
rect 85028 14952 85080 14958
rect 85028 14894 85080 14900
rect 84936 14408 84988 14414
rect 84936 14350 84988 14356
rect 84108 13932 84160 13938
rect 84108 13874 84160 13880
rect 84948 13870 84976 14350
rect 85040 14278 85068 14894
rect 85212 14816 85264 14822
rect 85212 14758 85264 14764
rect 85028 14272 85080 14278
rect 85028 14214 85080 14220
rect 84660 13864 84712 13870
rect 84660 13806 84712 13812
rect 84936 13864 84988 13870
rect 84936 13806 84988 13812
rect 84200 13524 84252 13530
rect 84200 13466 84252 13472
rect 84108 12844 84160 12850
rect 84108 12786 84160 12792
rect 84120 12442 84148 12786
rect 84108 12436 84160 12442
rect 84108 12378 84160 12384
rect 84016 12368 84068 12374
rect 84016 12310 84068 12316
rect 84028 11218 84056 12310
rect 84212 12238 84240 13466
rect 84476 13320 84528 13326
rect 84476 13262 84528 13268
rect 84488 12714 84516 13262
rect 84568 13252 84620 13258
rect 84568 13194 84620 13200
rect 84580 12986 84608 13194
rect 84568 12980 84620 12986
rect 84568 12922 84620 12928
rect 84476 12708 84528 12714
rect 84476 12650 84528 12656
rect 84568 12368 84620 12374
rect 84568 12310 84620 12316
rect 84108 12232 84160 12238
rect 84108 12174 84160 12180
rect 84200 12232 84252 12238
rect 84200 12174 84252 12180
rect 84120 11778 84148 12174
rect 84200 12096 84252 12102
rect 84200 12038 84252 12044
rect 84212 11898 84240 12038
rect 84200 11892 84252 11898
rect 84200 11834 84252 11840
rect 84292 11892 84344 11898
rect 84292 11834 84344 11840
rect 84304 11778 84332 11834
rect 84120 11750 84332 11778
rect 84384 11756 84436 11762
rect 84384 11698 84436 11704
rect 84292 11688 84344 11694
rect 84290 11656 84292 11665
rect 84344 11656 84346 11665
rect 84290 11591 84346 11600
rect 84292 11280 84344 11286
rect 84292 11222 84344 11228
rect 84016 11212 84068 11218
rect 84016 11154 84068 11160
rect 84108 11212 84160 11218
rect 84108 11154 84160 11160
rect 84014 11112 84070 11121
rect 84014 11047 84016 11056
rect 84068 11047 84070 11056
rect 84016 11018 84068 11024
rect 84120 11014 84148 11154
rect 84304 11014 84332 11222
rect 84108 11008 84160 11014
rect 84108 10950 84160 10956
rect 84292 11008 84344 11014
rect 84292 10950 84344 10956
rect 84120 10690 84148 10950
rect 84304 10713 84332 10950
rect 84290 10704 84346 10713
rect 84120 10674 84240 10690
rect 84120 10668 84252 10674
rect 84120 10662 84200 10668
rect 84290 10639 84346 10648
rect 84200 10610 84252 10616
rect 84304 10606 84332 10639
rect 84016 10600 84068 10606
rect 84292 10600 84344 10606
rect 84016 10542 84068 10548
rect 84198 10568 84254 10577
rect 84028 8906 84056 10542
rect 84292 10542 84344 10548
rect 84198 10503 84254 10512
rect 84212 10062 84240 10503
rect 84200 10056 84252 10062
rect 84200 9998 84252 10004
rect 84108 9376 84160 9382
rect 84396 9364 84424 11698
rect 84580 11506 84608 12310
rect 84672 11626 84700 13806
rect 85040 13802 85068 14214
rect 85028 13796 85080 13802
rect 85028 13738 85080 13744
rect 85040 12918 85068 13738
rect 85224 13530 85252 14758
rect 85672 14340 85724 14346
rect 85672 14282 85724 14288
rect 85212 13524 85264 13530
rect 85212 13466 85264 13472
rect 85028 12912 85080 12918
rect 85028 12854 85080 12860
rect 84660 11620 84712 11626
rect 84660 11562 84712 11568
rect 84752 11620 84804 11626
rect 84752 11562 84804 11568
rect 84764 11506 84792 11562
rect 84580 11478 84792 11506
rect 85040 11354 85068 12854
rect 85224 12850 85252 13466
rect 85212 12844 85264 12850
rect 85212 12786 85264 12792
rect 85120 12640 85172 12646
rect 85120 12582 85172 12588
rect 85580 12640 85632 12646
rect 85580 12582 85632 12588
rect 85132 12170 85160 12582
rect 85592 12306 85620 12582
rect 85212 12300 85264 12306
rect 85212 12242 85264 12248
rect 85580 12300 85632 12306
rect 85580 12242 85632 12248
rect 85120 12164 85172 12170
rect 85120 12106 85172 12112
rect 85224 11354 85252 12242
rect 85580 12164 85632 12170
rect 85580 12106 85632 12112
rect 85028 11348 85080 11354
rect 85028 11290 85080 11296
rect 85212 11348 85264 11354
rect 85212 11290 85264 11296
rect 84660 10668 84712 10674
rect 84660 10610 84712 10616
rect 84568 10600 84620 10606
rect 84568 10542 84620 10548
rect 84476 9716 84528 9722
rect 84476 9658 84528 9664
rect 84488 9586 84516 9658
rect 84476 9580 84528 9586
rect 84476 9522 84528 9528
rect 84160 9336 84424 9364
rect 84108 9318 84160 9324
rect 84016 8900 84068 8906
rect 84016 8842 84068 8848
rect 84292 8560 84344 8566
rect 84292 8502 84344 8508
rect 84200 8492 84252 8498
rect 84200 8434 84252 8440
rect 84212 8106 84240 8434
rect 84304 8294 84332 8502
rect 84292 8288 84344 8294
rect 84292 8230 84344 8236
rect 84212 8078 84332 8106
rect 84108 7948 84160 7954
rect 84108 7890 84160 7896
rect 84016 6996 84068 7002
rect 84016 6938 84068 6944
rect 84028 6662 84056 6938
rect 84120 6934 84148 7890
rect 84200 7268 84252 7274
rect 84200 7210 84252 7216
rect 84108 6928 84160 6934
rect 84108 6870 84160 6876
rect 84108 6724 84160 6730
rect 84108 6666 84160 6672
rect 84016 6656 84068 6662
rect 84016 6598 84068 6604
rect 84120 6390 84148 6666
rect 84108 6384 84160 6390
rect 84108 6326 84160 6332
rect 84016 5296 84068 5302
rect 84016 5238 84068 5244
rect 83568 4678 83780 4706
rect 83922 4720 83978 4729
rect 82728 4616 82780 4622
rect 82728 4558 82780 4564
rect 83372 4616 83424 4622
rect 83372 4558 83424 4564
rect 82452 4480 82504 4486
rect 82452 4422 82504 4428
rect 81992 4140 82044 4146
rect 81992 4082 82044 4088
rect 81992 3936 82044 3942
rect 81992 3878 82044 3884
rect 82004 3534 82032 3878
rect 82740 3534 82768 4558
rect 82979 3836 83287 3845
rect 82979 3834 82985 3836
rect 83041 3834 83065 3836
rect 83121 3834 83145 3836
rect 83201 3834 83225 3836
rect 83281 3834 83287 3836
rect 83041 3782 83043 3834
rect 83223 3782 83225 3834
rect 82979 3780 82985 3782
rect 83041 3780 83065 3782
rect 83121 3780 83145 3782
rect 83201 3780 83225 3782
rect 83281 3780 83287 3782
rect 82979 3771 83287 3780
rect 81716 3528 81768 3534
rect 81716 3470 81768 3476
rect 81992 3528 82044 3534
rect 81992 3470 82044 3476
rect 82728 3528 82780 3534
rect 82728 3470 82780 3476
rect 81440 3188 81492 3194
rect 81440 3130 81492 3136
rect 81532 3188 81584 3194
rect 81532 3130 81584 3136
rect 79876 3052 79928 3058
rect 79876 2994 79928 3000
rect 81728 2990 81756 3470
rect 82004 3194 82032 3470
rect 81992 3188 82044 3194
rect 81992 3130 82044 3136
rect 83384 2990 83412 4558
rect 83568 4146 83596 4678
rect 83922 4655 83978 4664
rect 83648 4616 83700 4622
rect 83648 4558 83700 4564
rect 83740 4616 83792 4622
rect 83740 4558 83792 4564
rect 83556 4140 83608 4146
rect 83556 4082 83608 4088
rect 83660 3602 83688 4558
rect 83752 4282 83780 4558
rect 83832 4548 83884 4554
rect 83832 4490 83884 4496
rect 83740 4276 83792 4282
rect 83740 4218 83792 4224
rect 83844 4146 83872 4490
rect 84028 4282 84056 5238
rect 84212 5114 84240 7210
rect 84304 5846 84332 8078
rect 84384 7744 84436 7750
rect 84384 7686 84436 7692
rect 84396 6798 84424 7686
rect 84476 7404 84528 7410
rect 84476 7346 84528 7352
rect 84488 7002 84516 7346
rect 84476 6996 84528 7002
rect 84476 6938 84528 6944
rect 84580 6798 84608 10542
rect 84672 9722 84700 10610
rect 85486 10568 85542 10577
rect 84844 10532 84896 10538
rect 85486 10503 85542 10512
rect 84844 10474 84896 10480
rect 84752 10464 84804 10470
rect 84752 10406 84804 10412
rect 84764 10130 84792 10406
rect 84752 10124 84804 10130
rect 84752 10066 84804 10072
rect 84856 10062 84884 10474
rect 85304 10464 85356 10470
rect 85304 10406 85356 10412
rect 85316 10266 85344 10406
rect 85304 10260 85356 10266
rect 85304 10202 85356 10208
rect 85396 10260 85448 10266
rect 85396 10202 85448 10208
rect 85408 10169 85436 10202
rect 85394 10160 85450 10169
rect 85500 10130 85528 10503
rect 85394 10095 85450 10104
rect 85488 10124 85540 10130
rect 85488 10066 85540 10072
rect 84844 10056 84896 10062
rect 84750 10024 84806 10033
rect 84844 9998 84896 10004
rect 84750 9959 84806 9968
rect 84764 9926 84792 9959
rect 84752 9920 84804 9926
rect 84752 9862 84804 9868
rect 84856 9722 84884 9998
rect 84660 9716 84712 9722
rect 84660 9658 84712 9664
rect 84844 9716 84896 9722
rect 84844 9658 84896 9664
rect 85592 9654 85620 12106
rect 85684 11898 85712 14282
rect 85856 14272 85908 14278
rect 85856 14214 85908 14220
rect 85868 13734 85896 14214
rect 85856 13728 85908 13734
rect 85856 13670 85908 13676
rect 85868 12306 85896 13670
rect 86224 13388 86276 13394
rect 86224 13330 86276 13336
rect 86236 12850 86264 13330
rect 86224 12844 86276 12850
rect 86224 12786 86276 12792
rect 86236 12374 86264 12786
rect 86328 12434 86356 16079
rect 86776 15360 86828 15366
rect 86776 15302 86828 15308
rect 86500 15020 86552 15026
rect 86500 14962 86552 14968
rect 86408 14272 86460 14278
rect 86408 14214 86460 14220
rect 86420 13326 86448 14214
rect 86408 13320 86460 13326
rect 86408 13262 86460 13268
rect 86512 13190 86540 14962
rect 86788 14958 86816 15302
rect 86776 14952 86828 14958
rect 86776 14894 86828 14900
rect 86788 14822 86816 14894
rect 86776 14816 86828 14822
rect 86776 14758 86828 14764
rect 86960 14816 87012 14822
rect 86960 14758 87012 14764
rect 86788 14414 86816 14758
rect 86972 14414 87000 14758
rect 86776 14408 86828 14414
rect 86776 14350 86828 14356
rect 86960 14408 87012 14414
rect 86960 14350 87012 14356
rect 86684 13320 86736 13326
rect 86684 13262 86736 13268
rect 86500 13184 86552 13190
rect 86500 13126 86552 13132
rect 86328 12406 86448 12434
rect 86224 12368 86276 12374
rect 86224 12310 86276 12316
rect 85856 12300 85908 12306
rect 85856 12242 85908 12248
rect 86224 12232 86276 12238
rect 86224 12174 86276 12180
rect 85672 11892 85724 11898
rect 85672 11834 85724 11840
rect 86132 11892 86184 11898
rect 86132 11834 86184 11840
rect 85948 11824 86000 11830
rect 85948 11766 86000 11772
rect 85960 11286 85988 11766
rect 86040 11552 86092 11558
rect 86040 11494 86092 11500
rect 85764 11280 85816 11286
rect 85762 11248 85764 11257
rect 85948 11280 86000 11286
rect 85816 11248 85818 11257
rect 85948 11222 86000 11228
rect 85762 11183 85818 11192
rect 86052 11150 86080 11494
rect 86040 11144 86092 11150
rect 86040 11086 86092 11092
rect 85764 10056 85816 10062
rect 85764 9998 85816 10004
rect 85580 9648 85632 9654
rect 85580 9590 85632 9596
rect 85396 9444 85448 9450
rect 85396 9386 85448 9392
rect 85408 8430 85436 9386
rect 85776 9382 85804 9998
rect 85948 9648 86000 9654
rect 85948 9590 86000 9596
rect 85764 9376 85816 9382
rect 85764 9318 85816 9324
rect 85672 9172 85724 9178
rect 85672 9114 85724 9120
rect 85486 8936 85542 8945
rect 85684 8906 85712 9114
rect 85486 8871 85542 8880
rect 85672 8900 85724 8906
rect 85500 8430 85528 8871
rect 85672 8842 85724 8848
rect 85396 8424 85448 8430
rect 85396 8366 85448 8372
rect 85488 8424 85540 8430
rect 85488 8366 85540 8372
rect 84660 8356 84712 8362
rect 84660 8298 84712 8304
rect 84672 7274 84700 8298
rect 84844 8084 84896 8090
rect 84844 8026 84896 8032
rect 84856 7818 84884 8026
rect 84844 7812 84896 7818
rect 84844 7754 84896 7760
rect 84660 7268 84712 7274
rect 84660 7210 84712 7216
rect 84384 6792 84436 6798
rect 84384 6734 84436 6740
rect 84568 6792 84620 6798
rect 84568 6734 84620 6740
rect 84752 6316 84804 6322
rect 84752 6258 84804 6264
rect 84384 6112 84436 6118
rect 84384 6054 84436 6060
rect 84292 5840 84344 5846
rect 84292 5782 84344 5788
rect 84212 5086 84332 5114
rect 84200 5024 84252 5030
rect 84200 4966 84252 4972
rect 84016 4276 84068 4282
rect 84016 4218 84068 4224
rect 83832 4140 83884 4146
rect 83832 4082 83884 4088
rect 84212 4010 84240 4966
rect 84304 4826 84332 5086
rect 84292 4820 84344 4826
rect 84292 4762 84344 4768
rect 84396 4758 84424 6054
rect 84764 5914 84792 6258
rect 84752 5908 84804 5914
rect 84752 5850 84804 5856
rect 84568 5160 84620 5166
rect 84568 5102 84620 5108
rect 84384 4752 84436 4758
rect 84384 4694 84436 4700
rect 84396 4622 84424 4694
rect 84384 4616 84436 4622
rect 84384 4558 84436 4564
rect 84580 4214 84608 5102
rect 84660 5024 84712 5030
rect 84660 4966 84712 4972
rect 84672 4622 84700 4966
rect 84660 4616 84712 4622
rect 84660 4558 84712 4564
rect 84672 4282 84700 4558
rect 84660 4276 84712 4282
rect 84660 4218 84712 4224
rect 84568 4208 84620 4214
rect 84568 4150 84620 4156
rect 84856 4146 84884 7754
rect 84934 7576 84990 7585
rect 85500 7546 85528 8366
rect 84934 7511 84990 7520
rect 85488 7540 85540 7546
rect 84948 5234 84976 7511
rect 85488 7482 85540 7488
rect 85028 7336 85080 7342
rect 85028 7278 85080 7284
rect 85040 6934 85068 7278
rect 85028 6928 85080 6934
rect 85028 6870 85080 6876
rect 85040 6322 85068 6870
rect 85028 6316 85080 6322
rect 85028 6258 85080 6264
rect 85488 6316 85540 6322
rect 85488 6258 85540 6264
rect 85396 5364 85448 5370
rect 85396 5306 85448 5312
rect 85408 5234 85436 5306
rect 84936 5228 84988 5234
rect 84936 5170 84988 5176
rect 85396 5228 85448 5234
rect 85396 5170 85448 5176
rect 84948 4758 84976 5170
rect 85120 5024 85172 5030
rect 85120 4966 85172 4972
rect 84936 4752 84988 4758
rect 84936 4694 84988 4700
rect 84844 4140 84896 4146
rect 84844 4082 84896 4088
rect 84200 4004 84252 4010
rect 84200 3946 84252 3952
rect 84856 3670 84884 4082
rect 84948 4010 84976 4694
rect 85132 4486 85160 4966
rect 85120 4480 85172 4486
rect 85120 4422 85172 4428
rect 85132 4282 85160 4422
rect 85120 4276 85172 4282
rect 85120 4218 85172 4224
rect 85500 4146 85528 6258
rect 85684 5234 85712 8842
rect 85960 7546 85988 9590
rect 86040 9036 86092 9042
rect 86040 8978 86092 8984
rect 85948 7540 86000 7546
rect 85948 7482 86000 7488
rect 86052 7410 86080 8978
rect 86144 7886 86172 11834
rect 86236 11558 86264 12174
rect 86224 11552 86276 11558
rect 86224 11494 86276 11500
rect 86236 11218 86264 11494
rect 86224 11212 86276 11218
rect 86224 11154 86276 11160
rect 86420 10062 86448 12406
rect 86512 10606 86540 13126
rect 86592 11076 86644 11082
rect 86696 11064 86724 13262
rect 86788 12782 86816 14350
rect 86972 14074 87000 14350
rect 86960 14068 87012 14074
rect 86960 14010 87012 14016
rect 86868 12844 86920 12850
rect 86972 12832 87000 14010
rect 87788 13252 87840 13258
rect 87788 13194 87840 13200
rect 87800 12986 87828 13194
rect 87788 12980 87840 12986
rect 87788 12922 87840 12928
rect 86920 12804 87000 12832
rect 87788 12844 87840 12850
rect 86868 12786 86920 12792
rect 87788 12786 87840 12792
rect 86776 12776 86828 12782
rect 86880 12753 86908 12786
rect 86776 12718 86828 12724
rect 86866 12744 86922 12753
rect 86644 11036 86724 11064
rect 86592 11018 86644 11024
rect 86500 10600 86552 10606
rect 86500 10542 86552 10548
rect 86408 10056 86460 10062
rect 86408 9998 86460 10004
rect 86132 7880 86184 7886
rect 86132 7822 86184 7828
rect 86040 7404 86092 7410
rect 86040 7346 86092 7352
rect 85764 6316 85816 6322
rect 85764 6258 85816 6264
rect 85776 6225 85804 6258
rect 85762 6216 85818 6225
rect 85762 6151 85818 6160
rect 85776 6118 85804 6151
rect 85764 6112 85816 6118
rect 85764 6054 85816 6060
rect 86052 5574 86080 7346
rect 86144 6254 86172 7822
rect 86132 6248 86184 6254
rect 86132 6190 86184 6196
rect 86144 5846 86172 6190
rect 86420 5914 86448 9998
rect 86500 9376 86552 9382
rect 86500 9318 86552 9324
rect 86592 9376 86644 9382
rect 86592 9318 86644 9324
rect 86512 8974 86540 9318
rect 86604 9178 86632 9318
rect 86592 9172 86644 9178
rect 86592 9114 86644 9120
rect 86500 8968 86552 8974
rect 86500 8910 86552 8916
rect 86684 8288 86736 8294
rect 86684 8230 86736 8236
rect 86696 8022 86724 8230
rect 86684 8016 86736 8022
rect 86684 7958 86736 7964
rect 86590 7576 86646 7585
rect 86590 7511 86592 7520
rect 86644 7511 86646 7520
rect 86592 7482 86644 7488
rect 86696 6798 86724 7958
rect 86684 6792 86736 6798
rect 86684 6734 86736 6740
rect 86408 5908 86460 5914
rect 86408 5850 86460 5856
rect 86132 5840 86184 5846
rect 86132 5782 86184 5788
rect 86040 5568 86092 5574
rect 86040 5510 86092 5516
rect 85672 5228 85724 5234
rect 85672 5170 85724 5176
rect 85488 4140 85540 4146
rect 85488 4082 85540 4088
rect 84936 4004 84988 4010
rect 84936 3946 84988 3952
rect 84844 3664 84896 3670
rect 84844 3606 84896 3612
rect 83648 3596 83700 3602
rect 83648 3538 83700 3544
rect 84948 3534 84976 3946
rect 85684 3602 85712 5170
rect 85856 4752 85908 4758
rect 85856 4694 85908 4700
rect 85868 4622 85896 4694
rect 85856 4616 85908 4622
rect 85856 4558 85908 4564
rect 86052 3738 86080 5510
rect 86144 4146 86172 5782
rect 86592 5772 86644 5778
rect 86592 5714 86644 5720
rect 86604 5234 86632 5714
rect 86592 5228 86644 5234
rect 86592 5170 86644 5176
rect 86604 4622 86632 5170
rect 86684 4684 86736 4690
rect 86788 4672 86816 12718
rect 86866 12679 86922 12688
rect 87800 12442 87828 12786
rect 87788 12436 87840 12442
rect 87788 12378 87840 12384
rect 86960 12096 87012 12102
rect 86960 12038 87012 12044
rect 86972 11694 87000 12038
rect 86960 11688 87012 11694
rect 86960 11630 87012 11636
rect 87696 11688 87748 11694
rect 87696 11630 87748 11636
rect 87708 11354 87736 11630
rect 87696 11348 87748 11354
rect 87696 11290 87748 11296
rect 86868 11212 86920 11218
rect 86868 11154 86920 11160
rect 86880 11014 86908 11154
rect 86868 11008 86920 11014
rect 86868 10950 86920 10956
rect 87892 10198 87920 16662
rect 92572 16584 92624 16590
rect 92572 16526 92624 16532
rect 92584 16250 92612 16526
rect 94697 16348 95005 16357
rect 94697 16346 94703 16348
rect 94759 16346 94783 16348
rect 94839 16346 94863 16348
rect 94919 16346 94943 16348
rect 94999 16346 95005 16348
rect 94759 16294 94761 16346
rect 94941 16294 94943 16346
rect 94697 16292 94703 16294
rect 94759 16292 94783 16294
rect 94839 16292 94863 16294
rect 94919 16292 94943 16294
rect 94999 16292 95005 16294
rect 94697 16283 95005 16292
rect 92572 16244 92624 16250
rect 92572 16186 92624 16192
rect 88248 15360 88300 15366
rect 88248 15302 88300 15308
rect 88984 15360 89036 15366
rect 88984 15302 89036 15308
rect 88260 14414 88288 15302
rect 88524 14544 88576 14550
rect 88524 14486 88576 14492
rect 88248 14408 88300 14414
rect 88248 14350 88300 14356
rect 88156 14272 88208 14278
rect 88156 14214 88208 14220
rect 88168 14113 88196 14214
rect 88154 14104 88210 14113
rect 88260 14074 88288 14350
rect 88154 14039 88210 14048
rect 88248 14068 88300 14074
rect 88248 14010 88300 14016
rect 87972 13864 88024 13870
rect 87972 13806 88024 13812
rect 87984 11694 88012 13806
rect 87972 11688 88024 11694
rect 87972 11630 88024 11636
rect 88156 11076 88208 11082
rect 88156 11018 88208 11024
rect 87880 10192 87932 10198
rect 87880 10134 87932 10140
rect 87788 10056 87840 10062
rect 87788 9998 87840 10004
rect 87696 9920 87748 9926
rect 87696 9862 87748 9868
rect 87708 9518 87736 9862
rect 87800 9654 87828 9998
rect 87788 9648 87840 9654
rect 87788 9590 87840 9596
rect 87236 9512 87288 9518
rect 87236 9454 87288 9460
rect 87696 9512 87748 9518
rect 87696 9454 87748 9460
rect 87248 9110 87276 9454
rect 87236 9104 87288 9110
rect 87236 9046 87288 9052
rect 87708 8974 87736 9454
rect 88064 9376 88116 9382
rect 88064 9318 88116 9324
rect 88076 9178 88104 9318
rect 88064 9172 88116 9178
rect 88064 9114 88116 9120
rect 88168 9042 88196 11018
rect 88536 10062 88564 14486
rect 88996 13870 89024 15302
rect 94697 15260 95005 15269
rect 94697 15258 94703 15260
rect 94759 15258 94783 15260
rect 94839 15258 94863 15260
rect 94919 15258 94943 15260
rect 94999 15258 95005 15260
rect 94759 15206 94761 15258
rect 94941 15206 94943 15258
rect 94697 15204 94703 15206
rect 94759 15204 94783 15206
rect 94839 15204 94863 15206
rect 94919 15204 94943 15206
rect 94999 15204 95005 15206
rect 94697 15195 95005 15204
rect 92664 14884 92716 14890
rect 92664 14826 92716 14832
rect 89076 14816 89128 14822
rect 89076 14758 89128 14764
rect 90456 14816 90508 14822
rect 90456 14758 90508 14764
rect 88984 13864 89036 13870
rect 88984 13806 89036 13812
rect 88996 13530 89024 13806
rect 88984 13524 89036 13530
rect 88984 13466 89036 13472
rect 88996 11694 89024 13466
rect 89088 13326 89116 14758
rect 89352 14408 89404 14414
rect 89352 14350 89404 14356
rect 89260 14340 89312 14346
rect 89260 14282 89312 14288
rect 89272 14006 89300 14282
rect 89260 14000 89312 14006
rect 89260 13942 89312 13948
rect 89364 13530 89392 14350
rect 89536 14272 89588 14278
rect 89536 14214 89588 14220
rect 89352 13524 89404 13530
rect 89352 13466 89404 13472
rect 89076 13320 89128 13326
rect 89076 13262 89128 13268
rect 89088 12782 89116 13262
rect 89364 12918 89392 13466
rect 89444 13252 89496 13258
rect 89444 13194 89496 13200
rect 89352 12912 89404 12918
rect 89456 12889 89484 13194
rect 89352 12854 89404 12860
rect 89442 12880 89498 12889
rect 89548 12850 89576 14214
rect 89812 14000 89864 14006
rect 89812 13942 89864 13948
rect 89824 13530 89852 13942
rect 89812 13524 89864 13530
rect 89812 13466 89864 13472
rect 89442 12815 89444 12824
rect 89496 12815 89498 12824
rect 89536 12844 89588 12850
rect 89444 12786 89496 12792
rect 89536 12786 89588 12792
rect 89076 12776 89128 12782
rect 89076 12718 89128 12724
rect 89088 11778 89116 12718
rect 89548 12238 89576 12786
rect 89628 12708 89680 12714
rect 89628 12650 89680 12656
rect 89536 12232 89588 12238
rect 89536 12174 89588 12180
rect 89168 12096 89220 12102
rect 89168 12038 89220 12044
rect 89180 11898 89208 12038
rect 89168 11892 89220 11898
rect 89168 11834 89220 11840
rect 89088 11762 89208 11778
rect 89088 11756 89220 11762
rect 89088 11750 89168 11756
rect 89168 11698 89220 11704
rect 88984 11688 89036 11694
rect 88984 11630 89036 11636
rect 89180 10674 89208 11698
rect 89640 11082 89668 12650
rect 90180 12640 90232 12646
rect 90180 12582 90232 12588
rect 89720 11620 89772 11626
rect 89720 11562 89772 11568
rect 89628 11076 89680 11082
rect 89628 11018 89680 11024
rect 88984 10668 89036 10674
rect 88984 10610 89036 10616
rect 89168 10668 89220 10674
rect 89168 10610 89220 10616
rect 88524 10056 88576 10062
rect 88524 9998 88576 10004
rect 88248 9580 88300 9586
rect 88248 9522 88300 9528
rect 88260 9382 88288 9522
rect 88248 9376 88300 9382
rect 88248 9318 88300 9324
rect 88156 9036 88208 9042
rect 88156 8978 88208 8984
rect 87696 8968 87748 8974
rect 87696 8910 87748 8916
rect 87880 8968 87932 8974
rect 87880 8910 87932 8916
rect 87236 7744 87288 7750
rect 87236 7686 87288 7692
rect 87144 7336 87196 7342
rect 87144 7278 87196 7284
rect 87156 6934 87184 7278
rect 87144 6928 87196 6934
rect 87144 6870 87196 6876
rect 87248 6866 87276 7686
rect 87892 6905 87920 8910
rect 88260 7041 88288 9318
rect 88432 9172 88484 9178
rect 88432 9114 88484 9120
rect 88444 9042 88472 9114
rect 88432 9036 88484 9042
rect 88432 8978 88484 8984
rect 88996 8634 89024 10610
rect 89732 9518 89760 11562
rect 89904 11008 89956 11014
rect 89904 10950 89956 10956
rect 89916 10742 89944 10950
rect 89904 10736 89956 10742
rect 89904 10678 89956 10684
rect 89812 10056 89864 10062
rect 89812 9998 89864 10004
rect 89720 9512 89772 9518
rect 89720 9454 89772 9460
rect 89824 9042 89852 9998
rect 89812 9036 89864 9042
rect 89812 8978 89864 8984
rect 89444 8968 89496 8974
rect 89444 8910 89496 8916
rect 89168 8832 89220 8838
rect 89168 8774 89220 8780
rect 88984 8628 89036 8634
rect 88984 8570 89036 8576
rect 88340 8560 88392 8566
rect 88340 8502 88392 8508
rect 88352 7478 88380 8502
rect 88432 7812 88484 7818
rect 88432 7754 88484 7760
rect 88340 7472 88392 7478
rect 88340 7414 88392 7420
rect 88444 7410 88472 7754
rect 89180 7478 89208 8774
rect 89260 8492 89312 8498
rect 89260 8434 89312 8440
rect 89272 7818 89300 8434
rect 89456 8430 89484 8910
rect 90192 8906 90220 12582
rect 90468 11150 90496 14758
rect 92676 14618 92704 14826
rect 92664 14612 92716 14618
rect 92664 14554 92716 14560
rect 91100 14272 91152 14278
rect 91100 14214 91152 14220
rect 92480 14272 92532 14278
rect 92480 14214 92532 14220
rect 90732 13932 90784 13938
rect 90732 13874 90784 13880
rect 90548 13728 90600 13734
rect 90548 13670 90600 13676
rect 90560 13326 90588 13670
rect 90548 13320 90600 13326
rect 90548 13262 90600 13268
rect 90560 12850 90588 13262
rect 90548 12844 90600 12850
rect 90548 12786 90600 12792
rect 90548 11824 90600 11830
rect 90548 11766 90600 11772
rect 90560 11354 90588 11766
rect 90548 11348 90600 11354
rect 90548 11290 90600 11296
rect 90456 11144 90508 11150
rect 90456 11086 90508 11092
rect 90468 10062 90496 11086
rect 90640 10736 90692 10742
rect 90640 10678 90692 10684
rect 90652 10266 90680 10678
rect 90744 10606 90772 13874
rect 91112 12170 91140 14214
rect 92492 13410 92520 14214
rect 92676 13938 92704 14554
rect 94697 14172 95005 14181
rect 94697 14170 94703 14172
rect 94759 14170 94783 14172
rect 94839 14170 94863 14172
rect 94919 14170 94943 14172
rect 94999 14170 95005 14172
rect 94759 14118 94761 14170
rect 94941 14118 94943 14170
rect 94697 14116 94703 14118
rect 94759 14116 94783 14118
rect 94839 14116 94863 14118
rect 94919 14116 94943 14118
rect 94999 14116 95005 14118
rect 94697 14107 95005 14116
rect 94044 14068 94096 14074
rect 94044 14010 94096 14016
rect 92664 13932 92716 13938
rect 92664 13874 92716 13880
rect 92664 13728 92716 13734
rect 92664 13670 92716 13676
rect 92492 13394 92612 13410
rect 92492 13388 92624 13394
rect 92492 13382 92572 13388
rect 92492 13297 92520 13382
rect 92572 13330 92624 13336
rect 92478 13288 92534 13297
rect 92676 13274 92704 13670
rect 92478 13223 92534 13232
rect 92584 13246 92704 13274
rect 93308 13252 93360 13258
rect 92584 13190 92612 13246
rect 93308 13194 93360 13200
rect 91836 13184 91888 13190
rect 91836 13126 91888 13132
rect 92572 13184 92624 13190
rect 92572 13126 92624 13132
rect 91100 12164 91152 12170
rect 91100 12106 91152 12112
rect 91112 11558 91140 12106
rect 91100 11552 91152 11558
rect 91100 11494 91152 11500
rect 91848 11354 91876 13126
rect 92480 12912 92532 12918
rect 92480 12854 92532 12860
rect 92112 12776 92164 12782
rect 92112 12718 92164 12724
rect 92124 11762 92152 12718
rect 92492 12306 92520 12854
rect 92584 12850 92612 13126
rect 93320 12986 93348 13194
rect 93308 12980 93360 12986
rect 93308 12922 93360 12928
rect 92572 12844 92624 12850
rect 92572 12786 92624 12792
rect 93308 12844 93360 12850
rect 93308 12786 93360 12792
rect 92940 12640 92992 12646
rect 92940 12582 92992 12588
rect 92480 12300 92532 12306
rect 92480 12242 92532 12248
rect 92112 11756 92164 11762
rect 92112 11698 92164 11704
rect 92296 11756 92348 11762
rect 92296 11698 92348 11704
rect 91836 11348 91888 11354
rect 91836 11290 91888 11296
rect 92124 10810 92152 11698
rect 92308 11354 92336 11698
rect 92480 11688 92532 11694
rect 92480 11630 92532 11636
rect 92296 11348 92348 11354
rect 92296 11290 92348 11296
rect 92492 11014 92520 11630
rect 92480 11008 92532 11014
rect 92480 10950 92532 10956
rect 92112 10804 92164 10810
rect 92112 10746 92164 10752
rect 92492 10606 92520 10950
rect 90732 10600 90784 10606
rect 90732 10542 90784 10548
rect 92480 10600 92532 10606
rect 92480 10542 92532 10548
rect 90640 10260 90692 10266
rect 90640 10202 90692 10208
rect 90456 10056 90508 10062
rect 90456 9998 90508 10004
rect 90732 9988 90784 9994
rect 90732 9930 90784 9936
rect 91100 9988 91152 9994
rect 91100 9930 91152 9936
rect 90640 9512 90692 9518
rect 90640 9454 90692 9460
rect 90180 8900 90232 8906
rect 90180 8842 90232 8848
rect 89720 8492 89772 8498
rect 89720 8434 89772 8440
rect 89444 8424 89496 8430
rect 89444 8366 89496 8372
rect 89456 7954 89484 8366
rect 89444 7948 89496 7954
rect 89444 7890 89496 7896
rect 89732 7886 89760 8434
rect 90180 8424 90232 8430
rect 90180 8366 90232 8372
rect 89812 8288 89864 8294
rect 89812 8230 89864 8236
rect 89720 7880 89772 7886
rect 89720 7822 89772 7828
rect 89260 7812 89312 7818
rect 89260 7754 89312 7760
rect 89628 7812 89680 7818
rect 89628 7754 89680 7760
rect 89168 7472 89220 7478
rect 89168 7414 89220 7420
rect 88432 7404 88484 7410
rect 88432 7346 88484 7352
rect 88246 7032 88302 7041
rect 88444 7002 88472 7346
rect 88892 7336 88944 7342
rect 88892 7278 88944 7284
rect 88246 6967 88302 6976
rect 88432 6996 88484 7002
rect 87972 6928 88024 6934
rect 87878 6896 87934 6905
rect 87236 6860 87288 6866
rect 87972 6870 88024 6876
rect 87878 6831 87934 6840
rect 87236 6802 87288 6808
rect 86960 6792 87012 6798
rect 86960 6734 87012 6740
rect 87420 6792 87472 6798
rect 87420 6734 87472 6740
rect 86972 6662 87000 6734
rect 86960 6656 87012 6662
rect 86960 6598 87012 6604
rect 87052 6656 87104 6662
rect 87052 6598 87104 6604
rect 87064 6390 87092 6598
rect 87052 6384 87104 6390
rect 87052 6326 87104 6332
rect 87432 6322 87460 6734
rect 86868 6316 86920 6322
rect 86868 6258 86920 6264
rect 87420 6316 87472 6322
rect 87420 6258 87472 6264
rect 86880 6225 86908 6258
rect 86866 6216 86922 6225
rect 86866 6151 86922 6160
rect 87604 6112 87656 6118
rect 87604 6054 87656 6060
rect 87696 6112 87748 6118
rect 87696 6054 87748 6060
rect 87616 5914 87644 6054
rect 87604 5908 87656 5914
rect 87604 5850 87656 5856
rect 87236 5840 87288 5846
rect 87236 5782 87288 5788
rect 86960 5704 87012 5710
rect 86960 5646 87012 5652
rect 86972 5370 87000 5646
rect 87248 5574 87276 5782
rect 87708 5692 87736 6054
rect 87984 5778 88012 6870
rect 88260 6866 88288 6967
rect 88432 6938 88484 6944
rect 88248 6860 88300 6866
rect 88248 6802 88300 6808
rect 88444 6322 88472 6938
rect 88904 6730 88932 7278
rect 89076 7268 89128 7274
rect 89076 7210 89128 7216
rect 89088 6798 89116 7210
rect 89442 6896 89498 6905
rect 89442 6831 89444 6840
rect 89496 6831 89498 6840
rect 89444 6802 89496 6808
rect 89640 6798 89668 7754
rect 89732 7274 89760 7822
rect 89720 7268 89772 7274
rect 89720 7210 89772 7216
rect 89824 7206 89852 8230
rect 90192 7342 90220 8366
rect 90456 7880 90508 7886
rect 90456 7822 90508 7828
rect 90468 7478 90496 7822
rect 90456 7472 90508 7478
rect 90456 7414 90508 7420
rect 90180 7336 90232 7342
rect 90180 7278 90232 7284
rect 89812 7200 89864 7206
rect 89812 7142 89864 7148
rect 89720 6996 89772 7002
rect 89720 6938 89772 6944
rect 89076 6792 89128 6798
rect 89076 6734 89128 6740
rect 89628 6792 89680 6798
rect 89628 6734 89680 6740
rect 88892 6724 88944 6730
rect 88892 6666 88944 6672
rect 88432 6316 88484 6322
rect 88432 6258 88484 6264
rect 88904 6254 88932 6666
rect 88892 6248 88944 6254
rect 88892 6190 88944 6196
rect 89732 5778 89760 6938
rect 89824 6934 89852 7142
rect 89902 7032 89958 7041
rect 90192 7002 90220 7278
rect 89902 6967 89958 6976
rect 90180 6996 90232 7002
rect 89812 6928 89864 6934
rect 89812 6870 89864 6876
rect 89824 5914 89852 6870
rect 89916 6798 89944 6967
rect 90180 6938 90232 6944
rect 89904 6792 89956 6798
rect 89904 6734 89956 6740
rect 89904 6248 89956 6254
rect 89904 6190 89956 6196
rect 89812 5908 89864 5914
rect 89812 5850 89864 5856
rect 87972 5772 88024 5778
rect 87972 5714 88024 5720
rect 89720 5772 89772 5778
rect 89720 5714 89772 5720
rect 87788 5704 87840 5710
rect 87708 5664 87788 5692
rect 87144 5568 87196 5574
rect 87144 5510 87196 5516
rect 87236 5568 87288 5574
rect 87236 5510 87288 5516
rect 86960 5364 87012 5370
rect 86960 5306 87012 5312
rect 86736 4644 86816 4672
rect 86684 4626 86736 4632
rect 86592 4616 86644 4622
rect 86592 4558 86644 4564
rect 86972 4146 87000 5306
rect 87052 5024 87104 5030
rect 87052 4966 87104 4972
rect 87064 4826 87092 4966
rect 87156 4826 87184 5510
rect 87708 5370 87736 5664
rect 87788 5646 87840 5652
rect 87696 5364 87748 5370
rect 87696 5306 87748 5312
rect 87708 5234 87736 5306
rect 87696 5228 87748 5234
rect 87696 5170 87748 5176
rect 87052 4820 87104 4826
rect 87052 4762 87104 4768
rect 87144 4820 87196 4826
rect 87144 4762 87196 4768
rect 87052 4480 87104 4486
rect 87052 4422 87104 4428
rect 86132 4140 86184 4146
rect 86132 4082 86184 4088
rect 86960 4140 87012 4146
rect 86960 4082 87012 4088
rect 86040 3732 86092 3738
rect 86040 3674 86092 3680
rect 85672 3596 85724 3602
rect 85672 3538 85724 3544
rect 84936 3528 84988 3534
rect 84936 3470 84988 3476
rect 84948 3194 84976 3470
rect 84936 3188 84988 3194
rect 84936 3130 84988 3136
rect 85684 3058 85712 3538
rect 85672 3052 85724 3058
rect 85672 2994 85724 3000
rect 86144 2990 86172 4082
rect 87064 3534 87092 4422
rect 87156 4282 87184 4762
rect 87708 4622 87736 5170
rect 87880 5024 87932 5030
rect 87984 5012 88012 5714
rect 89352 5704 89404 5710
rect 89352 5646 89404 5652
rect 89364 5030 89392 5646
rect 89916 5642 89944 6190
rect 89904 5636 89956 5642
rect 89904 5578 89956 5584
rect 87932 4984 88012 5012
rect 87880 4966 87932 4972
rect 87236 4616 87288 4622
rect 87236 4558 87288 4564
rect 87696 4616 87748 4622
rect 87696 4558 87748 4564
rect 87144 4276 87196 4282
rect 87144 4218 87196 4224
rect 87248 4146 87276 4558
rect 87984 4146 88012 4984
rect 88064 5024 88116 5030
rect 88064 4966 88116 4972
rect 88984 5024 89036 5030
rect 88984 4966 89036 4972
rect 89352 5024 89404 5030
rect 89352 4966 89404 4972
rect 88076 4826 88104 4966
rect 88064 4820 88116 4826
rect 88064 4762 88116 4768
rect 88524 4684 88576 4690
rect 88524 4626 88576 4632
rect 87236 4140 87288 4146
rect 87236 4082 87288 4088
rect 87972 4140 88024 4146
rect 87972 4082 88024 4088
rect 87248 3670 87276 4082
rect 88536 3738 88564 4626
rect 88616 4616 88668 4622
rect 88616 4558 88668 4564
rect 88628 4214 88656 4558
rect 88892 4548 88944 4554
rect 88892 4490 88944 4496
rect 88616 4208 88668 4214
rect 88616 4150 88668 4156
rect 88524 3732 88576 3738
rect 88524 3674 88576 3680
rect 87236 3664 87288 3670
rect 87236 3606 87288 3612
rect 88904 3602 88932 4490
rect 88996 3942 89024 4966
rect 89628 4548 89680 4554
rect 89628 4490 89680 4496
rect 89812 4548 89864 4554
rect 89812 4490 89864 4496
rect 89352 4480 89404 4486
rect 89352 4422 89404 4428
rect 89076 4004 89128 4010
rect 89076 3946 89128 3952
rect 88984 3936 89036 3942
rect 88984 3878 89036 3884
rect 88996 3670 89024 3878
rect 88984 3664 89036 3670
rect 88984 3606 89036 3612
rect 88892 3596 88944 3602
rect 88892 3538 88944 3544
rect 89088 3534 89116 3946
rect 89364 3602 89392 4422
rect 89640 4078 89668 4490
rect 89824 4214 89852 4490
rect 89812 4208 89864 4214
rect 89812 4150 89864 4156
rect 89628 4072 89680 4078
rect 89628 4014 89680 4020
rect 89352 3596 89404 3602
rect 89352 3538 89404 3544
rect 87052 3528 87104 3534
rect 87052 3470 87104 3476
rect 89076 3528 89128 3534
rect 89076 3470 89128 3476
rect 86868 3460 86920 3466
rect 86868 3402 86920 3408
rect 86880 3194 86908 3402
rect 86868 3188 86920 3194
rect 86868 3130 86920 3136
rect 81716 2984 81768 2990
rect 81716 2926 81768 2932
rect 83372 2984 83424 2990
rect 83372 2926 83424 2932
rect 86132 2984 86184 2990
rect 86132 2926 86184 2932
rect 82979 2748 83287 2757
rect 82979 2746 82985 2748
rect 83041 2746 83065 2748
rect 83121 2746 83145 2748
rect 83201 2746 83225 2748
rect 83281 2746 83287 2748
rect 83041 2694 83043 2746
rect 83223 2694 83225 2746
rect 82979 2692 82985 2694
rect 83041 2692 83065 2694
rect 83121 2692 83145 2694
rect 83201 2692 83225 2694
rect 83281 2692 83287 2694
rect 82979 2683 83287 2692
rect 86880 2650 86908 3130
rect 89088 2990 89116 3470
rect 89640 3126 89668 4014
rect 89916 4010 89944 5578
rect 90652 5370 90680 9454
rect 90744 7750 90772 9930
rect 91112 9382 91140 9930
rect 91192 9648 91244 9654
rect 91244 9596 91324 9602
rect 91192 9590 91324 9596
rect 91204 9574 91324 9590
rect 91296 9382 91324 9574
rect 92848 9580 92900 9586
rect 92848 9522 92900 9528
rect 91100 9376 91152 9382
rect 91100 9318 91152 9324
rect 91284 9376 91336 9382
rect 91284 9318 91336 9324
rect 92388 9376 92440 9382
rect 92388 9318 92440 9324
rect 92480 9376 92532 9382
rect 92480 9318 92532 9324
rect 91284 8968 91336 8974
rect 91284 8910 91336 8916
rect 91008 8832 91060 8838
rect 91008 8774 91060 8780
rect 91020 8430 91048 8774
rect 91008 8424 91060 8430
rect 91008 8366 91060 8372
rect 90824 7812 90876 7818
rect 90824 7754 90876 7760
rect 90732 7744 90784 7750
rect 90732 7686 90784 7692
rect 90744 6934 90772 7686
rect 90732 6928 90784 6934
rect 90732 6870 90784 6876
rect 90744 6662 90772 6870
rect 90732 6656 90784 6662
rect 90732 6598 90784 6604
rect 90836 6322 90864 7754
rect 91020 7410 91048 8366
rect 91192 8356 91244 8362
rect 91192 8298 91244 8304
rect 91204 7954 91232 8298
rect 91192 7948 91244 7954
rect 91192 7890 91244 7896
rect 91008 7404 91060 7410
rect 91008 7346 91060 7352
rect 90824 6316 90876 6322
rect 90824 6258 90876 6264
rect 90640 5364 90692 5370
rect 90640 5306 90692 5312
rect 90836 4706 90864 6258
rect 91020 6118 91048 7346
rect 91296 6322 91324 8910
rect 92400 6866 92428 9318
rect 92492 7954 92520 9318
rect 92860 8090 92888 9522
rect 92848 8084 92900 8090
rect 92848 8026 92900 8032
rect 92480 7948 92532 7954
rect 92480 7890 92532 7896
rect 92860 7546 92888 8026
rect 92848 7540 92900 7546
rect 92848 7482 92900 7488
rect 92756 7200 92808 7206
rect 92756 7142 92808 7148
rect 92388 6860 92440 6866
rect 92388 6802 92440 6808
rect 92768 6662 92796 7142
rect 92860 7002 92888 7482
rect 92952 7410 92980 12582
rect 93320 12442 93348 12786
rect 93308 12436 93360 12442
rect 93308 12378 93360 12384
rect 94056 12238 94084 14010
rect 94136 13728 94188 13734
rect 94136 13670 94188 13676
rect 94044 12232 94096 12238
rect 94044 12174 94096 12180
rect 93308 11756 93360 11762
rect 93308 11698 93360 11704
rect 93320 11354 93348 11698
rect 93400 11688 93452 11694
rect 93400 11630 93452 11636
rect 93308 11348 93360 11354
rect 93308 11290 93360 11296
rect 93320 10674 93348 11290
rect 93308 10668 93360 10674
rect 93308 10610 93360 10616
rect 93216 10600 93268 10606
rect 93216 10542 93268 10548
rect 93228 9042 93256 10542
rect 93216 9036 93268 9042
rect 93216 8978 93268 8984
rect 93124 8900 93176 8906
rect 93124 8842 93176 8848
rect 93032 7812 93084 7818
rect 93032 7754 93084 7760
rect 93044 7478 93072 7754
rect 93032 7472 93084 7478
rect 93032 7414 93084 7420
rect 92940 7404 92992 7410
rect 92940 7346 92992 7352
rect 92848 6996 92900 7002
rect 92848 6938 92900 6944
rect 92756 6656 92808 6662
rect 92756 6598 92808 6604
rect 91836 6384 91888 6390
rect 91836 6326 91888 6332
rect 91284 6316 91336 6322
rect 91284 6258 91336 6264
rect 91008 6112 91060 6118
rect 91008 6054 91060 6060
rect 91296 5778 91324 6258
rect 91848 6118 91876 6326
rect 92768 6118 92796 6598
rect 93044 6322 93072 7414
rect 93136 6730 93164 8842
rect 93412 8566 93440 11630
rect 93768 11144 93820 11150
rect 93768 11086 93820 11092
rect 93780 11014 93808 11086
rect 93768 11008 93820 11014
rect 93768 10950 93820 10956
rect 94148 10674 94176 13670
rect 94697 13084 95005 13093
rect 94697 13082 94703 13084
rect 94759 13082 94783 13084
rect 94839 13082 94863 13084
rect 94919 13082 94943 13084
rect 94999 13082 95005 13084
rect 94759 13030 94761 13082
rect 94941 13030 94943 13082
rect 94697 13028 94703 13030
rect 94759 13028 94783 13030
rect 94839 13028 94863 13030
rect 94919 13028 94943 13030
rect 94999 13028 95005 13030
rect 94697 13019 95005 13028
rect 94226 12472 94282 12481
rect 94226 12407 94228 12416
rect 94280 12407 94282 12416
rect 94228 12378 94280 12384
rect 94697 11996 95005 12005
rect 94697 11994 94703 11996
rect 94759 11994 94783 11996
rect 94839 11994 94863 11996
rect 94919 11994 94943 11996
rect 94999 11994 95005 11996
rect 94759 11942 94761 11994
rect 94941 11942 94943 11994
rect 94697 11940 94703 11942
rect 94759 11940 94783 11942
rect 94839 11940 94863 11942
rect 94919 11940 94943 11942
rect 94999 11940 95005 11942
rect 94697 11931 95005 11940
rect 94228 11076 94280 11082
rect 94228 11018 94280 11024
rect 94240 10810 94268 11018
rect 94697 10908 95005 10917
rect 94697 10906 94703 10908
rect 94759 10906 94783 10908
rect 94839 10906 94863 10908
rect 94919 10906 94943 10908
rect 94999 10906 95005 10908
rect 94759 10854 94761 10906
rect 94941 10854 94943 10906
rect 94697 10852 94703 10854
rect 94759 10852 94783 10854
rect 94839 10852 94863 10854
rect 94919 10852 94943 10854
rect 94999 10852 95005 10854
rect 94697 10843 95005 10852
rect 94228 10804 94280 10810
rect 94228 10746 94280 10752
rect 94136 10668 94188 10674
rect 94136 10610 94188 10616
rect 94148 10146 94176 10610
rect 93860 10124 93912 10130
rect 93860 10066 93912 10072
rect 94056 10118 94176 10146
rect 93768 9920 93820 9926
rect 93768 9862 93820 9868
rect 93780 9654 93808 9862
rect 93768 9648 93820 9654
rect 93768 9590 93820 9596
rect 93872 8974 93900 10066
rect 94056 9586 94084 10118
rect 94136 10056 94188 10062
rect 94136 9998 94188 10004
rect 94044 9580 94096 9586
rect 94044 9522 94096 9528
rect 93952 9512 94004 9518
rect 93952 9454 94004 9460
rect 93964 9178 93992 9454
rect 93952 9172 94004 9178
rect 93952 9114 94004 9120
rect 93860 8968 93912 8974
rect 93860 8910 93912 8916
rect 93400 8560 93452 8566
rect 93400 8502 93452 8508
rect 93584 8424 93636 8430
rect 93584 8366 93636 8372
rect 93596 8090 93624 8366
rect 93584 8084 93636 8090
rect 93584 8026 93636 8032
rect 93400 7880 93452 7886
rect 93400 7822 93452 7828
rect 93124 6724 93176 6730
rect 93124 6666 93176 6672
rect 93032 6316 93084 6322
rect 93032 6258 93084 6264
rect 91836 6112 91888 6118
rect 91836 6054 91888 6060
rect 92756 6112 92808 6118
rect 92756 6054 92808 6060
rect 91284 5772 91336 5778
rect 91284 5714 91336 5720
rect 91008 5364 91060 5370
rect 91008 5306 91060 5312
rect 91020 5030 91048 5306
rect 91296 5166 91324 5714
rect 91848 5710 91876 6054
rect 92768 5846 92796 6054
rect 92756 5840 92808 5846
rect 92756 5782 92808 5788
rect 91836 5704 91888 5710
rect 91836 5646 91888 5652
rect 91848 5370 91876 5646
rect 91836 5364 91888 5370
rect 91836 5306 91888 5312
rect 92020 5296 92072 5302
rect 92020 5238 92072 5244
rect 91284 5160 91336 5166
rect 91284 5102 91336 5108
rect 91008 5024 91060 5030
rect 91008 4966 91060 4972
rect 90836 4678 91048 4706
rect 90824 4616 90876 4622
rect 90824 4558 90876 4564
rect 90272 4480 90324 4486
rect 90272 4422 90324 4428
rect 90284 4282 90312 4422
rect 90272 4276 90324 4282
rect 90272 4218 90324 4224
rect 89996 4140 90048 4146
rect 89996 4082 90048 4088
rect 89904 4004 89956 4010
rect 89904 3946 89956 3952
rect 89916 3466 89944 3946
rect 90008 3738 90036 4082
rect 89996 3732 90048 3738
rect 89996 3674 90048 3680
rect 89904 3460 89956 3466
rect 89904 3402 89956 3408
rect 90836 3194 90864 4558
rect 90916 4480 90968 4486
rect 90916 4422 90968 4428
rect 90928 3738 90956 4422
rect 91020 3942 91048 4678
rect 92032 4622 92060 5238
rect 93044 5234 93072 6258
rect 93136 5914 93164 6666
rect 93214 6352 93270 6361
rect 93214 6287 93270 6296
rect 93124 5908 93176 5914
rect 93124 5850 93176 5856
rect 93228 5710 93256 6287
rect 93412 5914 93440 7822
rect 93768 6996 93820 7002
rect 93768 6938 93820 6944
rect 93780 5914 93808 6938
rect 93872 6798 93900 8910
rect 94056 6866 94084 9522
rect 94148 9110 94176 9998
rect 94228 9988 94280 9994
rect 94228 9930 94280 9936
rect 94240 9654 94268 9930
rect 94697 9820 95005 9829
rect 94697 9818 94703 9820
rect 94759 9818 94783 9820
rect 94839 9818 94863 9820
rect 94919 9818 94943 9820
rect 94999 9818 95005 9820
rect 94759 9766 94761 9818
rect 94941 9766 94943 9818
rect 94697 9764 94703 9766
rect 94759 9764 94783 9766
rect 94839 9764 94863 9766
rect 94919 9764 94943 9766
rect 94999 9764 95005 9766
rect 94697 9755 95005 9764
rect 94228 9648 94280 9654
rect 94228 9590 94280 9596
rect 94136 9104 94188 9110
rect 94136 9046 94188 9052
rect 94148 8362 94176 9046
rect 94697 8732 95005 8741
rect 94697 8730 94703 8732
rect 94759 8730 94783 8732
rect 94839 8730 94863 8732
rect 94919 8730 94943 8732
rect 94999 8730 95005 8732
rect 94759 8678 94761 8730
rect 94941 8678 94943 8730
rect 94697 8676 94703 8678
rect 94759 8676 94783 8678
rect 94839 8676 94863 8678
rect 94919 8676 94943 8678
rect 94999 8676 95005 8678
rect 94697 8667 95005 8676
rect 94136 8356 94188 8362
rect 94136 8298 94188 8304
rect 94044 6860 94096 6866
rect 94044 6802 94096 6808
rect 93860 6792 93912 6798
rect 93860 6734 93912 6740
rect 93400 5908 93452 5914
rect 93400 5850 93452 5856
rect 93768 5908 93820 5914
rect 93768 5850 93820 5856
rect 93216 5704 93268 5710
rect 93216 5646 93268 5652
rect 92388 5228 92440 5234
rect 92388 5170 92440 5176
rect 93032 5228 93084 5234
rect 93032 5170 93084 5176
rect 92020 4616 92072 4622
rect 92020 4558 92072 4564
rect 92032 4298 92060 4558
rect 92112 4548 92164 4554
rect 92296 4548 92348 4554
rect 92164 4508 92296 4536
rect 92112 4490 92164 4496
rect 92296 4490 92348 4496
rect 91940 4282 92060 4298
rect 91928 4276 92060 4282
rect 91980 4270 92060 4276
rect 91928 4218 91980 4224
rect 91008 3936 91060 3942
rect 91008 3878 91060 3884
rect 90916 3732 90968 3738
rect 90916 3674 90968 3680
rect 91020 3194 91048 3878
rect 91928 3528 91980 3534
rect 91928 3470 91980 3476
rect 90824 3188 90876 3194
rect 90824 3130 90876 3136
rect 91008 3188 91060 3194
rect 91008 3130 91060 3136
rect 89628 3120 89680 3126
rect 89628 3062 89680 3068
rect 91020 2990 91048 3130
rect 91940 2990 91968 3470
rect 92400 3194 92428 5170
rect 93124 4480 93176 4486
rect 93124 4422 93176 4428
rect 93136 4078 93164 4422
rect 93124 4072 93176 4078
rect 93124 4014 93176 4020
rect 93228 3738 93256 5646
rect 94056 5370 94084 6802
rect 94148 6458 94176 8298
rect 95148 7744 95200 7750
rect 95148 7686 95200 7692
rect 94697 7644 95005 7653
rect 94697 7642 94703 7644
rect 94759 7642 94783 7644
rect 94839 7642 94863 7644
rect 94919 7642 94943 7644
rect 94999 7642 95005 7644
rect 94759 7590 94761 7642
rect 94941 7590 94943 7642
rect 94697 7588 94703 7590
rect 94759 7588 94783 7590
rect 94839 7588 94863 7590
rect 94919 7588 94943 7590
rect 94999 7588 95005 7590
rect 94697 7579 95005 7588
rect 95160 7585 95188 7686
rect 95146 7576 95202 7585
rect 95146 7511 95202 7520
rect 94697 6556 95005 6565
rect 94697 6554 94703 6556
rect 94759 6554 94783 6556
rect 94839 6554 94863 6556
rect 94919 6554 94943 6556
rect 94999 6554 95005 6556
rect 94759 6502 94761 6554
rect 94941 6502 94943 6554
rect 94697 6500 94703 6502
rect 94759 6500 94783 6502
rect 94839 6500 94863 6502
rect 94919 6500 94943 6502
rect 94999 6500 95005 6502
rect 94697 6491 95005 6500
rect 94136 6452 94188 6458
rect 94136 6394 94188 6400
rect 94697 5468 95005 5477
rect 94697 5466 94703 5468
rect 94759 5466 94783 5468
rect 94839 5466 94863 5468
rect 94919 5466 94943 5468
rect 94999 5466 95005 5468
rect 94759 5414 94761 5466
rect 94941 5414 94943 5466
rect 94697 5412 94703 5414
rect 94759 5412 94783 5414
rect 94839 5412 94863 5414
rect 94919 5412 94943 5414
rect 94999 5412 95005 5414
rect 94697 5403 95005 5412
rect 93676 5364 93728 5370
rect 93676 5306 93728 5312
rect 94044 5364 94096 5370
rect 94044 5306 94096 5312
rect 93688 4486 93716 5306
rect 93676 4480 93728 4486
rect 93676 4422 93728 4428
rect 94228 4480 94280 4486
rect 94228 4422 94280 4428
rect 93216 3732 93268 3738
rect 93216 3674 93268 3680
rect 93688 3670 93716 4422
rect 94240 4078 94268 4422
rect 94697 4380 95005 4389
rect 94697 4378 94703 4380
rect 94759 4378 94783 4380
rect 94839 4378 94863 4380
rect 94919 4378 94943 4380
rect 94999 4378 95005 4380
rect 94759 4326 94761 4378
rect 94941 4326 94943 4378
rect 94697 4324 94703 4326
rect 94759 4324 94783 4326
rect 94839 4324 94863 4326
rect 94919 4324 94943 4326
rect 94999 4324 95005 4326
rect 94697 4315 95005 4324
rect 94228 4072 94280 4078
rect 94228 4014 94280 4020
rect 93676 3664 93728 3670
rect 93676 3606 93728 3612
rect 93768 3392 93820 3398
rect 93768 3334 93820 3340
rect 92388 3188 92440 3194
rect 92388 3130 92440 3136
rect 89076 2984 89128 2990
rect 89076 2926 89128 2932
rect 91008 2984 91060 2990
rect 91008 2926 91060 2932
rect 91928 2984 91980 2990
rect 91928 2926 91980 2932
rect 91020 2774 91048 2926
rect 90928 2746 91048 2774
rect 90928 2650 90956 2746
rect 93780 2689 93808 3334
rect 94697 3292 95005 3301
rect 94697 3290 94703 3292
rect 94759 3290 94783 3292
rect 94839 3290 94863 3292
rect 94919 3290 94943 3292
rect 94999 3290 95005 3292
rect 94759 3238 94761 3290
rect 94941 3238 94943 3290
rect 94697 3236 94703 3238
rect 94759 3236 94783 3238
rect 94839 3236 94863 3238
rect 94919 3236 94943 3238
rect 94999 3236 95005 3238
rect 94697 3227 95005 3236
rect 93766 2680 93822 2689
rect 75276 2644 75328 2650
rect 75276 2586 75328 2592
rect 78588 2644 78720 2650
rect 78640 2638 78720 2644
rect 78772 2644 78824 2650
rect 78588 2586 78640 2592
rect 78772 2586 78824 2592
rect 86868 2644 86920 2650
rect 86868 2586 86920 2592
rect 90916 2644 90968 2650
rect 93766 2615 93822 2624
rect 90916 2586 90968 2592
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 28448 2440 28500 2446
rect 28448 2382 28500 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 56324 2440 56376 2446
rect 56324 2382 56376 2388
rect 68376 2440 68428 2446
rect 68376 2382 68428 2388
rect 74816 2440 74868 2446
rect 74816 2382 74868 2388
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 20352 2304 20404 2310
rect 20352 2246 20404 2252
rect 28172 2304 28224 2310
rect 28172 2246 28224 2252
rect 4448 800 4476 2246
rect 12360 800 12388 2246
rect 20364 1170 20392 2246
rect 24386 2204 24694 2213
rect 24386 2202 24392 2204
rect 24448 2202 24472 2204
rect 24528 2202 24552 2204
rect 24608 2202 24632 2204
rect 24688 2202 24694 2204
rect 24448 2150 24450 2202
rect 24630 2150 24632 2202
rect 24386 2148 24392 2150
rect 24448 2148 24472 2150
rect 24528 2148 24552 2150
rect 24608 2148 24632 2150
rect 24688 2148 24694 2150
rect 24386 2139 24694 2148
rect 20272 1142 20392 1170
rect 20272 800 20300 1142
rect 28184 800 28212 2246
rect 36096 800 36124 2382
rect 75288 2378 75316 2586
rect 91468 2440 91520 2446
rect 91468 2382 91520 2388
rect 75276 2372 75328 2378
rect 75276 2314 75328 2320
rect 43996 2304 44048 2310
rect 43996 2246 44048 2252
rect 51908 2304 51960 2310
rect 51908 2246 51960 2252
rect 59820 2304 59872 2310
rect 59820 2246 59872 2252
rect 67732 2304 67784 2310
rect 67732 2246 67784 2252
rect 75644 2304 75696 2310
rect 75644 2246 75696 2252
rect 83556 2304 83608 2310
rect 83556 2246 83608 2252
rect 44008 800 44036 2246
rect 47823 2204 48131 2213
rect 47823 2202 47829 2204
rect 47885 2202 47909 2204
rect 47965 2202 47989 2204
rect 48045 2202 48069 2204
rect 48125 2202 48131 2204
rect 47885 2150 47887 2202
rect 48067 2150 48069 2202
rect 47823 2148 47829 2150
rect 47885 2148 47909 2150
rect 47965 2148 47989 2150
rect 48045 2148 48069 2150
rect 48125 2148 48131 2150
rect 47823 2139 48131 2148
rect 51920 800 51948 2246
rect 59832 800 59860 2246
rect 67744 800 67772 2246
rect 71260 2204 71568 2213
rect 71260 2202 71266 2204
rect 71322 2202 71346 2204
rect 71402 2202 71426 2204
rect 71482 2202 71506 2204
rect 71562 2202 71568 2204
rect 71322 2150 71324 2202
rect 71504 2150 71506 2202
rect 71260 2148 71266 2150
rect 71322 2148 71346 2150
rect 71402 2148 71426 2150
rect 71482 2148 71506 2150
rect 71562 2148 71568 2150
rect 71260 2139 71568 2148
rect 75656 800 75684 2246
rect 83568 800 83596 2246
rect 91480 800 91508 2382
rect 94697 2204 95005 2213
rect 94697 2202 94703 2204
rect 94759 2202 94783 2204
rect 94839 2202 94863 2204
rect 94919 2202 94943 2204
rect 94999 2202 95005 2204
rect 94759 2150 94761 2202
rect 94941 2150 94943 2202
rect 94697 2148 94703 2150
rect 94759 2148 94783 2150
rect 94839 2148 94863 2150
rect 94919 2148 94943 2150
rect 94999 2148 95005 2150
rect 94697 2139 95005 2148
rect 4434 0 4490 800
rect 12346 0 12402 800
rect 20258 0 20314 800
rect 28170 0 28226 800
rect 36082 0 36138 800
rect 43994 0 44050 800
rect 51906 0 51962 800
rect 59818 0 59874 800
rect 67730 0 67786 800
rect 75642 0 75698 800
rect 83554 0 83610 800
rect 91466 0 91522 800
<< via2 >>
rect 1582 16668 1584 16688
rect 1584 16668 1636 16688
rect 1636 16668 1638 16688
rect 1582 16632 1638 16668
rect 4802 13368 4858 13424
rect 1582 10004 1584 10024
rect 1584 10004 1636 10024
rect 1636 10004 1638 10024
rect 1582 9968 1638 10004
rect 7010 12724 7012 12744
rect 7012 12724 7064 12744
rect 7064 12724 7066 12744
rect 7010 12688 7066 12724
rect 8666 11600 8722 11656
rect 8482 11212 8538 11248
rect 8482 11192 8484 11212
rect 8484 11192 8536 11212
rect 8536 11192 8538 11212
rect 4066 3304 4122 3360
rect 12674 16890 12730 16892
rect 12754 16890 12810 16892
rect 12834 16890 12890 16892
rect 12914 16890 12970 16892
rect 12674 16838 12720 16890
rect 12720 16838 12730 16890
rect 12754 16838 12784 16890
rect 12784 16838 12796 16890
rect 12796 16838 12810 16890
rect 12834 16838 12848 16890
rect 12848 16838 12860 16890
rect 12860 16838 12890 16890
rect 12914 16838 12924 16890
rect 12924 16838 12970 16890
rect 12674 16836 12730 16838
rect 12754 16836 12810 16838
rect 12834 16836 12890 16838
rect 12914 16836 12970 16838
rect 20350 15988 20352 16008
rect 20352 15988 20404 16008
rect 20404 15988 20406 16008
rect 12674 15802 12730 15804
rect 12754 15802 12810 15804
rect 12834 15802 12890 15804
rect 12914 15802 12970 15804
rect 12674 15750 12720 15802
rect 12720 15750 12730 15802
rect 12754 15750 12784 15802
rect 12784 15750 12796 15802
rect 12796 15750 12810 15802
rect 12834 15750 12848 15802
rect 12848 15750 12860 15802
rect 12860 15750 12890 15802
rect 12914 15750 12924 15802
rect 12924 15750 12970 15802
rect 12674 15748 12730 15750
rect 12754 15748 12810 15750
rect 12834 15748 12890 15750
rect 12914 15748 12970 15750
rect 13910 15000 13966 15056
rect 12714 14884 12770 14920
rect 12714 14864 12716 14884
rect 12716 14864 12768 14884
rect 12768 14864 12770 14884
rect 12674 14714 12730 14716
rect 12754 14714 12810 14716
rect 12834 14714 12890 14716
rect 12914 14714 12970 14716
rect 12674 14662 12720 14714
rect 12720 14662 12730 14714
rect 12754 14662 12784 14714
rect 12784 14662 12796 14714
rect 12796 14662 12810 14714
rect 12834 14662 12848 14714
rect 12848 14662 12860 14714
rect 12860 14662 12890 14714
rect 12914 14662 12924 14714
rect 12924 14662 12970 14714
rect 12674 14660 12730 14662
rect 12754 14660 12810 14662
rect 12834 14660 12890 14662
rect 12914 14660 12970 14662
rect 13082 14340 13138 14376
rect 13082 14320 13084 14340
rect 13084 14320 13136 14340
rect 13136 14320 13138 14340
rect 13174 14048 13230 14104
rect 11978 13812 11980 13832
rect 11980 13812 12032 13832
rect 12032 13812 12034 13832
rect 11978 13776 12034 13812
rect 12674 13626 12730 13628
rect 12754 13626 12810 13628
rect 12834 13626 12890 13628
rect 12914 13626 12970 13628
rect 12674 13574 12720 13626
rect 12720 13574 12730 13626
rect 12754 13574 12784 13626
rect 12784 13574 12796 13626
rect 12796 13574 12810 13626
rect 12834 13574 12848 13626
rect 12848 13574 12860 13626
rect 12860 13574 12890 13626
rect 12914 13574 12924 13626
rect 12924 13574 12970 13626
rect 12674 13572 12730 13574
rect 12754 13572 12810 13574
rect 12834 13572 12890 13574
rect 12914 13572 12970 13574
rect 11886 10648 11942 10704
rect 9402 5072 9458 5128
rect 12674 12538 12730 12540
rect 12754 12538 12810 12540
rect 12834 12538 12890 12540
rect 12914 12538 12970 12540
rect 12674 12486 12720 12538
rect 12720 12486 12730 12538
rect 12754 12486 12784 12538
rect 12784 12486 12796 12538
rect 12796 12486 12810 12538
rect 12834 12486 12848 12538
rect 12848 12486 12860 12538
rect 12860 12486 12890 12538
rect 12914 12486 12924 12538
rect 12924 12486 12970 12538
rect 12674 12484 12730 12486
rect 12754 12484 12810 12486
rect 12834 12484 12890 12486
rect 12914 12484 12970 12486
rect 12990 11872 13046 11928
rect 12674 11450 12730 11452
rect 12754 11450 12810 11452
rect 12834 11450 12890 11452
rect 12914 11450 12970 11452
rect 12674 11398 12720 11450
rect 12720 11398 12730 11450
rect 12754 11398 12784 11450
rect 12784 11398 12796 11450
rect 12796 11398 12810 11450
rect 12834 11398 12848 11450
rect 12848 11398 12860 11450
rect 12860 11398 12890 11450
rect 12914 11398 12924 11450
rect 12924 11398 12970 11450
rect 12674 11396 12730 11398
rect 12754 11396 12810 11398
rect 12834 11396 12890 11398
rect 12914 11396 12970 11398
rect 12674 10362 12730 10364
rect 12754 10362 12810 10364
rect 12834 10362 12890 10364
rect 12914 10362 12970 10364
rect 12674 10310 12720 10362
rect 12720 10310 12730 10362
rect 12754 10310 12784 10362
rect 12784 10310 12796 10362
rect 12796 10310 12810 10362
rect 12834 10310 12848 10362
rect 12848 10310 12860 10362
rect 12860 10310 12890 10362
rect 12914 10310 12924 10362
rect 12924 10310 12970 10362
rect 12674 10308 12730 10310
rect 12754 10308 12810 10310
rect 12834 10308 12890 10310
rect 12914 10308 12970 10310
rect 12674 9274 12730 9276
rect 12754 9274 12810 9276
rect 12834 9274 12890 9276
rect 12914 9274 12970 9276
rect 12674 9222 12720 9274
rect 12720 9222 12730 9274
rect 12754 9222 12784 9274
rect 12784 9222 12796 9274
rect 12796 9222 12810 9274
rect 12834 9222 12848 9274
rect 12848 9222 12860 9274
rect 12860 9222 12890 9274
rect 12914 9222 12924 9274
rect 12924 9222 12970 9274
rect 12674 9220 12730 9222
rect 12754 9220 12810 9222
rect 12834 9220 12890 9222
rect 12914 9220 12970 9222
rect 12674 8186 12730 8188
rect 12754 8186 12810 8188
rect 12834 8186 12890 8188
rect 12914 8186 12970 8188
rect 12674 8134 12720 8186
rect 12720 8134 12730 8186
rect 12754 8134 12784 8186
rect 12784 8134 12796 8186
rect 12796 8134 12810 8186
rect 12834 8134 12848 8186
rect 12848 8134 12860 8186
rect 12860 8134 12890 8186
rect 12914 8134 12924 8186
rect 12924 8134 12970 8186
rect 12674 8132 12730 8134
rect 12754 8132 12810 8134
rect 12834 8132 12890 8134
rect 12914 8132 12970 8134
rect 20350 15952 20406 15988
rect 16946 15544 17002 15600
rect 15014 13912 15070 13968
rect 15382 11872 15438 11928
rect 14554 9444 14610 9480
rect 14554 9424 14556 9444
rect 14556 9424 14608 9444
rect 14608 9424 14610 9444
rect 13450 7928 13506 7984
rect 13174 7812 13230 7848
rect 13174 7792 13176 7812
rect 13176 7792 13228 7812
rect 13228 7792 13230 7812
rect 10874 4120 10930 4176
rect 12674 7098 12730 7100
rect 12754 7098 12810 7100
rect 12834 7098 12890 7100
rect 12914 7098 12970 7100
rect 12674 7046 12720 7098
rect 12720 7046 12730 7098
rect 12754 7046 12784 7098
rect 12784 7046 12796 7098
rect 12796 7046 12810 7098
rect 12834 7046 12848 7098
rect 12848 7046 12860 7098
rect 12860 7046 12890 7098
rect 12914 7046 12924 7098
rect 12924 7046 12970 7098
rect 12674 7044 12730 7046
rect 12754 7044 12810 7046
rect 12834 7044 12890 7046
rect 12914 7044 12970 7046
rect 12674 6010 12730 6012
rect 12754 6010 12810 6012
rect 12834 6010 12890 6012
rect 12914 6010 12970 6012
rect 12674 5958 12720 6010
rect 12720 5958 12730 6010
rect 12754 5958 12784 6010
rect 12784 5958 12796 6010
rect 12796 5958 12810 6010
rect 12834 5958 12848 6010
rect 12848 5958 12860 6010
rect 12860 5958 12890 6010
rect 12914 5958 12924 6010
rect 12924 5958 12970 6010
rect 12674 5956 12730 5958
rect 12754 5956 12810 5958
rect 12834 5956 12890 5958
rect 12914 5956 12970 5958
rect 12674 4922 12730 4924
rect 12754 4922 12810 4924
rect 12834 4922 12890 4924
rect 12914 4922 12970 4924
rect 12674 4870 12720 4922
rect 12720 4870 12730 4922
rect 12754 4870 12784 4922
rect 12784 4870 12796 4922
rect 12796 4870 12810 4922
rect 12834 4870 12848 4922
rect 12848 4870 12860 4922
rect 12860 4870 12890 4922
rect 12914 4870 12924 4922
rect 12924 4870 12970 4922
rect 12674 4868 12730 4870
rect 12754 4868 12810 4870
rect 12834 4868 12890 4870
rect 12914 4868 12970 4870
rect 15106 10240 15162 10296
rect 20442 13640 20498 13696
rect 16670 8336 16726 8392
rect 17130 8608 17186 8664
rect 17406 8472 17462 8528
rect 17682 8744 17738 8800
rect 17590 8356 17646 8392
rect 17590 8336 17592 8356
rect 17592 8336 17644 8356
rect 17644 8336 17646 8356
rect 18326 8744 18382 8800
rect 19338 11464 19394 11520
rect 19338 11092 19340 11112
rect 19340 11092 19392 11112
rect 19392 11092 19394 11112
rect 19338 11056 19394 11092
rect 19338 10956 19346 10976
rect 19346 10956 19394 10976
rect 19338 10920 19394 10956
rect 18694 9016 18750 9072
rect 19890 11328 19946 11384
rect 19798 10956 19800 10976
rect 19800 10956 19852 10976
rect 19852 10956 19854 10976
rect 19798 10920 19854 10956
rect 20718 9968 20774 10024
rect 19706 9696 19762 9752
rect 19890 9016 19946 9072
rect 20442 8608 20498 8664
rect 20626 8916 20628 8936
rect 20628 8916 20680 8936
rect 20680 8916 20682 8936
rect 20626 8880 20682 8916
rect 20718 8472 20774 8528
rect 20074 8336 20130 8392
rect 24392 17434 24448 17436
rect 24472 17434 24528 17436
rect 24552 17434 24608 17436
rect 24632 17434 24688 17436
rect 24392 17382 24438 17434
rect 24438 17382 24448 17434
rect 24472 17382 24502 17434
rect 24502 17382 24514 17434
rect 24514 17382 24528 17434
rect 24552 17382 24566 17434
rect 24566 17382 24578 17434
rect 24578 17382 24608 17434
rect 24632 17382 24642 17434
rect 24642 17382 24688 17434
rect 24392 17380 24448 17382
rect 24472 17380 24528 17382
rect 24552 17380 24608 17382
rect 24632 17380 24688 17382
rect 22098 13232 22154 13288
rect 24214 14048 24270 14104
rect 24392 16346 24448 16348
rect 24472 16346 24528 16348
rect 24552 16346 24608 16348
rect 24632 16346 24688 16348
rect 24392 16294 24438 16346
rect 24438 16294 24448 16346
rect 24472 16294 24502 16346
rect 24502 16294 24514 16346
rect 24514 16294 24528 16346
rect 24552 16294 24566 16346
rect 24566 16294 24578 16346
rect 24578 16294 24608 16346
rect 24632 16294 24642 16346
rect 24642 16294 24688 16346
rect 24392 16292 24448 16294
rect 24472 16292 24528 16294
rect 24552 16292 24608 16294
rect 24632 16292 24688 16294
rect 24392 15258 24448 15260
rect 24472 15258 24528 15260
rect 24552 15258 24608 15260
rect 24632 15258 24688 15260
rect 24392 15206 24438 15258
rect 24438 15206 24448 15258
rect 24472 15206 24502 15258
rect 24502 15206 24514 15258
rect 24514 15206 24528 15258
rect 24552 15206 24566 15258
rect 24566 15206 24578 15258
rect 24578 15206 24608 15258
rect 24632 15206 24642 15258
rect 24642 15206 24688 15258
rect 24392 15204 24448 15206
rect 24472 15204 24528 15206
rect 24552 15204 24608 15206
rect 24632 15204 24688 15206
rect 25594 14728 25650 14784
rect 24392 14170 24448 14172
rect 24472 14170 24528 14172
rect 24552 14170 24608 14172
rect 24632 14170 24688 14172
rect 24392 14118 24438 14170
rect 24438 14118 24448 14170
rect 24472 14118 24502 14170
rect 24502 14118 24514 14170
rect 24514 14118 24528 14170
rect 24552 14118 24566 14170
rect 24566 14118 24578 14170
rect 24578 14118 24608 14170
rect 24632 14118 24642 14170
rect 24642 14118 24688 14170
rect 24392 14116 24448 14118
rect 24472 14116 24528 14118
rect 24552 14116 24608 14118
rect 24632 14116 24688 14118
rect 24766 14048 24822 14104
rect 24392 13082 24448 13084
rect 24472 13082 24528 13084
rect 24552 13082 24608 13084
rect 24632 13082 24688 13084
rect 24392 13030 24438 13082
rect 24438 13030 24448 13082
rect 24472 13030 24502 13082
rect 24502 13030 24514 13082
rect 24514 13030 24528 13082
rect 24552 13030 24566 13082
rect 24566 13030 24578 13082
rect 24578 13030 24608 13082
rect 24632 13030 24642 13082
rect 24642 13030 24688 13082
rect 24392 13028 24448 13030
rect 24472 13028 24528 13030
rect 24552 13028 24608 13030
rect 24632 13028 24688 13030
rect 22558 11772 22560 11792
rect 22560 11772 22612 11792
rect 22612 11772 22614 11792
rect 22558 11736 22614 11772
rect 24030 12316 24032 12336
rect 24032 12316 24084 12336
rect 24084 12316 24086 12336
rect 24030 12280 24086 12316
rect 24392 11994 24448 11996
rect 24472 11994 24528 11996
rect 24552 11994 24608 11996
rect 24632 11994 24688 11996
rect 24392 11942 24438 11994
rect 24438 11942 24448 11994
rect 24472 11942 24502 11994
rect 24502 11942 24514 11994
rect 24514 11942 24528 11994
rect 24552 11942 24566 11994
rect 24566 11942 24578 11994
rect 24578 11942 24608 11994
rect 24632 11942 24642 11994
rect 24642 11942 24688 11994
rect 24392 11940 24448 11942
rect 24472 11940 24528 11942
rect 24552 11940 24608 11942
rect 24632 11940 24688 11942
rect 25410 11872 25466 11928
rect 22558 10376 22614 10432
rect 22006 10124 22062 10160
rect 22006 10104 22008 10124
rect 22008 10104 22060 10124
rect 22060 10104 22062 10124
rect 21914 9324 21916 9344
rect 21916 9324 21968 9344
rect 21968 9324 21970 9344
rect 21914 9288 21970 9324
rect 22190 9288 22246 9344
rect 21638 8744 21694 8800
rect 21454 8508 21456 8528
rect 21456 8508 21508 8528
rect 21508 8508 21510 8528
rect 21454 8472 21510 8508
rect 21914 8336 21970 8392
rect 20994 7420 20996 7440
rect 20996 7420 21048 7440
rect 21048 7420 21050 7440
rect 20994 7384 21050 7420
rect 22926 11076 22982 11112
rect 22926 11056 22928 11076
rect 22928 11056 22980 11076
rect 22980 11056 22982 11076
rect 24306 11056 24362 11112
rect 24392 10906 24448 10908
rect 24472 10906 24528 10908
rect 24552 10906 24608 10908
rect 24632 10906 24688 10908
rect 24392 10854 24438 10906
rect 24438 10854 24448 10906
rect 24472 10854 24502 10906
rect 24502 10854 24514 10906
rect 24514 10854 24528 10906
rect 24552 10854 24566 10906
rect 24566 10854 24578 10906
rect 24578 10854 24608 10906
rect 24632 10854 24642 10906
rect 24642 10854 24688 10906
rect 24392 10852 24448 10854
rect 24472 10852 24528 10854
rect 24552 10852 24608 10854
rect 24632 10852 24688 10854
rect 23938 10512 23994 10568
rect 24392 9818 24448 9820
rect 24472 9818 24528 9820
rect 24552 9818 24608 9820
rect 24632 9818 24688 9820
rect 24392 9766 24438 9818
rect 24438 9766 24448 9818
rect 24472 9766 24502 9818
rect 24502 9766 24514 9818
rect 24514 9766 24528 9818
rect 24552 9766 24566 9818
rect 24566 9766 24578 9818
rect 24578 9766 24608 9818
rect 24632 9766 24642 9818
rect 24642 9766 24688 9818
rect 24392 9764 24448 9766
rect 24472 9764 24528 9766
rect 24552 9764 24608 9766
rect 24632 9764 24688 9766
rect 23570 9696 23626 9752
rect 23386 9596 23388 9616
rect 23388 9596 23440 9616
rect 23440 9596 23442 9616
rect 23386 9560 23442 9596
rect 23386 9424 23442 9480
rect 23570 9424 23626 9480
rect 22650 8880 22706 8936
rect 22558 8744 22614 8800
rect 23202 9152 23258 9208
rect 23110 7284 23112 7304
rect 23112 7284 23164 7304
rect 23164 7284 23166 7304
rect 23110 7248 23166 7284
rect 19890 5908 19946 5944
rect 19890 5888 19892 5908
rect 19892 5888 19944 5908
rect 19944 5888 19946 5908
rect 24392 8730 24448 8732
rect 24472 8730 24528 8732
rect 24552 8730 24608 8732
rect 24632 8730 24688 8732
rect 24392 8678 24438 8730
rect 24438 8678 24448 8730
rect 24472 8678 24502 8730
rect 24502 8678 24514 8730
rect 24514 8678 24528 8730
rect 24552 8678 24566 8730
rect 24566 8678 24578 8730
rect 24578 8678 24608 8730
rect 24632 8678 24642 8730
rect 24642 8678 24688 8730
rect 24392 8676 24448 8678
rect 24472 8676 24528 8678
rect 24552 8676 24608 8678
rect 24632 8676 24688 8678
rect 23754 8492 23810 8528
rect 23754 8472 23756 8492
rect 23756 8472 23808 8492
rect 23808 8472 23810 8492
rect 24392 7642 24448 7644
rect 24472 7642 24528 7644
rect 24552 7642 24608 7644
rect 24632 7642 24688 7644
rect 24392 7590 24438 7642
rect 24438 7590 24448 7642
rect 24472 7590 24502 7642
rect 24502 7590 24514 7642
rect 24514 7590 24528 7642
rect 24552 7590 24566 7642
rect 24566 7590 24578 7642
rect 24578 7590 24608 7642
rect 24632 7590 24642 7642
rect 24642 7590 24688 7642
rect 24392 7588 24448 7590
rect 24472 7588 24528 7590
rect 24552 7588 24608 7590
rect 24632 7588 24688 7590
rect 23662 7148 23664 7168
rect 23664 7148 23716 7168
rect 23716 7148 23718 7168
rect 23662 7112 23718 7148
rect 22926 5752 22982 5808
rect 22650 5652 22652 5672
rect 22652 5652 22704 5672
rect 22704 5652 22706 5672
rect 22650 5616 22706 5652
rect 16394 4528 16450 4584
rect 27066 12280 27122 12336
rect 27434 11872 27490 11928
rect 27526 10684 27528 10704
rect 27528 10684 27580 10704
rect 27580 10684 27582 10704
rect 27526 10648 27582 10684
rect 28262 12960 28318 13016
rect 27894 12280 27950 12336
rect 28078 11328 28134 11384
rect 28998 12144 29054 12200
rect 29550 15272 29606 15328
rect 29642 14592 29698 14648
rect 29458 14456 29514 14512
rect 29642 13504 29698 13560
rect 29826 14184 29882 14240
rect 28630 11500 28632 11520
rect 28632 11500 28684 11520
rect 28684 11500 28686 11520
rect 28630 11464 28686 11500
rect 27802 11056 27858 11112
rect 27986 11056 28042 11112
rect 26606 9444 26662 9480
rect 26606 9424 26608 9444
rect 26608 9424 26660 9444
rect 26660 9424 26662 9444
rect 27066 10376 27122 10432
rect 27066 9968 27122 10024
rect 26790 9560 26846 9616
rect 27986 10512 28042 10568
rect 29182 11464 29238 11520
rect 28906 11192 28962 11248
rect 27526 9172 27582 9208
rect 27526 9152 27528 9172
rect 27528 9152 27580 9172
rect 27580 9152 27582 9172
rect 27526 8336 27582 8392
rect 24392 6554 24448 6556
rect 24472 6554 24528 6556
rect 24552 6554 24608 6556
rect 24632 6554 24688 6556
rect 24392 6502 24438 6554
rect 24438 6502 24448 6554
rect 24472 6502 24502 6554
rect 24502 6502 24514 6554
rect 24514 6502 24528 6554
rect 24552 6502 24566 6554
rect 24566 6502 24578 6554
rect 24578 6502 24608 6554
rect 24632 6502 24642 6554
rect 24642 6502 24688 6554
rect 24392 6500 24448 6502
rect 24472 6500 24528 6502
rect 24552 6500 24608 6502
rect 24632 6500 24688 6502
rect 24766 6296 24822 6352
rect 26146 6840 26202 6896
rect 25594 6724 25650 6760
rect 25594 6704 25596 6724
rect 25596 6704 25648 6724
rect 25648 6704 25650 6724
rect 24950 5616 25006 5672
rect 24392 5466 24448 5468
rect 24472 5466 24528 5468
rect 24552 5466 24608 5468
rect 24632 5466 24688 5468
rect 24392 5414 24438 5466
rect 24438 5414 24448 5466
rect 24472 5414 24502 5466
rect 24502 5414 24514 5466
rect 24514 5414 24528 5466
rect 24552 5414 24566 5466
rect 24566 5414 24578 5466
rect 24578 5414 24608 5466
rect 24632 5414 24642 5466
rect 24642 5414 24688 5466
rect 24392 5412 24448 5414
rect 24472 5412 24528 5414
rect 24552 5412 24608 5414
rect 24632 5412 24688 5414
rect 25134 5888 25190 5944
rect 24674 4972 24676 4992
rect 24676 4972 24728 4992
rect 24728 4972 24730 4992
rect 24674 4936 24730 4972
rect 24392 4378 24448 4380
rect 24472 4378 24528 4380
rect 24552 4378 24608 4380
rect 24632 4378 24688 4380
rect 24392 4326 24438 4378
rect 24438 4326 24448 4378
rect 24472 4326 24502 4378
rect 24502 4326 24514 4378
rect 24514 4326 24528 4378
rect 24552 4326 24566 4378
rect 24566 4326 24578 4378
rect 24578 4326 24608 4378
rect 24632 4326 24642 4378
rect 24642 4326 24688 4378
rect 24392 4324 24448 4326
rect 24472 4324 24528 4326
rect 24552 4324 24608 4326
rect 24632 4324 24688 4326
rect 12674 3834 12730 3836
rect 12754 3834 12810 3836
rect 12834 3834 12890 3836
rect 12914 3834 12970 3836
rect 12674 3782 12720 3834
rect 12720 3782 12730 3834
rect 12754 3782 12784 3834
rect 12784 3782 12796 3834
rect 12796 3782 12810 3834
rect 12834 3782 12848 3834
rect 12848 3782 12860 3834
rect 12860 3782 12890 3834
rect 12914 3782 12924 3834
rect 12924 3782 12970 3834
rect 12674 3780 12730 3782
rect 12754 3780 12810 3782
rect 12834 3780 12890 3782
rect 12914 3780 12970 3782
rect 12674 2746 12730 2748
rect 12754 2746 12810 2748
rect 12834 2746 12890 2748
rect 12914 2746 12970 2748
rect 12674 2694 12720 2746
rect 12720 2694 12730 2746
rect 12754 2694 12784 2746
rect 12784 2694 12796 2746
rect 12796 2694 12810 2746
rect 12834 2694 12848 2746
rect 12848 2694 12860 2746
rect 12860 2694 12890 2746
rect 12914 2694 12924 2746
rect 12924 2694 12970 2746
rect 12674 2692 12730 2694
rect 12754 2692 12810 2694
rect 12834 2692 12890 2694
rect 12914 2692 12970 2694
rect 28998 9696 29054 9752
rect 29826 12824 29882 12880
rect 30930 13504 30986 13560
rect 31114 13096 31170 13152
rect 30194 11872 30250 11928
rect 30010 11600 30066 11656
rect 31758 14592 31814 14648
rect 29826 10376 29882 10432
rect 29458 9696 29514 9752
rect 30194 9596 30196 9616
rect 30196 9596 30248 9616
rect 30248 9596 30250 9616
rect 30194 9560 30250 9596
rect 30470 10920 30526 10976
rect 31666 10920 31722 10976
rect 26698 6876 26700 6896
rect 26700 6876 26752 6896
rect 26752 6876 26754 6896
rect 26698 6840 26754 6876
rect 26422 6332 26424 6352
rect 26424 6332 26476 6352
rect 26476 6332 26478 6352
rect 26422 6296 26478 6332
rect 27066 5772 27122 5808
rect 27066 5752 27068 5772
rect 27068 5752 27120 5772
rect 27120 5752 27122 5772
rect 30286 9424 30342 9480
rect 32126 12280 32182 12336
rect 32586 12844 32642 12880
rect 32586 12824 32588 12844
rect 32588 12824 32640 12844
rect 32640 12824 32642 12844
rect 32402 12008 32458 12064
rect 32402 10240 32458 10296
rect 32678 11192 32734 11248
rect 33414 11500 33416 11520
rect 33416 11500 33468 11520
rect 33468 11500 33470 11520
rect 33414 11464 33470 11500
rect 32954 10532 33010 10568
rect 32954 10512 32956 10532
rect 32956 10512 33008 10532
rect 33008 10512 33010 10532
rect 32586 9424 32642 9480
rect 30470 6432 30526 6488
rect 31206 6876 31208 6896
rect 31208 6876 31260 6896
rect 31260 6876 31262 6896
rect 31206 6840 31262 6876
rect 32310 6296 32366 6352
rect 28262 5244 28264 5264
rect 28264 5244 28316 5264
rect 28316 5244 28318 5264
rect 28262 5208 28318 5244
rect 26422 4936 26478 4992
rect 24392 3290 24448 3292
rect 24472 3290 24528 3292
rect 24552 3290 24608 3292
rect 24632 3290 24688 3292
rect 24392 3238 24438 3290
rect 24438 3238 24448 3290
rect 24472 3238 24502 3290
rect 24502 3238 24514 3290
rect 24514 3238 24528 3290
rect 24552 3238 24566 3290
rect 24566 3238 24578 3290
rect 24578 3238 24608 3290
rect 24632 3238 24642 3290
rect 24642 3238 24688 3290
rect 24392 3236 24448 3238
rect 24472 3236 24528 3238
rect 24552 3236 24608 3238
rect 24632 3236 24688 3238
rect 32770 5636 32826 5672
rect 32770 5616 32772 5636
rect 32772 5616 32824 5636
rect 32824 5616 32826 5636
rect 33046 9152 33102 9208
rect 33322 9424 33378 9480
rect 33046 8472 33102 8528
rect 47829 17434 47885 17436
rect 47909 17434 47965 17436
rect 47989 17434 48045 17436
rect 48069 17434 48125 17436
rect 47829 17382 47875 17434
rect 47875 17382 47885 17434
rect 47909 17382 47939 17434
rect 47939 17382 47951 17434
rect 47951 17382 47965 17434
rect 47989 17382 48003 17434
rect 48003 17382 48015 17434
rect 48015 17382 48045 17434
rect 48069 17382 48079 17434
rect 48079 17382 48125 17434
rect 47829 17380 47885 17382
rect 47909 17380 47965 17382
rect 47989 17380 48045 17382
rect 48069 17380 48125 17382
rect 36111 16890 36167 16892
rect 36191 16890 36247 16892
rect 36271 16890 36327 16892
rect 36351 16890 36407 16892
rect 36111 16838 36157 16890
rect 36157 16838 36167 16890
rect 36191 16838 36221 16890
rect 36221 16838 36233 16890
rect 36233 16838 36247 16890
rect 36271 16838 36285 16890
rect 36285 16838 36297 16890
rect 36297 16838 36327 16890
rect 36351 16838 36361 16890
rect 36361 16838 36407 16890
rect 36111 16836 36167 16838
rect 36191 16836 36247 16838
rect 36271 16836 36327 16838
rect 36351 16836 36407 16838
rect 34886 15408 34942 15464
rect 35346 15408 35402 15464
rect 34702 15272 34758 15328
rect 35070 14728 35126 14784
rect 35070 14456 35126 14512
rect 35070 10376 35126 10432
rect 34518 9832 34574 9888
rect 33690 9152 33746 9208
rect 33874 8372 33876 8392
rect 33876 8372 33928 8392
rect 33928 8372 33930 8392
rect 33874 8336 33930 8372
rect 33138 7656 33194 7712
rect 33046 6568 33102 6624
rect 34518 8900 34574 8936
rect 34518 8880 34520 8900
rect 34520 8880 34572 8900
rect 34572 8880 34574 8900
rect 34334 8608 34390 8664
rect 36111 15802 36167 15804
rect 36191 15802 36247 15804
rect 36271 15802 36327 15804
rect 36351 15802 36407 15804
rect 36111 15750 36157 15802
rect 36157 15750 36167 15802
rect 36191 15750 36221 15802
rect 36221 15750 36233 15802
rect 36233 15750 36247 15802
rect 36271 15750 36285 15802
rect 36285 15750 36297 15802
rect 36297 15750 36327 15802
rect 36351 15750 36361 15802
rect 36361 15750 36407 15802
rect 36111 15748 36167 15750
rect 36191 15748 36247 15750
rect 36271 15748 36327 15750
rect 36351 15748 36407 15750
rect 35898 15544 35954 15600
rect 35806 15272 35862 15328
rect 35622 13640 35678 13696
rect 36111 14714 36167 14716
rect 36191 14714 36247 14716
rect 36271 14714 36327 14716
rect 36351 14714 36407 14716
rect 36111 14662 36157 14714
rect 36157 14662 36167 14714
rect 36191 14662 36221 14714
rect 36221 14662 36233 14714
rect 36233 14662 36247 14714
rect 36271 14662 36285 14714
rect 36285 14662 36297 14714
rect 36297 14662 36327 14714
rect 36351 14662 36361 14714
rect 36361 14662 36407 14714
rect 36111 14660 36167 14662
rect 36191 14660 36247 14662
rect 36271 14660 36327 14662
rect 36351 14660 36407 14662
rect 37094 14184 37150 14240
rect 36111 13626 36167 13628
rect 36191 13626 36247 13628
rect 36271 13626 36327 13628
rect 36351 13626 36407 13628
rect 36111 13574 36157 13626
rect 36157 13574 36167 13626
rect 36191 13574 36221 13626
rect 36221 13574 36233 13626
rect 36233 13574 36247 13626
rect 36271 13574 36285 13626
rect 36285 13574 36297 13626
rect 36297 13574 36327 13626
rect 36351 13574 36361 13626
rect 36361 13574 36407 13626
rect 36111 13572 36167 13574
rect 36191 13572 36247 13574
rect 36271 13572 36327 13574
rect 36351 13572 36407 13574
rect 36726 13640 36782 13696
rect 35530 12844 35586 12880
rect 35530 12824 35532 12844
rect 35532 12824 35584 12844
rect 35584 12824 35586 12844
rect 36111 12538 36167 12540
rect 36191 12538 36247 12540
rect 36271 12538 36327 12540
rect 36351 12538 36407 12540
rect 36111 12486 36157 12538
rect 36157 12486 36167 12538
rect 36191 12486 36221 12538
rect 36221 12486 36233 12538
rect 36233 12486 36247 12538
rect 36271 12486 36285 12538
rect 36285 12486 36297 12538
rect 36297 12486 36327 12538
rect 36351 12486 36361 12538
rect 36361 12486 36407 12538
rect 36111 12484 36167 12486
rect 36191 12484 36247 12486
rect 36271 12484 36327 12486
rect 36351 12484 36407 12486
rect 37462 13096 37518 13152
rect 36910 12144 36966 12200
rect 35714 11500 35716 11520
rect 35716 11500 35768 11520
rect 35768 11500 35770 11520
rect 35714 11464 35770 11500
rect 36111 11450 36167 11452
rect 36191 11450 36247 11452
rect 36271 11450 36327 11452
rect 36351 11450 36407 11452
rect 36111 11398 36157 11450
rect 36157 11398 36167 11450
rect 36191 11398 36221 11450
rect 36221 11398 36233 11450
rect 36233 11398 36247 11450
rect 36271 11398 36285 11450
rect 36285 11398 36297 11450
rect 36297 11398 36327 11450
rect 36351 11398 36361 11450
rect 36361 11398 36407 11450
rect 36111 11396 36167 11398
rect 36191 11396 36247 11398
rect 36271 11396 36327 11398
rect 36351 11396 36407 11398
rect 37002 11600 37058 11656
rect 36910 11056 36966 11112
rect 36542 10920 36598 10976
rect 36542 10376 36598 10432
rect 36111 10362 36167 10364
rect 36191 10362 36247 10364
rect 36271 10362 36327 10364
rect 36351 10362 36407 10364
rect 36111 10310 36157 10362
rect 36157 10310 36167 10362
rect 36191 10310 36221 10362
rect 36221 10310 36233 10362
rect 36233 10310 36247 10362
rect 36271 10310 36285 10362
rect 36285 10310 36297 10362
rect 36297 10310 36327 10362
rect 36351 10310 36361 10362
rect 36361 10310 36407 10362
rect 36111 10308 36167 10310
rect 36191 10308 36247 10310
rect 36271 10308 36327 10310
rect 36351 10308 36407 10310
rect 34426 7792 34482 7848
rect 36634 9832 36690 9888
rect 34886 9288 34942 9344
rect 35070 9152 35126 9208
rect 34702 6976 34758 7032
rect 34702 6432 34758 6488
rect 35162 8744 35218 8800
rect 35162 7792 35218 7848
rect 36818 9696 36874 9752
rect 35714 9152 35770 9208
rect 36111 9274 36167 9276
rect 36191 9274 36247 9276
rect 36271 9274 36327 9276
rect 36351 9274 36407 9276
rect 36111 9222 36157 9274
rect 36157 9222 36167 9274
rect 36191 9222 36221 9274
rect 36221 9222 36233 9274
rect 36233 9222 36247 9274
rect 36271 9222 36285 9274
rect 36285 9222 36297 9274
rect 36297 9222 36327 9274
rect 36351 9222 36361 9274
rect 36361 9222 36407 9274
rect 36111 9220 36167 9222
rect 36191 9220 36247 9222
rect 36271 9220 36327 9222
rect 36351 9220 36407 9222
rect 35530 8744 35586 8800
rect 36111 8186 36167 8188
rect 36191 8186 36247 8188
rect 36271 8186 36327 8188
rect 36351 8186 36407 8188
rect 36111 8134 36157 8186
rect 36157 8134 36167 8186
rect 36191 8134 36221 8186
rect 36221 8134 36233 8186
rect 36233 8134 36247 8186
rect 36271 8134 36285 8186
rect 36285 8134 36297 8186
rect 36297 8134 36327 8186
rect 36351 8134 36361 8186
rect 36361 8134 36407 8186
rect 36111 8132 36167 8134
rect 36191 8132 36247 8134
rect 36271 8132 36327 8134
rect 36351 8132 36407 8134
rect 36111 7098 36167 7100
rect 36191 7098 36247 7100
rect 36271 7098 36327 7100
rect 36351 7098 36407 7100
rect 36111 7046 36157 7098
rect 36157 7046 36167 7098
rect 36191 7046 36221 7098
rect 36221 7046 36233 7098
rect 36233 7046 36247 7098
rect 36271 7046 36285 7098
rect 36285 7046 36297 7098
rect 36297 7046 36327 7098
rect 36351 7046 36361 7098
rect 36361 7046 36407 7098
rect 36111 7044 36167 7046
rect 36191 7044 36247 7046
rect 36271 7044 36327 7046
rect 36351 7044 36407 7046
rect 35898 6976 35954 7032
rect 35806 6296 35862 6352
rect 35622 6196 35624 6216
rect 35624 6196 35676 6216
rect 35676 6196 35678 6216
rect 35622 6160 35678 6196
rect 36111 6010 36167 6012
rect 36191 6010 36247 6012
rect 36271 6010 36327 6012
rect 36351 6010 36407 6012
rect 36111 5958 36157 6010
rect 36157 5958 36167 6010
rect 36191 5958 36221 6010
rect 36221 5958 36233 6010
rect 36233 5958 36247 6010
rect 36271 5958 36285 6010
rect 36285 5958 36297 6010
rect 36297 5958 36327 6010
rect 36351 5958 36361 6010
rect 36361 5958 36407 6010
rect 36111 5956 36167 5958
rect 36191 5956 36247 5958
rect 36271 5956 36327 5958
rect 36351 5956 36407 5958
rect 36542 8200 36598 8256
rect 36726 6604 36728 6624
rect 36728 6604 36780 6624
rect 36780 6604 36782 6624
rect 36726 6568 36782 6604
rect 36542 5616 36598 5672
rect 38014 12960 38070 13016
rect 37830 12280 37886 12336
rect 40774 15988 40776 16008
rect 40776 15988 40828 16008
rect 40828 15988 40830 16008
rect 40774 15952 40830 15988
rect 40774 15544 40830 15600
rect 40958 14864 41014 14920
rect 40590 14476 40646 14512
rect 40590 14456 40592 14476
rect 40592 14456 40644 14476
rect 40644 14456 40646 14476
rect 39026 12416 39082 12472
rect 38934 12164 38990 12200
rect 38934 12144 38936 12164
rect 38936 12144 38988 12164
rect 38988 12144 38990 12164
rect 38658 11872 38714 11928
rect 38842 11600 38898 11656
rect 39578 11464 39634 11520
rect 38750 11328 38806 11384
rect 37738 10648 37794 10704
rect 37094 8628 37150 8664
rect 37094 8608 37096 8628
rect 37096 8608 37148 8628
rect 37148 8608 37150 8628
rect 37738 9832 37794 9888
rect 37830 8200 37886 8256
rect 37554 6296 37610 6352
rect 38106 8472 38162 8528
rect 38106 6840 38162 6896
rect 36111 4922 36167 4924
rect 36191 4922 36247 4924
rect 36271 4922 36327 4924
rect 36351 4922 36407 4924
rect 36111 4870 36157 4922
rect 36157 4870 36167 4922
rect 36191 4870 36221 4922
rect 36221 4870 36233 4922
rect 36233 4870 36247 4922
rect 36271 4870 36285 4922
rect 36285 4870 36297 4922
rect 36297 4870 36327 4922
rect 36351 4870 36361 4922
rect 36361 4870 36407 4922
rect 36111 4868 36167 4870
rect 36191 4868 36247 4870
rect 36271 4868 36327 4870
rect 36351 4868 36407 4870
rect 34426 4664 34482 4720
rect 36111 3834 36167 3836
rect 36191 3834 36247 3836
rect 36271 3834 36327 3836
rect 36351 3834 36407 3836
rect 36111 3782 36157 3834
rect 36157 3782 36167 3834
rect 36191 3782 36221 3834
rect 36221 3782 36233 3834
rect 36233 3782 36247 3834
rect 36271 3782 36285 3834
rect 36285 3782 36297 3834
rect 36297 3782 36327 3834
rect 36351 3782 36361 3834
rect 36361 3782 36407 3834
rect 36111 3780 36167 3782
rect 36191 3780 36247 3782
rect 36271 3780 36327 3782
rect 36351 3780 36407 3782
rect 38474 9016 38530 9072
rect 38842 9288 38898 9344
rect 38750 9016 38806 9072
rect 38934 9016 38990 9072
rect 38842 8880 38898 8936
rect 38566 6160 38622 6216
rect 40590 12552 40646 12608
rect 40222 11464 40278 11520
rect 40130 11056 40186 11112
rect 40498 10920 40554 10976
rect 41234 14592 41290 14648
rect 41418 14184 41474 14240
rect 42338 16496 42394 16552
rect 42246 14048 42302 14104
rect 41786 13096 41842 13152
rect 42430 15000 42486 15056
rect 41602 12008 41658 12064
rect 41418 11600 41474 11656
rect 39302 9696 39358 9752
rect 41142 10240 41198 10296
rect 39670 9016 39726 9072
rect 40222 9444 40278 9480
rect 40222 9424 40224 9444
rect 40224 9424 40276 9444
rect 40276 9424 40278 9444
rect 41142 9832 41198 9888
rect 41326 9832 41382 9888
rect 41234 9460 41236 9480
rect 41236 9460 41288 9480
rect 41288 9460 41290 9480
rect 40498 8608 40554 8664
rect 40774 8492 40830 8528
rect 40774 8472 40776 8492
rect 40776 8472 40828 8492
rect 40828 8472 40830 8492
rect 40406 8064 40462 8120
rect 40590 7112 40646 7168
rect 41234 9424 41290 9460
rect 41234 9172 41290 9208
rect 41234 9152 41236 9172
rect 41236 9152 41288 9172
rect 41288 9152 41290 9172
rect 41602 11328 41658 11384
rect 42338 12280 42394 12336
rect 44638 16088 44694 16144
rect 42890 13252 42946 13288
rect 42890 13232 42892 13252
rect 42892 13232 42944 13252
rect 42944 13232 42946 13252
rect 41786 11328 41842 11384
rect 42154 10920 42210 10976
rect 41786 10784 41842 10840
rect 42062 10260 42118 10296
rect 42062 10240 42064 10260
rect 42064 10240 42116 10260
rect 42116 10240 42118 10260
rect 42614 11736 42670 11792
rect 42890 11464 42946 11520
rect 44086 15680 44142 15736
rect 43810 14592 43866 14648
rect 43902 12008 43958 12064
rect 43994 11328 44050 11384
rect 44546 12164 44602 12200
rect 44546 12144 44548 12164
rect 44548 12144 44600 12164
rect 44600 12144 44602 12164
rect 46110 16496 46166 16552
rect 45742 13640 45798 13696
rect 44362 10240 44418 10296
rect 42706 9696 42762 9752
rect 41602 9152 41658 9208
rect 42430 8628 42486 8664
rect 42430 8608 42432 8628
rect 42432 8608 42484 8628
rect 42484 8608 42486 8628
rect 38198 4528 38254 4584
rect 42614 7656 42670 7712
rect 41878 7112 41934 7168
rect 42430 6704 42486 6760
rect 43442 9036 43498 9072
rect 43442 9016 43444 9036
rect 43444 9016 43496 9036
rect 43496 9016 43498 9036
rect 44822 9832 44878 9888
rect 43074 5344 43130 5400
rect 42982 4936 43038 4992
rect 45190 9832 45246 9888
rect 45006 9560 45062 9616
rect 45098 9424 45154 9480
rect 45466 8064 45522 8120
rect 45650 8084 45706 8120
rect 45650 8064 45652 8084
rect 45652 8064 45704 8084
rect 45704 8064 45706 8084
rect 45190 7792 45246 7848
rect 44178 5344 44234 5400
rect 47829 16346 47885 16348
rect 47909 16346 47965 16348
rect 47989 16346 48045 16348
rect 48069 16346 48125 16348
rect 47829 16294 47875 16346
rect 47875 16294 47885 16346
rect 47909 16294 47939 16346
rect 47939 16294 47951 16346
rect 47951 16294 47965 16346
rect 47989 16294 48003 16346
rect 48003 16294 48015 16346
rect 48015 16294 48045 16346
rect 48069 16294 48079 16346
rect 48079 16294 48125 16346
rect 47829 16292 47885 16294
rect 47909 16292 47965 16294
rect 47989 16292 48045 16294
rect 48069 16292 48125 16294
rect 47950 15680 48006 15736
rect 47829 15258 47885 15260
rect 47909 15258 47965 15260
rect 47989 15258 48045 15260
rect 48069 15258 48125 15260
rect 47829 15206 47875 15258
rect 47875 15206 47885 15258
rect 47909 15206 47939 15258
rect 47939 15206 47951 15258
rect 47951 15206 47965 15258
rect 47989 15206 48003 15258
rect 48003 15206 48015 15258
rect 48015 15206 48045 15258
rect 48069 15206 48079 15258
rect 48079 15206 48125 15258
rect 47829 15204 47885 15206
rect 47909 15204 47965 15206
rect 47989 15204 48045 15206
rect 48069 15204 48125 15206
rect 47030 14184 47086 14240
rect 48318 14320 48374 14376
rect 47829 14170 47885 14172
rect 47909 14170 47965 14172
rect 47989 14170 48045 14172
rect 48069 14170 48125 14172
rect 47829 14118 47875 14170
rect 47875 14118 47885 14170
rect 47909 14118 47939 14170
rect 47939 14118 47951 14170
rect 47951 14118 47965 14170
rect 47989 14118 48003 14170
rect 48003 14118 48015 14170
rect 48015 14118 48045 14170
rect 48069 14118 48079 14170
rect 48079 14118 48125 14170
rect 47829 14116 47885 14118
rect 47909 14116 47965 14118
rect 47989 14116 48045 14118
rect 48069 14116 48125 14118
rect 46754 12008 46810 12064
rect 47030 10784 47086 10840
rect 46570 9832 46626 9888
rect 47829 13082 47885 13084
rect 47909 13082 47965 13084
rect 47989 13082 48045 13084
rect 48069 13082 48125 13084
rect 47829 13030 47875 13082
rect 47875 13030 47885 13082
rect 47909 13030 47939 13082
rect 47939 13030 47951 13082
rect 47951 13030 47965 13082
rect 47989 13030 48003 13082
rect 48003 13030 48015 13082
rect 48015 13030 48045 13082
rect 48069 13030 48079 13082
rect 48079 13030 48125 13082
rect 47829 13028 47885 13030
rect 47909 13028 47965 13030
rect 47989 13028 48045 13030
rect 48069 13028 48125 13030
rect 48226 12688 48282 12744
rect 47829 11994 47885 11996
rect 47909 11994 47965 11996
rect 47989 11994 48045 11996
rect 48069 11994 48125 11996
rect 47829 11942 47875 11994
rect 47875 11942 47885 11994
rect 47909 11942 47939 11994
rect 47939 11942 47951 11994
rect 47951 11942 47965 11994
rect 47989 11942 48003 11994
rect 48003 11942 48015 11994
rect 48015 11942 48045 11994
rect 48069 11942 48079 11994
rect 48079 11942 48125 11994
rect 47829 11940 47885 11942
rect 47909 11940 47965 11942
rect 47989 11940 48045 11942
rect 48069 11940 48125 11942
rect 47829 10906 47885 10908
rect 47909 10906 47965 10908
rect 47989 10906 48045 10908
rect 48069 10906 48125 10908
rect 47829 10854 47875 10906
rect 47875 10854 47885 10906
rect 47909 10854 47939 10906
rect 47939 10854 47951 10906
rect 47951 10854 47965 10906
rect 47989 10854 48003 10906
rect 48003 10854 48015 10906
rect 48015 10854 48045 10906
rect 48069 10854 48079 10906
rect 48079 10854 48125 10906
rect 47829 10852 47885 10854
rect 47909 10852 47965 10854
rect 47989 10852 48045 10854
rect 48069 10852 48125 10854
rect 48778 15408 48834 15464
rect 50342 14864 50398 14920
rect 48962 11212 49018 11248
rect 48962 11192 48964 11212
rect 48964 11192 49016 11212
rect 49016 11192 49018 11212
rect 48410 10784 48466 10840
rect 47674 10512 47730 10568
rect 47829 9818 47885 9820
rect 47909 9818 47965 9820
rect 47989 9818 48045 9820
rect 48069 9818 48125 9820
rect 47829 9766 47875 9818
rect 47875 9766 47885 9818
rect 47909 9766 47939 9818
rect 47939 9766 47951 9818
rect 47951 9766 47965 9818
rect 47989 9766 48003 9818
rect 48003 9766 48015 9818
rect 48015 9766 48045 9818
rect 48069 9766 48079 9818
rect 48079 9766 48125 9818
rect 47829 9764 47885 9766
rect 47909 9764 47965 9766
rect 47989 9764 48045 9766
rect 48069 9764 48125 9766
rect 49330 10512 49386 10568
rect 46570 9288 46626 9344
rect 46570 8780 46572 8800
rect 46572 8780 46624 8800
rect 46624 8780 46626 8800
rect 46570 8744 46626 8780
rect 46570 8508 46572 8528
rect 46572 8508 46624 8528
rect 46624 8508 46626 8528
rect 46570 8472 46626 8508
rect 46570 7540 46626 7576
rect 46570 7520 46572 7540
rect 46572 7520 46624 7540
rect 46624 7520 46626 7540
rect 46754 9016 46810 9072
rect 47214 8744 47270 8800
rect 47398 8064 47454 8120
rect 47306 5636 47362 5672
rect 47306 5616 47308 5636
rect 47308 5616 47360 5636
rect 47360 5616 47362 5636
rect 45834 4528 45890 4584
rect 47582 9016 47638 9072
rect 47829 8730 47885 8732
rect 47909 8730 47965 8732
rect 47989 8730 48045 8732
rect 48069 8730 48125 8732
rect 47829 8678 47875 8730
rect 47875 8678 47885 8730
rect 47909 8678 47939 8730
rect 47939 8678 47951 8730
rect 47951 8678 47965 8730
rect 47989 8678 48003 8730
rect 48003 8678 48015 8730
rect 48015 8678 48045 8730
rect 48069 8678 48079 8730
rect 48079 8678 48125 8730
rect 47829 8676 47885 8678
rect 47909 8676 47965 8678
rect 47989 8676 48045 8678
rect 48069 8676 48125 8678
rect 48870 9324 48872 9344
rect 48872 9324 48924 9344
rect 48924 9324 48926 9344
rect 48870 9288 48926 9324
rect 48778 9016 48834 9072
rect 47829 7642 47885 7644
rect 47909 7642 47965 7644
rect 47989 7642 48045 7644
rect 48069 7642 48125 7644
rect 47829 7590 47875 7642
rect 47875 7590 47885 7642
rect 47909 7590 47939 7642
rect 47939 7590 47951 7642
rect 47951 7590 47965 7642
rect 47989 7590 48003 7642
rect 48003 7590 48015 7642
rect 48015 7590 48045 7642
rect 48069 7590 48079 7642
rect 48079 7590 48125 7642
rect 47829 7588 47885 7590
rect 47909 7588 47965 7590
rect 47989 7588 48045 7590
rect 48069 7588 48125 7590
rect 49882 11600 49938 11656
rect 49698 11192 49754 11248
rect 49514 10920 49570 10976
rect 49606 9288 49662 9344
rect 49514 8336 49570 8392
rect 50158 10804 50214 10840
rect 50158 10784 50160 10804
rect 50160 10784 50212 10804
rect 50212 10784 50214 10804
rect 51354 14320 51410 14376
rect 50618 11192 50674 11248
rect 50710 10920 50766 10976
rect 52366 15952 52422 16008
rect 53838 15000 53894 15056
rect 52090 13096 52146 13152
rect 51354 12144 51410 12200
rect 51170 11872 51226 11928
rect 52550 9832 52606 9888
rect 51078 7928 51134 7984
rect 49146 7112 49202 7168
rect 50342 6860 50398 6896
rect 51170 7828 51172 7848
rect 51172 7828 51224 7848
rect 51224 7828 51226 7848
rect 51170 7792 51226 7828
rect 51722 7792 51778 7848
rect 51078 7520 51134 7576
rect 50342 6840 50344 6860
rect 50344 6840 50396 6860
rect 50396 6840 50398 6860
rect 47829 6554 47885 6556
rect 47909 6554 47965 6556
rect 47989 6554 48045 6556
rect 48069 6554 48125 6556
rect 47829 6502 47875 6554
rect 47875 6502 47885 6554
rect 47909 6502 47939 6554
rect 47939 6502 47951 6554
rect 47951 6502 47965 6554
rect 47989 6502 48003 6554
rect 48003 6502 48015 6554
rect 48015 6502 48045 6554
rect 48069 6502 48079 6554
rect 48079 6502 48125 6554
rect 47829 6500 47885 6502
rect 47909 6500 47965 6502
rect 47989 6500 48045 6502
rect 48069 6500 48125 6502
rect 48226 6432 48282 6488
rect 48318 5752 48374 5808
rect 47490 5072 47546 5128
rect 47829 5466 47885 5468
rect 47909 5466 47965 5468
rect 47989 5466 48045 5468
rect 48069 5466 48125 5468
rect 47829 5414 47875 5466
rect 47875 5414 47885 5466
rect 47909 5414 47939 5466
rect 47939 5414 47951 5466
rect 47951 5414 47965 5466
rect 47989 5414 48003 5466
rect 48003 5414 48015 5466
rect 48015 5414 48045 5466
rect 48069 5414 48079 5466
rect 48079 5414 48125 5466
rect 47829 5412 47885 5414
rect 47909 5412 47965 5414
rect 47989 5412 48045 5414
rect 48069 5412 48125 5414
rect 47582 4936 47638 4992
rect 47490 4528 47546 4584
rect 49514 5908 49570 5944
rect 49514 5888 49516 5908
rect 49516 5888 49568 5908
rect 49568 5888 49570 5908
rect 51722 6432 51778 6488
rect 49974 6024 50030 6080
rect 47829 4378 47885 4380
rect 47909 4378 47965 4380
rect 47989 4378 48045 4380
rect 48069 4378 48125 4380
rect 47829 4326 47875 4378
rect 47875 4326 47885 4378
rect 47909 4326 47939 4378
rect 47939 4326 47951 4378
rect 47951 4326 47965 4378
rect 47989 4326 48003 4378
rect 48003 4326 48015 4378
rect 48015 4326 48045 4378
rect 48069 4326 48079 4378
rect 48079 4326 48125 4378
rect 47829 4324 47885 4326
rect 47909 4324 47965 4326
rect 47989 4324 48045 4326
rect 48069 4324 48125 4326
rect 50802 5908 50858 5944
rect 50802 5888 50804 5908
rect 50804 5888 50856 5908
rect 50856 5888 50858 5908
rect 50618 5072 50674 5128
rect 51170 4936 51226 4992
rect 51538 4936 51594 4992
rect 51998 4564 52000 4584
rect 52000 4564 52052 4584
rect 52052 4564 52054 4584
rect 51998 4528 52054 4564
rect 53286 10784 53342 10840
rect 53654 10784 53710 10840
rect 53286 10260 53342 10296
rect 53286 10240 53288 10260
rect 53288 10240 53340 10260
rect 53340 10240 53342 10260
rect 54850 13912 54906 13968
rect 54666 11228 54668 11248
rect 54668 11228 54720 11248
rect 54720 11228 54722 11248
rect 54666 11192 54722 11228
rect 53838 10920 53894 10976
rect 54482 10240 54538 10296
rect 53654 6196 53656 6216
rect 53656 6196 53708 6216
rect 53708 6196 53710 6216
rect 53654 6160 53710 6196
rect 54206 7112 54262 7168
rect 53838 6332 53840 6352
rect 53840 6332 53892 6352
rect 53892 6332 53894 6352
rect 53838 6296 53894 6332
rect 53654 5208 53710 5264
rect 36111 2746 36167 2748
rect 36191 2746 36247 2748
rect 36271 2746 36327 2748
rect 36351 2746 36407 2748
rect 36111 2694 36157 2746
rect 36157 2694 36167 2746
rect 36191 2694 36221 2746
rect 36221 2694 36233 2746
rect 36233 2694 36247 2746
rect 36271 2694 36285 2746
rect 36285 2694 36297 2746
rect 36297 2694 36327 2746
rect 36351 2694 36361 2746
rect 36361 2694 36407 2746
rect 36111 2692 36167 2694
rect 36191 2692 36247 2694
rect 36271 2692 36327 2694
rect 36351 2692 36407 2694
rect 47829 3290 47885 3292
rect 47909 3290 47965 3292
rect 47989 3290 48045 3292
rect 48069 3290 48125 3292
rect 47829 3238 47875 3290
rect 47875 3238 47885 3290
rect 47909 3238 47939 3290
rect 47939 3238 47951 3290
rect 47951 3238 47965 3290
rect 47989 3238 48003 3290
rect 48003 3238 48015 3290
rect 48015 3238 48045 3290
rect 48069 3238 48079 3290
rect 48079 3238 48125 3290
rect 47829 3236 47885 3238
rect 47909 3236 47965 3238
rect 47989 3236 48045 3238
rect 48069 3236 48125 3238
rect 55678 12960 55734 13016
rect 55678 12552 55734 12608
rect 56322 13232 56378 13288
rect 56138 12416 56194 12472
rect 56598 12044 56600 12064
rect 56600 12044 56652 12064
rect 56652 12044 56654 12064
rect 56598 12008 56654 12044
rect 56690 11756 56746 11792
rect 56690 11736 56692 11756
rect 56692 11736 56744 11756
rect 56744 11736 56746 11756
rect 56506 11620 56562 11656
rect 56506 11600 56508 11620
rect 56508 11600 56560 11620
rect 56560 11600 56562 11620
rect 56966 15544 57022 15600
rect 55402 10376 55458 10432
rect 55494 8880 55550 8936
rect 55402 8472 55458 8528
rect 56782 11056 56838 11112
rect 56046 9460 56048 9480
rect 56048 9460 56100 9480
rect 56100 9460 56102 9480
rect 56046 9424 56102 9460
rect 55218 6840 55274 6896
rect 54574 6024 54630 6080
rect 56046 5344 56102 5400
rect 57978 14048 58034 14104
rect 57702 12416 57758 12472
rect 57334 11092 57336 11112
rect 57336 11092 57388 11112
rect 57388 11092 57390 11112
rect 57334 11056 57390 11092
rect 59548 16890 59604 16892
rect 59628 16890 59684 16892
rect 59708 16890 59764 16892
rect 59788 16890 59844 16892
rect 59548 16838 59594 16890
rect 59594 16838 59604 16890
rect 59628 16838 59658 16890
rect 59658 16838 59670 16890
rect 59670 16838 59684 16890
rect 59708 16838 59722 16890
rect 59722 16838 59734 16890
rect 59734 16838 59764 16890
rect 59788 16838 59798 16890
rect 59798 16838 59844 16890
rect 59548 16836 59604 16838
rect 59628 16836 59684 16838
rect 59708 16836 59764 16838
rect 59788 16836 59844 16838
rect 57426 10104 57482 10160
rect 58254 10648 58310 10704
rect 57610 8900 57666 8936
rect 57610 8880 57612 8900
rect 57612 8880 57664 8900
rect 57664 8880 57666 8900
rect 57334 7792 57390 7848
rect 58070 7404 58126 7440
rect 58070 7384 58072 7404
rect 58072 7384 58124 7404
rect 58124 7384 58126 7404
rect 56966 6724 57022 6760
rect 56966 6704 56968 6724
rect 56968 6704 57020 6724
rect 57020 6704 57022 6724
rect 57150 5752 57206 5808
rect 56782 5072 56838 5128
rect 56690 4972 56692 4992
rect 56692 4972 56744 4992
rect 56744 4972 56746 4992
rect 56690 4936 56746 4972
rect 57334 4564 57336 4584
rect 57336 4564 57388 4584
rect 57388 4564 57390 4584
rect 57334 4528 57390 4564
rect 59082 15136 59138 15192
rect 58714 12008 58770 12064
rect 59548 15802 59604 15804
rect 59628 15802 59684 15804
rect 59708 15802 59764 15804
rect 59788 15802 59844 15804
rect 59548 15750 59594 15802
rect 59594 15750 59604 15802
rect 59628 15750 59658 15802
rect 59658 15750 59670 15802
rect 59670 15750 59684 15802
rect 59708 15750 59722 15802
rect 59722 15750 59734 15802
rect 59734 15750 59764 15802
rect 59788 15750 59798 15802
rect 59798 15750 59844 15802
rect 59548 15748 59604 15750
rect 59628 15748 59684 15750
rect 59708 15748 59764 15750
rect 59788 15748 59844 15750
rect 59174 13912 59230 13968
rect 59548 14714 59604 14716
rect 59628 14714 59684 14716
rect 59708 14714 59764 14716
rect 59788 14714 59844 14716
rect 59548 14662 59594 14714
rect 59594 14662 59604 14714
rect 59628 14662 59658 14714
rect 59658 14662 59670 14714
rect 59670 14662 59684 14714
rect 59708 14662 59722 14714
rect 59722 14662 59734 14714
rect 59734 14662 59764 14714
rect 59788 14662 59798 14714
rect 59798 14662 59844 14714
rect 59548 14660 59604 14662
rect 59628 14660 59684 14662
rect 59708 14660 59764 14662
rect 59788 14660 59844 14662
rect 59548 13626 59604 13628
rect 59628 13626 59684 13628
rect 59708 13626 59764 13628
rect 59788 13626 59844 13628
rect 59548 13574 59594 13626
rect 59594 13574 59604 13626
rect 59628 13574 59658 13626
rect 59658 13574 59670 13626
rect 59670 13574 59684 13626
rect 59708 13574 59722 13626
rect 59722 13574 59734 13626
rect 59734 13574 59764 13626
rect 59788 13574 59798 13626
rect 59798 13574 59844 13626
rect 59548 13572 59604 13574
rect 59628 13572 59684 13574
rect 59708 13572 59764 13574
rect 59788 13572 59844 13574
rect 59548 12538 59604 12540
rect 59628 12538 59684 12540
rect 59708 12538 59764 12540
rect 59788 12538 59844 12540
rect 59548 12486 59594 12538
rect 59594 12486 59604 12538
rect 59628 12486 59658 12538
rect 59658 12486 59670 12538
rect 59670 12486 59684 12538
rect 59708 12486 59722 12538
rect 59722 12486 59734 12538
rect 59734 12486 59764 12538
rect 59788 12486 59798 12538
rect 59798 12486 59844 12538
rect 59548 12484 59604 12486
rect 59628 12484 59684 12486
rect 59708 12484 59764 12486
rect 59788 12484 59844 12486
rect 59174 12144 59230 12200
rect 58898 11056 58954 11112
rect 59910 12280 59966 12336
rect 59548 11450 59604 11452
rect 59628 11450 59684 11452
rect 59708 11450 59764 11452
rect 59788 11450 59844 11452
rect 59548 11398 59594 11450
rect 59594 11398 59604 11450
rect 59628 11398 59658 11450
rect 59658 11398 59670 11450
rect 59670 11398 59684 11450
rect 59708 11398 59722 11450
rect 59722 11398 59734 11450
rect 59734 11398 59764 11450
rect 59788 11398 59798 11450
rect 59798 11398 59844 11450
rect 59548 11396 59604 11398
rect 59628 11396 59684 11398
rect 59708 11396 59764 11398
rect 59788 11396 59844 11398
rect 60186 12960 60242 13016
rect 60186 12552 60242 12608
rect 60370 13504 60426 13560
rect 59910 11056 59966 11112
rect 59548 10362 59604 10364
rect 59628 10362 59684 10364
rect 59708 10362 59764 10364
rect 59788 10362 59844 10364
rect 59548 10310 59594 10362
rect 59594 10310 59604 10362
rect 59628 10310 59658 10362
rect 59658 10310 59670 10362
rect 59670 10310 59684 10362
rect 59708 10310 59722 10362
rect 59722 10310 59734 10362
rect 59734 10310 59764 10362
rect 59788 10310 59798 10362
rect 59798 10310 59844 10362
rect 59548 10308 59604 10310
rect 59628 10308 59684 10310
rect 59708 10308 59764 10310
rect 59788 10308 59844 10310
rect 59358 10240 59414 10296
rect 59358 9696 59414 9752
rect 60370 11500 60372 11520
rect 60372 11500 60424 11520
rect 60424 11500 60426 11520
rect 60370 11464 60426 11500
rect 60094 11328 60150 11384
rect 60646 14184 60702 14240
rect 60646 13640 60702 13696
rect 61658 13912 61714 13968
rect 60646 12280 60702 12336
rect 60554 11736 60610 11792
rect 60738 11736 60794 11792
rect 61290 13096 61346 13152
rect 60922 11600 60978 11656
rect 64694 15408 64750 15464
rect 62026 12960 62082 13016
rect 61934 12144 61990 12200
rect 60370 9696 60426 9752
rect 59548 9274 59604 9276
rect 59628 9274 59684 9276
rect 59708 9274 59764 9276
rect 59788 9274 59844 9276
rect 59548 9222 59594 9274
rect 59594 9222 59604 9274
rect 59628 9222 59658 9274
rect 59658 9222 59670 9274
rect 59670 9222 59684 9274
rect 59708 9222 59722 9274
rect 59722 9222 59734 9274
rect 59734 9222 59764 9274
rect 59788 9222 59798 9274
rect 59798 9222 59844 9274
rect 59548 9220 59604 9222
rect 59628 9220 59684 9222
rect 59708 9220 59764 9222
rect 59788 9220 59844 9222
rect 60002 9152 60058 9208
rect 60002 8880 60058 8936
rect 58714 6432 58770 6488
rect 58806 5772 58862 5808
rect 58806 5752 58808 5772
rect 58808 5752 58860 5772
rect 58860 5752 58862 5772
rect 58806 5344 58862 5400
rect 59548 8186 59604 8188
rect 59628 8186 59684 8188
rect 59708 8186 59764 8188
rect 59788 8186 59844 8188
rect 59548 8134 59594 8186
rect 59594 8134 59604 8186
rect 59628 8134 59658 8186
rect 59658 8134 59670 8186
rect 59670 8134 59684 8186
rect 59708 8134 59722 8186
rect 59722 8134 59734 8186
rect 59734 8134 59764 8186
rect 59788 8134 59798 8186
rect 59798 8134 59844 8186
rect 59548 8132 59604 8134
rect 59628 8132 59684 8134
rect 59708 8132 59764 8134
rect 59788 8132 59844 8134
rect 59548 7098 59604 7100
rect 59628 7098 59684 7100
rect 59708 7098 59764 7100
rect 59788 7098 59844 7100
rect 59548 7046 59594 7098
rect 59594 7046 59604 7098
rect 59628 7046 59658 7098
rect 59658 7046 59670 7098
rect 59670 7046 59684 7098
rect 59708 7046 59722 7098
rect 59722 7046 59734 7098
rect 59734 7046 59764 7098
rect 59788 7046 59798 7098
rect 59798 7046 59844 7098
rect 59548 7044 59604 7046
rect 59628 7044 59684 7046
rect 59708 7044 59764 7046
rect 59788 7044 59844 7046
rect 59548 6010 59604 6012
rect 59628 6010 59684 6012
rect 59708 6010 59764 6012
rect 59788 6010 59844 6012
rect 59548 5958 59594 6010
rect 59594 5958 59604 6010
rect 59628 5958 59658 6010
rect 59658 5958 59670 6010
rect 59670 5958 59684 6010
rect 59708 5958 59722 6010
rect 59722 5958 59734 6010
rect 59734 5958 59764 6010
rect 59788 5958 59798 6010
rect 59798 5958 59844 6010
rect 59548 5956 59604 5958
rect 59628 5956 59684 5958
rect 59708 5956 59764 5958
rect 59788 5956 59844 5958
rect 59548 4922 59604 4924
rect 59628 4922 59684 4924
rect 59708 4922 59764 4924
rect 59788 4922 59844 4924
rect 59548 4870 59594 4922
rect 59594 4870 59604 4922
rect 59628 4870 59658 4922
rect 59658 4870 59670 4922
rect 59670 4870 59684 4922
rect 59708 4870 59722 4922
rect 59722 4870 59734 4922
rect 59734 4870 59764 4922
rect 59788 4870 59798 4922
rect 59798 4870 59844 4922
rect 59548 4868 59604 4870
rect 59628 4868 59684 4870
rect 59708 4868 59764 4870
rect 59788 4868 59844 4870
rect 61566 9968 61622 10024
rect 61014 8608 61070 8664
rect 60646 7520 60702 7576
rect 60738 5772 60794 5808
rect 60738 5752 60740 5772
rect 60740 5752 60792 5772
rect 60792 5752 60794 5772
rect 63038 12280 63094 12336
rect 63222 14048 63278 14104
rect 66074 14184 66130 14240
rect 64694 13676 64696 13696
rect 64696 13676 64748 13696
rect 64748 13676 64750 13696
rect 64694 13640 64750 13676
rect 66442 13912 66498 13968
rect 59548 3834 59604 3836
rect 59628 3834 59684 3836
rect 59708 3834 59764 3836
rect 59788 3834 59844 3836
rect 59548 3782 59594 3834
rect 59594 3782 59604 3834
rect 59628 3782 59658 3834
rect 59658 3782 59670 3834
rect 59670 3782 59684 3834
rect 59708 3782 59722 3834
rect 59722 3782 59734 3834
rect 59734 3782 59764 3834
rect 59788 3782 59798 3834
rect 59798 3782 59844 3834
rect 59548 3780 59604 3782
rect 59628 3780 59684 3782
rect 59708 3780 59764 3782
rect 59788 3780 59844 3782
rect 62578 7520 62634 7576
rect 63130 9444 63186 9480
rect 63130 9424 63132 9444
rect 63132 9424 63184 9444
rect 63184 9424 63186 9444
rect 63498 8608 63554 8664
rect 63314 7384 63370 7440
rect 63774 8472 63830 8528
rect 63682 8336 63738 8392
rect 64050 8336 64106 8392
rect 63590 4800 63646 4856
rect 64786 12144 64842 12200
rect 65062 11872 65118 11928
rect 64234 8916 64236 8936
rect 64236 8916 64288 8936
rect 64288 8916 64290 8936
rect 64234 8880 64290 8916
rect 65798 8744 65854 8800
rect 64510 8608 64566 8664
rect 59548 2746 59604 2748
rect 59628 2746 59684 2748
rect 59708 2746 59764 2748
rect 59788 2746 59844 2748
rect 59548 2694 59594 2746
rect 59594 2694 59604 2746
rect 59628 2694 59658 2746
rect 59658 2694 59670 2746
rect 59670 2694 59684 2746
rect 59708 2694 59722 2746
rect 59722 2694 59734 2746
rect 59734 2694 59764 2746
rect 59788 2694 59798 2746
rect 59798 2694 59844 2746
rect 59548 2692 59604 2694
rect 59628 2692 59684 2694
rect 59708 2692 59764 2694
rect 59788 2692 59844 2694
rect 65982 9696 66038 9752
rect 66718 13504 66774 13560
rect 66442 11328 66498 11384
rect 67178 12960 67234 13016
rect 67086 12008 67142 12064
rect 67086 9016 67142 9072
rect 66718 7792 66774 7848
rect 66626 7384 66682 7440
rect 67086 7112 67142 7168
rect 67454 14068 67510 14104
rect 67454 14048 67456 14068
rect 67456 14048 67508 14068
rect 67508 14048 67510 14068
rect 68466 14456 68522 14512
rect 68190 14356 68192 14376
rect 68192 14356 68244 14376
rect 68244 14356 68246 14376
rect 68190 14320 68246 14356
rect 67914 13096 67970 13152
rect 68466 13640 68522 13696
rect 68282 13504 68338 13560
rect 67546 12144 67602 12200
rect 67454 9424 67510 9480
rect 67638 9424 67694 9480
rect 67914 9832 67970 9888
rect 67822 9288 67878 9344
rect 68282 10784 68338 10840
rect 68466 10376 68522 10432
rect 68006 9424 68062 9480
rect 69570 12416 69626 12472
rect 71266 17434 71322 17436
rect 71346 17434 71402 17436
rect 71426 17434 71482 17436
rect 71506 17434 71562 17436
rect 71266 17382 71312 17434
rect 71312 17382 71322 17434
rect 71346 17382 71376 17434
rect 71376 17382 71388 17434
rect 71388 17382 71402 17434
rect 71426 17382 71440 17434
rect 71440 17382 71452 17434
rect 71452 17382 71482 17434
rect 71506 17382 71516 17434
rect 71516 17382 71562 17434
rect 71266 17380 71322 17382
rect 71346 17380 71402 17382
rect 71426 17380 71482 17382
rect 71506 17380 71562 17382
rect 71266 16346 71322 16348
rect 71346 16346 71402 16348
rect 71426 16346 71482 16348
rect 71506 16346 71562 16348
rect 71266 16294 71312 16346
rect 71312 16294 71322 16346
rect 71346 16294 71376 16346
rect 71376 16294 71388 16346
rect 71388 16294 71402 16346
rect 71426 16294 71440 16346
rect 71440 16294 71452 16346
rect 71452 16294 71482 16346
rect 71506 16294 71516 16346
rect 71516 16294 71562 16346
rect 71266 16292 71322 16294
rect 71346 16292 71402 16294
rect 71426 16292 71482 16294
rect 71506 16292 71562 16294
rect 69754 13368 69810 13424
rect 69478 12144 69534 12200
rect 68006 7384 68062 7440
rect 67178 6976 67234 7032
rect 66626 6432 66682 6488
rect 67822 6840 67878 6896
rect 68834 7520 68890 7576
rect 71266 15258 71322 15260
rect 71346 15258 71402 15260
rect 71426 15258 71482 15260
rect 71506 15258 71562 15260
rect 71266 15206 71312 15258
rect 71312 15206 71322 15258
rect 71346 15206 71376 15258
rect 71376 15206 71388 15258
rect 71388 15206 71402 15258
rect 71426 15206 71440 15258
rect 71440 15206 71452 15258
rect 71452 15206 71482 15258
rect 71506 15206 71516 15258
rect 71516 15206 71562 15258
rect 71266 15204 71322 15206
rect 71346 15204 71402 15206
rect 71426 15204 71482 15206
rect 71506 15204 71562 15206
rect 70674 13912 70730 13968
rect 71266 14170 71322 14172
rect 71346 14170 71402 14172
rect 71426 14170 71482 14172
rect 71506 14170 71562 14172
rect 71266 14118 71312 14170
rect 71312 14118 71322 14170
rect 71346 14118 71376 14170
rect 71376 14118 71388 14170
rect 71388 14118 71402 14170
rect 71426 14118 71440 14170
rect 71440 14118 71452 14170
rect 71452 14118 71482 14170
rect 71506 14118 71516 14170
rect 71516 14118 71562 14170
rect 71266 14116 71322 14118
rect 71346 14116 71402 14118
rect 71426 14116 71482 14118
rect 71506 14116 71562 14118
rect 71134 13368 71190 13424
rect 71266 13082 71322 13084
rect 71346 13082 71402 13084
rect 71426 13082 71482 13084
rect 71506 13082 71562 13084
rect 71266 13030 71312 13082
rect 71312 13030 71322 13082
rect 71346 13030 71376 13082
rect 71376 13030 71388 13082
rect 71388 13030 71402 13082
rect 71426 13030 71440 13082
rect 71440 13030 71452 13082
rect 71452 13030 71482 13082
rect 71506 13030 71516 13082
rect 71516 13030 71562 13082
rect 71266 13028 71322 13030
rect 71346 13028 71402 13030
rect 71426 13028 71482 13030
rect 71506 13028 71562 13030
rect 71686 12960 71742 13016
rect 69754 11600 69810 11656
rect 69570 10240 69626 10296
rect 70582 10784 70638 10840
rect 70306 9696 70362 9752
rect 70214 9424 70270 9480
rect 71134 12552 71190 12608
rect 71042 12416 71098 12472
rect 71318 12552 71374 12608
rect 71266 11994 71322 11996
rect 71346 11994 71402 11996
rect 71426 11994 71482 11996
rect 71506 11994 71562 11996
rect 71266 11942 71312 11994
rect 71312 11942 71322 11994
rect 71346 11942 71376 11994
rect 71376 11942 71388 11994
rect 71388 11942 71402 11994
rect 71426 11942 71440 11994
rect 71440 11942 71452 11994
rect 71452 11942 71482 11994
rect 71506 11942 71516 11994
rect 71516 11942 71562 11994
rect 71266 11940 71322 11942
rect 71346 11940 71402 11942
rect 71426 11940 71482 11942
rect 71506 11940 71562 11942
rect 71962 13096 72018 13152
rect 71134 11328 71190 11384
rect 71134 10956 71136 10976
rect 71136 10956 71188 10976
rect 71188 10956 71190 10976
rect 71134 10920 71190 10956
rect 71266 10906 71322 10908
rect 71346 10906 71402 10908
rect 71426 10906 71482 10908
rect 71506 10906 71562 10908
rect 71266 10854 71312 10906
rect 71312 10854 71322 10906
rect 71346 10854 71376 10906
rect 71376 10854 71388 10906
rect 71388 10854 71402 10906
rect 71426 10854 71440 10906
rect 71440 10854 71452 10906
rect 71452 10854 71482 10906
rect 71506 10854 71516 10906
rect 71516 10854 71562 10906
rect 71266 10852 71322 10854
rect 71346 10852 71402 10854
rect 71426 10852 71482 10854
rect 71506 10852 71562 10854
rect 70950 10376 71006 10432
rect 69570 7792 69626 7848
rect 69478 7248 69534 7304
rect 68834 7112 68890 7168
rect 69846 7112 69902 7168
rect 68742 6840 68798 6896
rect 69202 5752 69258 5808
rect 71266 9818 71322 9820
rect 71346 9818 71402 9820
rect 71426 9818 71482 9820
rect 71506 9818 71562 9820
rect 71266 9766 71312 9818
rect 71312 9766 71322 9818
rect 71346 9766 71376 9818
rect 71376 9766 71388 9818
rect 71388 9766 71402 9818
rect 71426 9766 71440 9818
rect 71440 9766 71452 9818
rect 71452 9766 71482 9818
rect 71506 9766 71516 9818
rect 71516 9766 71562 9818
rect 71266 9764 71322 9766
rect 71346 9764 71402 9766
rect 71426 9764 71482 9766
rect 71506 9764 71562 9766
rect 71134 9424 71190 9480
rect 72238 11192 72294 11248
rect 72606 14048 72662 14104
rect 73250 13504 73306 13560
rect 72422 12552 72478 12608
rect 72606 12280 72662 12336
rect 72514 12008 72570 12064
rect 72698 12164 72754 12200
rect 72698 12144 72700 12164
rect 72700 12144 72752 12164
rect 72752 12144 72754 12164
rect 72422 9288 72478 9344
rect 71870 9152 71926 9208
rect 71266 8730 71322 8732
rect 71346 8730 71402 8732
rect 71426 8730 71482 8732
rect 71506 8730 71562 8732
rect 71266 8678 71312 8730
rect 71312 8678 71322 8730
rect 71346 8678 71376 8730
rect 71376 8678 71388 8730
rect 71388 8678 71402 8730
rect 71426 8678 71440 8730
rect 71440 8678 71452 8730
rect 71452 8678 71482 8730
rect 71506 8678 71516 8730
rect 71516 8678 71562 8730
rect 71266 8676 71322 8678
rect 71346 8676 71402 8678
rect 71426 8676 71482 8678
rect 71506 8676 71562 8678
rect 71502 7928 71558 7984
rect 71266 7642 71322 7644
rect 71346 7642 71402 7644
rect 71426 7642 71482 7644
rect 71506 7642 71562 7644
rect 71266 7590 71312 7642
rect 71312 7590 71322 7642
rect 71346 7590 71376 7642
rect 71376 7590 71388 7642
rect 71388 7590 71402 7642
rect 71426 7590 71440 7642
rect 71440 7590 71452 7642
rect 71452 7590 71482 7642
rect 71506 7590 71516 7642
rect 71516 7590 71562 7642
rect 71266 7588 71322 7590
rect 71346 7588 71402 7590
rect 71426 7588 71482 7590
rect 71506 7588 71562 7590
rect 71870 7112 71926 7168
rect 71870 6840 71926 6896
rect 73802 13932 73858 13968
rect 73802 13912 73804 13932
rect 73804 13912 73856 13932
rect 73856 13912 73858 13932
rect 75274 14884 75330 14920
rect 75274 14864 75276 14884
rect 75276 14864 75328 14884
rect 75328 14864 75330 14884
rect 73618 12008 73674 12064
rect 74630 12280 74686 12336
rect 72882 10104 72938 10160
rect 73986 9424 74042 9480
rect 75734 13640 75790 13696
rect 82985 16890 83041 16892
rect 83065 16890 83121 16892
rect 83145 16890 83201 16892
rect 83225 16890 83281 16892
rect 82985 16838 83031 16890
rect 83031 16838 83041 16890
rect 83065 16838 83095 16890
rect 83095 16838 83107 16890
rect 83107 16838 83121 16890
rect 83145 16838 83159 16890
rect 83159 16838 83171 16890
rect 83171 16838 83201 16890
rect 83225 16838 83235 16890
rect 83235 16838 83281 16890
rect 82985 16836 83041 16838
rect 83065 16836 83121 16838
rect 83145 16836 83201 16838
rect 83225 16836 83281 16838
rect 75182 12416 75238 12472
rect 74722 11636 74724 11656
rect 74724 11636 74776 11656
rect 74776 11636 74778 11656
rect 74722 11600 74778 11636
rect 75182 11192 75238 11248
rect 75458 11328 75514 11384
rect 76378 12180 76380 12200
rect 76380 12180 76432 12200
rect 76432 12180 76434 12200
rect 76378 12144 76434 12180
rect 76194 11872 76250 11928
rect 76102 10240 76158 10296
rect 75458 9424 75514 9480
rect 72606 7248 72662 7304
rect 72790 6704 72846 6760
rect 73526 7284 73528 7304
rect 73528 7284 73580 7304
rect 73580 7284 73582 7304
rect 73526 7248 73582 7284
rect 71266 6554 71322 6556
rect 71346 6554 71402 6556
rect 71426 6554 71482 6556
rect 71506 6554 71562 6556
rect 71266 6502 71312 6554
rect 71312 6502 71322 6554
rect 71346 6502 71376 6554
rect 71376 6502 71388 6554
rect 71388 6502 71402 6554
rect 71426 6502 71440 6554
rect 71440 6502 71452 6554
rect 71452 6502 71482 6554
rect 71506 6502 71516 6554
rect 71516 6502 71562 6554
rect 71266 6500 71322 6502
rect 71346 6500 71402 6502
rect 71426 6500 71482 6502
rect 71506 6500 71562 6502
rect 71266 5466 71322 5468
rect 71346 5466 71402 5468
rect 71426 5466 71482 5468
rect 71506 5466 71562 5468
rect 71266 5414 71312 5466
rect 71312 5414 71322 5466
rect 71346 5414 71376 5466
rect 71376 5414 71388 5466
rect 71388 5414 71402 5466
rect 71426 5414 71440 5466
rect 71440 5414 71452 5466
rect 71452 5414 71482 5466
rect 71506 5414 71516 5466
rect 71516 5414 71562 5466
rect 71266 5412 71322 5414
rect 71346 5412 71402 5414
rect 71426 5412 71482 5414
rect 71506 5412 71562 5414
rect 71778 5480 71834 5536
rect 71962 6432 72018 6488
rect 71266 4378 71322 4380
rect 71346 4378 71402 4380
rect 71426 4378 71482 4380
rect 71506 4378 71562 4380
rect 71266 4326 71312 4378
rect 71312 4326 71322 4378
rect 71346 4326 71376 4378
rect 71376 4326 71388 4378
rect 71388 4326 71402 4378
rect 71426 4326 71440 4378
rect 71440 4326 71452 4378
rect 71452 4326 71482 4378
rect 71506 4326 71516 4378
rect 71516 4326 71562 4378
rect 71266 4324 71322 4326
rect 71346 4324 71402 4326
rect 71426 4324 71482 4326
rect 71506 4324 71562 4326
rect 74538 7928 74594 7984
rect 74078 5888 74134 5944
rect 71266 3290 71322 3292
rect 71346 3290 71402 3292
rect 71426 3290 71482 3292
rect 71506 3290 71562 3292
rect 71266 3238 71312 3290
rect 71312 3238 71322 3290
rect 71346 3238 71376 3290
rect 71376 3238 71388 3290
rect 71388 3238 71402 3290
rect 71426 3238 71440 3290
rect 71440 3238 71452 3290
rect 71452 3238 71482 3290
rect 71506 3238 71516 3290
rect 71516 3238 71562 3290
rect 71266 3236 71322 3238
rect 71346 3236 71402 3238
rect 71426 3236 71482 3238
rect 71506 3236 71562 3238
rect 75918 6976 75974 7032
rect 74998 6568 75054 6624
rect 75274 5516 75276 5536
rect 75276 5516 75328 5536
rect 75328 5516 75330 5536
rect 75274 5480 75330 5516
rect 75458 6060 75460 6080
rect 75460 6060 75512 6080
rect 75512 6060 75514 6080
rect 75458 6024 75514 6060
rect 75550 5208 75606 5264
rect 77022 13368 77078 13424
rect 77022 13096 77078 13152
rect 77114 12960 77170 13016
rect 77206 11192 77262 11248
rect 76286 6568 76342 6624
rect 76562 6604 76564 6624
rect 76564 6604 76616 6624
rect 76616 6604 76618 6624
rect 76286 5908 76342 5944
rect 76286 5888 76288 5908
rect 76288 5888 76340 5908
rect 76340 5888 76342 5908
rect 76562 6568 76618 6604
rect 77850 15408 77906 15464
rect 78678 15036 78680 15056
rect 78680 15036 78732 15056
rect 78732 15036 78734 15056
rect 78678 15000 78734 15036
rect 82174 15952 82230 16008
rect 77482 13368 77538 13424
rect 77574 12300 77630 12336
rect 77574 12280 77576 12300
rect 77576 12280 77628 12300
rect 77628 12280 77630 12300
rect 77942 11872 77998 11928
rect 78586 11192 78642 11248
rect 79046 11872 79102 11928
rect 79414 13096 79470 13152
rect 77666 10376 77722 10432
rect 77298 6740 77300 6760
rect 77300 6740 77352 6760
rect 77352 6740 77354 6760
rect 76746 6024 76802 6080
rect 77298 6704 77354 6740
rect 76838 5228 76894 5264
rect 76838 5208 76840 5228
rect 76840 5208 76892 5228
rect 76892 5208 76894 5228
rect 77850 5908 77906 5944
rect 77850 5888 77852 5908
rect 77852 5888 77904 5908
rect 77904 5888 77906 5908
rect 80702 13776 80758 13832
rect 79966 10104 80022 10160
rect 78862 8880 78918 8936
rect 77574 4120 77630 4176
rect 79782 8472 79838 8528
rect 79874 8336 79930 8392
rect 79966 6568 80022 6624
rect 80058 5516 80060 5536
rect 80060 5516 80112 5536
rect 80112 5516 80114 5536
rect 80058 5480 80114 5516
rect 80518 8916 80520 8936
rect 80520 8916 80572 8936
rect 80572 8916 80574 8936
rect 80518 8880 80574 8916
rect 81438 11736 81494 11792
rect 82985 15802 83041 15804
rect 83065 15802 83121 15804
rect 83145 15802 83201 15804
rect 83225 15802 83281 15804
rect 82985 15750 83031 15802
rect 83031 15750 83041 15802
rect 83065 15750 83095 15802
rect 83095 15750 83107 15802
rect 83107 15750 83121 15802
rect 83145 15750 83159 15802
rect 83159 15750 83171 15802
rect 83171 15750 83201 15802
rect 83225 15750 83235 15802
rect 83235 15750 83281 15802
rect 82985 15748 83041 15750
rect 83065 15748 83121 15750
rect 83145 15748 83201 15750
rect 83225 15748 83281 15750
rect 81622 11600 81678 11656
rect 82985 14714 83041 14716
rect 83065 14714 83121 14716
rect 83145 14714 83201 14716
rect 83225 14714 83281 14716
rect 82985 14662 83031 14714
rect 83031 14662 83041 14714
rect 83065 14662 83095 14714
rect 83095 14662 83107 14714
rect 83107 14662 83121 14714
rect 83145 14662 83159 14714
rect 83159 14662 83171 14714
rect 83171 14662 83201 14714
rect 83225 14662 83235 14714
rect 83235 14662 83281 14714
rect 82985 14660 83041 14662
rect 83065 14660 83121 14662
rect 83145 14660 83201 14662
rect 83225 14660 83281 14662
rect 82985 13626 83041 13628
rect 83065 13626 83121 13628
rect 83145 13626 83201 13628
rect 83225 13626 83281 13628
rect 82985 13574 83031 13626
rect 83031 13574 83041 13626
rect 83065 13574 83095 13626
rect 83095 13574 83107 13626
rect 83107 13574 83121 13626
rect 83145 13574 83159 13626
rect 83159 13574 83171 13626
rect 83171 13574 83201 13626
rect 83225 13574 83235 13626
rect 83235 13574 83281 13626
rect 82985 13572 83041 13574
rect 83065 13572 83121 13574
rect 83145 13572 83201 13574
rect 83225 13572 83281 13574
rect 82266 13096 82322 13152
rect 82985 12538 83041 12540
rect 83065 12538 83121 12540
rect 83145 12538 83201 12540
rect 83225 12538 83281 12540
rect 82985 12486 83031 12538
rect 83031 12486 83041 12538
rect 83065 12486 83095 12538
rect 83095 12486 83107 12538
rect 83107 12486 83121 12538
rect 83145 12486 83159 12538
rect 83159 12486 83171 12538
rect 83171 12486 83201 12538
rect 83225 12486 83235 12538
rect 83235 12486 83281 12538
rect 82985 12484 83041 12486
rect 83065 12484 83121 12486
rect 83145 12484 83201 12486
rect 83225 12484 83281 12486
rect 82542 11600 82598 11656
rect 82985 11450 83041 11452
rect 83065 11450 83121 11452
rect 83145 11450 83201 11452
rect 83225 11450 83281 11452
rect 82985 11398 83031 11450
rect 83031 11398 83041 11450
rect 83065 11398 83095 11450
rect 83095 11398 83107 11450
rect 83107 11398 83121 11450
rect 83145 11398 83159 11450
rect 83159 11398 83171 11450
rect 83171 11398 83201 11450
rect 83225 11398 83235 11450
rect 83235 11398 83281 11450
rect 82985 11396 83041 11398
rect 83065 11396 83121 11398
rect 83145 11396 83201 11398
rect 83225 11396 83281 11398
rect 81806 10104 81862 10160
rect 82985 10362 83041 10364
rect 83065 10362 83121 10364
rect 83145 10362 83201 10364
rect 83225 10362 83281 10364
rect 82985 10310 83031 10362
rect 83031 10310 83041 10362
rect 83065 10310 83095 10362
rect 83095 10310 83107 10362
rect 83107 10310 83121 10362
rect 83145 10310 83159 10362
rect 83159 10310 83171 10362
rect 83171 10310 83201 10362
rect 83225 10310 83235 10362
rect 83235 10310 83281 10362
rect 82985 10308 83041 10310
rect 83065 10308 83121 10310
rect 83145 10308 83201 10310
rect 83225 10308 83281 10310
rect 81530 9560 81586 9616
rect 80794 8472 80850 8528
rect 80334 6740 80336 6760
rect 80336 6740 80388 6760
rect 80388 6740 80390 6760
rect 80334 6704 80390 6740
rect 80334 6568 80390 6624
rect 81254 5752 81310 5808
rect 82985 9274 83041 9276
rect 83065 9274 83121 9276
rect 83145 9274 83201 9276
rect 83225 9274 83281 9276
rect 82985 9222 83031 9274
rect 83031 9222 83041 9274
rect 83065 9222 83095 9274
rect 83095 9222 83107 9274
rect 83107 9222 83121 9274
rect 83145 9222 83159 9274
rect 83159 9222 83171 9274
rect 83171 9222 83201 9274
rect 83225 9222 83235 9274
rect 83235 9222 83281 9274
rect 82985 9220 83041 9222
rect 83065 9220 83121 9222
rect 83145 9220 83201 9222
rect 83225 9220 83281 9222
rect 81714 6724 81770 6760
rect 81714 6704 81716 6724
rect 81716 6704 81768 6724
rect 81768 6704 81770 6724
rect 81438 5616 81494 5672
rect 81622 5516 81624 5536
rect 81624 5516 81676 5536
rect 81676 5516 81678 5536
rect 81622 5480 81678 5516
rect 82985 8186 83041 8188
rect 83065 8186 83121 8188
rect 83145 8186 83201 8188
rect 83225 8186 83281 8188
rect 82985 8134 83031 8186
rect 83031 8134 83041 8186
rect 83065 8134 83095 8186
rect 83095 8134 83107 8186
rect 83107 8134 83121 8186
rect 83145 8134 83159 8186
rect 83159 8134 83171 8186
rect 83171 8134 83201 8186
rect 83225 8134 83235 8186
rect 83235 8134 83281 8186
rect 82985 8132 83041 8134
rect 83065 8132 83121 8134
rect 83145 8132 83201 8134
rect 83225 8132 83281 8134
rect 82985 7098 83041 7100
rect 83065 7098 83121 7100
rect 83145 7098 83201 7100
rect 83225 7098 83281 7100
rect 82985 7046 83031 7098
rect 83031 7046 83041 7098
rect 83065 7046 83095 7098
rect 83095 7046 83107 7098
rect 83107 7046 83121 7098
rect 83145 7046 83159 7098
rect 83159 7046 83171 7098
rect 83171 7046 83201 7098
rect 83225 7046 83235 7098
rect 83235 7046 83281 7098
rect 82985 7044 83041 7046
rect 83065 7044 83121 7046
rect 83145 7044 83201 7046
rect 83225 7044 83281 7046
rect 83738 11756 83794 11792
rect 83738 11736 83740 11756
rect 83740 11736 83792 11756
rect 83792 11736 83794 11756
rect 83554 7520 83610 7576
rect 83830 9988 83886 10024
rect 83830 9968 83832 9988
rect 83832 9968 83884 9988
rect 83884 9968 83886 9988
rect 82726 5888 82782 5944
rect 82985 6010 83041 6012
rect 83065 6010 83121 6012
rect 83145 6010 83201 6012
rect 83225 6010 83281 6012
rect 82985 5958 83031 6010
rect 83031 5958 83041 6010
rect 83065 5958 83095 6010
rect 83095 5958 83107 6010
rect 83107 5958 83121 6010
rect 83145 5958 83159 6010
rect 83159 5958 83171 6010
rect 83171 5958 83201 6010
rect 83225 5958 83235 6010
rect 83235 5958 83281 6010
rect 82985 5956 83041 5958
rect 83065 5956 83121 5958
rect 83145 5956 83201 5958
rect 83225 5956 83281 5958
rect 82985 4922 83041 4924
rect 83065 4922 83121 4924
rect 83145 4922 83201 4924
rect 83225 4922 83281 4924
rect 82985 4870 83031 4922
rect 83031 4870 83041 4922
rect 83065 4870 83095 4922
rect 83095 4870 83107 4922
rect 83107 4870 83121 4922
rect 83145 4870 83159 4922
rect 83159 4870 83171 4922
rect 83171 4870 83201 4922
rect 83225 4870 83235 4922
rect 83235 4870 83281 4922
rect 82985 4868 83041 4870
rect 83065 4868 83121 4870
rect 83145 4868 83201 4870
rect 83225 4868 83281 4870
rect 94703 17434 94759 17436
rect 94783 17434 94839 17436
rect 94863 17434 94919 17436
rect 94943 17434 94999 17436
rect 94703 17382 94749 17434
rect 94749 17382 94759 17434
rect 94783 17382 94813 17434
rect 94813 17382 94825 17434
rect 94825 17382 94839 17434
rect 94863 17382 94877 17434
rect 94877 17382 94889 17434
rect 94889 17382 94919 17434
rect 94943 17382 94953 17434
rect 94953 17382 94999 17434
rect 94703 17380 94759 17382
rect 94783 17380 94839 17382
rect 94863 17380 94919 17382
rect 94943 17380 94999 17382
rect 94226 16788 94282 16824
rect 94226 16768 94228 16788
rect 94228 16768 94280 16788
rect 94280 16768 94282 16788
rect 86314 16088 86370 16144
rect 84290 11636 84292 11656
rect 84292 11636 84344 11656
rect 84344 11636 84346 11656
rect 84290 11600 84346 11636
rect 84014 11076 84070 11112
rect 84014 11056 84016 11076
rect 84016 11056 84068 11076
rect 84068 11056 84070 11076
rect 84290 10648 84346 10704
rect 84198 10512 84254 10568
rect 82985 3834 83041 3836
rect 83065 3834 83121 3836
rect 83145 3834 83201 3836
rect 83225 3834 83281 3836
rect 82985 3782 83031 3834
rect 83031 3782 83041 3834
rect 83065 3782 83095 3834
rect 83095 3782 83107 3834
rect 83107 3782 83121 3834
rect 83145 3782 83159 3834
rect 83159 3782 83171 3834
rect 83171 3782 83201 3834
rect 83225 3782 83235 3834
rect 83235 3782 83281 3834
rect 82985 3780 83041 3782
rect 83065 3780 83121 3782
rect 83145 3780 83201 3782
rect 83225 3780 83281 3782
rect 83922 4664 83978 4720
rect 85486 10512 85542 10568
rect 85394 10104 85450 10160
rect 84750 9968 84806 10024
rect 85762 11228 85764 11248
rect 85764 11228 85816 11248
rect 85816 11228 85818 11248
rect 85762 11192 85818 11228
rect 85486 8880 85542 8936
rect 84934 7520 84990 7576
rect 85762 6160 85818 6216
rect 86590 7540 86646 7576
rect 86590 7520 86592 7540
rect 86592 7520 86644 7540
rect 86644 7520 86646 7540
rect 86866 12688 86922 12744
rect 94703 16346 94759 16348
rect 94783 16346 94839 16348
rect 94863 16346 94919 16348
rect 94943 16346 94999 16348
rect 94703 16294 94749 16346
rect 94749 16294 94759 16346
rect 94783 16294 94813 16346
rect 94813 16294 94825 16346
rect 94825 16294 94839 16346
rect 94863 16294 94877 16346
rect 94877 16294 94889 16346
rect 94889 16294 94919 16346
rect 94943 16294 94953 16346
rect 94953 16294 94999 16346
rect 94703 16292 94759 16294
rect 94783 16292 94839 16294
rect 94863 16292 94919 16294
rect 94943 16292 94999 16294
rect 88154 14048 88210 14104
rect 94703 15258 94759 15260
rect 94783 15258 94839 15260
rect 94863 15258 94919 15260
rect 94943 15258 94999 15260
rect 94703 15206 94749 15258
rect 94749 15206 94759 15258
rect 94783 15206 94813 15258
rect 94813 15206 94825 15258
rect 94825 15206 94839 15258
rect 94863 15206 94877 15258
rect 94877 15206 94889 15258
rect 94889 15206 94919 15258
rect 94943 15206 94953 15258
rect 94953 15206 94999 15258
rect 94703 15204 94759 15206
rect 94783 15204 94839 15206
rect 94863 15204 94919 15206
rect 94943 15204 94999 15206
rect 89442 12844 89498 12880
rect 89442 12824 89444 12844
rect 89444 12824 89496 12844
rect 89496 12824 89498 12844
rect 94703 14170 94759 14172
rect 94783 14170 94839 14172
rect 94863 14170 94919 14172
rect 94943 14170 94999 14172
rect 94703 14118 94749 14170
rect 94749 14118 94759 14170
rect 94783 14118 94813 14170
rect 94813 14118 94825 14170
rect 94825 14118 94839 14170
rect 94863 14118 94877 14170
rect 94877 14118 94889 14170
rect 94889 14118 94919 14170
rect 94943 14118 94953 14170
rect 94953 14118 94999 14170
rect 94703 14116 94759 14118
rect 94783 14116 94839 14118
rect 94863 14116 94919 14118
rect 94943 14116 94999 14118
rect 92478 13232 92534 13288
rect 88246 6976 88302 7032
rect 87878 6840 87934 6896
rect 86866 6160 86922 6216
rect 89442 6860 89498 6896
rect 89442 6840 89444 6860
rect 89444 6840 89496 6860
rect 89496 6840 89498 6860
rect 89902 6976 89958 7032
rect 82985 2746 83041 2748
rect 83065 2746 83121 2748
rect 83145 2746 83201 2748
rect 83225 2746 83281 2748
rect 82985 2694 83031 2746
rect 83031 2694 83041 2746
rect 83065 2694 83095 2746
rect 83095 2694 83107 2746
rect 83107 2694 83121 2746
rect 83145 2694 83159 2746
rect 83159 2694 83171 2746
rect 83171 2694 83201 2746
rect 83225 2694 83235 2746
rect 83235 2694 83281 2746
rect 82985 2692 83041 2694
rect 83065 2692 83121 2694
rect 83145 2692 83201 2694
rect 83225 2692 83281 2694
rect 94703 13082 94759 13084
rect 94783 13082 94839 13084
rect 94863 13082 94919 13084
rect 94943 13082 94999 13084
rect 94703 13030 94749 13082
rect 94749 13030 94759 13082
rect 94783 13030 94813 13082
rect 94813 13030 94825 13082
rect 94825 13030 94839 13082
rect 94863 13030 94877 13082
rect 94877 13030 94889 13082
rect 94889 13030 94919 13082
rect 94943 13030 94953 13082
rect 94953 13030 94999 13082
rect 94703 13028 94759 13030
rect 94783 13028 94839 13030
rect 94863 13028 94919 13030
rect 94943 13028 94999 13030
rect 94226 12436 94282 12472
rect 94226 12416 94228 12436
rect 94228 12416 94280 12436
rect 94280 12416 94282 12436
rect 94703 11994 94759 11996
rect 94783 11994 94839 11996
rect 94863 11994 94919 11996
rect 94943 11994 94999 11996
rect 94703 11942 94749 11994
rect 94749 11942 94759 11994
rect 94783 11942 94813 11994
rect 94813 11942 94825 11994
rect 94825 11942 94839 11994
rect 94863 11942 94877 11994
rect 94877 11942 94889 11994
rect 94889 11942 94919 11994
rect 94943 11942 94953 11994
rect 94953 11942 94999 11994
rect 94703 11940 94759 11942
rect 94783 11940 94839 11942
rect 94863 11940 94919 11942
rect 94943 11940 94999 11942
rect 94703 10906 94759 10908
rect 94783 10906 94839 10908
rect 94863 10906 94919 10908
rect 94943 10906 94999 10908
rect 94703 10854 94749 10906
rect 94749 10854 94759 10906
rect 94783 10854 94813 10906
rect 94813 10854 94825 10906
rect 94825 10854 94839 10906
rect 94863 10854 94877 10906
rect 94877 10854 94889 10906
rect 94889 10854 94919 10906
rect 94943 10854 94953 10906
rect 94953 10854 94999 10906
rect 94703 10852 94759 10854
rect 94783 10852 94839 10854
rect 94863 10852 94919 10854
rect 94943 10852 94999 10854
rect 93214 6296 93270 6352
rect 94703 9818 94759 9820
rect 94783 9818 94839 9820
rect 94863 9818 94919 9820
rect 94943 9818 94999 9820
rect 94703 9766 94749 9818
rect 94749 9766 94759 9818
rect 94783 9766 94813 9818
rect 94813 9766 94825 9818
rect 94825 9766 94839 9818
rect 94863 9766 94877 9818
rect 94877 9766 94889 9818
rect 94889 9766 94919 9818
rect 94943 9766 94953 9818
rect 94953 9766 94999 9818
rect 94703 9764 94759 9766
rect 94783 9764 94839 9766
rect 94863 9764 94919 9766
rect 94943 9764 94999 9766
rect 94703 8730 94759 8732
rect 94783 8730 94839 8732
rect 94863 8730 94919 8732
rect 94943 8730 94999 8732
rect 94703 8678 94749 8730
rect 94749 8678 94759 8730
rect 94783 8678 94813 8730
rect 94813 8678 94825 8730
rect 94825 8678 94839 8730
rect 94863 8678 94877 8730
rect 94877 8678 94889 8730
rect 94889 8678 94919 8730
rect 94943 8678 94953 8730
rect 94953 8678 94999 8730
rect 94703 8676 94759 8678
rect 94783 8676 94839 8678
rect 94863 8676 94919 8678
rect 94943 8676 94999 8678
rect 94703 7642 94759 7644
rect 94783 7642 94839 7644
rect 94863 7642 94919 7644
rect 94943 7642 94999 7644
rect 94703 7590 94749 7642
rect 94749 7590 94759 7642
rect 94783 7590 94813 7642
rect 94813 7590 94825 7642
rect 94825 7590 94839 7642
rect 94863 7590 94877 7642
rect 94877 7590 94889 7642
rect 94889 7590 94919 7642
rect 94943 7590 94953 7642
rect 94953 7590 94999 7642
rect 94703 7588 94759 7590
rect 94783 7588 94839 7590
rect 94863 7588 94919 7590
rect 94943 7588 94999 7590
rect 95146 7520 95202 7576
rect 94703 6554 94759 6556
rect 94783 6554 94839 6556
rect 94863 6554 94919 6556
rect 94943 6554 94999 6556
rect 94703 6502 94749 6554
rect 94749 6502 94759 6554
rect 94783 6502 94813 6554
rect 94813 6502 94825 6554
rect 94825 6502 94839 6554
rect 94863 6502 94877 6554
rect 94877 6502 94889 6554
rect 94889 6502 94919 6554
rect 94943 6502 94953 6554
rect 94953 6502 94999 6554
rect 94703 6500 94759 6502
rect 94783 6500 94839 6502
rect 94863 6500 94919 6502
rect 94943 6500 94999 6502
rect 94703 5466 94759 5468
rect 94783 5466 94839 5468
rect 94863 5466 94919 5468
rect 94943 5466 94999 5468
rect 94703 5414 94749 5466
rect 94749 5414 94759 5466
rect 94783 5414 94813 5466
rect 94813 5414 94825 5466
rect 94825 5414 94839 5466
rect 94863 5414 94877 5466
rect 94877 5414 94889 5466
rect 94889 5414 94919 5466
rect 94943 5414 94953 5466
rect 94953 5414 94999 5466
rect 94703 5412 94759 5414
rect 94783 5412 94839 5414
rect 94863 5412 94919 5414
rect 94943 5412 94999 5414
rect 94703 4378 94759 4380
rect 94783 4378 94839 4380
rect 94863 4378 94919 4380
rect 94943 4378 94999 4380
rect 94703 4326 94749 4378
rect 94749 4326 94759 4378
rect 94783 4326 94813 4378
rect 94813 4326 94825 4378
rect 94825 4326 94839 4378
rect 94863 4326 94877 4378
rect 94877 4326 94889 4378
rect 94889 4326 94919 4378
rect 94943 4326 94953 4378
rect 94953 4326 94999 4378
rect 94703 4324 94759 4326
rect 94783 4324 94839 4326
rect 94863 4324 94919 4326
rect 94943 4324 94999 4326
rect 94703 3290 94759 3292
rect 94783 3290 94839 3292
rect 94863 3290 94919 3292
rect 94943 3290 94999 3292
rect 94703 3238 94749 3290
rect 94749 3238 94759 3290
rect 94783 3238 94813 3290
rect 94813 3238 94825 3290
rect 94825 3238 94839 3290
rect 94863 3238 94877 3290
rect 94877 3238 94889 3290
rect 94889 3238 94919 3290
rect 94943 3238 94953 3290
rect 94953 3238 94999 3290
rect 94703 3236 94759 3238
rect 94783 3236 94839 3238
rect 94863 3236 94919 3238
rect 94943 3236 94999 3238
rect 93766 2624 93822 2680
rect 24392 2202 24448 2204
rect 24472 2202 24528 2204
rect 24552 2202 24608 2204
rect 24632 2202 24688 2204
rect 24392 2150 24438 2202
rect 24438 2150 24448 2202
rect 24472 2150 24502 2202
rect 24502 2150 24514 2202
rect 24514 2150 24528 2202
rect 24552 2150 24566 2202
rect 24566 2150 24578 2202
rect 24578 2150 24608 2202
rect 24632 2150 24642 2202
rect 24642 2150 24688 2202
rect 24392 2148 24448 2150
rect 24472 2148 24528 2150
rect 24552 2148 24608 2150
rect 24632 2148 24688 2150
rect 47829 2202 47885 2204
rect 47909 2202 47965 2204
rect 47989 2202 48045 2204
rect 48069 2202 48125 2204
rect 47829 2150 47875 2202
rect 47875 2150 47885 2202
rect 47909 2150 47939 2202
rect 47939 2150 47951 2202
rect 47951 2150 47965 2202
rect 47989 2150 48003 2202
rect 48003 2150 48015 2202
rect 48015 2150 48045 2202
rect 48069 2150 48079 2202
rect 48079 2150 48125 2202
rect 47829 2148 47885 2150
rect 47909 2148 47965 2150
rect 47989 2148 48045 2150
rect 48069 2148 48125 2150
rect 71266 2202 71322 2204
rect 71346 2202 71402 2204
rect 71426 2202 71482 2204
rect 71506 2202 71562 2204
rect 71266 2150 71312 2202
rect 71312 2150 71322 2202
rect 71346 2150 71376 2202
rect 71376 2150 71388 2202
rect 71388 2150 71402 2202
rect 71426 2150 71440 2202
rect 71440 2150 71452 2202
rect 71452 2150 71482 2202
rect 71506 2150 71516 2202
rect 71516 2150 71562 2202
rect 71266 2148 71322 2150
rect 71346 2148 71402 2150
rect 71426 2148 71482 2150
rect 71506 2148 71562 2150
rect 94703 2202 94759 2204
rect 94783 2202 94839 2204
rect 94863 2202 94919 2204
rect 94943 2202 94999 2204
rect 94703 2150 94749 2202
rect 94749 2150 94759 2202
rect 94783 2150 94813 2202
rect 94813 2150 94825 2202
rect 94825 2150 94839 2202
rect 94863 2150 94877 2202
rect 94877 2150 94889 2202
rect 94889 2150 94919 2202
rect 94943 2150 94953 2202
rect 94953 2150 94999 2202
rect 94703 2148 94759 2150
rect 94783 2148 94839 2150
rect 94863 2148 94919 2150
rect 94943 2148 94999 2150
<< metal3 >>
rect 24382 17440 24698 17441
rect 24382 17376 24388 17440
rect 24452 17376 24468 17440
rect 24532 17376 24548 17440
rect 24612 17376 24628 17440
rect 24692 17376 24698 17440
rect 24382 17375 24698 17376
rect 47819 17440 48135 17441
rect 47819 17376 47825 17440
rect 47889 17376 47905 17440
rect 47969 17376 47985 17440
rect 48049 17376 48065 17440
rect 48129 17376 48135 17440
rect 47819 17375 48135 17376
rect 71256 17440 71572 17441
rect 71256 17376 71262 17440
rect 71326 17376 71342 17440
rect 71406 17376 71422 17440
rect 71486 17376 71502 17440
rect 71566 17376 71572 17440
rect 71256 17375 71572 17376
rect 94693 17440 95009 17441
rect 94693 17376 94699 17440
rect 94763 17376 94779 17440
rect 94843 17376 94859 17440
rect 94923 17376 94939 17440
rect 95003 17376 95009 17440
rect 94693 17375 95009 17376
rect 95200 17280 96000 17400
rect 12664 16896 12980 16897
rect 12664 16832 12670 16896
rect 12734 16832 12750 16896
rect 12814 16832 12830 16896
rect 12894 16832 12910 16896
rect 12974 16832 12980 16896
rect 12664 16831 12980 16832
rect 36101 16896 36417 16897
rect 36101 16832 36107 16896
rect 36171 16832 36187 16896
rect 36251 16832 36267 16896
rect 36331 16832 36347 16896
rect 36411 16832 36417 16896
rect 36101 16831 36417 16832
rect 59538 16896 59854 16897
rect 59538 16832 59544 16896
rect 59608 16832 59624 16896
rect 59688 16832 59704 16896
rect 59768 16832 59784 16896
rect 59848 16832 59854 16896
rect 59538 16831 59854 16832
rect 82975 16896 83291 16897
rect 82975 16832 82981 16896
rect 83045 16832 83061 16896
rect 83125 16832 83141 16896
rect 83205 16832 83221 16896
rect 83285 16832 83291 16896
rect 82975 16831 83291 16832
rect 94221 16826 94287 16829
rect 95374 16826 95434 17280
rect 94221 16824 95434 16826
rect 94221 16768 94226 16824
rect 94282 16768 95434 16824
rect 94221 16766 95434 16768
rect 94221 16763 94287 16766
rect 0 16690 800 16720
rect 1577 16690 1643 16693
rect 0 16688 1643 16690
rect 0 16632 1582 16688
rect 1638 16632 1643 16688
rect 0 16630 1643 16632
rect 0 16600 800 16630
rect 1577 16627 1643 16630
rect 42333 16554 42399 16557
rect 46105 16554 46171 16557
rect 42333 16552 46171 16554
rect 42333 16496 42338 16552
rect 42394 16496 46110 16552
rect 46166 16496 46171 16552
rect 42333 16494 46171 16496
rect 42333 16491 42399 16494
rect 46105 16491 46171 16494
rect 24382 16352 24698 16353
rect 24382 16288 24388 16352
rect 24452 16288 24468 16352
rect 24532 16288 24548 16352
rect 24612 16288 24628 16352
rect 24692 16288 24698 16352
rect 24382 16287 24698 16288
rect 47819 16352 48135 16353
rect 47819 16288 47825 16352
rect 47889 16288 47905 16352
rect 47969 16288 47985 16352
rect 48049 16288 48065 16352
rect 48129 16288 48135 16352
rect 47819 16287 48135 16288
rect 71256 16352 71572 16353
rect 71256 16288 71262 16352
rect 71326 16288 71342 16352
rect 71406 16288 71422 16352
rect 71486 16288 71502 16352
rect 71566 16288 71572 16352
rect 71256 16287 71572 16288
rect 94693 16352 95009 16353
rect 94693 16288 94699 16352
rect 94763 16288 94779 16352
rect 94843 16288 94859 16352
rect 94923 16288 94939 16352
rect 95003 16288 95009 16352
rect 94693 16287 95009 16288
rect 44633 16146 44699 16149
rect 86309 16146 86375 16149
rect 44633 16144 86375 16146
rect 44633 16088 44638 16144
rect 44694 16088 86314 16144
rect 86370 16088 86375 16144
rect 44633 16086 86375 16088
rect 44633 16083 44699 16086
rect 86309 16083 86375 16086
rect 20345 16010 20411 16013
rect 40769 16010 40835 16013
rect 20345 16008 40835 16010
rect 20345 15952 20350 16008
rect 20406 15952 40774 16008
rect 40830 15952 40835 16008
rect 20345 15950 40835 15952
rect 20345 15947 20411 15950
rect 40769 15947 40835 15950
rect 52361 16010 52427 16013
rect 82169 16010 82235 16013
rect 52361 16008 82235 16010
rect 52361 15952 52366 16008
rect 52422 15952 82174 16008
rect 82230 15952 82235 16008
rect 52361 15950 82235 15952
rect 52361 15947 52427 15950
rect 82169 15947 82235 15950
rect 12664 15808 12980 15809
rect 12664 15744 12670 15808
rect 12734 15744 12750 15808
rect 12814 15744 12830 15808
rect 12894 15744 12910 15808
rect 12974 15744 12980 15808
rect 12664 15743 12980 15744
rect 36101 15808 36417 15809
rect 36101 15744 36107 15808
rect 36171 15744 36187 15808
rect 36251 15744 36267 15808
rect 36331 15744 36347 15808
rect 36411 15744 36417 15808
rect 36101 15743 36417 15744
rect 59538 15808 59854 15809
rect 59538 15744 59544 15808
rect 59608 15744 59624 15808
rect 59688 15744 59704 15808
rect 59768 15744 59784 15808
rect 59848 15744 59854 15808
rect 59538 15743 59854 15744
rect 82975 15808 83291 15809
rect 82975 15744 82981 15808
rect 83045 15744 83061 15808
rect 83125 15744 83141 15808
rect 83205 15744 83221 15808
rect 83285 15744 83291 15808
rect 82975 15743 83291 15744
rect 44081 15738 44147 15741
rect 47945 15738 48011 15741
rect 44081 15736 48011 15738
rect 44081 15680 44086 15736
rect 44142 15680 47950 15736
rect 48006 15680 48011 15736
rect 44081 15678 48011 15680
rect 44081 15675 44147 15678
rect 47945 15675 48011 15678
rect 16941 15602 17007 15605
rect 35893 15602 35959 15605
rect 16941 15600 35959 15602
rect 16941 15544 16946 15600
rect 17002 15544 35898 15600
rect 35954 15544 35959 15600
rect 16941 15542 35959 15544
rect 16941 15539 17007 15542
rect 35893 15539 35959 15542
rect 40769 15602 40835 15605
rect 56961 15602 57027 15605
rect 40769 15600 57027 15602
rect 40769 15544 40774 15600
rect 40830 15544 56966 15600
rect 57022 15544 57027 15600
rect 40769 15542 57027 15544
rect 40769 15539 40835 15542
rect 56961 15539 57027 15542
rect 34881 15466 34947 15469
rect 35341 15466 35407 15469
rect 48773 15466 48839 15469
rect 34881 15464 48839 15466
rect 34881 15408 34886 15464
rect 34942 15408 35346 15464
rect 35402 15408 48778 15464
rect 48834 15408 48839 15464
rect 34881 15406 48839 15408
rect 34881 15403 34947 15406
rect 35341 15403 35407 15406
rect 48773 15403 48839 15406
rect 64689 15466 64755 15469
rect 77845 15466 77911 15469
rect 64689 15464 77911 15466
rect 64689 15408 64694 15464
rect 64750 15408 77850 15464
rect 77906 15408 77911 15464
rect 64689 15406 77911 15408
rect 64689 15403 64755 15406
rect 77845 15403 77911 15406
rect 29545 15330 29611 15333
rect 34697 15330 34763 15333
rect 35801 15330 35867 15333
rect 29545 15328 35910 15330
rect 29545 15272 29550 15328
rect 29606 15272 34702 15328
rect 34758 15272 35806 15328
rect 35862 15272 35910 15328
rect 29545 15270 35910 15272
rect 29545 15267 29611 15270
rect 34697 15267 34763 15270
rect 35801 15267 35910 15270
rect 24382 15264 24698 15265
rect 24382 15200 24388 15264
rect 24452 15200 24468 15264
rect 24532 15200 24548 15264
rect 24612 15200 24628 15264
rect 24692 15200 24698 15264
rect 24382 15199 24698 15200
rect 35850 15194 35910 15267
rect 47819 15264 48135 15265
rect 47819 15200 47825 15264
rect 47889 15200 47905 15264
rect 47969 15200 47985 15264
rect 48049 15200 48065 15264
rect 48129 15200 48135 15264
rect 47819 15199 48135 15200
rect 71256 15264 71572 15265
rect 71256 15200 71262 15264
rect 71326 15200 71342 15264
rect 71406 15200 71422 15264
rect 71486 15200 71502 15264
rect 71566 15200 71572 15264
rect 71256 15199 71572 15200
rect 94693 15264 95009 15265
rect 94693 15200 94699 15264
rect 94763 15200 94779 15264
rect 94843 15200 94859 15264
rect 94923 15200 94939 15264
rect 95003 15200 95009 15264
rect 94693 15199 95009 15200
rect 59077 15194 59143 15197
rect 35850 15134 46306 15194
rect 13905 15058 13971 15061
rect 42425 15058 42491 15061
rect 13905 15056 42491 15058
rect 13905 15000 13910 15056
rect 13966 15000 42430 15056
rect 42486 15000 42491 15056
rect 13905 14998 42491 15000
rect 46246 15058 46306 15134
rect 51030 15192 59143 15194
rect 51030 15136 59082 15192
rect 59138 15136 59143 15192
rect 51030 15134 59143 15136
rect 51030 15058 51090 15134
rect 59077 15131 59143 15134
rect 46246 14998 51090 15058
rect 53833 15058 53899 15061
rect 78673 15058 78739 15061
rect 53833 15056 78739 15058
rect 53833 15000 53838 15056
rect 53894 15000 78678 15056
rect 78734 15000 78739 15056
rect 53833 14998 78739 15000
rect 13905 14995 13971 14998
rect 42425 14995 42491 14998
rect 53833 14995 53899 14998
rect 78673 14995 78739 14998
rect 12709 14922 12775 14925
rect 40953 14922 41019 14925
rect 12709 14920 41019 14922
rect 12709 14864 12714 14920
rect 12770 14864 40958 14920
rect 41014 14864 41019 14920
rect 12709 14862 41019 14864
rect 12709 14859 12775 14862
rect 40953 14859 41019 14862
rect 50337 14922 50403 14925
rect 75269 14922 75335 14925
rect 50337 14920 75335 14922
rect 50337 14864 50342 14920
rect 50398 14864 75274 14920
rect 75330 14864 75335 14920
rect 50337 14862 75335 14864
rect 50337 14859 50403 14862
rect 75269 14859 75335 14862
rect 25589 14786 25655 14789
rect 35065 14786 35131 14789
rect 25589 14784 35131 14786
rect 25589 14728 25594 14784
rect 25650 14728 35070 14784
rect 35126 14728 35131 14784
rect 25589 14726 35131 14728
rect 25589 14723 25655 14726
rect 35065 14723 35131 14726
rect 12664 14720 12980 14721
rect 12664 14656 12670 14720
rect 12734 14656 12750 14720
rect 12814 14656 12830 14720
rect 12894 14656 12910 14720
rect 12974 14656 12980 14720
rect 12664 14655 12980 14656
rect 36101 14720 36417 14721
rect 36101 14656 36107 14720
rect 36171 14656 36187 14720
rect 36251 14656 36267 14720
rect 36331 14656 36347 14720
rect 36411 14656 36417 14720
rect 36101 14655 36417 14656
rect 59538 14720 59854 14721
rect 59538 14656 59544 14720
rect 59608 14656 59624 14720
rect 59688 14656 59704 14720
rect 59768 14656 59784 14720
rect 59848 14656 59854 14720
rect 59538 14655 59854 14656
rect 82975 14720 83291 14721
rect 82975 14656 82981 14720
rect 83045 14656 83061 14720
rect 83125 14656 83141 14720
rect 83205 14656 83221 14720
rect 83285 14656 83291 14720
rect 82975 14655 83291 14656
rect 29637 14650 29703 14653
rect 31753 14650 31819 14653
rect 29637 14648 31819 14650
rect 29637 14592 29642 14648
rect 29698 14592 31758 14648
rect 31814 14592 31819 14648
rect 29637 14590 31819 14592
rect 29637 14587 29703 14590
rect 31753 14587 31819 14590
rect 41229 14650 41295 14653
rect 43805 14650 43871 14653
rect 41229 14648 43871 14650
rect 41229 14592 41234 14648
rect 41290 14592 43810 14648
rect 43866 14592 43871 14648
rect 41229 14590 43871 14592
rect 41229 14587 41295 14590
rect 43805 14587 43871 14590
rect 29453 14514 29519 14517
rect 35065 14514 35131 14517
rect 29453 14512 35131 14514
rect 29453 14456 29458 14512
rect 29514 14456 35070 14512
rect 35126 14456 35131 14512
rect 29453 14454 35131 14456
rect 29453 14451 29519 14454
rect 35065 14451 35131 14454
rect 40585 14514 40651 14517
rect 68461 14514 68527 14517
rect 40585 14512 68527 14514
rect 40585 14456 40590 14512
rect 40646 14456 68466 14512
rect 68522 14456 68527 14512
rect 40585 14454 68527 14456
rect 40585 14451 40651 14454
rect 68461 14451 68527 14454
rect 13077 14378 13143 14381
rect 48313 14378 48379 14381
rect 13077 14376 48379 14378
rect 13077 14320 13082 14376
rect 13138 14320 48318 14376
rect 48374 14320 48379 14376
rect 13077 14318 48379 14320
rect 13077 14315 13143 14318
rect 48313 14315 48379 14318
rect 51349 14378 51415 14381
rect 68185 14378 68251 14381
rect 51349 14376 68251 14378
rect 51349 14320 51354 14376
rect 51410 14320 68190 14376
rect 68246 14320 68251 14376
rect 51349 14318 68251 14320
rect 51349 14315 51415 14318
rect 68185 14315 68251 14318
rect 29821 14242 29887 14245
rect 37089 14242 37155 14245
rect 29821 14240 37155 14242
rect 29821 14184 29826 14240
rect 29882 14184 37094 14240
rect 37150 14184 37155 14240
rect 29821 14182 37155 14184
rect 29821 14179 29887 14182
rect 37089 14179 37155 14182
rect 41413 14242 41479 14245
rect 47025 14242 47091 14245
rect 41413 14240 47091 14242
rect 41413 14184 41418 14240
rect 41474 14184 47030 14240
rect 47086 14184 47091 14240
rect 41413 14182 47091 14184
rect 41413 14179 41479 14182
rect 47025 14179 47091 14182
rect 60641 14242 60707 14245
rect 66069 14242 66135 14245
rect 60641 14240 66135 14242
rect 60641 14184 60646 14240
rect 60702 14184 66074 14240
rect 66130 14184 66135 14240
rect 60641 14182 66135 14184
rect 60641 14179 60707 14182
rect 66069 14179 66135 14182
rect 24382 14176 24698 14177
rect 24382 14112 24388 14176
rect 24452 14112 24468 14176
rect 24532 14112 24548 14176
rect 24612 14112 24628 14176
rect 24692 14112 24698 14176
rect 24382 14111 24698 14112
rect 47819 14176 48135 14177
rect 47819 14112 47825 14176
rect 47889 14112 47905 14176
rect 47969 14112 47985 14176
rect 48049 14112 48065 14176
rect 48129 14112 48135 14176
rect 47819 14111 48135 14112
rect 71256 14176 71572 14177
rect 71256 14112 71262 14176
rect 71326 14112 71342 14176
rect 71406 14112 71422 14176
rect 71486 14112 71502 14176
rect 71566 14112 71572 14176
rect 71256 14111 71572 14112
rect 94693 14176 95009 14177
rect 94693 14112 94699 14176
rect 94763 14112 94779 14176
rect 94843 14112 94859 14176
rect 94923 14112 94939 14176
rect 95003 14112 95009 14176
rect 94693 14111 95009 14112
rect 13169 14106 13235 14109
rect 24209 14106 24275 14109
rect 13169 14104 24275 14106
rect 13169 14048 13174 14104
rect 13230 14048 24214 14104
rect 24270 14048 24275 14104
rect 13169 14046 24275 14048
rect 13169 14043 13235 14046
rect 24209 14043 24275 14046
rect 24761 14106 24827 14109
rect 42241 14106 42307 14109
rect 24761 14104 42307 14106
rect 24761 14048 24766 14104
rect 24822 14048 42246 14104
rect 42302 14048 42307 14104
rect 24761 14046 42307 14048
rect 24761 14043 24827 14046
rect 42241 14043 42307 14046
rect 57973 14106 58039 14109
rect 63217 14106 63283 14109
rect 67449 14106 67515 14109
rect 57973 14104 61946 14106
rect 57973 14048 57978 14104
rect 58034 14048 61946 14104
rect 57973 14046 61946 14048
rect 57973 14043 58039 14046
rect 15009 13970 15075 13973
rect 54845 13970 54911 13973
rect 15009 13968 54911 13970
rect 15009 13912 15014 13968
rect 15070 13912 54850 13968
rect 54906 13912 54911 13968
rect 15009 13910 54911 13912
rect 15009 13907 15075 13910
rect 54845 13907 54911 13910
rect 59169 13970 59235 13973
rect 61653 13970 61719 13973
rect 59169 13968 61719 13970
rect 59169 13912 59174 13968
rect 59230 13912 61658 13968
rect 61714 13912 61719 13968
rect 59169 13910 61719 13912
rect 61886 13970 61946 14046
rect 63217 14104 67515 14106
rect 63217 14048 63222 14104
rect 63278 14048 67454 14104
rect 67510 14048 67515 14104
rect 63217 14046 67515 14048
rect 63217 14043 63283 14046
rect 67449 14043 67515 14046
rect 72601 14106 72667 14109
rect 88149 14106 88215 14109
rect 72601 14104 88215 14106
rect 72601 14048 72606 14104
rect 72662 14048 88154 14104
rect 88210 14048 88215 14104
rect 72601 14046 88215 14048
rect 72601 14043 72667 14046
rect 88149 14043 88215 14046
rect 66437 13970 66503 13973
rect 61886 13968 66503 13970
rect 61886 13912 66442 13968
rect 66498 13912 66503 13968
rect 61886 13910 66503 13912
rect 59169 13907 59235 13910
rect 61653 13907 61719 13910
rect 66437 13907 66503 13910
rect 70669 13970 70735 13973
rect 73797 13970 73863 13973
rect 70669 13968 73863 13970
rect 70669 13912 70674 13968
rect 70730 13912 73802 13968
rect 73858 13912 73863 13968
rect 70669 13910 73863 13912
rect 70669 13907 70735 13910
rect 73797 13907 73863 13910
rect 11973 13834 12039 13837
rect 80697 13834 80763 13837
rect 11973 13832 80763 13834
rect 11973 13776 11978 13832
rect 12034 13776 80702 13832
rect 80758 13776 80763 13832
rect 11973 13774 80763 13776
rect 11973 13771 12039 13774
rect 80697 13771 80763 13774
rect 20437 13698 20503 13701
rect 35617 13698 35683 13701
rect 20437 13696 35683 13698
rect 20437 13640 20442 13696
rect 20498 13640 35622 13696
rect 35678 13640 35683 13696
rect 20437 13638 35683 13640
rect 20437 13635 20503 13638
rect 35617 13635 35683 13638
rect 36721 13698 36787 13701
rect 45737 13698 45803 13701
rect 36721 13696 45803 13698
rect 36721 13640 36726 13696
rect 36782 13640 45742 13696
rect 45798 13640 45803 13696
rect 36721 13638 45803 13640
rect 36721 13635 36787 13638
rect 45737 13635 45803 13638
rect 60641 13698 60707 13701
rect 64689 13698 64755 13701
rect 60641 13696 64755 13698
rect 60641 13640 60646 13696
rect 60702 13640 64694 13696
rect 64750 13640 64755 13696
rect 60641 13638 64755 13640
rect 60641 13635 60707 13638
rect 64689 13635 64755 13638
rect 68461 13698 68527 13701
rect 75729 13698 75795 13701
rect 68461 13696 75795 13698
rect 68461 13640 68466 13696
rect 68522 13640 75734 13696
rect 75790 13640 75795 13696
rect 68461 13638 75795 13640
rect 68461 13635 68527 13638
rect 75729 13635 75795 13638
rect 12664 13632 12980 13633
rect 12664 13568 12670 13632
rect 12734 13568 12750 13632
rect 12814 13568 12830 13632
rect 12894 13568 12910 13632
rect 12974 13568 12980 13632
rect 12664 13567 12980 13568
rect 36101 13632 36417 13633
rect 36101 13568 36107 13632
rect 36171 13568 36187 13632
rect 36251 13568 36267 13632
rect 36331 13568 36347 13632
rect 36411 13568 36417 13632
rect 36101 13567 36417 13568
rect 59538 13632 59854 13633
rect 59538 13568 59544 13632
rect 59608 13568 59624 13632
rect 59688 13568 59704 13632
rect 59768 13568 59784 13632
rect 59848 13568 59854 13632
rect 59538 13567 59854 13568
rect 82975 13632 83291 13633
rect 82975 13568 82981 13632
rect 83045 13568 83061 13632
rect 83125 13568 83141 13632
rect 83205 13568 83221 13632
rect 83285 13568 83291 13632
rect 82975 13567 83291 13568
rect 29637 13562 29703 13565
rect 30925 13562 30991 13565
rect 29637 13560 30991 13562
rect 29637 13504 29642 13560
rect 29698 13504 30930 13560
rect 30986 13504 30991 13560
rect 29637 13502 30991 13504
rect 29637 13499 29703 13502
rect 30925 13499 30991 13502
rect 60365 13562 60431 13565
rect 66713 13562 66779 13565
rect 60365 13560 66779 13562
rect 60365 13504 60370 13560
rect 60426 13504 66718 13560
rect 66774 13504 66779 13560
rect 60365 13502 66779 13504
rect 60365 13499 60431 13502
rect 66713 13499 66779 13502
rect 68277 13562 68343 13565
rect 73245 13562 73311 13565
rect 68277 13560 73311 13562
rect 68277 13504 68282 13560
rect 68338 13504 73250 13560
rect 73306 13504 73311 13560
rect 68277 13502 73311 13504
rect 68277 13499 68343 13502
rect 73245 13499 73311 13502
rect 4797 13426 4863 13429
rect 69749 13426 69815 13429
rect 4797 13424 69815 13426
rect 4797 13368 4802 13424
rect 4858 13368 69754 13424
rect 69810 13368 69815 13424
rect 4797 13366 69815 13368
rect 4797 13363 4863 13366
rect 69749 13363 69815 13366
rect 71129 13426 71195 13429
rect 77017 13426 77083 13429
rect 77477 13426 77543 13429
rect 71129 13424 77543 13426
rect 71129 13368 71134 13424
rect 71190 13368 77022 13424
rect 77078 13368 77482 13424
rect 77538 13368 77543 13424
rect 71129 13366 77543 13368
rect 71129 13363 71195 13366
rect 77017 13363 77083 13366
rect 77477 13363 77543 13366
rect 22093 13290 22159 13293
rect 42885 13290 42951 13293
rect 56317 13290 56383 13293
rect 92473 13290 92539 13293
rect 22093 13288 42951 13290
rect 22093 13232 22098 13288
rect 22154 13232 42890 13288
rect 42946 13232 42951 13288
rect 22093 13230 42951 13232
rect 22093 13227 22159 13230
rect 42885 13227 42951 13230
rect 43118 13230 51090 13290
rect 31109 13154 31175 13157
rect 37457 13154 37523 13157
rect 31109 13152 37523 13154
rect 31109 13096 31114 13152
rect 31170 13096 37462 13152
rect 37518 13096 37523 13152
rect 31109 13094 37523 13096
rect 31109 13091 31175 13094
rect 37457 13091 37523 13094
rect 41781 13154 41847 13157
rect 43118 13154 43178 13230
rect 41781 13152 43178 13154
rect 41781 13096 41786 13152
rect 41842 13096 43178 13152
rect 41781 13094 43178 13096
rect 51030 13154 51090 13230
rect 56317 13288 92539 13290
rect 56317 13232 56322 13288
rect 56378 13232 92478 13288
rect 92534 13232 92539 13288
rect 56317 13230 92539 13232
rect 56317 13227 56383 13230
rect 92473 13227 92539 13230
rect 52085 13154 52151 13157
rect 60222 13154 60228 13156
rect 51030 13152 60228 13154
rect 51030 13096 52090 13152
rect 52146 13096 60228 13152
rect 51030 13094 60228 13096
rect 41781 13091 41847 13094
rect 52085 13091 52151 13094
rect 60222 13092 60228 13094
rect 60292 13092 60298 13156
rect 61285 13154 61351 13157
rect 67909 13154 67975 13157
rect 61285 13152 67975 13154
rect 61285 13096 61290 13152
rect 61346 13096 67914 13152
rect 67970 13096 67975 13152
rect 61285 13094 67975 13096
rect 61285 13091 61351 13094
rect 67909 13091 67975 13094
rect 71957 13154 72023 13157
rect 77017 13154 77083 13157
rect 71957 13152 77083 13154
rect 71957 13096 71962 13152
rect 72018 13096 77022 13152
rect 77078 13096 77083 13152
rect 71957 13094 77083 13096
rect 71957 13091 72023 13094
rect 77017 13091 77083 13094
rect 79409 13154 79475 13157
rect 82261 13154 82327 13157
rect 79409 13152 82327 13154
rect 79409 13096 79414 13152
rect 79470 13096 82266 13152
rect 82322 13096 82327 13152
rect 79409 13094 82327 13096
rect 79409 13091 79475 13094
rect 82261 13091 82327 13094
rect 24382 13088 24698 13089
rect 24382 13024 24388 13088
rect 24452 13024 24468 13088
rect 24532 13024 24548 13088
rect 24612 13024 24628 13088
rect 24692 13024 24698 13088
rect 24382 13023 24698 13024
rect 47819 13088 48135 13089
rect 47819 13024 47825 13088
rect 47889 13024 47905 13088
rect 47969 13024 47985 13088
rect 48049 13024 48065 13088
rect 48129 13024 48135 13088
rect 47819 13023 48135 13024
rect 71256 13088 71572 13089
rect 71256 13024 71262 13088
rect 71326 13024 71342 13088
rect 71406 13024 71422 13088
rect 71486 13024 71502 13088
rect 71566 13024 71572 13088
rect 71256 13023 71572 13024
rect 94693 13088 95009 13089
rect 94693 13024 94699 13088
rect 94763 13024 94779 13088
rect 94843 13024 94859 13088
rect 94923 13024 94939 13088
rect 95003 13024 95009 13088
rect 94693 13023 95009 13024
rect 28257 13018 28323 13021
rect 38009 13018 38075 13021
rect 28257 13016 38075 13018
rect 28257 12960 28262 13016
rect 28318 12960 38014 13016
rect 38070 12960 38075 13016
rect 28257 12958 38075 12960
rect 28257 12955 28323 12958
rect 38009 12955 38075 12958
rect 55673 13018 55739 13021
rect 60181 13018 60247 13021
rect 55673 13016 60247 13018
rect 55673 12960 55678 13016
rect 55734 12960 60186 13016
rect 60242 12960 60247 13016
rect 55673 12958 60247 12960
rect 55673 12955 55739 12958
rect 60181 12955 60247 12958
rect 62021 13018 62087 13021
rect 67173 13018 67239 13021
rect 62021 13016 67239 13018
rect 62021 12960 62026 13016
rect 62082 12960 67178 13016
rect 67234 12960 67239 13016
rect 62021 12958 67239 12960
rect 62021 12955 62087 12958
rect 67173 12955 67239 12958
rect 71681 13018 71747 13021
rect 77109 13018 77175 13021
rect 71681 13016 77175 13018
rect 71681 12960 71686 13016
rect 71742 12960 77114 13016
rect 77170 12960 77175 13016
rect 71681 12958 77175 12960
rect 71681 12955 71747 12958
rect 77109 12955 77175 12958
rect 29821 12882 29887 12885
rect 32581 12882 32647 12885
rect 29821 12880 32647 12882
rect 29821 12824 29826 12880
rect 29882 12824 32586 12880
rect 32642 12824 32647 12880
rect 29821 12822 32647 12824
rect 29821 12819 29887 12822
rect 32581 12819 32647 12822
rect 35525 12882 35591 12885
rect 89437 12882 89503 12885
rect 35525 12880 89503 12882
rect 35525 12824 35530 12880
rect 35586 12824 89442 12880
rect 89498 12824 89503 12880
rect 35525 12822 89503 12824
rect 35525 12819 35591 12822
rect 89437 12819 89503 12822
rect 7005 12746 7071 12749
rect 48221 12746 48287 12749
rect 7005 12744 48287 12746
rect 7005 12688 7010 12744
rect 7066 12688 48226 12744
rect 48282 12688 48287 12744
rect 7005 12686 48287 12688
rect 7005 12683 7071 12686
rect 48221 12683 48287 12686
rect 55814 12686 60060 12746
rect 40585 12610 40651 12613
rect 55673 12610 55739 12613
rect 40585 12608 55739 12610
rect 40585 12552 40590 12608
rect 40646 12552 55678 12608
rect 55734 12552 55739 12608
rect 40585 12550 55739 12552
rect 40585 12547 40651 12550
rect 55673 12547 55739 12550
rect 12664 12544 12980 12545
rect 12664 12480 12670 12544
rect 12734 12480 12750 12544
rect 12814 12480 12830 12544
rect 12894 12480 12910 12544
rect 12974 12480 12980 12544
rect 12664 12479 12980 12480
rect 36101 12544 36417 12545
rect 36101 12480 36107 12544
rect 36171 12480 36187 12544
rect 36251 12480 36267 12544
rect 36331 12480 36347 12544
rect 36411 12480 36417 12544
rect 36101 12479 36417 12480
rect 39021 12474 39087 12477
rect 55814 12474 55874 12686
rect 59538 12544 59854 12545
rect 59538 12480 59544 12544
rect 59608 12480 59624 12544
rect 59688 12480 59704 12544
rect 59768 12480 59784 12544
rect 59848 12480 59854 12544
rect 59538 12479 59854 12480
rect 39021 12472 55874 12474
rect 39021 12416 39026 12472
rect 39082 12416 55874 12472
rect 39021 12414 55874 12416
rect 56133 12474 56199 12477
rect 57697 12474 57763 12477
rect 56133 12472 57763 12474
rect 56133 12416 56138 12472
rect 56194 12416 57702 12472
rect 57758 12416 57763 12472
rect 56133 12414 57763 12416
rect 60000 12474 60060 12686
rect 60222 12684 60228 12748
rect 60292 12746 60298 12748
rect 86861 12746 86927 12749
rect 60292 12744 86927 12746
rect 60292 12688 86866 12744
rect 86922 12688 86927 12744
rect 60292 12686 86927 12688
rect 60292 12684 60298 12686
rect 86861 12683 86927 12686
rect 60181 12610 60247 12613
rect 71129 12610 71195 12613
rect 60181 12608 71195 12610
rect 60181 12552 60186 12608
rect 60242 12552 71134 12608
rect 71190 12552 71195 12608
rect 60181 12550 71195 12552
rect 60181 12547 60247 12550
rect 71129 12547 71195 12550
rect 71313 12610 71379 12613
rect 72417 12610 72483 12613
rect 71313 12608 72483 12610
rect 71313 12552 71318 12608
rect 71374 12552 72422 12608
rect 72478 12552 72483 12608
rect 71313 12550 72483 12552
rect 71313 12547 71379 12550
rect 72417 12547 72483 12550
rect 82975 12544 83291 12545
rect 82975 12480 82981 12544
rect 83045 12480 83061 12544
rect 83125 12480 83141 12544
rect 83205 12480 83221 12544
rect 83285 12480 83291 12544
rect 82975 12479 83291 12480
rect 69565 12474 69631 12477
rect 60000 12472 69631 12474
rect 60000 12416 69570 12472
rect 69626 12416 69631 12472
rect 60000 12414 69631 12416
rect 39021 12411 39087 12414
rect 56133 12411 56199 12414
rect 57697 12411 57763 12414
rect 69565 12411 69631 12414
rect 71037 12474 71103 12477
rect 75177 12474 75243 12477
rect 71037 12472 75243 12474
rect 71037 12416 71042 12472
rect 71098 12416 75182 12472
rect 75238 12416 75243 12472
rect 71037 12414 75243 12416
rect 71037 12411 71103 12414
rect 75177 12411 75243 12414
rect 94221 12474 94287 12477
rect 95200 12474 96000 12504
rect 94221 12472 96000 12474
rect 94221 12416 94226 12472
rect 94282 12416 96000 12472
rect 94221 12414 96000 12416
rect 94221 12411 94287 12414
rect 95200 12384 96000 12414
rect 24025 12338 24091 12341
rect 27061 12338 27127 12341
rect 24025 12336 27127 12338
rect 24025 12280 24030 12336
rect 24086 12280 27066 12336
rect 27122 12280 27127 12336
rect 24025 12278 27127 12280
rect 24025 12275 24091 12278
rect 27061 12275 27127 12278
rect 27889 12338 27955 12341
rect 32121 12338 32187 12341
rect 37825 12338 37891 12341
rect 27889 12336 32187 12338
rect 27889 12280 27894 12336
rect 27950 12280 32126 12336
rect 32182 12280 32187 12336
rect 27889 12278 32187 12280
rect 27889 12275 27955 12278
rect 32121 12275 32187 12278
rect 32262 12336 37891 12338
rect 32262 12280 37830 12336
rect 37886 12280 37891 12336
rect 32262 12278 37891 12280
rect 28993 12202 29059 12205
rect 32262 12202 32322 12278
rect 37825 12275 37891 12278
rect 42333 12338 42399 12341
rect 59905 12338 59971 12341
rect 42333 12336 59971 12338
rect 42333 12280 42338 12336
rect 42394 12280 59910 12336
rect 59966 12280 59971 12336
rect 42333 12278 59971 12280
rect 42333 12275 42399 12278
rect 59905 12275 59971 12278
rect 60641 12338 60707 12341
rect 63033 12338 63099 12341
rect 60641 12336 63099 12338
rect 60641 12280 60646 12336
rect 60702 12280 63038 12336
rect 63094 12280 63099 12336
rect 60641 12278 63099 12280
rect 60641 12275 60707 12278
rect 63033 12275 63099 12278
rect 72601 12338 72667 12341
rect 74625 12338 74691 12341
rect 77569 12338 77635 12341
rect 72601 12336 77635 12338
rect 72601 12280 72606 12336
rect 72662 12280 74630 12336
rect 74686 12280 77574 12336
rect 77630 12280 77635 12336
rect 72601 12278 77635 12280
rect 72601 12275 72667 12278
rect 74625 12275 74691 12278
rect 77569 12275 77635 12278
rect 28993 12200 32322 12202
rect 28993 12144 28998 12200
rect 29054 12144 32322 12200
rect 28993 12142 32322 12144
rect 36905 12202 36971 12205
rect 38929 12202 38995 12205
rect 36905 12200 38995 12202
rect 36905 12144 36910 12200
rect 36966 12144 38934 12200
rect 38990 12144 38995 12200
rect 36905 12142 38995 12144
rect 28993 12139 29059 12142
rect 36905 12139 36971 12142
rect 38929 12139 38995 12142
rect 44541 12202 44607 12205
rect 51349 12202 51415 12205
rect 44541 12200 51415 12202
rect 44541 12144 44546 12200
rect 44602 12144 51354 12200
rect 51410 12144 51415 12200
rect 44541 12142 51415 12144
rect 44541 12139 44607 12142
rect 51349 12139 51415 12142
rect 59169 12202 59235 12205
rect 61929 12202 61995 12205
rect 59169 12200 61995 12202
rect 59169 12144 59174 12200
rect 59230 12144 61934 12200
rect 61990 12144 61995 12200
rect 59169 12142 61995 12144
rect 59169 12139 59235 12142
rect 61929 12139 61995 12142
rect 64781 12202 64847 12205
rect 67541 12202 67607 12205
rect 64781 12200 67607 12202
rect 64781 12144 64786 12200
rect 64842 12144 67546 12200
rect 67602 12144 67607 12200
rect 64781 12142 67607 12144
rect 64781 12139 64847 12142
rect 67541 12139 67607 12142
rect 69473 12202 69539 12205
rect 72693 12202 72759 12205
rect 76373 12202 76439 12205
rect 69473 12200 72434 12202
rect 69473 12144 69478 12200
rect 69534 12144 72434 12200
rect 69473 12142 72434 12144
rect 69473 12139 69539 12142
rect 32397 12066 32463 12069
rect 41597 12066 41663 12069
rect 32397 12064 41663 12066
rect 32397 12008 32402 12064
rect 32458 12008 41602 12064
rect 41658 12008 41663 12064
rect 32397 12006 41663 12008
rect 32397 12003 32463 12006
rect 41597 12003 41663 12006
rect 43897 12066 43963 12069
rect 46749 12066 46815 12069
rect 43897 12064 46815 12066
rect 43897 12008 43902 12064
rect 43958 12008 46754 12064
rect 46810 12008 46815 12064
rect 43897 12006 46815 12008
rect 43897 12003 43963 12006
rect 46749 12003 46815 12006
rect 56593 12066 56659 12069
rect 58709 12066 58775 12069
rect 67081 12066 67147 12069
rect 56593 12064 67147 12066
rect 56593 12008 56598 12064
rect 56654 12008 58714 12064
rect 58770 12008 67086 12064
rect 67142 12008 67147 12064
rect 56593 12006 67147 12008
rect 56593 12003 56659 12006
rect 58709 12003 58775 12006
rect 67081 12003 67147 12006
rect 24382 12000 24698 12001
rect 24382 11936 24388 12000
rect 24452 11936 24468 12000
rect 24532 11936 24548 12000
rect 24612 11936 24628 12000
rect 24692 11936 24698 12000
rect 24382 11935 24698 11936
rect 47819 12000 48135 12001
rect 47819 11936 47825 12000
rect 47889 11936 47905 12000
rect 47969 11936 47985 12000
rect 48049 11936 48065 12000
rect 48129 11936 48135 12000
rect 47819 11935 48135 11936
rect 71256 12000 71572 12001
rect 71256 11936 71262 12000
rect 71326 11936 71342 12000
rect 71406 11936 71422 12000
rect 71486 11936 71502 12000
rect 71566 11936 71572 12000
rect 71256 11935 71572 11936
rect 12985 11930 13051 11933
rect 15377 11930 15443 11933
rect 12985 11928 15443 11930
rect 12985 11872 12990 11928
rect 13046 11872 15382 11928
rect 15438 11872 15443 11928
rect 12985 11870 15443 11872
rect 12985 11867 13051 11870
rect 15377 11867 15443 11870
rect 25405 11930 25471 11933
rect 27429 11930 27495 11933
rect 25405 11928 27495 11930
rect 25405 11872 25410 11928
rect 25466 11872 27434 11928
rect 27490 11872 27495 11928
rect 25405 11870 27495 11872
rect 25405 11867 25471 11870
rect 27429 11867 27495 11870
rect 30189 11930 30255 11933
rect 38653 11930 38719 11933
rect 30189 11928 38719 11930
rect 30189 11872 30194 11928
rect 30250 11872 38658 11928
rect 38714 11872 38719 11928
rect 30189 11870 38719 11872
rect 30189 11867 30255 11870
rect 38653 11867 38719 11870
rect 51165 11930 51231 11933
rect 65057 11930 65123 11933
rect 51165 11928 65123 11930
rect 51165 11872 51170 11928
rect 51226 11872 65062 11928
rect 65118 11872 65123 11928
rect 51165 11870 65123 11872
rect 72374 11930 72434 12142
rect 72693 12200 76439 12202
rect 72693 12144 72698 12200
rect 72754 12144 76378 12200
rect 76434 12144 76439 12200
rect 72693 12142 76439 12144
rect 72693 12139 72759 12142
rect 76373 12139 76439 12142
rect 72509 12066 72575 12069
rect 73613 12066 73679 12069
rect 72509 12064 73679 12066
rect 72509 12008 72514 12064
rect 72570 12008 73618 12064
rect 73674 12008 73679 12064
rect 72509 12006 73679 12008
rect 72509 12003 72575 12006
rect 73613 12003 73679 12006
rect 94693 12000 95009 12001
rect 94693 11936 94699 12000
rect 94763 11936 94779 12000
rect 94843 11936 94859 12000
rect 94923 11936 94939 12000
rect 95003 11936 95009 12000
rect 94693 11935 95009 11936
rect 76189 11930 76255 11933
rect 72374 11928 76255 11930
rect 72374 11872 76194 11928
rect 76250 11872 76255 11928
rect 72374 11870 76255 11872
rect 51165 11867 51231 11870
rect 65057 11867 65123 11870
rect 76189 11867 76255 11870
rect 77937 11930 78003 11933
rect 79041 11930 79107 11933
rect 77937 11928 79107 11930
rect 77937 11872 77942 11928
rect 77998 11872 79046 11928
rect 79102 11872 79107 11928
rect 77937 11870 79107 11872
rect 77937 11867 78003 11870
rect 79041 11867 79107 11870
rect 22553 11794 22619 11797
rect 42609 11794 42675 11797
rect 22553 11792 42675 11794
rect 22553 11736 22558 11792
rect 22614 11736 42614 11792
rect 42670 11736 42675 11792
rect 22553 11734 42675 11736
rect 22553 11731 22619 11734
rect 42609 11731 42675 11734
rect 56685 11794 56751 11797
rect 60549 11794 60615 11797
rect 56685 11792 60615 11794
rect 56685 11736 56690 11792
rect 56746 11736 60554 11792
rect 60610 11736 60615 11792
rect 56685 11734 60615 11736
rect 56685 11731 56751 11734
rect 60549 11731 60615 11734
rect 60733 11794 60799 11797
rect 81433 11794 81499 11797
rect 83733 11794 83799 11797
rect 60733 11792 83799 11794
rect 60733 11736 60738 11792
rect 60794 11736 81438 11792
rect 81494 11736 83738 11792
rect 83794 11736 83799 11792
rect 60733 11734 83799 11736
rect 60733 11731 60799 11734
rect 81433 11731 81499 11734
rect 83733 11731 83799 11734
rect 8661 11658 8727 11661
rect 30005 11658 30071 11661
rect 36997 11658 37063 11661
rect 8661 11656 30071 11658
rect 8661 11600 8666 11656
rect 8722 11600 30010 11656
rect 30066 11600 30071 11656
rect 8661 11598 30071 11600
rect 8661 11595 8727 11598
rect 30005 11595 30071 11598
rect 30192 11656 37063 11658
rect 30192 11600 37002 11656
rect 37058 11600 37063 11656
rect 30192 11598 37063 11600
rect 19333 11522 19399 11525
rect 28625 11522 28691 11525
rect 19333 11520 28691 11522
rect 19333 11464 19338 11520
rect 19394 11464 28630 11520
rect 28686 11464 28691 11520
rect 19333 11462 28691 11464
rect 19333 11459 19399 11462
rect 28625 11459 28691 11462
rect 29177 11522 29243 11525
rect 30192 11522 30252 11598
rect 36997 11595 37063 11598
rect 38837 11658 38903 11661
rect 41413 11658 41479 11661
rect 38837 11656 41479 11658
rect 38837 11600 38842 11656
rect 38898 11600 41418 11656
rect 41474 11600 41479 11656
rect 38837 11598 41479 11600
rect 38837 11595 38903 11598
rect 41413 11595 41479 11598
rect 49877 11658 49943 11661
rect 56501 11658 56567 11661
rect 60917 11658 60983 11661
rect 49877 11656 60983 11658
rect 49877 11600 49882 11656
rect 49938 11600 56506 11656
rect 56562 11600 60922 11656
rect 60978 11600 60983 11656
rect 49877 11598 60983 11600
rect 49877 11595 49943 11598
rect 56501 11595 56567 11598
rect 60917 11595 60983 11598
rect 69749 11658 69815 11661
rect 74717 11658 74783 11661
rect 81617 11658 81683 11661
rect 82537 11658 82603 11661
rect 84285 11658 84351 11661
rect 69749 11656 74783 11658
rect 69749 11600 69754 11656
rect 69810 11600 74722 11656
rect 74778 11600 74783 11656
rect 69749 11598 74783 11600
rect 69749 11595 69815 11598
rect 74717 11595 74783 11598
rect 80010 11656 84351 11658
rect 80010 11600 81622 11656
rect 81678 11600 82542 11656
rect 82598 11600 84290 11656
rect 84346 11600 84351 11656
rect 80010 11598 84351 11600
rect 29177 11520 30252 11522
rect 29177 11464 29182 11520
rect 29238 11464 30252 11520
rect 29177 11462 30252 11464
rect 33409 11522 33475 11525
rect 35709 11522 35775 11525
rect 33409 11520 35775 11522
rect 33409 11464 33414 11520
rect 33470 11464 35714 11520
rect 35770 11464 35775 11520
rect 33409 11462 35775 11464
rect 29177 11459 29243 11462
rect 33409 11459 33475 11462
rect 35709 11459 35775 11462
rect 39573 11522 39639 11525
rect 40217 11522 40283 11525
rect 42885 11522 42951 11525
rect 39573 11520 42951 11522
rect 39573 11464 39578 11520
rect 39634 11464 40222 11520
rect 40278 11464 42890 11520
rect 42946 11464 42951 11520
rect 39573 11462 42951 11464
rect 39573 11459 39639 11462
rect 40217 11459 40283 11462
rect 42885 11459 42951 11462
rect 60365 11522 60431 11525
rect 80010 11522 80070 11598
rect 81617 11595 81683 11598
rect 82537 11595 82603 11598
rect 84285 11595 84351 11598
rect 60365 11520 80070 11522
rect 60365 11464 60370 11520
rect 60426 11464 80070 11520
rect 60365 11462 80070 11464
rect 60365 11459 60431 11462
rect 12664 11456 12980 11457
rect 12664 11392 12670 11456
rect 12734 11392 12750 11456
rect 12814 11392 12830 11456
rect 12894 11392 12910 11456
rect 12974 11392 12980 11456
rect 12664 11391 12980 11392
rect 36101 11456 36417 11457
rect 36101 11392 36107 11456
rect 36171 11392 36187 11456
rect 36251 11392 36267 11456
rect 36331 11392 36347 11456
rect 36411 11392 36417 11456
rect 36101 11391 36417 11392
rect 59538 11456 59854 11457
rect 59538 11392 59544 11456
rect 59608 11392 59624 11456
rect 59688 11392 59704 11456
rect 59768 11392 59784 11456
rect 59848 11392 59854 11456
rect 59538 11391 59854 11392
rect 82975 11456 83291 11457
rect 82975 11392 82981 11456
rect 83045 11392 83061 11456
rect 83125 11392 83141 11456
rect 83205 11392 83221 11456
rect 83285 11392 83291 11456
rect 82975 11391 83291 11392
rect 19885 11386 19951 11389
rect 28073 11386 28139 11389
rect 19885 11384 28139 11386
rect 19885 11328 19890 11384
rect 19946 11328 28078 11384
rect 28134 11328 28139 11384
rect 19885 11326 28139 11328
rect 19885 11323 19951 11326
rect 28073 11323 28139 11326
rect 38745 11386 38811 11389
rect 41597 11386 41663 11389
rect 38745 11384 41663 11386
rect 38745 11328 38750 11384
rect 38806 11328 41602 11384
rect 41658 11328 41663 11384
rect 38745 11326 41663 11328
rect 38745 11323 38811 11326
rect 41597 11323 41663 11326
rect 41781 11386 41847 11389
rect 43989 11386 44055 11389
rect 41781 11384 44055 11386
rect 41781 11328 41786 11384
rect 41842 11328 43994 11384
rect 44050 11328 44055 11384
rect 41781 11326 44055 11328
rect 41781 11323 41847 11326
rect 43989 11323 44055 11326
rect 60089 11386 60155 11389
rect 66437 11386 66503 11389
rect 60089 11384 66503 11386
rect 60089 11328 60094 11384
rect 60150 11328 66442 11384
rect 66498 11328 66503 11384
rect 60089 11326 66503 11328
rect 60089 11323 60155 11326
rect 66437 11323 66503 11326
rect 71129 11386 71195 11389
rect 75453 11386 75519 11389
rect 71129 11384 75519 11386
rect 71129 11328 71134 11384
rect 71190 11328 75458 11384
rect 75514 11328 75519 11384
rect 71129 11326 75519 11328
rect 71129 11323 71195 11326
rect 75453 11323 75519 11326
rect 8477 11250 8543 11253
rect 28901 11250 28967 11253
rect 8477 11248 28967 11250
rect 8477 11192 8482 11248
rect 8538 11192 28906 11248
rect 28962 11192 28967 11248
rect 8477 11190 28967 11192
rect 8477 11187 8543 11190
rect 28901 11187 28967 11190
rect 32673 11250 32739 11253
rect 48957 11250 49023 11253
rect 32673 11248 49023 11250
rect 32673 11192 32678 11248
rect 32734 11192 48962 11248
rect 49018 11192 49023 11248
rect 32673 11190 49023 11192
rect 32673 11187 32739 11190
rect 48957 11187 49023 11190
rect 49693 11250 49759 11253
rect 50613 11250 50679 11253
rect 49693 11248 50679 11250
rect 49693 11192 49698 11248
rect 49754 11192 50618 11248
rect 50674 11192 50679 11248
rect 49693 11190 50679 11192
rect 49693 11187 49759 11190
rect 50613 11187 50679 11190
rect 54661 11250 54727 11253
rect 72233 11250 72299 11253
rect 54661 11248 72299 11250
rect 54661 11192 54666 11248
rect 54722 11192 72238 11248
rect 72294 11192 72299 11248
rect 54661 11190 72299 11192
rect 54661 11187 54727 11190
rect 72233 11187 72299 11190
rect 75177 11250 75243 11253
rect 77201 11250 77267 11253
rect 75177 11248 77267 11250
rect 75177 11192 75182 11248
rect 75238 11192 77206 11248
rect 77262 11192 77267 11248
rect 75177 11190 77267 11192
rect 75177 11187 75243 11190
rect 77201 11187 77267 11190
rect 78581 11250 78647 11253
rect 85757 11250 85823 11253
rect 78581 11248 85823 11250
rect 78581 11192 78586 11248
rect 78642 11192 85762 11248
rect 85818 11192 85823 11248
rect 78581 11190 85823 11192
rect 78581 11187 78647 11190
rect 85757 11187 85823 11190
rect 19333 11114 19399 11117
rect 22921 11114 22987 11117
rect 19333 11112 22987 11114
rect 19333 11056 19338 11112
rect 19394 11056 22926 11112
rect 22982 11056 22987 11112
rect 19333 11054 22987 11056
rect 19333 11051 19399 11054
rect 22921 11051 22987 11054
rect 24301 11114 24367 11117
rect 27797 11114 27863 11117
rect 24301 11112 27863 11114
rect 24301 11056 24306 11112
rect 24362 11056 27802 11112
rect 27858 11056 27863 11112
rect 24301 11054 27863 11056
rect 24301 11051 24367 11054
rect 27797 11051 27863 11054
rect 27981 11114 28047 11117
rect 36905 11114 36971 11117
rect 27981 11112 36971 11114
rect 27981 11056 27986 11112
rect 28042 11056 36910 11112
rect 36966 11056 36971 11112
rect 27981 11054 36971 11056
rect 27981 11051 28047 11054
rect 36905 11051 36971 11054
rect 40125 11114 40191 11117
rect 56777 11114 56843 11117
rect 57329 11114 57395 11117
rect 40125 11112 57395 11114
rect 40125 11056 40130 11112
rect 40186 11056 56782 11112
rect 56838 11056 57334 11112
rect 57390 11056 57395 11112
rect 40125 11054 57395 11056
rect 40125 11051 40191 11054
rect 56777 11051 56843 11054
rect 57329 11051 57395 11054
rect 58893 11114 58959 11117
rect 59302 11114 59308 11116
rect 58893 11112 59308 11114
rect 58893 11056 58898 11112
rect 58954 11056 59308 11112
rect 58893 11054 59308 11056
rect 58893 11051 58959 11054
rect 59302 11052 59308 11054
rect 59372 11052 59378 11116
rect 59905 11114 59971 11117
rect 84009 11114 84075 11117
rect 59905 11112 84075 11114
rect 59905 11056 59910 11112
rect 59966 11056 84014 11112
rect 84070 11056 84075 11112
rect 59905 11054 84075 11056
rect 59905 11051 59971 11054
rect 84009 11051 84075 11054
rect 19333 10978 19399 10981
rect 19793 10978 19859 10981
rect 19333 10976 19859 10978
rect 19333 10920 19338 10976
rect 19394 10920 19798 10976
rect 19854 10920 19859 10976
rect 19333 10918 19859 10920
rect 19333 10915 19399 10918
rect 19793 10915 19859 10918
rect 30465 10978 30531 10981
rect 31661 10978 31727 10981
rect 36537 10978 36603 10981
rect 30465 10976 36603 10978
rect 30465 10920 30470 10976
rect 30526 10920 31666 10976
rect 31722 10920 36542 10976
rect 36598 10920 36603 10976
rect 30465 10918 36603 10920
rect 30465 10915 30531 10918
rect 31661 10915 31727 10918
rect 36537 10915 36603 10918
rect 40493 10978 40559 10981
rect 42149 10978 42215 10981
rect 40493 10976 42215 10978
rect 40493 10920 40498 10976
rect 40554 10920 42154 10976
rect 42210 10920 42215 10976
rect 40493 10918 42215 10920
rect 40493 10915 40559 10918
rect 42149 10915 42215 10918
rect 49509 10978 49575 10981
rect 50705 10978 50771 10981
rect 49509 10976 50771 10978
rect 49509 10920 49514 10976
rect 49570 10920 50710 10976
rect 50766 10920 50771 10976
rect 49509 10918 50771 10920
rect 49509 10915 49575 10918
rect 50705 10915 50771 10918
rect 53833 10978 53899 10981
rect 71129 10978 71195 10981
rect 53833 10976 71195 10978
rect 53833 10920 53838 10976
rect 53894 10920 71134 10976
rect 71190 10920 71195 10976
rect 53833 10918 71195 10920
rect 53833 10915 53899 10918
rect 71129 10915 71195 10918
rect 24382 10912 24698 10913
rect 24382 10848 24388 10912
rect 24452 10848 24468 10912
rect 24532 10848 24548 10912
rect 24612 10848 24628 10912
rect 24692 10848 24698 10912
rect 24382 10847 24698 10848
rect 47819 10912 48135 10913
rect 47819 10848 47825 10912
rect 47889 10848 47905 10912
rect 47969 10848 47985 10912
rect 48049 10848 48065 10912
rect 48129 10848 48135 10912
rect 47819 10847 48135 10848
rect 71256 10912 71572 10913
rect 71256 10848 71262 10912
rect 71326 10848 71342 10912
rect 71406 10848 71422 10912
rect 71486 10848 71502 10912
rect 71566 10848 71572 10912
rect 71256 10847 71572 10848
rect 94693 10912 95009 10913
rect 94693 10848 94699 10912
rect 94763 10848 94779 10912
rect 94843 10848 94859 10912
rect 94923 10848 94939 10912
rect 95003 10848 95009 10912
rect 94693 10847 95009 10848
rect 41781 10842 41847 10845
rect 47025 10842 47091 10845
rect 26926 10782 41430 10842
rect 11881 10706 11947 10709
rect 26926 10706 26986 10782
rect 11881 10704 26986 10706
rect 11881 10648 11886 10704
rect 11942 10648 26986 10704
rect 11881 10646 26986 10648
rect 27521 10706 27587 10709
rect 37733 10706 37799 10709
rect 27521 10704 37799 10706
rect 27521 10648 27526 10704
rect 27582 10648 37738 10704
rect 37794 10648 37799 10704
rect 27521 10646 37799 10648
rect 41370 10706 41430 10782
rect 41781 10840 47091 10842
rect 41781 10784 41786 10840
rect 41842 10784 47030 10840
rect 47086 10784 47091 10840
rect 41781 10782 47091 10784
rect 41781 10779 41847 10782
rect 47025 10779 47091 10782
rect 48405 10842 48471 10845
rect 50153 10842 50219 10845
rect 48405 10840 50219 10842
rect 48405 10784 48410 10840
rect 48466 10784 50158 10840
rect 50214 10784 50219 10840
rect 48405 10782 50219 10784
rect 48405 10779 48471 10782
rect 50153 10779 50219 10782
rect 53281 10842 53347 10845
rect 53649 10842 53715 10845
rect 53281 10840 53715 10842
rect 53281 10784 53286 10840
rect 53342 10784 53654 10840
rect 53710 10784 53715 10840
rect 53281 10782 53715 10784
rect 53281 10779 53347 10782
rect 53649 10779 53715 10782
rect 68277 10842 68343 10845
rect 70577 10842 70643 10845
rect 68277 10840 70643 10842
rect 68277 10784 68282 10840
rect 68338 10784 70582 10840
rect 70638 10784 70643 10840
rect 68277 10782 70643 10784
rect 68277 10779 68343 10782
rect 70577 10779 70643 10782
rect 58249 10706 58315 10709
rect 84285 10706 84351 10709
rect 41370 10704 84351 10706
rect 41370 10648 58254 10704
rect 58310 10648 84290 10704
rect 84346 10648 84351 10704
rect 41370 10646 84351 10648
rect 11881 10643 11947 10646
rect 27521 10643 27587 10646
rect 37733 10643 37799 10646
rect 58249 10643 58315 10646
rect 84285 10643 84351 10646
rect 23933 10570 23999 10573
rect 27981 10570 28047 10573
rect 23933 10568 28047 10570
rect 23933 10512 23938 10568
rect 23994 10512 27986 10568
rect 28042 10512 28047 10568
rect 23933 10510 28047 10512
rect 23933 10507 23999 10510
rect 27981 10507 28047 10510
rect 32949 10570 33015 10573
rect 47669 10570 47735 10573
rect 32949 10568 47735 10570
rect 32949 10512 32954 10568
rect 33010 10512 47674 10568
rect 47730 10512 47735 10568
rect 32949 10510 47735 10512
rect 32949 10507 33015 10510
rect 47669 10507 47735 10510
rect 49325 10570 49391 10573
rect 84193 10570 84259 10573
rect 85481 10570 85547 10573
rect 49325 10568 85547 10570
rect 49325 10512 49330 10568
rect 49386 10512 84198 10568
rect 84254 10512 85486 10568
rect 85542 10512 85547 10568
rect 49325 10510 85547 10512
rect 49325 10507 49391 10510
rect 84193 10507 84259 10510
rect 85481 10507 85547 10510
rect 22553 10434 22619 10437
rect 27061 10434 27127 10437
rect 22553 10432 27127 10434
rect 22553 10376 22558 10432
rect 22614 10376 27066 10432
rect 27122 10376 27127 10432
rect 22553 10374 27127 10376
rect 22553 10371 22619 10374
rect 27061 10371 27127 10374
rect 29821 10434 29887 10437
rect 35065 10434 35131 10437
rect 29821 10432 35131 10434
rect 29821 10376 29826 10432
rect 29882 10376 35070 10432
rect 35126 10376 35131 10432
rect 29821 10374 35131 10376
rect 29821 10371 29887 10374
rect 35065 10371 35131 10374
rect 36537 10434 36603 10437
rect 55397 10434 55463 10437
rect 36537 10432 55463 10434
rect 36537 10376 36542 10432
rect 36598 10376 55402 10432
rect 55458 10376 55463 10432
rect 36537 10374 55463 10376
rect 36537 10371 36603 10374
rect 55397 10371 55463 10374
rect 68461 10434 68527 10437
rect 70945 10434 71011 10437
rect 77661 10434 77727 10437
rect 68461 10432 77727 10434
rect 68461 10376 68466 10432
rect 68522 10376 70950 10432
rect 71006 10376 77666 10432
rect 77722 10376 77727 10432
rect 68461 10374 77727 10376
rect 68461 10371 68527 10374
rect 70945 10371 71011 10374
rect 77661 10371 77727 10374
rect 12664 10368 12980 10369
rect 12664 10304 12670 10368
rect 12734 10304 12750 10368
rect 12814 10304 12830 10368
rect 12894 10304 12910 10368
rect 12974 10304 12980 10368
rect 12664 10303 12980 10304
rect 36101 10368 36417 10369
rect 36101 10304 36107 10368
rect 36171 10304 36187 10368
rect 36251 10304 36267 10368
rect 36331 10304 36347 10368
rect 36411 10304 36417 10368
rect 36101 10303 36417 10304
rect 59538 10368 59854 10369
rect 59538 10304 59544 10368
rect 59608 10304 59624 10368
rect 59688 10304 59704 10368
rect 59768 10304 59784 10368
rect 59848 10304 59854 10368
rect 59538 10303 59854 10304
rect 82975 10368 83291 10369
rect 82975 10304 82981 10368
rect 83045 10304 83061 10368
rect 83125 10304 83141 10368
rect 83205 10304 83221 10368
rect 83285 10304 83291 10368
rect 82975 10303 83291 10304
rect 15101 10298 15167 10301
rect 32397 10298 32463 10301
rect 15101 10296 32463 10298
rect 15101 10240 15106 10296
rect 15162 10240 32402 10296
rect 32458 10240 32463 10296
rect 15101 10238 32463 10240
rect 15101 10235 15167 10238
rect 32397 10235 32463 10238
rect 41137 10298 41203 10301
rect 42057 10298 42123 10301
rect 44357 10298 44423 10301
rect 41137 10296 44423 10298
rect 41137 10240 41142 10296
rect 41198 10240 42062 10296
rect 42118 10240 44362 10296
rect 44418 10240 44423 10296
rect 41137 10238 44423 10240
rect 41137 10235 41203 10238
rect 42057 10235 42123 10238
rect 44357 10235 44423 10238
rect 53281 10298 53347 10301
rect 54477 10298 54543 10301
rect 59353 10298 59419 10301
rect 53281 10296 54543 10298
rect 53281 10240 53286 10296
rect 53342 10240 54482 10296
rect 54538 10240 54543 10296
rect 53281 10238 54543 10240
rect 53281 10235 53347 10238
rect 54477 10235 54543 10238
rect 57286 10296 59419 10298
rect 57286 10240 59358 10296
rect 59414 10240 59419 10296
rect 57286 10238 59419 10240
rect 22001 10162 22067 10165
rect 57286 10162 57346 10238
rect 59353 10235 59419 10238
rect 69565 10298 69631 10301
rect 76097 10298 76163 10301
rect 69565 10296 76163 10298
rect 69565 10240 69570 10296
rect 69626 10240 76102 10296
rect 76158 10240 76163 10296
rect 69565 10238 76163 10240
rect 69565 10235 69631 10238
rect 76097 10235 76163 10238
rect 22001 10160 57346 10162
rect 22001 10104 22006 10160
rect 22062 10104 57346 10160
rect 22001 10102 57346 10104
rect 57421 10162 57487 10165
rect 72877 10162 72943 10165
rect 57421 10160 72943 10162
rect 57421 10104 57426 10160
rect 57482 10104 72882 10160
rect 72938 10104 72943 10160
rect 57421 10102 72943 10104
rect 22001 10099 22067 10102
rect 57421 10099 57487 10102
rect 72877 10099 72943 10102
rect 79961 10162 80027 10165
rect 81801 10162 81867 10165
rect 85389 10162 85455 10165
rect 79961 10160 85455 10162
rect 79961 10104 79966 10160
rect 80022 10104 81806 10160
rect 81862 10104 85394 10160
rect 85450 10104 85455 10160
rect 79961 10102 85455 10104
rect 79961 10099 80027 10102
rect 81801 10099 81867 10102
rect 85389 10099 85455 10102
rect 0 10026 800 10056
rect 1577 10026 1643 10029
rect 0 10024 1643 10026
rect 0 9968 1582 10024
rect 1638 9968 1643 10024
rect 0 9966 1643 9968
rect 0 9936 800 9966
rect 1577 9963 1643 9966
rect 20713 10026 20779 10029
rect 27061 10026 27127 10029
rect 61561 10026 61627 10029
rect 20713 10024 26986 10026
rect 20713 9968 20718 10024
rect 20774 9968 26986 10024
rect 20713 9966 26986 9968
rect 20713 9963 20779 9966
rect 26926 9890 26986 9966
rect 27061 10024 61627 10026
rect 27061 9968 27066 10024
rect 27122 9968 61566 10024
rect 61622 9968 61627 10024
rect 27061 9966 61627 9968
rect 27061 9963 27127 9966
rect 61561 9963 61627 9966
rect 83825 10026 83891 10029
rect 84745 10026 84811 10029
rect 83825 10024 84811 10026
rect 83825 9968 83830 10024
rect 83886 9968 84750 10024
rect 84806 9968 84811 10024
rect 83825 9966 84811 9968
rect 83825 9963 83891 9966
rect 84745 9963 84811 9966
rect 34513 9890 34579 9893
rect 36629 9890 36695 9893
rect 26926 9830 31770 9890
rect 24382 9824 24698 9825
rect 24382 9760 24388 9824
rect 24452 9760 24468 9824
rect 24532 9760 24548 9824
rect 24612 9760 24628 9824
rect 24692 9760 24698 9824
rect 24382 9759 24698 9760
rect 19701 9754 19767 9757
rect 23565 9754 23631 9757
rect 19701 9752 23631 9754
rect 19701 9696 19706 9752
rect 19762 9696 23570 9752
rect 23626 9696 23631 9752
rect 19701 9694 23631 9696
rect 19701 9691 19767 9694
rect 23565 9691 23631 9694
rect 28993 9754 29059 9757
rect 29453 9754 29519 9757
rect 28993 9752 29519 9754
rect 28993 9696 28998 9752
rect 29054 9696 29458 9752
rect 29514 9696 29519 9752
rect 28993 9694 29519 9696
rect 31710 9754 31770 9830
rect 34513 9888 36695 9890
rect 34513 9832 34518 9888
rect 34574 9832 36634 9888
rect 36690 9832 36695 9888
rect 34513 9830 36695 9832
rect 34513 9827 34579 9830
rect 36629 9827 36695 9830
rect 37733 9890 37799 9893
rect 41137 9890 41203 9893
rect 37733 9888 41203 9890
rect 37733 9832 37738 9888
rect 37794 9832 41142 9888
rect 41198 9832 41203 9888
rect 37733 9830 41203 9832
rect 37733 9827 37799 9830
rect 41137 9827 41203 9830
rect 41321 9890 41387 9893
rect 44817 9890 44883 9893
rect 41321 9888 44883 9890
rect 41321 9832 41326 9888
rect 41382 9832 44822 9888
rect 44878 9832 44883 9888
rect 41321 9830 44883 9832
rect 41321 9827 41387 9830
rect 44817 9827 44883 9830
rect 45185 9890 45251 9893
rect 46565 9890 46631 9893
rect 45185 9888 46631 9890
rect 45185 9832 45190 9888
rect 45246 9832 46570 9888
rect 46626 9832 46631 9888
rect 45185 9830 46631 9832
rect 45185 9827 45251 9830
rect 46565 9827 46631 9830
rect 52545 9890 52611 9893
rect 67909 9890 67975 9893
rect 52545 9888 67975 9890
rect 52545 9832 52550 9888
rect 52606 9832 67914 9888
rect 67970 9832 67975 9888
rect 52545 9830 67975 9832
rect 52545 9827 52611 9830
rect 67909 9827 67975 9830
rect 47819 9824 48135 9825
rect 47819 9760 47825 9824
rect 47889 9760 47905 9824
rect 47969 9760 47985 9824
rect 48049 9760 48065 9824
rect 48129 9760 48135 9824
rect 47819 9759 48135 9760
rect 71256 9824 71572 9825
rect 71256 9760 71262 9824
rect 71326 9760 71342 9824
rect 71406 9760 71422 9824
rect 71486 9760 71502 9824
rect 71566 9760 71572 9824
rect 71256 9759 71572 9760
rect 94693 9824 95009 9825
rect 94693 9760 94699 9824
rect 94763 9760 94779 9824
rect 94843 9760 94859 9824
rect 94923 9760 94939 9824
rect 95003 9760 95009 9824
rect 94693 9759 95009 9760
rect 36813 9754 36879 9757
rect 31710 9752 36879 9754
rect 31710 9696 36818 9752
rect 36874 9696 36879 9752
rect 31710 9694 36879 9696
rect 28993 9691 29059 9694
rect 29453 9691 29519 9694
rect 36813 9691 36879 9694
rect 39297 9754 39363 9757
rect 42701 9754 42767 9757
rect 39297 9752 42767 9754
rect 39297 9696 39302 9752
rect 39358 9696 42706 9752
rect 42762 9696 42767 9752
rect 39297 9694 42767 9696
rect 39297 9691 39363 9694
rect 42701 9691 42767 9694
rect 59353 9754 59419 9757
rect 60365 9754 60431 9757
rect 65977 9754 66043 9757
rect 70301 9754 70367 9757
rect 59353 9752 70367 9754
rect 59353 9696 59358 9752
rect 59414 9696 60370 9752
rect 60426 9696 65982 9752
rect 66038 9696 70306 9752
rect 70362 9696 70367 9752
rect 59353 9694 70367 9696
rect 59353 9691 59419 9694
rect 60365 9691 60431 9694
rect 65977 9691 66043 9694
rect 70301 9691 70367 9694
rect 23381 9618 23447 9621
rect 26785 9618 26851 9621
rect 23381 9616 26851 9618
rect 23381 9560 23386 9616
rect 23442 9560 26790 9616
rect 26846 9560 26851 9616
rect 23381 9558 26851 9560
rect 23381 9555 23447 9558
rect 26785 9555 26851 9558
rect 30189 9618 30255 9621
rect 45001 9618 45067 9621
rect 81525 9618 81591 9621
rect 30189 9616 45067 9618
rect 30189 9560 30194 9616
rect 30250 9560 45006 9616
rect 45062 9560 45067 9616
rect 30189 9558 45067 9560
rect 30189 9555 30255 9558
rect 45001 9555 45067 9558
rect 60690 9616 81591 9618
rect 60690 9560 81530 9616
rect 81586 9560 81591 9616
rect 60690 9558 81591 9560
rect 14549 9482 14615 9485
rect 23381 9482 23447 9485
rect 14549 9480 23447 9482
rect 14549 9424 14554 9480
rect 14610 9424 23386 9480
rect 23442 9424 23447 9480
rect 14549 9422 23447 9424
rect 14549 9419 14615 9422
rect 23381 9419 23447 9422
rect 23565 9482 23631 9485
rect 26601 9482 26667 9485
rect 23565 9480 26667 9482
rect 23565 9424 23570 9480
rect 23626 9424 26606 9480
rect 26662 9424 26667 9480
rect 23565 9422 26667 9424
rect 23565 9419 23631 9422
rect 26601 9419 26667 9422
rect 30281 9482 30347 9485
rect 32581 9482 32647 9485
rect 30281 9480 32647 9482
rect 30281 9424 30286 9480
rect 30342 9424 32586 9480
rect 32642 9424 32647 9480
rect 30281 9422 32647 9424
rect 30281 9419 30347 9422
rect 32581 9419 32647 9422
rect 33317 9482 33383 9485
rect 40217 9482 40283 9485
rect 33317 9480 40283 9482
rect 33317 9424 33322 9480
rect 33378 9424 40222 9480
rect 40278 9424 40283 9480
rect 33317 9422 40283 9424
rect 33317 9419 33383 9422
rect 40217 9419 40283 9422
rect 41229 9482 41295 9485
rect 45093 9482 45159 9485
rect 41229 9480 45159 9482
rect 41229 9424 41234 9480
rect 41290 9424 45098 9480
rect 45154 9424 45159 9480
rect 41229 9422 45159 9424
rect 41229 9419 41295 9422
rect 45093 9419 45159 9422
rect 56041 9482 56107 9485
rect 60690 9482 60750 9558
rect 81525 9555 81591 9558
rect 56041 9480 60750 9482
rect 56041 9424 56046 9480
rect 56102 9424 60750 9480
rect 56041 9422 60750 9424
rect 63125 9482 63191 9485
rect 67449 9482 67515 9485
rect 63125 9480 67515 9482
rect 63125 9424 63130 9480
rect 63186 9424 67454 9480
rect 67510 9424 67515 9480
rect 63125 9422 67515 9424
rect 56041 9419 56107 9422
rect 63125 9419 63191 9422
rect 67449 9419 67515 9422
rect 67633 9482 67699 9485
rect 68001 9482 68067 9485
rect 67633 9480 68067 9482
rect 67633 9424 67638 9480
rect 67694 9424 68006 9480
rect 68062 9424 68067 9480
rect 67633 9422 68067 9424
rect 67633 9419 67699 9422
rect 68001 9419 68067 9422
rect 70209 9482 70275 9485
rect 71129 9482 71195 9485
rect 70209 9480 71195 9482
rect 70209 9424 70214 9480
rect 70270 9424 71134 9480
rect 71190 9424 71195 9480
rect 70209 9422 71195 9424
rect 70209 9419 70275 9422
rect 71129 9419 71195 9422
rect 73981 9482 74047 9485
rect 75453 9482 75519 9485
rect 73981 9480 75519 9482
rect 73981 9424 73986 9480
rect 74042 9424 75458 9480
rect 75514 9424 75519 9480
rect 73981 9422 75519 9424
rect 73981 9419 74047 9422
rect 75453 9419 75519 9422
rect 21909 9346 21975 9349
rect 22185 9346 22251 9349
rect 21909 9344 22251 9346
rect 21909 9288 21914 9344
rect 21970 9288 22190 9344
rect 22246 9288 22251 9344
rect 21909 9286 22251 9288
rect 32584 9346 32644 9419
rect 34881 9346 34947 9349
rect 32584 9344 34947 9346
rect 32584 9288 34886 9344
rect 34942 9288 34947 9344
rect 32584 9286 34947 9288
rect 21909 9283 21975 9286
rect 22185 9283 22251 9286
rect 34881 9283 34947 9286
rect 38837 9346 38903 9349
rect 46565 9346 46631 9349
rect 38837 9344 46631 9346
rect 38837 9288 38842 9344
rect 38898 9288 46570 9344
rect 46626 9288 46631 9344
rect 38837 9286 46631 9288
rect 38837 9283 38903 9286
rect 46565 9283 46631 9286
rect 48865 9346 48931 9349
rect 49601 9346 49667 9349
rect 48865 9344 49667 9346
rect 48865 9288 48870 9344
rect 48926 9288 49606 9344
rect 49662 9288 49667 9344
rect 48865 9286 49667 9288
rect 48865 9283 48931 9286
rect 49601 9283 49667 9286
rect 67817 9346 67883 9349
rect 72417 9346 72483 9349
rect 67817 9344 72483 9346
rect 67817 9288 67822 9344
rect 67878 9288 72422 9344
rect 72478 9288 72483 9344
rect 67817 9286 72483 9288
rect 67817 9283 67883 9286
rect 72417 9283 72483 9286
rect 12664 9280 12980 9281
rect 12664 9216 12670 9280
rect 12734 9216 12750 9280
rect 12814 9216 12830 9280
rect 12894 9216 12910 9280
rect 12974 9216 12980 9280
rect 12664 9215 12980 9216
rect 36101 9280 36417 9281
rect 36101 9216 36107 9280
rect 36171 9216 36187 9280
rect 36251 9216 36267 9280
rect 36331 9216 36347 9280
rect 36411 9216 36417 9280
rect 36101 9215 36417 9216
rect 59538 9280 59854 9281
rect 59538 9216 59544 9280
rect 59608 9216 59624 9280
rect 59688 9216 59704 9280
rect 59768 9216 59784 9280
rect 59848 9216 59854 9280
rect 59538 9215 59854 9216
rect 82975 9280 83291 9281
rect 82975 9216 82981 9280
rect 83045 9216 83061 9280
rect 83125 9216 83141 9280
rect 83205 9216 83221 9280
rect 83285 9216 83291 9280
rect 82975 9215 83291 9216
rect 23197 9210 23263 9213
rect 27521 9210 27587 9213
rect 23197 9208 27587 9210
rect 23197 9152 23202 9208
rect 23258 9152 27526 9208
rect 27582 9152 27587 9208
rect 23197 9150 27587 9152
rect 23197 9147 23263 9150
rect 27521 9147 27587 9150
rect 33041 9210 33107 9213
rect 33685 9210 33751 9213
rect 33041 9208 33751 9210
rect 33041 9152 33046 9208
rect 33102 9152 33690 9208
rect 33746 9152 33751 9208
rect 33041 9150 33751 9152
rect 33041 9147 33107 9150
rect 33685 9147 33751 9150
rect 35065 9210 35131 9213
rect 35709 9210 35775 9213
rect 35065 9208 35775 9210
rect 35065 9152 35070 9208
rect 35126 9152 35714 9208
rect 35770 9152 35775 9208
rect 35065 9150 35775 9152
rect 35065 9147 35131 9150
rect 35709 9147 35775 9150
rect 41229 9210 41295 9213
rect 41597 9210 41663 9213
rect 41229 9208 41663 9210
rect 41229 9152 41234 9208
rect 41290 9152 41602 9208
rect 41658 9152 41663 9208
rect 41229 9150 41663 9152
rect 41229 9147 41295 9150
rect 41597 9147 41663 9150
rect 59997 9210 60063 9213
rect 71865 9210 71931 9213
rect 59997 9208 71931 9210
rect 59997 9152 60002 9208
rect 60058 9152 71870 9208
rect 71926 9152 71931 9208
rect 59997 9150 71931 9152
rect 59997 9147 60063 9150
rect 71865 9147 71931 9150
rect 18689 9074 18755 9077
rect 19885 9074 19951 9077
rect 38469 9074 38535 9077
rect 38745 9074 38811 9077
rect 18689 9072 38811 9074
rect 18689 9016 18694 9072
rect 18750 9016 19890 9072
rect 19946 9016 38474 9072
rect 38530 9016 38750 9072
rect 38806 9016 38811 9072
rect 18689 9014 38811 9016
rect 18689 9011 18755 9014
rect 19885 9011 19951 9014
rect 38469 9011 38535 9014
rect 38745 9011 38811 9014
rect 38929 9074 38995 9077
rect 39665 9074 39731 9077
rect 43437 9074 43503 9077
rect 46749 9074 46815 9077
rect 38929 9072 46815 9074
rect 38929 9016 38934 9072
rect 38990 9016 39670 9072
rect 39726 9016 43442 9072
rect 43498 9016 46754 9072
rect 46810 9016 46815 9072
rect 38929 9014 46815 9016
rect 38929 9011 38995 9014
rect 39665 9011 39731 9014
rect 43437 9011 43503 9014
rect 46749 9011 46815 9014
rect 47577 9074 47643 9077
rect 48773 9074 48839 9077
rect 67081 9074 67147 9077
rect 47577 9072 67147 9074
rect 47577 9016 47582 9072
rect 47638 9016 48778 9072
rect 48834 9016 67086 9072
rect 67142 9016 67147 9072
rect 47577 9014 67147 9016
rect 47577 9011 47643 9014
rect 48773 9011 48839 9014
rect 67081 9011 67147 9014
rect 20621 8938 20687 8941
rect 22645 8938 22711 8941
rect 20621 8936 22711 8938
rect 20621 8880 20626 8936
rect 20682 8880 22650 8936
rect 22706 8880 22711 8936
rect 20621 8878 22711 8880
rect 20621 8875 20687 8878
rect 22645 8875 22711 8878
rect 34513 8938 34579 8941
rect 38837 8938 38903 8941
rect 55489 8938 55555 8941
rect 34513 8936 38903 8938
rect 34513 8880 34518 8936
rect 34574 8880 38842 8936
rect 38898 8880 38903 8936
rect 34513 8878 38903 8880
rect 34513 8875 34579 8878
rect 38837 8875 38903 8878
rect 41370 8936 55555 8938
rect 41370 8880 55494 8936
rect 55550 8880 55555 8936
rect 41370 8878 55555 8880
rect 17677 8802 17743 8805
rect 18321 8802 18387 8805
rect 21633 8802 21699 8805
rect 22553 8802 22619 8805
rect 17677 8800 22619 8802
rect 17677 8744 17682 8800
rect 17738 8744 18326 8800
rect 18382 8744 21638 8800
rect 21694 8744 22558 8800
rect 22614 8744 22619 8800
rect 17677 8742 22619 8744
rect 17677 8739 17743 8742
rect 18321 8739 18387 8742
rect 21633 8739 21699 8742
rect 22553 8739 22619 8742
rect 35157 8802 35223 8805
rect 35525 8802 35591 8805
rect 41370 8802 41430 8878
rect 55489 8875 55555 8878
rect 57605 8938 57671 8941
rect 59997 8938 60063 8941
rect 57605 8936 60063 8938
rect 57605 8880 57610 8936
rect 57666 8880 60002 8936
rect 60058 8880 60063 8936
rect 57605 8878 60063 8880
rect 57605 8875 57671 8878
rect 59997 8875 60063 8878
rect 64229 8938 64295 8941
rect 78857 8938 78923 8941
rect 64229 8936 78923 8938
rect 64229 8880 64234 8936
rect 64290 8880 78862 8936
rect 78918 8880 78923 8936
rect 64229 8878 78923 8880
rect 64229 8875 64295 8878
rect 78857 8875 78923 8878
rect 80513 8938 80579 8941
rect 85481 8938 85547 8941
rect 80513 8936 85547 8938
rect 80513 8880 80518 8936
rect 80574 8880 85486 8936
rect 85542 8880 85547 8936
rect 80513 8878 85547 8880
rect 80513 8875 80579 8878
rect 85481 8875 85547 8878
rect 35157 8800 41430 8802
rect 35157 8744 35162 8800
rect 35218 8744 35530 8800
rect 35586 8744 41430 8800
rect 35157 8742 41430 8744
rect 46565 8802 46631 8805
rect 47209 8802 47275 8805
rect 46565 8800 47275 8802
rect 46565 8744 46570 8800
rect 46626 8744 47214 8800
rect 47270 8744 47275 8800
rect 46565 8742 47275 8744
rect 35157 8739 35223 8742
rect 35525 8739 35591 8742
rect 46565 8739 46631 8742
rect 47209 8739 47275 8742
rect 59302 8740 59308 8804
rect 59372 8802 59378 8804
rect 65793 8802 65859 8805
rect 59372 8800 65859 8802
rect 59372 8744 65798 8800
rect 65854 8744 65859 8800
rect 59372 8742 65859 8744
rect 59372 8740 59378 8742
rect 65793 8739 65859 8742
rect 24382 8736 24698 8737
rect 24382 8672 24388 8736
rect 24452 8672 24468 8736
rect 24532 8672 24548 8736
rect 24612 8672 24628 8736
rect 24692 8672 24698 8736
rect 24382 8671 24698 8672
rect 47819 8736 48135 8737
rect 47819 8672 47825 8736
rect 47889 8672 47905 8736
rect 47969 8672 47985 8736
rect 48049 8672 48065 8736
rect 48129 8672 48135 8736
rect 47819 8671 48135 8672
rect 71256 8736 71572 8737
rect 71256 8672 71262 8736
rect 71326 8672 71342 8736
rect 71406 8672 71422 8736
rect 71486 8672 71502 8736
rect 71566 8672 71572 8736
rect 71256 8671 71572 8672
rect 94693 8736 95009 8737
rect 94693 8672 94699 8736
rect 94763 8672 94779 8736
rect 94843 8672 94859 8736
rect 94923 8672 94939 8736
rect 95003 8672 95009 8736
rect 94693 8671 95009 8672
rect 17125 8666 17191 8669
rect 20437 8666 20503 8669
rect 17125 8664 20503 8666
rect 17125 8608 17130 8664
rect 17186 8608 20442 8664
rect 20498 8608 20503 8664
rect 17125 8606 20503 8608
rect 17125 8603 17191 8606
rect 20437 8603 20503 8606
rect 34329 8666 34395 8669
rect 37089 8666 37155 8669
rect 34329 8664 37155 8666
rect 34329 8608 34334 8664
rect 34390 8608 37094 8664
rect 37150 8608 37155 8664
rect 34329 8606 37155 8608
rect 34329 8603 34395 8606
rect 37089 8603 37155 8606
rect 40493 8666 40559 8669
rect 42425 8666 42491 8669
rect 40493 8664 42491 8666
rect 40493 8608 40498 8664
rect 40554 8608 42430 8664
rect 42486 8608 42491 8664
rect 40493 8606 42491 8608
rect 40493 8603 40559 8606
rect 42425 8603 42491 8606
rect 61009 8666 61075 8669
rect 63493 8666 63559 8669
rect 64505 8666 64571 8669
rect 61009 8664 64571 8666
rect 61009 8608 61014 8664
rect 61070 8608 63498 8664
rect 63554 8608 64510 8664
rect 64566 8608 64571 8664
rect 61009 8606 64571 8608
rect 61009 8603 61075 8606
rect 63493 8603 63559 8606
rect 64505 8603 64571 8606
rect 17401 8530 17467 8533
rect 20713 8530 20779 8533
rect 17401 8528 20779 8530
rect 17401 8472 17406 8528
rect 17462 8472 20718 8528
rect 20774 8472 20779 8528
rect 17401 8470 20779 8472
rect 17401 8467 17467 8470
rect 20713 8467 20779 8470
rect 21449 8530 21515 8533
rect 23749 8530 23815 8533
rect 21449 8528 23815 8530
rect 21449 8472 21454 8528
rect 21510 8472 23754 8528
rect 23810 8472 23815 8528
rect 21449 8470 23815 8472
rect 21449 8467 21515 8470
rect 23749 8467 23815 8470
rect 33041 8530 33107 8533
rect 38101 8530 38167 8533
rect 33041 8528 38167 8530
rect 33041 8472 33046 8528
rect 33102 8472 38106 8528
rect 38162 8472 38167 8528
rect 33041 8470 38167 8472
rect 33041 8467 33107 8470
rect 38101 8467 38167 8470
rect 40769 8530 40835 8533
rect 46565 8530 46631 8533
rect 40769 8528 46631 8530
rect 40769 8472 40774 8528
rect 40830 8472 46570 8528
rect 46626 8472 46631 8528
rect 40769 8470 46631 8472
rect 40769 8467 40835 8470
rect 46565 8467 46631 8470
rect 55397 8530 55463 8533
rect 63534 8530 63540 8532
rect 55397 8528 63540 8530
rect 55397 8472 55402 8528
rect 55458 8472 63540 8528
rect 55397 8470 63540 8472
rect 55397 8467 55463 8470
rect 63534 8468 63540 8470
rect 63604 8530 63610 8532
rect 63769 8530 63835 8533
rect 79777 8530 79843 8533
rect 80789 8530 80855 8533
rect 63604 8528 80855 8530
rect 63604 8472 63774 8528
rect 63830 8472 79782 8528
rect 79838 8472 80794 8528
rect 80850 8472 80855 8528
rect 63604 8470 80855 8472
rect 63604 8468 63610 8470
rect 63769 8467 63835 8470
rect 79777 8467 79843 8470
rect 80789 8467 80855 8470
rect 16665 8394 16731 8397
rect 17585 8394 17651 8397
rect 16665 8392 17651 8394
rect 16665 8336 16670 8392
rect 16726 8336 17590 8392
rect 17646 8336 17651 8392
rect 16665 8334 17651 8336
rect 16665 8331 16731 8334
rect 17585 8331 17651 8334
rect 20069 8394 20135 8397
rect 21909 8394 21975 8397
rect 27521 8394 27587 8397
rect 20069 8392 27587 8394
rect 20069 8336 20074 8392
rect 20130 8336 21914 8392
rect 21970 8336 27526 8392
rect 27582 8336 27587 8392
rect 20069 8334 27587 8336
rect 20069 8331 20135 8334
rect 21909 8331 21975 8334
rect 27521 8331 27587 8334
rect 33869 8394 33935 8397
rect 49509 8394 49575 8397
rect 33869 8392 49575 8394
rect 33869 8336 33874 8392
rect 33930 8336 49514 8392
rect 49570 8336 49575 8392
rect 33869 8334 49575 8336
rect 33869 8331 33935 8334
rect 49509 8331 49575 8334
rect 63677 8394 63743 8397
rect 64045 8394 64111 8397
rect 79869 8394 79935 8397
rect 63677 8392 79935 8394
rect 63677 8336 63682 8392
rect 63738 8336 64050 8392
rect 64106 8336 79874 8392
rect 79930 8336 79935 8392
rect 63677 8334 79935 8336
rect 63677 8331 63743 8334
rect 64045 8331 64111 8334
rect 79869 8331 79935 8334
rect 36537 8258 36603 8261
rect 37825 8258 37891 8261
rect 36537 8256 37891 8258
rect 36537 8200 36542 8256
rect 36598 8200 37830 8256
rect 37886 8200 37891 8256
rect 36537 8198 37891 8200
rect 36537 8195 36603 8198
rect 37825 8195 37891 8198
rect 12664 8192 12980 8193
rect 12664 8128 12670 8192
rect 12734 8128 12750 8192
rect 12814 8128 12830 8192
rect 12894 8128 12910 8192
rect 12974 8128 12980 8192
rect 12664 8127 12980 8128
rect 36101 8192 36417 8193
rect 36101 8128 36107 8192
rect 36171 8128 36187 8192
rect 36251 8128 36267 8192
rect 36331 8128 36347 8192
rect 36411 8128 36417 8192
rect 36101 8127 36417 8128
rect 59538 8192 59854 8193
rect 59538 8128 59544 8192
rect 59608 8128 59624 8192
rect 59688 8128 59704 8192
rect 59768 8128 59784 8192
rect 59848 8128 59854 8192
rect 59538 8127 59854 8128
rect 82975 8192 83291 8193
rect 82975 8128 82981 8192
rect 83045 8128 83061 8192
rect 83125 8128 83141 8192
rect 83205 8128 83221 8192
rect 83285 8128 83291 8192
rect 82975 8127 83291 8128
rect 40401 8122 40467 8125
rect 45461 8122 45527 8125
rect 40401 8120 45527 8122
rect 40401 8064 40406 8120
rect 40462 8064 45466 8120
rect 45522 8064 45527 8120
rect 40401 8062 45527 8064
rect 40401 8059 40467 8062
rect 45461 8059 45527 8062
rect 45645 8122 45711 8125
rect 47393 8122 47459 8125
rect 45645 8120 47459 8122
rect 45645 8064 45650 8120
rect 45706 8064 47398 8120
rect 47454 8064 47459 8120
rect 45645 8062 47459 8064
rect 45645 8059 45711 8062
rect 47393 8059 47459 8062
rect 13445 7986 13511 7989
rect 51073 7986 51139 7989
rect 13445 7984 51139 7986
rect 13445 7928 13450 7984
rect 13506 7928 51078 7984
rect 51134 7928 51139 7984
rect 13445 7926 51139 7928
rect 13445 7923 13511 7926
rect 51073 7923 51139 7926
rect 71497 7986 71563 7989
rect 74533 7986 74599 7989
rect 71497 7984 74599 7986
rect 71497 7928 71502 7984
rect 71558 7928 74538 7984
rect 74594 7928 74599 7984
rect 71497 7926 74599 7928
rect 71497 7923 71563 7926
rect 74533 7923 74599 7926
rect 13169 7850 13235 7853
rect 34421 7850 34487 7853
rect 13169 7848 34487 7850
rect 13169 7792 13174 7848
rect 13230 7792 34426 7848
rect 34482 7792 34487 7848
rect 13169 7790 34487 7792
rect 13169 7787 13235 7790
rect 34421 7787 34487 7790
rect 35157 7850 35223 7853
rect 45185 7850 45251 7853
rect 35157 7848 45251 7850
rect 35157 7792 35162 7848
rect 35218 7792 45190 7848
rect 45246 7792 45251 7848
rect 35157 7790 45251 7792
rect 35157 7787 35223 7790
rect 45185 7787 45251 7790
rect 51165 7850 51231 7853
rect 51717 7850 51783 7853
rect 57329 7850 57395 7853
rect 51165 7848 57395 7850
rect 51165 7792 51170 7848
rect 51226 7792 51722 7848
rect 51778 7792 57334 7848
rect 57390 7792 57395 7848
rect 51165 7790 57395 7792
rect 51165 7787 51231 7790
rect 51717 7787 51783 7790
rect 57329 7787 57395 7790
rect 66713 7850 66779 7853
rect 69565 7850 69631 7853
rect 66713 7848 69631 7850
rect 66713 7792 66718 7848
rect 66774 7792 69570 7848
rect 69626 7792 69631 7848
rect 66713 7790 69631 7792
rect 66713 7787 66779 7790
rect 69565 7787 69631 7790
rect 33133 7714 33199 7717
rect 42609 7714 42675 7717
rect 33133 7712 42675 7714
rect 33133 7656 33138 7712
rect 33194 7656 42614 7712
rect 42670 7656 42675 7712
rect 33133 7654 42675 7656
rect 33133 7651 33199 7654
rect 42609 7651 42675 7654
rect 24382 7648 24698 7649
rect 24382 7584 24388 7648
rect 24452 7584 24468 7648
rect 24532 7584 24548 7648
rect 24612 7584 24628 7648
rect 24692 7584 24698 7648
rect 24382 7583 24698 7584
rect 47819 7648 48135 7649
rect 47819 7584 47825 7648
rect 47889 7584 47905 7648
rect 47969 7584 47985 7648
rect 48049 7584 48065 7648
rect 48129 7584 48135 7648
rect 47819 7583 48135 7584
rect 71256 7648 71572 7649
rect 71256 7584 71262 7648
rect 71326 7584 71342 7648
rect 71406 7584 71422 7648
rect 71486 7584 71502 7648
rect 71566 7584 71572 7648
rect 71256 7583 71572 7584
rect 94693 7648 95009 7649
rect 94693 7584 94699 7648
rect 94763 7584 94779 7648
rect 94843 7584 94859 7648
rect 94923 7584 94939 7648
rect 95003 7584 95009 7648
rect 94693 7583 95009 7584
rect 95200 7581 96000 7608
rect 46565 7578 46631 7581
rect 26926 7576 46631 7578
rect 26926 7520 46570 7576
rect 46626 7520 46631 7576
rect 26926 7518 46631 7520
rect 20989 7442 21055 7445
rect 26926 7442 26986 7518
rect 46565 7515 46631 7518
rect 51073 7578 51139 7581
rect 60641 7578 60707 7581
rect 62573 7578 62639 7581
rect 68829 7578 68895 7581
rect 83549 7578 83615 7581
rect 84929 7578 84995 7581
rect 86585 7578 86651 7581
rect 51073 7576 70410 7578
rect 51073 7520 51078 7576
rect 51134 7520 60646 7576
rect 60702 7520 62578 7576
rect 62634 7520 68834 7576
rect 68890 7520 70410 7576
rect 51073 7518 70410 7520
rect 51073 7515 51139 7518
rect 60641 7515 60707 7518
rect 62573 7515 62639 7518
rect 68829 7515 68895 7518
rect 58065 7442 58131 7445
rect 20989 7440 26986 7442
rect 20989 7384 20994 7440
rect 21050 7384 26986 7440
rect 20989 7382 26986 7384
rect 27478 7440 58131 7442
rect 27478 7384 58070 7440
rect 58126 7384 58131 7440
rect 27478 7382 58131 7384
rect 20989 7379 21055 7382
rect 23105 7306 23171 7309
rect 27478 7306 27538 7382
rect 58065 7379 58131 7382
rect 63309 7442 63375 7445
rect 66621 7442 66687 7445
rect 68001 7442 68067 7445
rect 63309 7440 68067 7442
rect 63309 7384 63314 7440
rect 63370 7384 66626 7440
rect 66682 7384 68006 7440
rect 68062 7384 68067 7440
rect 63309 7382 68067 7384
rect 63309 7379 63375 7382
rect 66621 7379 66687 7382
rect 68001 7379 68067 7382
rect 69473 7306 69539 7309
rect 23105 7304 27538 7306
rect 23105 7248 23110 7304
rect 23166 7248 27538 7304
rect 23105 7246 27538 7248
rect 31710 7304 69539 7306
rect 31710 7248 69478 7304
rect 69534 7248 69539 7304
rect 31710 7246 69539 7248
rect 70350 7306 70410 7518
rect 83549 7576 86651 7578
rect 83549 7520 83554 7576
rect 83610 7520 84934 7576
rect 84990 7520 86590 7576
rect 86646 7520 86651 7576
rect 83549 7518 86651 7520
rect 83549 7515 83615 7518
rect 84929 7515 84995 7518
rect 86585 7515 86651 7518
rect 95141 7576 96000 7581
rect 95141 7520 95146 7576
rect 95202 7520 96000 7576
rect 95141 7515 96000 7520
rect 95200 7488 96000 7515
rect 72601 7306 72667 7309
rect 73521 7306 73587 7309
rect 70350 7304 73587 7306
rect 70350 7248 72606 7304
rect 72662 7248 73526 7304
rect 73582 7248 73587 7304
rect 70350 7246 73587 7248
rect 23105 7243 23171 7246
rect 23657 7170 23723 7173
rect 31710 7170 31770 7246
rect 69473 7243 69539 7246
rect 72601 7243 72667 7246
rect 73521 7243 73587 7246
rect 23657 7168 31770 7170
rect 23657 7112 23662 7168
rect 23718 7112 31770 7168
rect 23657 7110 31770 7112
rect 40585 7170 40651 7173
rect 41873 7170 41939 7173
rect 40585 7168 41939 7170
rect 40585 7112 40590 7168
rect 40646 7112 41878 7168
rect 41934 7112 41939 7168
rect 40585 7110 41939 7112
rect 23657 7107 23723 7110
rect 40585 7107 40651 7110
rect 41873 7107 41939 7110
rect 49141 7170 49207 7173
rect 54201 7170 54267 7173
rect 49141 7168 54267 7170
rect 49141 7112 49146 7168
rect 49202 7112 54206 7168
rect 54262 7112 54267 7168
rect 49141 7110 54267 7112
rect 49141 7107 49207 7110
rect 54201 7107 54267 7110
rect 67081 7170 67147 7173
rect 68829 7170 68895 7173
rect 67081 7168 68895 7170
rect 67081 7112 67086 7168
rect 67142 7112 68834 7168
rect 68890 7112 68895 7168
rect 67081 7110 68895 7112
rect 67081 7107 67147 7110
rect 68829 7107 68895 7110
rect 69841 7170 69907 7173
rect 71865 7170 71931 7173
rect 69841 7168 71931 7170
rect 69841 7112 69846 7168
rect 69902 7112 71870 7168
rect 71926 7112 71931 7168
rect 69841 7110 71931 7112
rect 69841 7107 69907 7110
rect 71865 7107 71931 7110
rect 12664 7104 12980 7105
rect 12664 7040 12670 7104
rect 12734 7040 12750 7104
rect 12814 7040 12830 7104
rect 12894 7040 12910 7104
rect 12974 7040 12980 7104
rect 12664 7039 12980 7040
rect 36101 7104 36417 7105
rect 36101 7040 36107 7104
rect 36171 7040 36187 7104
rect 36251 7040 36267 7104
rect 36331 7040 36347 7104
rect 36411 7040 36417 7104
rect 36101 7039 36417 7040
rect 59538 7104 59854 7105
rect 59538 7040 59544 7104
rect 59608 7040 59624 7104
rect 59688 7040 59704 7104
rect 59768 7040 59784 7104
rect 59848 7040 59854 7104
rect 59538 7039 59854 7040
rect 82975 7104 83291 7105
rect 82975 7040 82981 7104
rect 83045 7040 83061 7104
rect 83125 7040 83141 7104
rect 83205 7040 83221 7104
rect 83285 7040 83291 7104
rect 82975 7039 83291 7040
rect 34697 7034 34763 7037
rect 35893 7034 35959 7037
rect 34697 7032 35959 7034
rect 34697 6976 34702 7032
rect 34758 6976 35898 7032
rect 35954 6976 35959 7032
rect 34697 6974 35959 6976
rect 34697 6971 34763 6974
rect 35893 6971 35959 6974
rect 67173 7034 67239 7037
rect 75913 7034 75979 7037
rect 67173 7032 75979 7034
rect 67173 6976 67178 7032
rect 67234 6976 75918 7032
rect 75974 6976 75979 7032
rect 67173 6974 75979 6976
rect 67173 6971 67239 6974
rect 75913 6971 75979 6974
rect 88241 7034 88307 7037
rect 89897 7034 89963 7037
rect 88241 7032 89963 7034
rect 88241 6976 88246 7032
rect 88302 6976 89902 7032
rect 89958 6976 89963 7032
rect 88241 6974 89963 6976
rect 88241 6971 88307 6974
rect 89897 6971 89963 6974
rect 26141 6898 26207 6901
rect 26693 6898 26759 6901
rect 26141 6896 26759 6898
rect 26141 6840 26146 6896
rect 26202 6840 26698 6896
rect 26754 6840 26759 6896
rect 26141 6838 26759 6840
rect 26141 6835 26207 6838
rect 26693 6835 26759 6838
rect 31201 6898 31267 6901
rect 38101 6898 38167 6901
rect 31201 6896 38167 6898
rect 31201 6840 31206 6896
rect 31262 6840 38106 6896
rect 38162 6840 38167 6896
rect 31201 6838 38167 6840
rect 31201 6835 31267 6838
rect 38101 6835 38167 6838
rect 50337 6898 50403 6901
rect 55213 6898 55279 6901
rect 50337 6896 55279 6898
rect 50337 6840 50342 6896
rect 50398 6840 55218 6896
rect 55274 6840 55279 6896
rect 50337 6838 55279 6840
rect 50337 6835 50403 6838
rect 55213 6835 55279 6838
rect 67817 6898 67883 6901
rect 68737 6898 68803 6901
rect 67817 6896 68803 6898
rect 67817 6840 67822 6896
rect 67878 6840 68742 6896
rect 68798 6840 68803 6896
rect 67817 6838 68803 6840
rect 67817 6835 67883 6838
rect 68737 6835 68803 6838
rect 71865 6898 71931 6901
rect 87873 6898 87939 6901
rect 89437 6898 89503 6901
rect 71865 6896 89503 6898
rect 71865 6840 71870 6896
rect 71926 6840 87878 6896
rect 87934 6840 89442 6896
rect 89498 6840 89503 6896
rect 71865 6838 89503 6840
rect 71865 6835 71931 6838
rect 87873 6835 87939 6838
rect 89437 6835 89503 6838
rect 25589 6762 25655 6765
rect 42425 6762 42491 6765
rect 25589 6760 42491 6762
rect 25589 6704 25594 6760
rect 25650 6704 42430 6760
rect 42486 6704 42491 6760
rect 25589 6702 42491 6704
rect 25589 6699 25655 6702
rect 42425 6699 42491 6702
rect 56961 6762 57027 6765
rect 72785 6762 72851 6765
rect 77293 6762 77359 6765
rect 56961 6760 71698 6762
rect 56961 6704 56966 6760
rect 57022 6704 71698 6760
rect 56961 6702 71698 6704
rect 56961 6699 57027 6702
rect 33041 6626 33107 6629
rect 36721 6626 36787 6629
rect 33041 6624 36787 6626
rect 33041 6568 33046 6624
rect 33102 6568 36726 6624
rect 36782 6568 36787 6624
rect 33041 6566 36787 6568
rect 33041 6563 33107 6566
rect 36721 6563 36787 6566
rect 24382 6560 24698 6561
rect 24382 6496 24388 6560
rect 24452 6496 24468 6560
rect 24532 6496 24548 6560
rect 24612 6496 24628 6560
rect 24692 6496 24698 6560
rect 24382 6495 24698 6496
rect 47819 6560 48135 6561
rect 47819 6496 47825 6560
rect 47889 6496 47905 6560
rect 47969 6496 47985 6560
rect 48049 6496 48065 6560
rect 48129 6496 48135 6560
rect 47819 6495 48135 6496
rect 71256 6560 71572 6561
rect 71256 6496 71262 6560
rect 71326 6496 71342 6560
rect 71406 6496 71422 6560
rect 71486 6496 71502 6560
rect 71566 6496 71572 6560
rect 71256 6495 71572 6496
rect 30465 6490 30531 6493
rect 34697 6490 34763 6493
rect 30465 6488 34763 6490
rect 30465 6432 30470 6488
rect 30526 6432 34702 6488
rect 34758 6432 34763 6488
rect 30465 6430 34763 6432
rect 30465 6427 30531 6430
rect 34697 6427 34763 6430
rect 48221 6490 48287 6493
rect 51717 6490 51783 6493
rect 48221 6488 51783 6490
rect 48221 6432 48226 6488
rect 48282 6432 51722 6488
rect 51778 6432 51783 6488
rect 48221 6430 51783 6432
rect 48221 6427 48287 6430
rect 51717 6427 51783 6430
rect 58709 6490 58775 6493
rect 66621 6490 66687 6493
rect 58709 6488 66687 6490
rect 58709 6432 58714 6488
rect 58770 6432 66626 6488
rect 66682 6432 66687 6488
rect 58709 6430 66687 6432
rect 71638 6490 71698 6702
rect 72785 6760 77359 6762
rect 72785 6704 72790 6760
rect 72846 6704 77298 6760
rect 77354 6704 77359 6760
rect 72785 6702 77359 6704
rect 72785 6699 72851 6702
rect 77293 6699 77359 6702
rect 80329 6762 80395 6765
rect 81709 6762 81775 6765
rect 80329 6760 81775 6762
rect 80329 6704 80334 6760
rect 80390 6704 81714 6760
rect 81770 6704 81775 6760
rect 80329 6702 81775 6704
rect 80329 6699 80395 6702
rect 81709 6699 81775 6702
rect 74993 6626 75059 6629
rect 76281 6626 76347 6629
rect 76557 6626 76623 6629
rect 74993 6624 76623 6626
rect 74993 6568 74998 6624
rect 75054 6568 76286 6624
rect 76342 6568 76562 6624
rect 76618 6568 76623 6624
rect 74993 6566 76623 6568
rect 74993 6563 75059 6566
rect 76281 6563 76347 6566
rect 76557 6563 76623 6566
rect 79961 6626 80027 6629
rect 80329 6626 80395 6629
rect 79961 6624 80395 6626
rect 79961 6568 79966 6624
rect 80022 6568 80334 6624
rect 80390 6568 80395 6624
rect 79961 6566 80395 6568
rect 79961 6563 80027 6566
rect 80329 6563 80395 6566
rect 94693 6560 95009 6561
rect 94693 6496 94699 6560
rect 94763 6496 94779 6560
rect 94843 6496 94859 6560
rect 94923 6496 94939 6560
rect 95003 6496 95009 6560
rect 94693 6495 95009 6496
rect 71957 6490 72023 6493
rect 71638 6488 72023 6490
rect 71638 6432 71962 6488
rect 72018 6432 72023 6488
rect 71638 6430 72023 6432
rect 58709 6427 58775 6430
rect 66621 6427 66687 6430
rect 71957 6427 72023 6430
rect 24761 6354 24827 6357
rect 26417 6354 26483 6357
rect 24761 6352 26483 6354
rect 24761 6296 24766 6352
rect 24822 6296 26422 6352
rect 26478 6296 26483 6352
rect 24761 6294 26483 6296
rect 24761 6291 24827 6294
rect 26417 6291 26483 6294
rect 32305 6354 32371 6357
rect 35801 6354 35867 6357
rect 32305 6352 35867 6354
rect 32305 6296 32310 6352
rect 32366 6296 35806 6352
rect 35862 6296 35867 6352
rect 32305 6294 35867 6296
rect 32305 6291 32371 6294
rect 35801 6291 35867 6294
rect 37549 6354 37615 6357
rect 53833 6354 53899 6357
rect 93209 6354 93275 6357
rect 37549 6352 53899 6354
rect 37549 6296 37554 6352
rect 37610 6296 53838 6352
rect 53894 6296 53899 6352
rect 37549 6294 53899 6296
rect 37549 6291 37615 6294
rect 53833 6291 53899 6294
rect 60690 6352 93275 6354
rect 60690 6296 93214 6352
rect 93270 6296 93275 6352
rect 60690 6294 93275 6296
rect 35617 6218 35683 6221
rect 38561 6218 38627 6221
rect 35617 6216 38627 6218
rect 35617 6160 35622 6216
rect 35678 6160 38566 6216
rect 38622 6160 38627 6216
rect 35617 6158 38627 6160
rect 35617 6155 35683 6158
rect 38561 6155 38627 6158
rect 53649 6218 53715 6221
rect 60690 6218 60750 6294
rect 93209 6291 93275 6294
rect 53649 6216 60750 6218
rect 53649 6160 53654 6216
rect 53710 6160 60750 6216
rect 53649 6158 60750 6160
rect 85757 6218 85823 6221
rect 86861 6218 86927 6221
rect 85757 6216 86927 6218
rect 85757 6160 85762 6216
rect 85818 6160 86866 6216
rect 86922 6160 86927 6216
rect 85757 6158 86927 6160
rect 53649 6155 53715 6158
rect 85757 6155 85823 6158
rect 86861 6155 86927 6158
rect 49969 6082 50035 6085
rect 54569 6082 54635 6085
rect 49969 6080 54635 6082
rect 49969 6024 49974 6080
rect 50030 6024 54574 6080
rect 54630 6024 54635 6080
rect 49969 6022 54635 6024
rect 49969 6019 50035 6022
rect 54569 6019 54635 6022
rect 75453 6082 75519 6085
rect 76741 6082 76807 6085
rect 75453 6080 76807 6082
rect 75453 6024 75458 6080
rect 75514 6024 76746 6080
rect 76802 6024 76807 6080
rect 75453 6022 76807 6024
rect 75453 6019 75519 6022
rect 76741 6019 76807 6022
rect 12664 6016 12980 6017
rect 12664 5952 12670 6016
rect 12734 5952 12750 6016
rect 12814 5952 12830 6016
rect 12894 5952 12910 6016
rect 12974 5952 12980 6016
rect 12664 5951 12980 5952
rect 36101 6016 36417 6017
rect 36101 5952 36107 6016
rect 36171 5952 36187 6016
rect 36251 5952 36267 6016
rect 36331 5952 36347 6016
rect 36411 5952 36417 6016
rect 36101 5951 36417 5952
rect 59538 6016 59854 6017
rect 59538 5952 59544 6016
rect 59608 5952 59624 6016
rect 59688 5952 59704 6016
rect 59768 5952 59784 6016
rect 59848 5952 59854 6016
rect 59538 5951 59854 5952
rect 82975 6016 83291 6017
rect 82975 5952 82981 6016
rect 83045 5952 83061 6016
rect 83125 5952 83141 6016
rect 83205 5952 83221 6016
rect 83285 5952 83291 6016
rect 82975 5951 83291 5952
rect 19885 5946 19951 5949
rect 25129 5946 25195 5949
rect 19885 5944 25195 5946
rect 19885 5888 19890 5944
rect 19946 5888 25134 5944
rect 25190 5888 25195 5944
rect 19885 5886 25195 5888
rect 19885 5883 19951 5886
rect 25129 5883 25195 5886
rect 49509 5946 49575 5949
rect 50797 5946 50863 5949
rect 49509 5944 50863 5946
rect 49509 5888 49514 5944
rect 49570 5888 50802 5944
rect 50858 5888 50863 5944
rect 49509 5886 50863 5888
rect 49509 5883 49575 5886
rect 50797 5883 50863 5886
rect 74073 5946 74139 5949
rect 76281 5946 76347 5949
rect 74073 5944 76347 5946
rect 74073 5888 74078 5944
rect 74134 5888 76286 5944
rect 76342 5888 76347 5944
rect 74073 5886 76347 5888
rect 74073 5883 74139 5886
rect 76281 5883 76347 5886
rect 77845 5946 77911 5949
rect 82721 5946 82787 5949
rect 77845 5944 82787 5946
rect 77845 5888 77850 5944
rect 77906 5888 82726 5944
rect 82782 5888 82787 5944
rect 77845 5886 82787 5888
rect 77845 5883 77911 5886
rect 82721 5883 82787 5886
rect 22921 5810 22987 5813
rect 27061 5810 27127 5813
rect 22921 5808 27127 5810
rect 22921 5752 22926 5808
rect 22982 5752 27066 5808
rect 27122 5752 27127 5808
rect 22921 5750 27127 5752
rect 22921 5747 22987 5750
rect 27061 5747 27127 5750
rect 48313 5810 48379 5813
rect 57145 5810 57211 5813
rect 48313 5808 57211 5810
rect 48313 5752 48318 5808
rect 48374 5752 57150 5808
rect 57206 5752 57211 5808
rect 48313 5750 57211 5752
rect 48313 5747 48379 5750
rect 57145 5747 57211 5750
rect 58801 5810 58867 5813
rect 60733 5810 60799 5813
rect 58801 5808 60799 5810
rect 58801 5752 58806 5808
rect 58862 5752 60738 5808
rect 60794 5752 60799 5808
rect 58801 5750 60799 5752
rect 58801 5747 58867 5750
rect 60733 5747 60799 5750
rect 69197 5810 69263 5813
rect 81249 5810 81315 5813
rect 69197 5808 81315 5810
rect 69197 5752 69202 5808
rect 69258 5752 81254 5808
rect 81310 5752 81315 5808
rect 69197 5750 81315 5752
rect 69197 5747 69263 5750
rect 81249 5747 81315 5750
rect 22645 5674 22711 5677
rect 24945 5674 25011 5677
rect 22645 5672 25011 5674
rect 22645 5616 22650 5672
rect 22706 5616 24950 5672
rect 25006 5616 25011 5672
rect 22645 5614 25011 5616
rect 22645 5611 22711 5614
rect 24945 5611 25011 5614
rect 32765 5674 32831 5677
rect 36537 5674 36603 5677
rect 32765 5672 36603 5674
rect 32765 5616 32770 5672
rect 32826 5616 36542 5672
rect 36598 5616 36603 5672
rect 32765 5614 36603 5616
rect 32765 5611 32831 5614
rect 36537 5611 36603 5614
rect 47301 5674 47367 5677
rect 81433 5674 81499 5677
rect 47301 5672 81499 5674
rect 47301 5616 47306 5672
rect 47362 5616 81438 5672
rect 81494 5616 81499 5672
rect 47301 5614 81499 5616
rect 47301 5611 47367 5614
rect 81433 5611 81499 5614
rect 71773 5538 71839 5541
rect 75269 5538 75335 5541
rect 71773 5536 75335 5538
rect 71773 5480 71778 5536
rect 71834 5480 75274 5536
rect 75330 5480 75335 5536
rect 71773 5478 75335 5480
rect 71773 5475 71839 5478
rect 75269 5475 75335 5478
rect 80053 5538 80119 5541
rect 81617 5538 81683 5541
rect 80053 5536 81683 5538
rect 80053 5480 80058 5536
rect 80114 5480 81622 5536
rect 81678 5480 81683 5536
rect 80053 5478 81683 5480
rect 80053 5475 80119 5478
rect 81617 5475 81683 5478
rect 24382 5472 24698 5473
rect 24382 5408 24388 5472
rect 24452 5408 24468 5472
rect 24532 5408 24548 5472
rect 24612 5408 24628 5472
rect 24692 5408 24698 5472
rect 24382 5407 24698 5408
rect 47819 5472 48135 5473
rect 47819 5408 47825 5472
rect 47889 5408 47905 5472
rect 47969 5408 47985 5472
rect 48049 5408 48065 5472
rect 48129 5408 48135 5472
rect 47819 5407 48135 5408
rect 71256 5472 71572 5473
rect 71256 5408 71262 5472
rect 71326 5408 71342 5472
rect 71406 5408 71422 5472
rect 71486 5408 71502 5472
rect 71566 5408 71572 5472
rect 71256 5407 71572 5408
rect 94693 5472 95009 5473
rect 94693 5408 94699 5472
rect 94763 5408 94779 5472
rect 94843 5408 94859 5472
rect 94923 5408 94939 5472
rect 95003 5408 95009 5472
rect 94693 5407 95009 5408
rect 43069 5402 43135 5405
rect 44173 5402 44239 5405
rect 43069 5400 44239 5402
rect 43069 5344 43074 5400
rect 43130 5344 44178 5400
rect 44234 5344 44239 5400
rect 43069 5342 44239 5344
rect 43069 5339 43135 5342
rect 44173 5339 44239 5342
rect 56041 5402 56107 5405
rect 58801 5402 58867 5405
rect 56041 5400 58867 5402
rect 56041 5344 56046 5400
rect 56102 5344 58806 5400
rect 58862 5344 58867 5400
rect 56041 5342 58867 5344
rect 56041 5339 56107 5342
rect 58801 5339 58867 5342
rect 28257 5266 28323 5269
rect 53649 5266 53715 5269
rect 28257 5264 53715 5266
rect 28257 5208 28262 5264
rect 28318 5208 53654 5264
rect 53710 5208 53715 5264
rect 28257 5206 53715 5208
rect 28257 5203 28323 5206
rect 53649 5203 53715 5206
rect 75545 5266 75611 5269
rect 76833 5266 76899 5269
rect 75545 5264 76899 5266
rect 75545 5208 75550 5264
rect 75606 5208 76838 5264
rect 76894 5208 76899 5264
rect 75545 5206 76899 5208
rect 75545 5203 75611 5206
rect 76833 5203 76899 5206
rect 9397 5130 9463 5133
rect 47485 5130 47551 5133
rect 9397 5128 47551 5130
rect 9397 5072 9402 5128
rect 9458 5072 47490 5128
rect 47546 5072 47551 5128
rect 9397 5070 47551 5072
rect 9397 5067 9463 5070
rect 47485 5067 47551 5070
rect 50613 5130 50679 5133
rect 56777 5130 56843 5133
rect 50613 5128 56843 5130
rect 50613 5072 50618 5128
rect 50674 5072 56782 5128
rect 56838 5072 56843 5128
rect 50613 5070 56843 5072
rect 50613 5067 50679 5070
rect 56777 5067 56843 5070
rect 24669 4994 24735 4997
rect 26417 4994 26483 4997
rect 24669 4992 26483 4994
rect 24669 4936 24674 4992
rect 24730 4936 26422 4992
rect 26478 4936 26483 4992
rect 24669 4934 26483 4936
rect 24669 4931 24735 4934
rect 26417 4931 26483 4934
rect 42977 4994 43043 4997
rect 47577 4994 47643 4997
rect 42977 4992 47643 4994
rect 42977 4936 42982 4992
rect 43038 4936 47582 4992
rect 47638 4936 47643 4992
rect 42977 4934 47643 4936
rect 42977 4931 43043 4934
rect 47577 4931 47643 4934
rect 51165 4994 51231 4997
rect 51533 4994 51599 4997
rect 56685 4994 56751 4997
rect 51165 4992 56751 4994
rect 51165 4936 51170 4992
rect 51226 4936 51538 4992
rect 51594 4936 56690 4992
rect 56746 4936 56751 4992
rect 51165 4934 56751 4936
rect 51165 4931 51231 4934
rect 51533 4931 51599 4934
rect 56685 4931 56751 4934
rect 12664 4928 12980 4929
rect 12664 4864 12670 4928
rect 12734 4864 12750 4928
rect 12814 4864 12830 4928
rect 12894 4864 12910 4928
rect 12974 4864 12980 4928
rect 12664 4863 12980 4864
rect 36101 4928 36417 4929
rect 36101 4864 36107 4928
rect 36171 4864 36187 4928
rect 36251 4864 36267 4928
rect 36331 4864 36347 4928
rect 36411 4864 36417 4928
rect 36101 4863 36417 4864
rect 59538 4928 59854 4929
rect 59538 4864 59544 4928
rect 59608 4864 59624 4928
rect 59688 4864 59704 4928
rect 59768 4864 59784 4928
rect 59848 4864 59854 4928
rect 59538 4863 59854 4864
rect 82975 4928 83291 4929
rect 82975 4864 82981 4928
rect 83045 4864 83061 4928
rect 83125 4864 83141 4928
rect 83205 4864 83221 4928
rect 83285 4864 83291 4928
rect 82975 4863 83291 4864
rect 63585 4860 63651 4861
rect 63534 4796 63540 4860
rect 63604 4858 63651 4860
rect 63604 4856 63696 4858
rect 63646 4800 63696 4856
rect 63604 4798 63696 4800
rect 63604 4796 63651 4798
rect 63585 4795 63651 4796
rect 34421 4722 34487 4725
rect 83917 4722 83983 4725
rect 34421 4720 83983 4722
rect 34421 4664 34426 4720
rect 34482 4664 83922 4720
rect 83978 4664 83983 4720
rect 34421 4662 83983 4664
rect 34421 4659 34487 4662
rect 83917 4659 83983 4662
rect 16389 4586 16455 4589
rect 38193 4586 38259 4589
rect 16389 4584 38259 4586
rect 16389 4528 16394 4584
rect 16450 4528 38198 4584
rect 38254 4528 38259 4584
rect 16389 4526 38259 4528
rect 16389 4523 16455 4526
rect 38193 4523 38259 4526
rect 45829 4586 45895 4589
rect 47485 4586 47551 4589
rect 45829 4584 47551 4586
rect 45829 4528 45834 4584
rect 45890 4528 47490 4584
rect 47546 4528 47551 4584
rect 45829 4526 47551 4528
rect 45829 4523 45895 4526
rect 47485 4523 47551 4526
rect 51993 4586 52059 4589
rect 57329 4586 57395 4589
rect 51993 4584 57395 4586
rect 51993 4528 51998 4584
rect 52054 4528 57334 4584
rect 57390 4528 57395 4584
rect 51993 4526 57395 4528
rect 51993 4523 52059 4526
rect 57329 4523 57395 4526
rect 24382 4384 24698 4385
rect 24382 4320 24388 4384
rect 24452 4320 24468 4384
rect 24532 4320 24548 4384
rect 24612 4320 24628 4384
rect 24692 4320 24698 4384
rect 24382 4319 24698 4320
rect 47819 4384 48135 4385
rect 47819 4320 47825 4384
rect 47889 4320 47905 4384
rect 47969 4320 47985 4384
rect 48049 4320 48065 4384
rect 48129 4320 48135 4384
rect 47819 4319 48135 4320
rect 71256 4384 71572 4385
rect 71256 4320 71262 4384
rect 71326 4320 71342 4384
rect 71406 4320 71422 4384
rect 71486 4320 71502 4384
rect 71566 4320 71572 4384
rect 71256 4319 71572 4320
rect 94693 4384 95009 4385
rect 94693 4320 94699 4384
rect 94763 4320 94779 4384
rect 94843 4320 94859 4384
rect 94923 4320 94939 4384
rect 95003 4320 95009 4384
rect 94693 4319 95009 4320
rect 10869 4178 10935 4181
rect 77569 4178 77635 4181
rect 10869 4176 77635 4178
rect 10869 4120 10874 4176
rect 10930 4120 77574 4176
rect 77630 4120 77635 4176
rect 10869 4118 77635 4120
rect 10869 4115 10935 4118
rect 77569 4115 77635 4118
rect 12664 3840 12980 3841
rect 12664 3776 12670 3840
rect 12734 3776 12750 3840
rect 12814 3776 12830 3840
rect 12894 3776 12910 3840
rect 12974 3776 12980 3840
rect 12664 3775 12980 3776
rect 36101 3840 36417 3841
rect 36101 3776 36107 3840
rect 36171 3776 36187 3840
rect 36251 3776 36267 3840
rect 36331 3776 36347 3840
rect 36411 3776 36417 3840
rect 36101 3775 36417 3776
rect 59538 3840 59854 3841
rect 59538 3776 59544 3840
rect 59608 3776 59624 3840
rect 59688 3776 59704 3840
rect 59768 3776 59784 3840
rect 59848 3776 59854 3840
rect 59538 3775 59854 3776
rect 82975 3840 83291 3841
rect 82975 3776 82981 3840
rect 83045 3776 83061 3840
rect 83125 3776 83141 3840
rect 83205 3776 83221 3840
rect 83285 3776 83291 3840
rect 82975 3775 83291 3776
rect 0 3362 800 3392
rect 4061 3362 4127 3365
rect 0 3360 4127 3362
rect 0 3304 4066 3360
rect 4122 3304 4127 3360
rect 0 3302 4127 3304
rect 0 3272 800 3302
rect 4061 3299 4127 3302
rect 24382 3296 24698 3297
rect 24382 3232 24388 3296
rect 24452 3232 24468 3296
rect 24532 3232 24548 3296
rect 24612 3232 24628 3296
rect 24692 3232 24698 3296
rect 24382 3231 24698 3232
rect 47819 3296 48135 3297
rect 47819 3232 47825 3296
rect 47889 3232 47905 3296
rect 47969 3232 47985 3296
rect 48049 3232 48065 3296
rect 48129 3232 48135 3296
rect 47819 3231 48135 3232
rect 71256 3296 71572 3297
rect 71256 3232 71262 3296
rect 71326 3232 71342 3296
rect 71406 3232 71422 3296
rect 71486 3232 71502 3296
rect 71566 3232 71572 3296
rect 71256 3231 71572 3232
rect 94693 3296 95009 3297
rect 94693 3232 94699 3296
rect 94763 3232 94779 3296
rect 94843 3232 94859 3296
rect 94923 3232 94939 3296
rect 95003 3232 95009 3296
rect 94693 3231 95009 3232
rect 12664 2752 12980 2753
rect 12664 2688 12670 2752
rect 12734 2688 12750 2752
rect 12814 2688 12830 2752
rect 12894 2688 12910 2752
rect 12974 2688 12980 2752
rect 12664 2687 12980 2688
rect 36101 2752 36417 2753
rect 36101 2688 36107 2752
rect 36171 2688 36187 2752
rect 36251 2688 36267 2752
rect 36331 2688 36347 2752
rect 36411 2688 36417 2752
rect 36101 2687 36417 2688
rect 59538 2752 59854 2753
rect 59538 2688 59544 2752
rect 59608 2688 59624 2752
rect 59688 2688 59704 2752
rect 59768 2688 59784 2752
rect 59848 2688 59854 2752
rect 59538 2687 59854 2688
rect 82975 2752 83291 2753
rect 82975 2688 82981 2752
rect 83045 2688 83061 2752
rect 83125 2688 83141 2752
rect 83205 2688 83221 2752
rect 83285 2688 83291 2752
rect 82975 2687 83291 2688
rect 93761 2682 93827 2685
rect 95200 2682 96000 2712
rect 93761 2680 96000 2682
rect 93761 2624 93766 2680
rect 93822 2624 96000 2680
rect 93761 2622 96000 2624
rect 93761 2619 93827 2622
rect 95200 2592 96000 2622
rect 24382 2208 24698 2209
rect 24382 2144 24388 2208
rect 24452 2144 24468 2208
rect 24532 2144 24548 2208
rect 24612 2144 24628 2208
rect 24692 2144 24698 2208
rect 24382 2143 24698 2144
rect 47819 2208 48135 2209
rect 47819 2144 47825 2208
rect 47889 2144 47905 2208
rect 47969 2144 47985 2208
rect 48049 2144 48065 2208
rect 48129 2144 48135 2208
rect 47819 2143 48135 2144
rect 71256 2208 71572 2209
rect 71256 2144 71262 2208
rect 71326 2144 71342 2208
rect 71406 2144 71422 2208
rect 71486 2144 71502 2208
rect 71566 2144 71572 2208
rect 71256 2143 71572 2144
rect 94693 2208 95009 2209
rect 94693 2144 94699 2208
rect 94763 2144 94779 2208
rect 94843 2144 94859 2208
rect 94923 2144 94939 2208
rect 95003 2144 95009 2208
rect 94693 2143 95009 2144
<< via3 >>
rect 24388 17436 24452 17440
rect 24388 17380 24392 17436
rect 24392 17380 24448 17436
rect 24448 17380 24452 17436
rect 24388 17376 24452 17380
rect 24468 17436 24532 17440
rect 24468 17380 24472 17436
rect 24472 17380 24528 17436
rect 24528 17380 24532 17436
rect 24468 17376 24532 17380
rect 24548 17436 24612 17440
rect 24548 17380 24552 17436
rect 24552 17380 24608 17436
rect 24608 17380 24612 17436
rect 24548 17376 24612 17380
rect 24628 17436 24692 17440
rect 24628 17380 24632 17436
rect 24632 17380 24688 17436
rect 24688 17380 24692 17436
rect 24628 17376 24692 17380
rect 47825 17436 47889 17440
rect 47825 17380 47829 17436
rect 47829 17380 47885 17436
rect 47885 17380 47889 17436
rect 47825 17376 47889 17380
rect 47905 17436 47969 17440
rect 47905 17380 47909 17436
rect 47909 17380 47965 17436
rect 47965 17380 47969 17436
rect 47905 17376 47969 17380
rect 47985 17436 48049 17440
rect 47985 17380 47989 17436
rect 47989 17380 48045 17436
rect 48045 17380 48049 17436
rect 47985 17376 48049 17380
rect 48065 17436 48129 17440
rect 48065 17380 48069 17436
rect 48069 17380 48125 17436
rect 48125 17380 48129 17436
rect 48065 17376 48129 17380
rect 71262 17436 71326 17440
rect 71262 17380 71266 17436
rect 71266 17380 71322 17436
rect 71322 17380 71326 17436
rect 71262 17376 71326 17380
rect 71342 17436 71406 17440
rect 71342 17380 71346 17436
rect 71346 17380 71402 17436
rect 71402 17380 71406 17436
rect 71342 17376 71406 17380
rect 71422 17436 71486 17440
rect 71422 17380 71426 17436
rect 71426 17380 71482 17436
rect 71482 17380 71486 17436
rect 71422 17376 71486 17380
rect 71502 17436 71566 17440
rect 71502 17380 71506 17436
rect 71506 17380 71562 17436
rect 71562 17380 71566 17436
rect 71502 17376 71566 17380
rect 94699 17436 94763 17440
rect 94699 17380 94703 17436
rect 94703 17380 94759 17436
rect 94759 17380 94763 17436
rect 94699 17376 94763 17380
rect 94779 17436 94843 17440
rect 94779 17380 94783 17436
rect 94783 17380 94839 17436
rect 94839 17380 94843 17436
rect 94779 17376 94843 17380
rect 94859 17436 94923 17440
rect 94859 17380 94863 17436
rect 94863 17380 94919 17436
rect 94919 17380 94923 17436
rect 94859 17376 94923 17380
rect 94939 17436 95003 17440
rect 94939 17380 94943 17436
rect 94943 17380 94999 17436
rect 94999 17380 95003 17436
rect 94939 17376 95003 17380
rect 12670 16892 12734 16896
rect 12670 16836 12674 16892
rect 12674 16836 12730 16892
rect 12730 16836 12734 16892
rect 12670 16832 12734 16836
rect 12750 16892 12814 16896
rect 12750 16836 12754 16892
rect 12754 16836 12810 16892
rect 12810 16836 12814 16892
rect 12750 16832 12814 16836
rect 12830 16892 12894 16896
rect 12830 16836 12834 16892
rect 12834 16836 12890 16892
rect 12890 16836 12894 16892
rect 12830 16832 12894 16836
rect 12910 16892 12974 16896
rect 12910 16836 12914 16892
rect 12914 16836 12970 16892
rect 12970 16836 12974 16892
rect 12910 16832 12974 16836
rect 36107 16892 36171 16896
rect 36107 16836 36111 16892
rect 36111 16836 36167 16892
rect 36167 16836 36171 16892
rect 36107 16832 36171 16836
rect 36187 16892 36251 16896
rect 36187 16836 36191 16892
rect 36191 16836 36247 16892
rect 36247 16836 36251 16892
rect 36187 16832 36251 16836
rect 36267 16892 36331 16896
rect 36267 16836 36271 16892
rect 36271 16836 36327 16892
rect 36327 16836 36331 16892
rect 36267 16832 36331 16836
rect 36347 16892 36411 16896
rect 36347 16836 36351 16892
rect 36351 16836 36407 16892
rect 36407 16836 36411 16892
rect 36347 16832 36411 16836
rect 59544 16892 59608 16896
rect 59544 16836 59548 16892
rect 59548 16836 59604 16892
rect 59604 16836 59608 16892
rect 59544 16832 59608 16836
rect 59624 16892 59688 16896
rect 59624 16836 59628 16892
rect 59628 16836 59684 16892
rect 59684 16836 59688 16892
rect 59624 16832 59688 16836
rect 59704 16892 59768 16896
rect 59704 16836 59708 16892
rect 59708 16836 59764 16892
rect 59764 16836 59768 16892
rect 59704 16832 59768 16836
rect 59784 16892 59848 16896
rect 59784 16836 59788 16892
rect 59788 16836 59844 16892
rect 59844 16836 59848 16892
rect 59784 16832 59848 16836
rect 82981 16892 83045 16896
rect 82981 16836 82985 16892
rect 82985 16836 83041 16892
rect 83041 16836 83045 16892
rect 82981 16832 83045 16836
rect 83061 16892 83125 16896
rect 83061 16836 83065 16892
rect 83065 16836 83121 16892
rect 83121 16836 83125 16892
rect 83061 16832 83125 16836
rect 83141 16892 83205 16896
rect 83141 16836 83145 16892
rect 83145 16836 83201 16892
rect 83201 16836 83205 16892
rect 83141 16832 83205 16836
rect 83221 16892 83285 16896
rect 83221 16836 83225 16892
rect 83225 16836 83281 16892
rect 83281 16836 83285 16892
rect 83221 16832 83285 16836
rect 24388 16348 24452 16352
rect 24388 16292 24392 16348
rect 24392 16292 24448 16348
rect 24448 16292 24452 16348
rect 24388 16288 24452 16292
rect 24468 16348 24532 16352
rect 24468 16292 24472 16348
rect 24472 16292 24528 16348
rect 24528 16292 24532 16348
rect 24468 16288 24532 16292
rect 24548 16348 24612 16352
rect 24548 16292 24552 16348
rect 24552 16292 24608 16348
rect 24608 16292 24612 16348
rect 24548 16288 24612 16292
rect 24628 16348 24692 16352
rect 24628 16292 24632 16348
rect 24632 16292 24688 16348
rect 24688 16292 24692 16348
rect 24628 16288 24692 16292
rect 47825 16348 47889 16352
rect 47825 16292 47829 16348
rect 47829 16292 47885 16348
rect 47885 16292 47889 16348
rect 47825 16288 47889 16292
rect 47905 16348 47969 16352
rect 47905 16292 47909 16348
rect 47909 16292 47965 16348
rect 47965 16292 47969 16348
rect 47905 16288 47969 16292
rect 47985 16348 48049 16352
rect 47985 16292 47989 16348
rect 47989 16292 48045 16348
rect 48045 16292 48049 16348
rect 47985 16288 48049 16292
rect 48065 16348 48129 16352
rect 48065 16292 48069 16348
rect 48069 16292 48125 16348
rect 48125 16292 48129 16348
rect 48065 16288 48129 16292
rect 71262 16348 71326 16352
rect 71262 16292 71266 16348
rect 71266 16292 71322 16348
rect 71322 16292 71326 16348
rect 71262 16288 71326 16292
rect 71342 16348 71406 16352
rect 71342 16292 71346 16348
rect 71346 16292 71402 16348
rect 71402 16292 71406 16348
rect 71342 16288 71406 16292
rect 71422 16348 71486 16352
rect 71422 16292 71426 16348
rect 71426 16292 71482 16348
rect 71482 16292 71486 16348
rect 71422 16288 71486 16292
rect 71502 16348 71566 16352
rect 71502 16292 71506 16348
rect 71506 16292 71562 16348
rect 71562 16292 71566 16348
rect 71502 16288 71566 16292
rect 94699 16348 94763 16352
rect 94699 16292 94703 16348
rect 94703 16292 94759 16348
rect 94759 16292 94763 16348
rect 94699 16288 94763 16292
rect 94779 16348 94843 16352
rect 94779 16292 94783 16348
rect 94783 16292 94839 16348
rect 94839 16292 94843 16348
rect 94779 16288 94843 16292
rect 94859 16348 94923 16352
rect 94859 16292 94863 16348
rect 94863 16292 94919 16348
rect 94919 16292 94923 16348
rect 94859 16288 94923 16292
rect 94939 16348 95003 16352
rect 94939 16292 94943 16348
rect 94943 16292 94999 16348
rect 94999 16292 95003 16348
rect 94939 16288 95003 16292
rect 12670 15804 12734 15808
rect 12670 15748 12674 15804
rect 12674 15748 12730 15804
rect 12730 15748 12734 15804
rect 12670 15744 12734 15748
rect 12750 15804 12814 15808
rect 12750 15748 12754 15804
rect 12754 15748 12810 15804
rect 12810 15748 12814 15804
rect 12750 15744 12814 15748
rect 12830 15804 12894 15808
rect 12830 15748 12834 15804
rect 12834 15748 12890 15804
rect 12890 15748 12894 15804
rect 12830 15744 12894 15748
rect 12910 15804 12974 15808
rect 12910 15748 12914 15804
rect 12914 15748 12970 15804
rect 12970 15748 12974 15804
rect 12910 15744 12974 15748
rect 36107 15804 36171 15808
rect 36107 15748 36111 15804
rect 36111 15748 36167 15804
rect 36167 15748 36171 15804
rect 36107 15744 36171 15748
rect 36187 15804 36251 15808
rect 36187 15748 36191 15804
rect 36191 15748 36247 15804
rect 36247 15748 36251 15804
rect 36187 15744 36251 15748
rect 36267 15804 36331 15808
rect 36267 15748 36271 15804
rect 36271 15748 36327 15804
rect 36327 15748 36331 15804
rect 36267 15744 36331 15748
rect 36347 15804 36411 15808
rect 36347 15748 36351 15804
rect 36351 15748 36407 15804
rect 36407 15748 36411 15804
rect 36347 15744 36411 15748
rect 59544 15804 59608 15808
rect 59544 15748 59548 15804
rect 59548 15748 59604 15804
rect 59604 15748 59608 15804
rect 59544 15744 59608 15748
rect 59624 15804 59688 15808
rect 59624 15748 59628 15804
rect 59628 15748 59684 15804
rect 59684 15748 59688 15804
rect 59624 15744 59688 15748
rect 59704 15804 59768 15808
rect 59704 15748 59708 15804
rect 59708 15748 59764 15804
rect 59764 15748 59768 15804
rect 59704 15744 59768 15748
rect 59784 15804 59848 15808
rect 59784 15748 59788 15804
rect 59788 15748 59844 15804
rect 59844 15748 59848 15804
rect 59784 15744 59848 15748
rect 82981 15804 83045 15808
rect 82981 15748 82985 15804
rect 82985 15748 83041 15804
rect 83041 15748 83045 15804
rect 82981 15744 83045 15748
rect 83061 15804 83125 15808
rect 83061 15748 83065 15804
rect 83065 15748 83121 15804
rect 83121 15748 83125 15804
rect 83061 15744 83125 15748
rect 83141 15804 83205 15808
rect 83141 15748 83145 15804
rect 83145 15748 83201 15804
rect 83201 15748 83205 15804
rect 83141 15744 83205 15748
rect 83221 15804 83285 15808
rect 83221 15748 83225 15804
rect 83225 15748 83281 15804
rect 83281 15748 83285 15804
rect 83221 15744 83285 15748
rect 24388 15260 24452 15264
rect 24388 15204 24392 15260
rect 24392 15204 24448 15260
rect 24448 15204 24452 15260
rect 24388 15200 24452 15204
rect 24468 15260 24532 15264
rect 24468 15204 24472 15260
rect 24472 15204 24528 15260
rect 24528 15204 24532 15260
rect 24468 15200 24532 15204
rect 24548 15260 24612 15264
rect 24548 15204 24552 15260
rect 24552 15204 24608 15260
rect 24608 15204 24612 15260
rect 24548 15200 24612 15204
rect 24628 15260 24692 15264
rect 24628 15204 24632 15260
rect 24632 15204 24688 15260
rect 24688 15204 24692 15260
rect 24628 15200 24692 15204
rect 47825 15260 47889 15264
rect 47825 15204 47829 15260
rect 47829 15204 47885 15260
rect 47885 15204 47889 15260
rect 47825 15200 47889 15204
rect 47905 15260 47969 15264
rect 47905 15204 47909 15260
rect 47909 15204 47965 15260
rect 47965 15204 47969 15260
rect 47905 15200 47969 15204
rect 47985 15260 48049 15264
rect 47985 15204 47989 15260
rect 47989 15204 48045 15260
rect 48045 15204 48049 15260
rect 47985 15200 48049 15204
rect 48065 15260 48129 15264
rect 48065 15204 48069 15260
rect 48069 15204 48125 15260
rect 48125 15204 48129 15260
rect 48065 15200 48129 15204
rect 71262 15260 71326 15264
rect 71262 15204 71266 15260
rect 71266 15204 71322 15260
rect 71322 15204 71326 15260
rect 71262 15200 71326 15204
rect 71342 15260 71406 15264
rect 71342 15204 71346 15260
rect 71346 15204 71402 15260
rect 71402 15204 71406 15260
rect 71342 15200 71406 15204
rect 71422 15260 71486 15264
rect 71422 15204 71426 15260
rect 71426 15204 71482 15260
rect 71482 15204 71486 15260
rect 71422 15200 71486 15204
rect 71502 15260 71566 15264
rect 71502 15204 71506 15260
rect 71506 15204 71562 15260
rect 71562 15204 71566 15260
rect 71502 15200 71566 15204
rect 94699 15260 94763 15264
rect 94699 15204 94703 15260
rect 94703 15204 94759 15260
rect 94759 15204 94763 15260
rect 94699 15200 94763 15204
rect 94779 15260 94843 15264
rect 94779 15204 94783 15260
rect 94783 15204 94839 15260
rect 94839 15204 94843 15260
rect 94779 15200 94843 15204
rect 94859 15260 94923 15264
rect 94859 15204 94863 15260
rect 94863 15204 94919 15260
rect 94919 15204 94923 15260
rect 94859 15200 94923 15204
rect 94939 15260 95003 15264
rect 94939 15204 94943 15260
rect 94943 15204 94999 15260
rect 94999 15204 95003 15260
rect 94939 15200 95003 15204
rect 12670 14716 12734 14720
rect 12670 14660 12674 14716
rect 12674 14660 12730 14716
rect 12730 14660 12734 14716
rect 12670 14656 12734 14660
rect 12750 14716 12814 14720
rect 12750 14660 12754 14716
rect 12754 14660 12810 14716
rect 12810 14660 12814 14716
rect 12750 14656 12814 14660
rect 12830 14716 12894 14720
rect 12830 14660 12834 14716
rect 12834 14660 12890 14716
rect 12890 14660 12894 14716
rect 12830 14656 12894 14660
rect 12910 14716 12974 14720
rect 12910 14660 12914 14716
rect 12914 14660 12970 14716
rect 12970 14660 12974 14716
rect 12910 14656 12974 14660
rect 36107 14716 36171 14720
rect 36107 14660 36111 14716
rect 36111 14660 36167 14716
rect 36167 14660 36171 14716
rect 36107 14656 36171 14660
rect 36187 14716 36251 14720
rect 36187 14660 36191 14716
rect 36191 14660 36247 14716
rect 36247 14660 36251 14716
rect 36187 14656 36251 14660
rect 36267 14716 36331 14720
rect 36267 14660 36271 14716
rect 36271 14660 36327 14716
rect 36327 14660 36331 14716
rect 36267 14656 36331 14660
rect 36347 14716 36411 14720
rect 36347 14660 36351 14716
rect 36351 14660 36407 14716
rect 36407 14660 36411 14716
rect 36347 14656 36411 14660
rect 59544 14716 59608 14720
rect 59544 14660 59548 14716
rect 59548 14660 59604 14716
rect 59604 14660 59608 14716
rect 59544 14656 59608 14660
rect 59624 14716 59688 14720
rect 59624 14660 59628 14716
rect 59628 14660 59684 14716
rect 59684 14660 59688 14716
rect 59624 14656 59688 14660
rect 59704 14716 59768 14720
rect 59704 14660 59708 14716
rect 59708 14660 59764 14716
rect 59764 14660 59768 14716
rect 59704 14656 59768 14660
rect 59784 14716 59848 14720
rect 59784 14660 59788 14716
rect 59788 14660 59844 14716
rect 59844 14660 59848 14716
rect 59784 14656 59848 14660
rect 82981 14716 83045 14720
rect 82981 14660 82985 14716
rect 82985 14660 83041 14716
rect 83041 14660 83045 14716
rect 82981 14656 83045 14660
rect 83061 14716 83125 14720
rect 83061 14660 83065 14716
rect 83065 14660 83121 14716
rect 83121 14660 83125 14716
rect 83061 14656 83125 14660
rect 83141 14716 83205 14720
rect 83141 14660 83145 14716
rect 83145 14660 83201 14716
rect 83201 14660 83205 14716
rect 83141 14656 83205 14660
rect 83221 14716 83285 14720
rect 83221 14660 83225 14716
rect 83225 14660 83281 14716
rect 83281 14660 83285 14716
rect 83221 14656 83285 14660
rect 24388 14172 24452 14176
rect 24388 14116 24392 14172
rect 24392 14116 24448 14172
rect 24448 14116 24452 14172
rect 24388 14112 24452 14116
rect 24468 14172 24532 14176
rect 24468 14116 24472 14172
rect 24472 14116 24528 14172
rect 24528 14116 24532 14172
rect 24468 14112 24532 14116
rect 24548 14172 24612 14176
rect 24548 14116 24552 14172
rect 24552 14116 24608 14172
rect 24608 14116 24612 14172
rect 24548 14112 24612 14116
rect 24628 14172 24692 14176
rect 24628 14116 24632 14172
rect 24632 14116 24688 14172
rect 24688 14116 24692 14172
rect 24628 14112 24692 14116
rect 47825 14172 47889 14176
rect 47825 14116 47829 14172
rect 47829 14116 47885 14172
rect 47885 14116 47889 14172
rect 47825 14112 47889 14116
rect 47905 14172 47969 14176
rect 47905 14116 47909 14172
rect 47909 14116 47965 14172
rect 47965 14116 47969 14172
rect 47905 14112 47969 14116
rect 47985 14172 48049 14176
rect 47985 14116 47989 14172
rect 47989 14116 48045 14172
rect 48045 14116 48049 14172
rect 47985 14112 48049 14116
rect 48065 14172 48129 14176
rect 48065 14116 48069 14172
rect 48069 14116 48125 14172
rect 48125 14116 48129 14172
rect 48065 14112 48129 14116
rect 71262 14172 71326 14176
rect 71262 14116 71266 14172
rect 71266 14116 71322 14172
rect 71322 14116 71326 14172
rect 71262 14112 71326 14116
rect 71342 14172 71406 14176
rect 71342 14116 71346 14172
rect 71346 14116 71402 14172
rect 71402 14116 71406 14172
rect 71342 14112 71406 14116
rect 71422 14172 71486 14176
rect 71422 14116 71426 14172
rect 71426 14116 71482 14172
rect 71482 14116 71486 14172
rect 71422 14112 71486 14116
rect 71502 14172 71566 14176
rect 71502 14116 71506 14172
rect 71506 14116 71562 14172
rect 71562 14116 71566 14172
rect 71502 14112 71566 14116
rect 94699 14172 94763 14176
rect 94699 14116 94703 14172
rect 94703 14116 94759 14172
rect 94759 14116 94763 14172
rect 94699 14112 94763 14116
rect 94779 14172 94843 14176
rect 94779 14116 94783 14172
rect 94783 14116 94839 14172
rect 94839 14116 94843 14172
rect 94779 14112 94843 14116
rect 94859 14172 94923 14176
rect 94859 14116 94863 14172
rect 94863 14116 94919 14172
rect 94919 14116 94923 14172
rect 94859 14112 94923 14116
rect 94939 14172 95003 14176
rect 94939 14116 94943 14172
rect 94943 14116 94999 14172
rect 94999 14116 95003 14172
rect 94939 14112 95003 14116
rect 12670 13628 12734 13632
rect 12670 13572 12674 13628
rect 12674 13572 12730 13628
rect 12730 13572 12734 13628
rect 12670 13568 12734 13572
rect 12750 13628 12814 13632
rect 12750 13572 12754 13628
rect 12754 13572 12810 13628
rect 12810 13572 12814 13628
rect 12750 13568 12814 13572
rect 12830 13628 12894 13632
rect 12830 13572 12834 13628
rect 12834 13572 12890 13628
rect 12890 13572 12894 13628
rect 12830 13568 12894 13572
rect 12910 13628 12974 13632
rect 12910 13572 12914 13628
rect 12914 13572 12970 13628
rect 12970 13572 12974 13628
rect 12910 13568 12974 13572
rect 36107 13628 36171 13632
rect 36107 13572 36111 13628
rect 36111 13572 36167 13628
rect 36167 13572 36171 13628
rect 36107 13568 36171 13572
rect 36187 13628 36251 13632
rect 36187 13572 36191 13628
rect 36191 13572 36247 13628
rect 36247 13572 36251 13628
rect 36187 13568 36251 13572
rect 36267 13628 36331 13632
rect 36267 13572 36271 13628
rect 36271 13572 36327 13628
rect 36327 13572 36331 13628
rect 36267 13568 36331 13572
rect 36347 13628 36411 13632
rect 36347 13572 36351 13628
rect 36351 13572 36407 13628
rect 36407 13572 36411 13628
rect 36347 13568 36411 13572
rect 59544 13628 59608 13632
rect 59544 13572 59548 13628
rect 59548 13572 59604 13628
rect 59604 13572 59608 13628
rect 59544 13568 59608 13572
rect 59624 13628 59688 13632
rect 59624 13572 59628 13628
rect 59628 13572 59684 13628
rect 59684 13572 59688 13628
rect 59624 13568 59688 13572
rect 59704 13628 59768 13632
rect 59704 13572 59708 13628
rect 59708 13572 59764 13628
rect 59764 13572 59768 13628
rect 59704 13568 59768 13572
rect 59784 13628 59848 13632
rect 59784 13572 59788 13628
rect 59788 13572 59844 13628
rect 59844 13572 59848 13628
rect 59784 13568 59848 13572
rect 82981 13628 83045 13632
rect 82981 13572 82985 13628
rect 82985 13572 83041 13628
rect 83041 13572 83045 13628
rect 82981 13568 83045 13572
rect 83061 13628 83125 13632
rect 83061 13572 83065 13628
rect 83065 13572 83121 13628
rect 83121 13572 83125 13628
rect 83061 13568 83125 13572
rect 83141 13628 83205 13632
rect 83141 13572 83145 13628
rect 83145 13572 83201 13628
rect 83201 13572 83205 13628
rect 83141 13568 83205 13572
rect 83221 13628 83285 13632
rect 83221 13572 83225 13628
rect 83225 13572 83281 13628
rect 83281 13572 83285 13628
rect 83221 13568 83285 13572
rect 60228 13092 60292 13156
rect 24388 13084 24452 13088
rect 24388 13028 24392 13084
rect 24392 13028 24448 13084
rect 24448 13028 24452 13084
rect 24388 13024 24452 13028
rect 24468 13084 24532 13088
rect 24468 13028 24472 13084
rect 24472 13028 24528 13084
rect 24528 13028 24532 13084
rect 24468 13024 24532 13028
rect 24548 13084 24612 13088
rect 24548 13028 24552 13084
rect 24552 13028 24608 13084
rect 24608 13028 24612 13084
rect 24548 13024 24612 13028
rect 24628 13084 24692 13088
rect 24628 13028 24632 13084
rect 24632 13028 24688 13084
rect 24688 13028 24692 13084
rect 24628 13024 24692 13028
rect 47825 13084 47889 13088
rect 47825 13028 47829 13084
rect 47829 13028 47885 13084
rect 47885 13028 47889 13084
rect 47825 13024 47889 13028
rect 47905 13084 47969 13088
rect 47905 13028 47909 13084
rect 47909 13028 47965 13084
rect 47965 13028 47969 13084
rect 47905 13024 47969 13028
rect 47985 13084 48049 13088
rect 47985 13028 47989 13084
rect 47989 13028 48045 13084
rect 48045 13028 48049 13084
rect 47985 13024 48049 13028
rect 48065 13084 48129 13088
rect 48065 13028 48069 13084
rect 48069 13028 48125 13084
rect 48125 13028 48129 13084
rect 48065 13024 48129 13028
rect 71262 13084 71326 13088
rect 71262 13028 71266 13084
rect 71266 13028 71322 13084
rect 71322 13028 71326 13084
rect 71262 13024 71326 13028
rect 71342 13084 71406 13088
rect 71342 13028 71346 13084
rect 71346 13028 71402 13084
rect 71402 13028 71406 13084
rect 71342 13024 71406 13028
rect 71422 13084 71486 13088
rect 71422 13028 71426 13084
rect 71426 13028 71482 13084
rect 71482 13028 71486 13084
rect 71422 13024 71486 13028
rect 71502 13084 71566 13088
rect 71502 13028 71506 13084
rect 71506 13028 71562 13084
rect 71562 13028 71566 13084
rect 71502 13024 71566 13028
rect 94699 13084 94763 13088
rect 94699 13028 94703 13084
rect 94703 13028 94759 13084
rect 94759 13028 94763 13084
rect 94699 13024 94763 13028
rect 94779 13084 94843 13088
rect 94779 13028 94783 13084
rect 94783 13028 94839 13084
rect 94839 13028 94843 13084
rect 94779 13024 94843 13028
rect 94859 13084 94923 13088
rect 94859 13028 94863 13084
rect 94863 13028 94919 13084
rect 94919 13028 94923 13084
rect 94859 13024 94923 13028
rect 94939 13084 95003 13088
rect 94939 13028 94943 13084
rect 94943 13028 94999 13084
rect 94999 13028 95003 13084
rect 94939 13024 95003 13028
rect 12670 12540 12734 12544
rect 12670 12484 12674 12540
rect 12674 12484 12730 12540
rect 12730 12484 12734 12540
rect 12670 12480 12734 12484
rect 12750 12540 12814 12544
rect 12750 12484 12754 12540
rect 12754 12484 12810 12540
rect 12810 12484 12814 12540
rect 12750 12480 12814 12484
rect 12830 12540 12894 12544
rect 12830 12484 12834 12540
rect 12834 12484 12890 12540
rect 12890 12484 12894 12540
rect 12830 12480 12894 12484
rect 12910 12540 12974 12544
rect 12910 12484 12914 12540
rect 12914 12484 12970 12540
rect 12970 12484 12974 12540
rect 12910 12480 12974 12484
rect 36107 12540 36171 12544
rect 36107 12484 36111 12540
rect 36111 12484 36167 12540
rect 36167 12484 36171 12540
rect 36107 12480 36171 12484
rect 36187 12540 36251 12544
rect 36187 12484 36191 12540
rect 36191 12484 36247 12540
rect 36247 12484 36251 12540
rect 36187 12480 36251 12484
rect 36267 12540 36331 12544
rect 36267 12484 36271 12540
rect 36271 12484 36327 12540
rect 36327 12484 36331 12540
rect 36267 12480 36331 12484
rect 36347 12540 36411 12544
rect 36347 12484 36351 12540
rect 36351 12484 36407 12540
rect 36407 12484 36411 12540
rect 36347 12480 36411 12484
rect 59544 12540 59608 12544
rect 59544 12484 59548 12540
rect 59548 12484 59604 12540
rect 59604 12484 59608 12540
rect 59544 12480 59608 12484
rect 59624 12540 59688 12544
rect 59624 12484 59628 12540
rect 59628 12484 59684 12540
rect 59684 12484 59688 12540
rect 59624 12480 59688 12484
rect 59704 12540 59768 12544
rect 59704 12484 59708 12540
rect 59708 12484 59764 12540
rect 59764 12484 59768 12540
rect 59704 12480 59768 12484
rect 59784 12540 59848 12544
rect 59784 12484 59788 12540
rect 59788 12484 59844 12540
rect 59844 12484 59848 12540
rect 59784 12480 59848 12484
rect 60228 12684 60292 12748
rect 82981 12540 83045 12544
rect 82981 12484 82985 12540
rect 82985 12484 83041 12540
rect 83041 12484 83045 12540
rect 82981 12480 83045 12484
rect 83061 12540 83125 12544
rect 83061 12484 83065 12540
rect 83065 12484 83121 12540
rect 83121 12484 83125 12540
rect 83061 12480 83125 12484
rect 83141 12540 83205 12544
rect 83141 12484 83145 12540
rect 83145 12484 83201 12540
rect 83201 12484 83205 12540
rect 83141 12480 83205 12484
rect 83221 12540 83285 12544
rect 83221 12484 83225 12540
rect 83225 12484 83281 12540
rect 83281 12484 83285 12540
rect 83221 12480 83285 12484
rect 24388 11996 24452 12000
rect 24388 11940 24392 11996
rect 24392 11940 24448 11996
rect 24448 11940 24452 11996
rect 24388 11936 24452 11940
rect 24468 11996 24532 12000
rect 24468 11940 24472 11996
rect 24472 11940 24528 11996
rect 24528 11940 24532 11996
rect 24468 11936 24532 11940
rect 24548 11996 24612 12000
rect 24548 11940 24552 11996
rect 24552 11940 24608 11996
rect 24608 11940 24612 11996
rect 24548 11936 24612 11940
rect 24628 11996 24692 12000
rect 24628 11940 24632 11996
rect 24632 11940 24688 11996
rect 24688 11940 24692 11996
rect 24628 11936 24692 11940
rect 47825 11996 47889 12000
rect 47825 11940 47829 11996
rect 47829 11940 47885 11996
rect 47885 11940 47889 11996
rect 47825 11936 47889 11940
rect 47905 11996 47969 12000
rect 47905 11940 47909 11996
rect 47909 11940 47965 11996
rect 47965 11940 47969 11996
rect 47905 11936 47969 11940
rect 47985 11996 48049 12000
rect 47985 11940 47989 11996
rect 47989 11940 48045 11996
rect 48045 11940 48049 11996
rect 47985 11936 48049 11940
rect 48065 11996 48129 12000
rect 48065 11940 48069 11996
rect 48069 11940 48125 11996
rect 48125 11940 48129 11996
rect 48065 11936 48129 11940
rect 71262 11996 71326 12000
rect 71262 11940 71266 11996
rect 71266 11940 71322 11996
rect 71322 11940 71326 11996
rect 71262 11936 71326 11940
rect 71342 11996 71406 12000
rect 71342 11940 71346 11996
rect 71346 11940 71402 11996
rect 71402 11940 71406 11996
rect 71342 11936 71406 11940
rect 71422 11996 71486 12000
rect 71422 11940 71426 11996
rect 71426 11940 71482 11996
rect 71482 11940 71486 11996
rect 71422 11936 71486 11940
rect 71502 11996 71566 12000
rect 71502 11940 71506 11996
rect 71506 11940 71562 11996
rect 71562 11940 71566 11996
rect 71502 11936 71566 11940
rect 94699 11996 94763 12000
rect 94699 11940 94703 11996
rect 94703 11940 94759 11996
rect 94759 11940 94763 11996
rect 94699 11936 94763 11940
rect 94779 11996 94843 12000
rect 94779 11940 94783 11996
rect 94783 11940 94839 11996
rect 94839 11940 94843 11996
rect 94779 11936 94843 11940
rect 94859 11996 94923 12000
rect 94859 11940 94863 11996
rect 94863 11940 94919 11996
rect 94919 11940 94923 11996
rect 94859 11936 94923 11940
rect 94939 11996 95003 12000
rect 94939 11940 94943 11996
rect 94943 11940 94999 11996
rect 94999 11940 95003 11996
rect 94939 11936 95003 11940
rect 12670 11452 12734 11456
rect 12670 11396 12674 11452
rect 12674 11396 12730 11452
rect 12730 11396 12734 11452
rect 12670 11392 12734 11396
rect 12750 11452 12814 11456
rect 12750 11396 12754 11452
rect 12754 11396 12810 11452
rect 12810 11396 12814 11452
rect 12750 11392 12814 11396
rect 12830 11452 12894 11456
rect 12830 11396 12834 11452
rect 12834 11396 12890 11452
rect 12890 11396 12894 11452
rect 12830 11392 12894 11396
rect 12910 11452 12974 11456
rect 12910 11396 12914 11452
rect 12914 11396 12970 11452
rect 12970 11396 12974 11452
rect 12910 11392 12974 11396
rect 36107 11452 36171 11456
rect 36107 11396 36111 11452
rect 36111 11396 36167 11452
rect 36167 11396 36171 11452
rect 36107 11392 36171 11396
rect 36187 11452 36251 11456
rect 36187 11396 36191 11452
rect 36191 11396 36247 11452
rect 36247 11396 36251 11452
rect 36187 11392 36251 11396
rect 36267 11452 36331 11456
rect 36267 11396 36271 11452
rect 36271 11396 36327 11452
rect 36327 11396 36331 11452
rect 36267 11392 36331 11396
rect 36347 11452 36411 11456
rect 36347 11396 36351 11452
rect 36351 11396 36407 11452
rect 36407 11396 36411 11452
rect 36347 11392 36411 11396
rect 59544 11452 59608 11456
rect 59544 11396 59548 11452
rect 59548 11396 59604 11452
rect 59604 11396 59608 11452
rect 59544 11392 59608 11396
rect 59624 11452 59688 11456
rect 59624 11396 59628 11452
rect 59628 11396 59684 11452
rect 59684 11396 59688 11452
rect 59624 11392 59688 11396
rect 59704 11452 59768 11456
rect 59704 11396 59708 11452
rect 59708 11396 59764 11452
rect 59764 11396 59768 11452
rect 59704 11392 59768 11396
rect 59784 11452 59848 11456
rect 59784 11396 59788 11452
rect 59788 11396 59844 11452
rect 59844 11396 59848 11452
rect 59784 11392 59848 11396
rect 82981 11452 83045 11456
rect 82981 11396 82985 11452
rect 82985 11396 83041 11452
rect 83041 11396 83045 11452
rect 82981 11392 83045 11396
rect 83061 11452 83125 11456
rect 83061 11396 83065 11452
rect 83065 11396 83121 11452
rect 83121 11396 83125 11452
rect 83061 11392 83125 11396
rect 83141 11452 83205 11456
rect 83141 11396 83145 11452
rect 83145 11396 83201 11452
rect 83201 11396 83205 11452
rect 83141 11392 83205 11396
rect 83221 11452 83285 11456
rect 83221 11396 83225 11452
rect 83225 11396 83281 11452
rect 83281 11396 83285 11452
rect 83221 11392 83285 11396
rect 59308 11052 59372 11116
rect 24388 10908 24452 10912
rect 24388 10852 24392 10908
rect 24392 10852 24448 10908
rect 24448 10852 24452 10908
rect 24388 10848 24452 10852
rect 24468 10908 24532 10912
rect 24468 10852 24472 10908
rect 24472 10852 24528 10908
rect 24528 10852 24532 10908
rect 24468 10848 24532 10852
rect 24548 10908 24612 10912
rect 24548 10852 24552 10908
rect 24552 10852 24608 10908
rect 24608 10852 24612 10908
rect 24548 10848 24612 10852
rect 24628 10908 24692 10912
rect 24628 10852 24632 10908
rect 24632 10852 24688 10908
rect 24688 10852 24692 10908
rect 24628 10848 24692 10852
rect 47825 10908 47889 10912
rect 47825 10852 47829 10908
rect 47829 10852 47885 10908
rect 47885 10852 47889 10908
rect 47825 10848 47889 10852
rect 47905 10908 47969 10912
rect 47905 10852 47909 10908
rect 47909 10852 47965 10908
rect 47965 10852 47969 10908
rect 47905 10848 47969 10852
rect 47985 10908 48049 10912
rect 47985 10852 47989 10908
rect 47989 10852 48045 10908
rect 48045 10852 48049 10908
rect 47985 10848 48049 10852
rect 48065 10908 48129 10912
rect 48065 10852 48069 10908
rect 48069 10852 48125 10908
rect 48125 10852 48129 10908
rect 48065 10848 48129 10852
rect 71262 10908 71326 10912
rect 71262 10852 71266 10908
rect 71266 10852 71322 10908
rect 71322 10852 71326 10908
rect 71262 10848 71326 10852
rect 71342 10908 71406 10912
rect 71342 10852 71346 10908
rect 71346 10852 71402 10908
rect 71402 10852 71406 10908
rect 71342 10848 71406 10852
rect 71422 10908 71486 10912
rect 71422 10852 71426 10908
rect 71426 10852 71482 10908
rect 71482 10852 71486 10908
rect 71422 10848 71486 10852
rect 71502 10908 71566 10912
rect 71502 10852 71506 10908
rect 71506 10852 71562 10908
rect 71562 10852 71566 10908
rect 71502 10848 71566 10852
rect 94699 10908 94763 10912
rect 94699 10852 94703 10908
rect 94703 10852 94759 10908
rect 94759 10852 94763 10908
rect 94699 10848 94763 10852
rect 94779 10908 94843 10912
rect 94779 10852 94783 10908
rect 94783 10852 94839 10908
rect 94839 10852 94843 10908
rect 94779 10848 94843 10852
rect 94859 10908 94923 10912
rect 94859 10852 94863 10908
rect 94863 10852 94919 10908
rect 94919 10852 94923 10908
rect 94859 10848 94923 10852
rect 94939 10908 95003 10912
rect 94939 10852 94943 10908
rect 94943 10852 94999 10908
rect 94999 10852 95003 10908
rect 94939 10848 95003 10852
rect 12670 10364 12734 10368
rect 12670 10308 12674 10364
rect 12674 10308 12730 10364
rect 12730 10308 12734 10364
rect 12670 10304 12734 10308
rect 12750 10364 12814 10368
rect 12750 10308 12754 10364
rect 12754 10308 12810 10364
rect 12810 10308 12814 10364
rect 12750 10304 12814 10308
rect 12830 10364 12894 10368
rect 12830 10308 12834 10364
rect 12834 10308 12890 10364
rect 12890 10308 12894 10364
rect 12830 10304 12894 10308
rect 12910 10364 12974 10368
rect 12910 10308 12914 10364
rect 12914 10308 12970 10364
rect 12970 10308 12974 10364
rect 12910 10304 12974 10308
rect 36107 10364 36171 10368
rect 36107 10308 36111 10364
rect 36111 10308 36167 10364
rect 36167 10308 36171 10364
rect 36107 10304 36171 10308
rect 36187 10364 36251 10368
rect 36187 10308 36191 10364
rect 36191 10308 36247 10364
rect 36247 10308 36251 10364
rect 36187 10304 36251 10308
rect 36267 10364 36331 10368
rect 36267 10308 36271 10364
rect 36271 10308 36327 10364
rect 36327 10308 36331 10364
rect 36267 10304 36331 10308
rect 36347 10364 36411 10368
rect 36347 10308 36351 10364
rect 36351 10308 36407 10364
rect 36407 10308 36411 10364
rect 36347 10304 36411 10308
rect 59544 10364 59608 10368
rect 59544 10308 59548 10364
rect 59548 10308 59604 10364
rect 59604 10308 59608 10364
rect 59544 10304 59608 10308
rect 59624 10364 59688 10368
rect 59624 10308 59628 10364
rect 59628 10308 59684 10364
rect 59684 10308 59688 10364
rect 59624 10304 59688 10308
rect 59704 10364 59768 10368
rect 59704 10308 59708 10364
rect 59708 10308 59764 10364
rect 59764 10308 59768 10364
rect 59704 10304 59768 10308
rect 59784 10364 59848 10368
rect 59784 10308 59788 10364
rect 59788 10308 59844 10364
rect 59844 10308 59848 10364
rect 59784 10304 59848 10308
rect 82981 10364 83045 10368
rect 82981 10308 82985 10364
rect 82985 10308 83041 10364
rect 83041 10308 83045 10364
rect 82981 10304 83045 10308
rect 83061 10364 83125 10368
rect 83061 10308 83065 10364
rect 83065 10308 83121 10364
rect 83121 10308 83125 10364
rect 83061 10304 83125 10308
rect 83141 10364 83205 10368
rect 83141 10308 83145 10364
rect 83145 10308 83201 10364
rect 83201 10308 83205 10364
rect 83141 10304 83205 10308
rect 83221 10364 83285 10368
rect 83221 10308 83225 10364
rect 83225 10308 83281 10364
rect 83281 10308 83285 10364
rect 83221 10304 83285 10308
rect 24388 9820 24452 9824
rect 24388 9764 24392 9820
rect 24392 9764 24448 9820
rect 24448 9764 24452 9820
rect 24388 9760 24452 9764
rect 24468 9820 24532 9824
rect 24468 9764 24472 9820
rect 24472 9764 24528 9820
rect 24528 9764 24532 9820
rect 24468 9760 24532 9764
rect 24548 9820 24612 9824
rect 24548 9764 24552 9820
rect 24552 9764 24608 9820
rect 24608 9764 24612 9820
rect 24548 9760 24612 9764
rect 24628 9820 24692 9824
rect 24628 9764 24632 9820
rect 24632 9764 24688 9820
rect 24688 9764 24692 9820
rect 24628 9760 24692 9764
rect 47825 9820 47889 9824
rect 47825 9764 47829 9820
rect 47829 9764 47885 9820
rect 47885 9764 47889 9820
rect 47825 9760 47889 9764
rect 47905 9820 47969 9824
rect 47905 9764 47909 9820
rect 47909 9764 47965 9820
rect 47965 9764 47969 9820
rect 47905 9760 47969 9764
rect 47985 9820 48049 9824
rect 47985 9764 47989 9820
rect 47989 9764 48045 9820
rect 48045 9764 48049 9820
rect 47985 9760 48049 9764
rect 48065 9820 48129 9824
rect 48065 9764 48069 9820
rect 48069 9764 48125 9820
rect 48125 9764 48129 9820
rect 48065 9760 48129 9764
rect 71262 9820 71326 9824
rect 71262 9764 71266 9820
rect 71266 9764 71322 9820
rect 71322 9764 71326 9820
rect 71262 9760 71326 9764
rect 71342 9820 71406 9824
rect 71342 9764 71346 9820
rect 71346 9764 71402 9820
rect 71402 9764 71406 9820
rect 71342 9760 71406 9764
rect 71422 9820 71486 9824
rect 71422 9764 71426 9820
rect 71426 9764 71482 9820
rect 71482 9764 71486 9820
rect 71422 9760 71486 9764
rect 71502 9820 71566 9824
rect 71502 9764 71506 9820
rect 71506 9764 71562 9820
rect 71562 9764 71566 9820
rect 71502 9760 71566 9764
rect 94699 9820 94763 9824
rect 94699 9764 94703 9820
rect 94703 9764 94759 9820
rect 94759 9764 94763 9820
rect 94699 9760 94763 9764
rect 94779 9820 94843 9824
rect 94779 9764 94783 9820
rect 94783 9764 94839 9820
rect 94839 9764 94843 9820
rect 94779 9760 94843 9764
rect 94859 9820 94923 9824
rect 94859 9764 94863 9820
rect 94863 9764 94919 9820
rect 94919 9764 94923 9820
rect 94859 9760 94923 9764
rect 94939 9820 95003 9824
rect 94939 9764 94943 9820
rect 94943 9764 94999 9820
rect 94999 9764 95003 9820
rect 94939 9760 95003 9764
rect 12670 9276 12734 9280
rect 12670 9220 12674 9276
rect 12674 9220 12730 9276
rect 12730 9220 12734 9276
rect 12670 9216 12734 9220
rect 12750 9276 12814 9280
rect 12750 9220 12754 9276
rect 12754 9220 12810 9276
rect 12810 9220 12814 9276
rect 12750 9216 12814 9220
rect 12830 9276 12894 9280
rect 12830 9220 12834 9276
rect 12834 9220 12890 9276
rect 12890 9220 12894 9276
rect 12830 9216 12894 9220
rect 12910 9276 12974 9280
rect 12910 9220 12914 9276
rect 12914 9220 12970 9276
rect 12970 9220 12974 9276
rect 12910 9216 12974 9220
rect 36107 9276 36171 9280
rect 36107 9220 36111 9276
rect 36111 9220 36167 9276
rect 36167 9220 36171 9276
rect 36107 9216 36171 9220
rect 36187 9276 36251 9280
rect 36187 9220 36191 9276
rect 36191 9220 36247 9276
rect 36247 9220 36251 9276
rect 36187 9216 36251 9220
rect 36267 9276 36331 9280
rect 36267 9220 36271 9276
rect 36271 9220 36327 9276
rect 36327 9220 36331 9276
rect 36267 9216 36331 9220
rect 36347 9276 36411 9280
rect 36347 9220 36351 9276
rect 36351 9220 36407 9276
rect 36407 9220 36411 9276
rect 36347 9216 36411 9220
rect 59544 9276 59608 9280
rect 59544 9220 59548 9276
rect 59548 9220 59604 9276
rect 59604 9220 59608 9276
rect 59544 9216 59608 9220
rect 59624 9276 59688 9280
rect 59624 9220 59628 9276
rect 59628 9220 59684 9276
rect 59684 9220 59688 9276
rect 59624 9216 59688 9220
rect 59704 9276 59768 9280
rect 59704 9220 59708 9276
rect 59708 9220 59764 9276
rect 59764 9220 59768 9276
rect 59704 9216 59768 9220
rect 59784 9276 59848 9280
rect 59784 9220 59788 9276
rect 59788 9220 59844 9276
rect 59844 9220 59848 9276
rect 59784 9216 59848 9220
rect 82981 9276 83045 9280
rect 82981 9220 82985 9276
rect 82985 9220 83041 9276
rect 83041 9220 83045 9276
rect 82981 9216 83045 9220
rect 83061 9276 83125 9280
rect 83061 9220 83065 9276
rect 83065 9220 83121 9276
rect 83121 9220 83125 9276
rect 83061 9216 83125 9220
rect 83141 9276 83205 9280
rect 83141 9220 83145 9276
rect 83145 9220 83201 9276
rect 83201 9220 83205 9276
rect 83141 9216 83205 9220
rect 83221 9276 83285 9280
rect 83221 9220 83225 9276
rect 83225 9220 83281 9276
rect 83281 9220 83285 9276
rect 83221 9216 83285 9220
rect 59308 8740 59372 8804
rect 24388 8732 24452 8736
rect 24388 8676 24392 8732
rect 24392 8676 24448 8732
rect 24448 8676 24452 8732
rect 24388 8672 24452 8676
rect 24468 8732 24532 8736
rect 24468 8676 24472 8732
rect 24472 8676 24528 8732
rect 24528 8676 24532 8732
rect 24468 8672 24532 8676
rect 24548 8732 24612 8736
rect 24548 8676 24552 8732
rect 24552 8676 24608 8732
rect 24608 8676 24612 8732
rect 24548 8672 24612 8676
rect 24628 8732 24692 8736
rect 24628 8676 24632 8732
rect 24632 8676 24688 8732
rect 24688 8676 24692 8732
rect 24628 8672 24692 8676
rect 47825 8732 47889 8736
rect 47825 8676 47829 8732
rect 47829 8676 47885 8732
rect 47885 8676 47889 8732
rect 47825 8672 47889 8676
rect 47905 8732 47969 8736
rect 47905 8676 47909 8732
rect 47909 8676 47965 8732
rect 47965 8676 47969 8732
rect 47905 8672 47969 8676
rect 47985 8732 48049 8736
rect 47985 8676 47989 8732
rect 47989 8676 48045 8732
rect 48045 8676 48049 8732
rect 47985 8672 48049 8676
rect 48065 8732 48129 8736
rect 48065 8676 48069 8732
rect 48069 8676 48125 8732
rect 48125 8676 48129 8732
rect 48065 8672 48129 8676
rect 71262 8732 71326 8736
rect 71262 8676 71266 8732
rect 71266 8676 71322 8732
rect 71322 8676 71326 8732
rect 71262 8672 71326 8676
rect 71342 8732 71406 8736
rect 71342 8676 71346 8732
rect 71346 8676 71402 8732
rect 71402 8676 71406 8732
rect 71342 8672 71406 8676
rect 71422 8732 71486 8736
rect 71422 8676 71426 8732
rect 71426 8676 71482 8732
rect 71482 8676 71486 8732
rect 71422 8672 71486 8676
rect 71502 8732 71566 8736
rect 71502 8676 71506 8732
rect 71506 8676 71562 8732
rect 71562 8676 71566 8732
rect 71502 8672 71566 8676
rect 94699 8732 94763 8736
rect 94699 8676 94703 8732
rect 94703 8676 94759 8732
rect 94759 8676 94763 8732
rect 94699 8672 94763 8676
rect 94779 8732 94843 8736
rect 94779 8676 94783 8732
rect 94783 8676 94839 8732
rect 94839 8676 94843 8732
rect 94779 8672 94843 8676
rect 94859 8732 94923 8736
rect 94859 8676 94863 8732
rect 94863 8676 94919 8732
rect 94919 8676 94923 8732
rect 94859 8672 94923 8676
rect 94939 8732 95003 8736
rect 94939 8676 94943 8732
rect 94943 8676 94999 8732
rect 94999 8676 95003 8732
rect 94939 8672 95003 8676
rect 63540 8468 63604 8532
rect 12670 8188 12734 8192
rect 12670 8132 12674 8188
rect 12674 8132 12730 8188
rect 12730 8132 12734 8188
rect 12670 8128 12734 8132
rect 12750 8188 12814 8192
rect 12750 8132 12754 8188
rect 12754 8132 12810 8188
rect 12810 8132 12814 8188
rect 12750 8128 12814 8132
rect 12830 8188 12894 8192
rect 12830 8132 12834 8188
rect 12834 8132 12890 8188
rect 12890 8132 12894 8188
rect 12830 8128 12894 8132
rect 12910 8188 12974 8192
rect 12910 8132 12914 8188
rect 12914 8132 12970 8188
rect 12970 8132 12974 8188
rect 12910 8128 12974 8132
rect 36107 8188 36171 8192
rect 36107 8132 36111 8188
rect 36111 8132 36167 8188
rect 36167 8132 36171 8188
rect 36107 8128 36171 8132
rect 36187 8188 36251 8192
rect 36187 8132 36191 8188
rect 36191 8132 36247 8188
rect 36247 8132 36251 8188
rect 36187 8128 36251 8132
rect 36267 8188 36331 8192
rect 36267 8132 36271 8188
rect 36271 8132 36327 8188
rect 36327 8132 36331 8188
rect 36267 8128 36331 8132
rect 36347 8188 36411 8192
rect 36347 8132 36351 8188
rect 36351 8132 36407 8188
rect 36407 8132 36411 8188
rect 36347 8128 36411 8132
rect 59544 8188 59608 8192
rect 59544 8132 59548 8188
rect 59548 8132 59604 8188
rect 59604 8132 59608 8188
rect 59544 8128 59608 8132
rect 59624 8188 59688 8192
rect 59624 8132 59628 8188
rect 59628 8132 59684 8188
rect 59684 8132 59688 8188
rect 59624 8128 59688 8132
rect 59704 8188 59768 8192
rect 59704 8132 59708 8188
rect 59708 8132 59764 8188
rect 59764 8132 59768 8188
rect 59704 8128 59768 8132
rect 59784 8188 59848 8192
rect 59784 8132 59788 8188
rect 59788 8132 59844 8188
rect 59844 8132 59848 8188
rect 59784 8128 59848 8132
rect 82981 8188 83045 8192
rect 82981 8132 82985 8188
rect 82985 8132 83041 8188
rect 83041 8132 83045 8188
rect 82981 8128 83045 8132
rect 83061 8188 83125 8192
rect 83061 8132 83065 8188
rect 83065 8132 83121 8188
rect 83121 8132 83125 8188
rect 83061 8128 83125 8132
rect 83141 8188 83205 8192
rect 83141 8132 83145 8188
rect 83145 8132 83201 8188
rect 83201 8132 83205 8188
rect 83141 8128 83205 8132
rect 83221 8188 83285 8192
rect 83221 8132 83225 8188
rect 83225 8132 83281 8188
rect 83281 8132 83285 8188
rect 83221 8128 83285 8132
rect 24388 7644 24452 7648
rect 24388 7588 24392 7644
rect 24392 7588 24448 7644
rect 24448 7588 24452 7644
rect 24388 7584 24452 7588
rect 24468 7644 24532 7648
rect 24468 7588 24472 7644
rect 24472 7588 24528 7644
rect 24528 7588 24532 7644
rect 24468 7584 24532 7588
rect 24548 7644 24612 7648
rect 24548 7588 24552 7644
rect 24552 7588 24608 7644
rect 24608 7588 24612 7644
rect 24548 7584 24612 7588
rect 24628 7644 24692 7648
rect 24628 7588 24632 7644
rect 24632 7588 24688 7644
rect 24688 7588 24692 7644
rect 24628 7584 24692 7588
rect 47825 7644 47889 7648
rect 47825 7588 47829 7644
rect 47829 7588 47885 7644
rect 47885 7588 47889 7644
rect 47825 7584 47889 7588
rect 47905 7644 47969 7648
rect 47905 7588 47909 7644
rect 47909 7588 47965 7644
rect 47965 7588 47969 7644
rect 47905 7584 47969 7588
rect 47985 7644 48049 7648
rect 47985 7588 47989 7644
rect 47989 7588 48045 7644
rect 48045 7588 48049 7644
rect 47985 7584 48049 7588
rect 48065 7644 48129 7648
rect 48065 7588 48069 7644
rect 48069 7588 48125 7644
rect 48125 7588 48129 7644
rect 48065 7584 48129 7588
rect 71262 7644 71326 7648
rect 71262 7588 71266 7644
rect 71266 7588 71322 7644
rect 71322 7588 71326 7644
rect 71262 7584 71326 7588
rect 71342 7644 71406 7648
rect 71342 7588 71346 7644
rect 71346 7588 71402 7644
rect 71402 7588 71406 7644
rect 71342 7584 71406 7588
rect 71422 7644 71486 7648
rect 71422 7588 71426 7644
rect 71426 7588 71482 7644
rect 71482 7588 71486 7644
rect 71422 7584 71486 7588
rect 71502 7644 71566 7648
rect 71502 7588 71506 7644
rect 71506 7588 71562 7644
rect 71562 7588 71566 7644
rect 71502 7584 71566 7588
rect 94699 7644 94763 7648
rect 94699 7588 94703 7644
rect 94703 7588 94759 7644
rect 94759 7588 94763 7644
rect 94699 7584 94763 7588
rect 94779 7644 94843 7648
rect 94779 7588 94783 7644
rect 94783 7588 94839 7644
rect 94839 7588 94843 7644
rect 94779 7584 94843 7588
rect 94859 7644 94923 7648
rect 94859 7588 94863 7644
rect 94863 7588 94919 7644
rect 94919 7588 94923 7644
rect 94859 7584 94923 7588
rect 94939 7644 95003 7648
rect 94939 7588 94943 7644
rect 94943 7588 94999 7644
rect 94999 7588 95003 7644
rect 94939 7584 95003 7588
rect 12670 7100 12734 7104
rect 12670 7044 12674 7100
rect 12674 7044 12730 7100
rect 12730 7044 12734 7100
rect 12670 7040 12734 7044
rect 12750 7100 12814 7104
rect 12750 7044 12754 7100
rect 12754 7044 12810 7100
rect 12810 7044 12814 7100
rect 12750 7040 12814 7044
rect 12830 7100 12894 7104
rect 12830 7044 12834 7100
rect 12834 7044 12890 7100
rect 12890 7044 12894 7100
rect 12830 7040 12894 7044
rect 12910 7100 12974 7104
rect 12910 7044 12914 7100
rect 12914 7044 12970 7100
rect 12970 7044 12974 7100
rect 12910 7040 12974 7044
rect 36107 7100 36171 7104
rect 36107 7044 36111 7100
rect 36111 7044 36167 7100
rect 36167 7044 36171 7100
rect 36107 7040 36171 7044
rect 36187 7100 36251 7104
rect 36187 7044 36191 7100
rect 36191 7044 36247 7100
rect 36247 7044 36251 7100
rect 36187 7040 36251 7044
rect 36267 7100 36331 7104
rect 36267 7044 36271 7100
rect 36271 7044 36327 7100
rect 36327 7044 36331 7100
rect 36267 7040 36331 7044
rect 36347 7100 36411 7104
rect 36347 7044 36351 7100
rect 36351 7044 36407 7100
rect 36407 7044 36411 7100
rect 36347 7040 36411 7044
rect 59544 7100 59608 7104
rect 59544 7044 59548 7100
rect 59548 7044 59604 7100
rect 59604 7044 59608 7100
rect 59544 7040 59608 7044
rect 59624 7100 59688 7104
rect 59624 7044 59628 7100
rect 59628 7044 59684 7100
rect 59684 7044 59688 7100
rect 59624 7040 59688 7044
rect 59704 7100 59768 7104
rect 59704 7044 59708 7100
rect 59708 7044 59764 7100
rect 59764 7044 59768 7100
rect 59704 7040 59768 7044
rect 59784 7100 59848 7104
rect 59784 7044 59788 7100
rect 59788 7044 59844 7100
rect 59844 7044 59848 7100
rect 59784 7040 59848 7044
rect 82981 7100 83045 7104
rect 82981 7044 82985 7100
rect 82985 7044 83041 7100
rect 83041 7044 83045 7100
rect 82981 7040 83045 7044
rect 83061 7100 83125 7104
rect 83061 7044 83065 7100
rect 83065 7044 83121 7100
rect 83121 7044 83125 7100
rect 83061 7040 83125 7044
rect 83141 7100 83205 7104
rect 83141 7044 83145 7100
rect 83145 7044 83201 7100
rect 83201 7044 83205 7100
rect 83141 7040 83205 7044
rect 83221 7100 83285 7104
rect 83221 7044 83225 7100
rect 83225 7044 83281 7100
rect 83281 7044 83285 7100
rect 83221 7040 83285 7044
rect 24388 6556 24452 6560
rect 24388 6500 24392 6556
rect 24392 6500 24448 6556
rect 24448 6500 24452 6556
rect 24388 6496 24452 6500
rect 24468 6556 24532 6560
rect 24468 6500 24472 6556
rect 24472 6500 24528 6556
rect 24528 6500 24532 6556
rect 24468 6496 24532 6500
rect 24548 6556 24612 6560
rect 24548 6500 24552 6556
rect 24552 6500 24608 6556
rect 24608 6500 24612 6556
rect 24548 6496 24612 6500
rect 24628 6556 24692 6560
rect 24628 6500 24632 6556
rect 24632 6500 24688 6556
rect 24688 6500 24692 6556
rect 24628 6496 24692 6500
rect 47825 6556 47889 6560
rect 47825 6500 47829 6556
rect 47829 6500 47885 6556
rect 47885 6500 47889 6556
rect 47825 6496 47889 6500
rect 47905 6556 47969 6560
rect 47905 6500 47909 6556
rect 47909 6500 47965 6556
rect 47965 6500 47969 6556
rect 47905 6496 47969 6500
rect 47985 6556 48049 6560
rect 47985 6500 47989 6556
rect 47989 6500 48045 6556
rect 48045 6500 48049 6556
rect 47985 6496 48049 6500
rect 48065 6556 48129 6560
rect 48065 6500 48069 6556
rect 48069 6500 48125 6556
rect 48125 6500 48129 6556
rect 48065 6496 48129 6500
rect 71262 6556 71326 6560
rect 71262 6500 71266 6556
rect 71266 6500 71322 6556
rect 71322 6500 71326 6556
rect 71262 6496 71326 6500
rect 71342 6556 71406 6560
rect 71342 6500 71346 6556
rect 71346 6500 71402 6556
rect 71402 6500 71406 6556
rect 71342 6496 71406 6500
rect 71422 6556 71486 6560
rect 71422 6500 71426 6556
rect 71426 6500 71482 6556
rect 71482 6500 71486 6556
rect 71422 6496 71486 6500
rect 71502 6556 71566 6560
rect 71502 6500 71506 6556
rect 71506 6500 71562 6556
rect 71562 6500 71566 6556
rect 71502 6496 71566 6500
rect 94699 6556 94763 6560
rect 94699 6500 94703 6556
rect 94703 6500 94759 6556
rect 94759 6500 94763 6556
rect 94699 6496 94763 6500
rect 94779 6556 94843 6560
rect 94779 6500 94783 6556
rect 94783 6500 94839 6556
rect 94839 6500 94843 6556
rect 94779 6496 94843 6500
rect 94859 6556 94923 6560
rect 94859 6500 94863 6556
rect 94863 6500 94919 6556
rect 94919 6500 94923 6556
rect 94859 6496 94923 6500
rect 94939 6556 95003 6560
rect 94939 6500 94943 6556
rect 94943 6500 94999 6556
rect 94999 6500 95003 6556
rect 94939 6496 95003 6500
rect 12670 6012 12734 6016
rect 12670 5956 12674 6012
rect 12674 5956 12730 6012
rect 12730 5956 12734 6012
rect 12670 5952 12734 5956
rect 12750 6012 12814 6016
rect 12750 5956 12754 6012
rect 12754 5956 12810 6012
rect 12810 5956 12814 6012
rect 12750 5952 12814 5956
rect 12830 6012 12894 6016
rect 12830 5956 12834 6012
rect 12834 5956 12890 6012
rect 12890 5956 12894 6012
rect 12830 5952 12894 5956
rect 12910 6012 12974 6016
rect 12910 5956 12914 6012
rect 12914 5956 12970 6012
rect 12970 5956 12974 6012
rect 12910 5952 12974 5956
rect 36107 6012 36171 6016
rect 36107 5956 36111 6012
rect 36111 5956 36167 6012
rect 36167 5956 36171 6012
rect 36107 5952 36171 5956
rect 36187 6012 36251 6016
rect 36187 5956 36191 6012
rect 36191 5956 36247 6012
rect 36247 5956 36251 6012
rect 36187 5952 36251 5956
rect 36267 6012 36331 6016
rect 36267 5956 36271 6012
rect 36271 5956 36327 6012
rect 36327 5956 36331 6012
rect 36267 5952 36331 5956
rect 36347 6012 36411 6016
rect 36347 5956 36351 6012
rect 36351 5956 36407 6012
rect 36407 5956 36411 6012
rect 36347 5952 36411 5956
rect 59544 6012 59608 6016
rect 59544 5956 59548 6012
rect 59548 5956 59604 6012
rect 59604 5956 59608 6012
rect 59544 5952 59608 5956
rect 59624 6012 59688 6016
rect 59624 5956 59628 6012
rect 59628 5956 59684 6012
rect 59684 5956 59688 6012
rect 59624 5952 59688 5956
rect 59704 6012 59768 6016
rect 59704 5956 59708 6012
rect 59708 5956 59764 6012
rect 59764 5956 59768 6012
rect 59704 5952 59768 5956
rect 59784 6012 59848 6016
rect 59784 5956 59788 6012
rect 59788 5956 59844 6012
rect 59844 5956 59848 6012
rect 59784 5952 59848 5956
rect 82981 6012 83045 6016
rect 82981 5956 82985 6012
rect 82985 5956 83041 6012
rect 83041 5956 83045 6012
rect 82981 5952 83045 5956
rect 83061 6012 83125 6016
rect 83061 5956 83065 6012
rect 83065 5956 83121 6012
rect 83121 5956 83125 6012
rect 83061 5952 83125 5956
rect 83141 6012 83205 6016
rect 83141 5956 83145 6012
rect 83145 5956 83201 6012
rect 83201 5956 83205 6012
rect 83141 5952 83205 5956
rect 83221 6012 83285 6016
rect 83221 5956 83225 6012
rect 83225 5956 83281 6012
rect 83281 5956 83285 6012
rect 83221 5952 83285 5956
rect 24388 5468 24452 5472
rect 24388 5412 24392 5468
rect 24392 5412 24448 5468
rect 24448 5412 24452 5468
rect 24388 5408 24452 5412
rect 24468 5468 24532 5472
rect 24468 5412 24472 5468
rect 24472 5412 24528 5468
rect 24528 5412 24532 5468
rect 24468 5408 24532 5412
rect 24548 5468 24612 5472
rect 24548 5412 24552 5468
rect 24552 5412 24608 5468
rect 24608 5412 24612 5468
rect 24548 5408 24612 5412
rect 24628 5468 24692 5472
rect 24628 5412 24632 5468
rect 24632 5412 24688 5468
rect 24688 5412 24692 5468
rect 24628 5408 24692 5412
rect 47825 5468 47889 5472
rect 47825 5412 47829 5468
rect 47829 5412 47885 5468
rect 47885 5412 47889 5468
rect 47825 5408 47889 5412
rect 47905 5468 47969 5472
rect 47905 5412 47909 5468
rect 47909 5412 47965 5468
rect 47965 5412 47969 5468
rect 47905 5408 47969 5412
rect 47985 5468 48049 5472
rect 47985 5412 47989 5468
rect 47989 5412 48045 5468
rect 48045 5412 48049 5468
rect 47985 5408 48049 5412
rect 48065 5468 48129 5472
rect 48065 5412 48069 5468
rect 48069 5412 48125 5468
rect 48125 5412 48129 5468
rect 48065 5408 48129 5412
rect 71262 5468 71326 5472
rect 71262 5412 71266 5468
rect 71266 5412 71322 5468
rect 71322 5412 71326 5468
rect 71262 5408 71326 5412
rect 71342 5468 71406 5472
rect 71342 5412 71346 5468
rect 71346 5412 71402 5468
rect 71402 5412 71406 5468
rect 71342 5408 71406 5412
rect 71422 5468 71486 5472
rect 71422 5412 71426 5468
rect 71426 5412 71482 5468
rect 71482 5412 71486 5468
rect 71422 5408 71486 5412
rect 71502 5468 71566 5472
rect 71502 5412 71506 5468
rect 71506 5412 71562 5468
rect 71562 5412 71566 5468
rect 71502 5408 71566 5412
rect 94699 5468 94763 5472
rect 94699 5412 94703 5468
rect 94703 5412 94759 5468
rect 94759 5412 94763 5468
rect 94699 5408 94763 5412
rect 94779 5468 94843 5472
rect 94779 5412 94783 5468
rect 94783 5412 94839 5468
rect 94839 5412 94843 5468
rect 94779 5408 94843 5412
rect 94859 5468 94923 5472
rect 94859 5412 94863 5468
rect 94863 5412 94919 5468
rect 94919 5412 94923 5468
rect 94859 5408 94923 5412
rect 94939 5468 95003 5472
rect 94939 5412 94943 5468
rect 94943 5412 94999 5468
rect 94999 5412 95003 5468
rect 94939 5408 95003 5412
rect 12670 4924 12734 4928
rect 12670 4868 12674 4924
rect 12674 4868 12730 4924
rect 12730 4868 12734 4924
rect 12670 4864 12734 4868
rect 12750 4924 12814 4928
rect 12750 4868 12754 4924
rect 12754 4868 12810 4924
rect 12810 4868 12814 4924
rect 12750 4864 12814 4868
rect 12830 4924 12894 4928
rect 12830 4868 12834 4924
rect 12834 4868 12890 4924
rect 12890 4868 12894 4924
rect 12830 4864 12894 4868
rect 12910 4924 12974 4928
rect 12910 4868 12914 4924
rect 12914 4868 12970 4924
rect 12970 4868 12974 4924
rect 12910 4864 12974 4868
rect 36107 4924 36171 4928
rect 36107 4868 36111 4924
rect 36111 4868 36167 4924
rect 36167 4868 36171 4924
rect 36107 4864 36171 4868
rect 36187 4924 36251 4928
rect 36187 4868 36191 4924
rect 36191 4868 36247 4924
rect 36247 4868 36251 4924
rect 36187 4864 36251 4868
rect 36267 4924 36331 4928
rect 36267 4868 36271 4924
rect 36271 4868 36327 4924
rect 36327 4868 36331 4924
rect 36267 4864 36331 4868
rect 36347 4924 36411 4928
rect 36347 4868 36351 4924
rect 36351 4868 36407 4924
rect 36407 4868 36411 4924
rect 36347 4864 36411 4868
rect 59544 4924 59608 4928
rect 59544 4868 59548 4924
rect 59548 4868 59604 4924
rect 59604 4868 59608 4924
rect 59544 4864 59608 4868
rect 59624 4924 59688 4928
rect 59624 4868 59628 4924
rect 59628 4868 59684 4924
rect 59684 4868 59688 4924
rect 59624 4864 59688 4868
rect 59704 4924 59768 4928
rect 59704 4868 59708 4924
rect 59708 4868 59764 4924
rect 59764 4868 59768 4924
rect 59704 4864 59768 4868
rect 59784 4924 59848 4928
rect 59784 4868 59788 4924
rect 59788 4868 59844 4924
rect 59844 4868 59848 4924
rect 59784 4864 59848 4868
rect 82981 4924 83045 4928
rect 82981 4868 82985 4924
rect 82985 4868 83041 4924
rect 83041 4868 83045 4924
rect 82981 4864 83045 4868
rect 83061 4924 83125 4928
rect 83061 4868 83065 4924
rect 83065 4868 83121 4924
rect 83121 4868 83125 4924
rect 83061 4864 83125 4868
rect 83141 4924 83205 4928
rect 83141 4868 83145 4924
rect 83145 4868 83201 4924
rect 83201 4868 83205 4924
rect 83141 4864 83205 4868
rect 83221 4924 83285 4928
rect 83221 4868 83225 4924
rect 83225 4868 83281 4924
rect 83281 4868 83285 4924
rect 83221 4864 83285 4868
rect 63540 4856 63604 4860
rect 63540 4800 63590 4856
rect 63590 4800 63604 4856
rect 63540 4796 63604 4800
rect 24388 4380 24452 4384
rect 24388 4324 24392 4380
rect 24392 4324 24448 4380
rect 24448 4324 24452 4380
rect 24388 4320 24452 4324
rect 24468 4380 24532 4384
rect 24468 4324 24472 4380
rect 24472 4324 24528 4380
rect 24528 4324 24532 4380
rect 24468 4320 24532 4324
rect 24548 4380 24612 4384
rect 24548 4324 24552 4380
rect 24552 4324 24608 4380
rect 24608 4324 24612 4380
rect 24548 4320 24612 4324
rect 24628 4380 24692 4384
rect 24628 4324 24632 4380
rect 24632 4324 24688 4380
rect 24688 4324 24692 4380
rect 24628 4320 24692 4324
rect 47825 4380 47889 4384
rect 47825 4324 47829 4380
rect 47829 4324 47885 4380
rect 47885 4324 47889 4380
rect 47825 4320 47889 4324
rect 47905 4380 47969 4384
rect 47905 4324 47909 4380
rect 47909 4324 47965 4380
rect 47965 4324 47969 4380
rect 47905 4320 47969 4324
rect 47985 4380 48049 4384
rect 47985 4324 47989 4380
rect 47989 4324 48045 4380
rect 48045 4324 48049 4380
rect 47985 4320 48049 4324
rect 48065 4380 48129 4384
rect 48065 4324 48069 4380
rect 48069 4324 48125 4380
rect 48125 4324 48129 4380
rect 48065 4320 48129 4324
rect 71262 4380 71326 4384
rect 71262 4324 71266 4380
rect 71266 4324 71322 4380
rect 71322 4324 71326 4380
rect 71262 4320 71326 4324
rect 71342 4380 71406 4384
rect 71342 4324 71346 4380
rect 71346 4324 71402 4380
rect 71402 4324 71406 4380
rect 71342 4320 71406 4324
rect 71422 4380 71486 4384
rect 71422 4324 71426 4380
rect 71426 4324 71482 4380
rect 71482 4324 71486 4380
rect 71422 4320 71486 4324
rect 71502 4380 71566 4384
rect 71502 4324 71506 4380
rect 71506 4324 71562 4380
rect 71562 4324 71566 4380
rect 71502 4320 71566 4324
rect 94699 4380 94763 4384
rect 94699 4324 94703 4380
rect 94703 4324 94759 4380
rect 94759 4324 94763 4380
rect 94699 4320 94763 4324
rect 94779 4380 94843 4384
rect 94779 4324 94783 4380
rect 94783 4324 94839 4380
rect 94839 4324 94843 4380
rect 94779 4320 94843 4324
rect 94859 4380 94923 4384
rect 94859 4324 94863 4380
rect 94863 4324 94919 4380
rect 94919 4324 94923 4380
rect 94859 4320 94923 4324
rect 94939 4380 95003 4384
rect 94939 4324 94943 4380
rect 94943 4324 94999 4380
rect 94999 4324 95003 4380
rect 94939 4320 95003 4324
rect 12670 3836 12734 3840
rect 12670 3780 12674 3836
rect 12674 3780 12730 3836
rect 12730 3780 12734 3836
rect 12670 3776 12734 3780
rect 12750 3836 12814 3840
rect 12750 3780 12754 3836
rect 12754 3780 12810 3836
rect 12810 3780 12814 3836
rect 12750 3776 12814 3780
rect 12830 3836 12894 3840
rect 12830 3780 12834 3836
rect 12834 3780 12890 3836
rect 12890 3780 12894 3836
rect 12830 3776 12894 3780
rect 12910 3836 12974 3840
rect 12910 3780 12914 3836
rect 12914 3780 12970 3836
rect 12970 3780 12974 3836
rect 12910 3776 12974 3780
rect 36107 3836 36171 3840
rect 36107 3780 36111 3836
rect 36111 3780 36167 3836
rect 36167 3780 36171 3836
rect 36107 3776 36171 3780
rect 36187 3836 36251 3840
rect 36187 3780 36191 3836
rect 36191 3780 36247 3836
rect 36247 3780 36251 3836
rect 36187 3776 36251 3780
rect 36267 3836 36331 3840
rect 36267 3780 36271 3836
rect 36271 3780 36327 3836
rect 36327 3780 36331 3836
rect 36267 3776 36331 3780
rect 36347 3836 36411 3840
rect 36347 3780 36351 3836
rect 36351 3780 36407 3836
rect 36407 3780 36411 3836
rect 36347 3776 36411 3780
rect 59544 3836 59608 3840
rect 59544 3780 59548 3836
rect 59548 3780 59604 3836
rect 59604 3780 59608 3836
rect 59544 3776 59608 3780
rect 59624 3836 59688 3840
rect 59624 3780 59628 3836
rect 59628 3780 59684 3836
rect 59684 3780 59688 3836
rect 59624 3776 59688 3780
rect 59704 3836 59768 3840
rect 59704 3780 59708 3836
rect 59708 3780 59764 3836
rect 59764 3780 59768 3836
rect 59704 3776 59768 3780
rect 59784 3836 59848 3840
rect 59784 3780 59788 3836
rect 59788 3780 59844 3836
rect 59844 3780 59848 3836
rect 59784 3776 59848 3780
rect 82981 3836 83045 3840
rect 82981 3780 82985 3836
rect 82985 3780 83041 3836
rect 83041 3780 83045 3836
rect 82981 3776 83045 3780
rect 83061 3836 83125 3840
rect 83061 3780 83065 3836
rect 83065 3780 83121 3836
rect 83121 3780 83125 3836
rect 83061 3776 83125 3780
rect 83141 3836 83205 3840
rect 83141 3780 83145 3836
rect 83145 3780 83201 3836
rect 83201 3780 83205 3836
rect 83141 3776 83205 3780
rect 83221 3836 83285 3840
rect 83221 3780 83225 3836
rect 83225 3780 83281 3836
rect 83281 3780 83285 3836
rect 83221 3776 83285 3780
rect 24388 3292 24452 3296
rect 24388 3236 24392 3292
rect 24392 3236 24448 3292
rect 24448 3236 24452 3292
rect 24388 3232 24452 3236
rect 24468 3292 24532 3296
rect 24468 3236 24472 3292
rect 24472 3236 24528 3292
rect 24528 3236 24532 3292
rect 24468 3232 24532 3236
rect 24548 3292 24612 3296
rect 24548 3236 24552 3292
rect 24552 3236 24608 3292
rect 24608 3236 24612 3292
rect 24548 3232 24612 3236
rect 24628 3292 24692 3296
rect 24628 3236 24632 3292
rect 24632 3236 24688 3292
rect 24688 3236 24692 3292
rect 24628 3232 24692 3236
rect 47825 3292 47889 3296
rect 47825 3236 47829 3292
rect 47829 3236 47885 3292
rect 47885 3236 47889 3292
rect 47825 3232 47889 3236
rect 47905 3292 47969 3296
rect 47905 3236 47909 3292
rect 47909 3236 47965 3292
rect 47965 3236 47969 3292
rect 47905 3232 47969 3236
rect 47985 3292 48049 3296
rect 47985 3236 47989 3292
rect 47989 3236 48045 3292
rect 48045 3236 48049 3292
rect 47985 3232 48049 3236
rect 48065 3292 48129 3296
rect 48065 3236 48069 3292
rect 48069 3236 48125 3292
rect 48125 3236 48129 3292
rect 48065 3232 48129 3236
rect 71262 3292 71326 3296
rect 71262 3236 71266 3292
rect 71266 3236 71322 3292
rect 71322 3236 71326 3292
rect 71262 3232 71326 3236
rect 71342 3292 71406 3296
rect 71342 3236 71346 3292
rect 71346 3236 71402 3292
rect 71402 3236 71406 3292
rect 71342 3232 71406 3236
rect 71422 3292 71486 3296
rect 71422 3236 71426 3292
rect 71426 3236 71482 3292
rect 71482 3236 71486 3292
rect 71422 3232 71486 3236
rect 71502 3292 71566 3296
rect 71502 3236 71506 3292
rect 71506 3236 71562 3292
rect 71562 3236 71566 3292
rect 71502 3232 71566 3236
rect 94699 3292 94763 3296
rect 94699 3236 94703 3292
rect 94703 3236 94759 3292
rect 94759 3236 94763 3292
rect 94699 3232 94763 3236
rect 94779 3292 94843 3296
rect 94779 3236 94783 3292
rect 94783 3236 94839 3292
rect 94839 3236 94843 3292
rect 94779 3232 94843 3236
rect 94859 3292 94923 3296
rect 94859 3236 94863 3292
rect 94863 3236 94919 3292
rect 94919 3236 94923 3292
rect 94859 3232 94923 3236
rect 94939 3292 95003 3296
rect 94939 3236 94943 3292
rect 94943 3236 94999 3292
rect 94999 3236 95003 3292
rect 94939 3232 95003 3236
rect 12670 2748 12734 2752
rect 12670 2692 12674 2748
rect 12674 2692 12730 2748
rect 12730 2692 12734 2748
rect 12670 2688 12734 2692
rect 12750 2748 12814 2752
rect 12750 2692 12754 2748
rect 12754 2692 12810 2748
rect 12810 2692 12814 2748
rect 12750 2688 12814 2692
rect 12830 2748 12894 2752
rect 12830 2692 12834 2748
rect 12834 2692 12890 2748
rect 12890 2692 12894 2748
rect 12830 2688 12894 2692
rect 12910 2748 12974 2752
rect 12910 2692 12914 2748
rect 12914 2692 12970 2748
rect 12970 2692 12974 2748
rect 12910 2688 12974 2692
rect 36107 2748 36171 2752
rect 36107 2692 36111 2748
rect 36111 2692 36167 2748
rect 36167 2692 36171 2748
rect 36107 2688 36171 2692
rect 36187 2748 36251 2752
rect 36187 2692 36191 2748
rect 36191 2692 36247 2748
rect 36247 2692 36251 2748
rect 36187 2688 36251 2692
rect 36267 2748 36331 2752
rect 36267 2692 36271 2748
rect 36271 2692 36327 2748
rect 36327 2692 36331 2748
rect 36267 2688 36331 2692
rect 36347 2748 36411 2752
rect 36347 2692 36351 2748
rect 36351 2692 36407 2748
rect 36407 2692 36411 2748
rect 36347 2688 36411 2692
rect 59544 2748 59608 2752
rect 59544 2692 59548 2748
rect 59548 2692 59604 2748
rect 59604 2692 59608 2748
rect 59544 2688 59608 2692
rect 59624 2748 59688 2752
rect 59624 2692 59628 2748
rect 59628 2692 59684 2748
rect 59684 2692 59688 2748
rect 59624 2688 59688 2692
rect 59704 2748 59768 2752
rect 59704 2692 59708 2748
rect 59708 2692 59764 2748
rect 59764 2692 59768 2748
rect 59704 2688 59768 2692
rect 59784 2748 59848 2752
rect 59784 2692 59788 2748
rect 59788 2692 59844 2748
rect 59844 2692 59848 2748
rect 59784 2688 59848 2692
rect 82981 2748 83045 2752
rect 82981 2692 82985 2748
rect 82985 2692 83041 2748
rect 83041 2692 83045 2748
rect 82981 2688 83045 2692
rect 83061 2748 83125 2752
rect 83061 2692 83065 2748
rect 83065 2692 83121 2748
rect 83121 2692 83125 2748
rect 83061 2688 83125 2692
rect 83141 2748 83205 2752
rect 83141 2692 83145 2748
rect 83145 2692 83201 2748
rect 83201 2692 83205 2748
rect 83141 2688 83205 2692
rect 83221 2748 83285 2752
rect 83221 2692 83225 2748
rect 83225 2692 83281 2748
rect 83281 2692 83285 2748
rect 83221 2688 83285 2692
rect 24388 2204 24452 2208
rect 24388 2148 24392 2204
rect 24392 2148 24448 2204
rect 24448 2148 24452 2204
rect 24388 2144 24452 2148
rect 24468 2204 24532 2208
rect 24468 2148 24472 2204
rect 24472 2148 24528 2204
rect 24528 2148 24532 2204
rect 24468 2144 24532 2148
rect 24548 2204 24612 2208
rect 24548 2148 24552 2204
rect 24552 2148 24608 2204
rect 24608 2148 24612 2204
rect 24548 2144 24612 2148
rect 24628 2204 24692 2208
rect 24628 2148 24632 2204
rect 24632 2148 24688 2204
rect 24688 2148 24692 2204
rect 24628 2144 24692 2148
rect 47825 2204 47889 2208
rect 47825 2148 47829 2204
rect 47829 2148 47885 2204
rect 47885 2148 47889 2204
rect 47825 2144 47889 2148
rect 47905 2204 47969 2208
rect 47905 2148 47909 2204
rect 47909 2148 47965 2204
rect 47965 2148 47969 2204
rect 47905 2144 47969 2148
rect 47985 2204 48049 2208
rect 47985 2148 47989 2204
rect 47989 2148 48045 2204
rect 48045 2148 48049 2204
rect 47985 2144 48049 2148
rect 48065 2204 48129 2208
rect 48065 2148 48069 2204
rect 48069 2148 48125 2204
rect 48125 2148 48129 2204
rect 48065 2144 48129 2148
rect 71262 2204 71326 2208
rect 71262 2148 71266 2204
rect 71266 2148 71322 2204
rect 71322 2148 71326 2204
rect 71262 2144 71326 2148
rect 71342 2204 71406 2208
rect 71342 2148 71346 2204
rect 71346 2148 71402 2204
rect 71402 2148 71406 2204
rect 71342 2144 71406 2148
rect 71422 2204 71486 2208
rect 71422 2148 71426 2204
rect 71426 2148 71482 2204
rect 71482 2148 71486 2204
rect 71422 2144 71486 2148
rect 71502 2204 71566 2208
rect 71502 2148 71506 2204
rect 71506 2148 71562 2204
rect 71562 2148 71566 2204
rect 71502 2144 71566 2148
rect 94699 2204 94763 2208
rect 94699 2148 94703 2204
rect 94703 2148 94759 2204
rect 94759 2148 94763 2204
rect 94699 2144 94763 2148
rect 94779 2204 94843 2208
rect 94779 2148 94783 2204
rect 94783 2148 94839 2204
rect 94839 2148 94843 2204
rect 94779 2144 94843 2148
rect 94859 2204 94923 2208
rect 94859 2148 94863 2204
rect 94863 2148 94919 2204
rect 94919 2148 94923 2204
rect 94859 2144 94923 2148
rect 94939 2204 95003 2208
rect 94939 2148 94943 2204
rect 94943 2148 94999 2204
rect 94999 2148 95003 2204
rect 94939 2144 95003 2148
<< metal4 >>
rect 12662 16896 12982 17456
rect 12662 16832 12670 16896
rect 12734 16832 12750 16896
rect 12814 16832 12830 16896
rect 12894 16832 12910 16896
rect 12974 16832 12982 16896
rect 12662 15808 12982 16832
rect 12662 15744 12670 15808
rect 12734 15744 12750 15808
rect 12814 15744 12830 15808
rect 12894 15744 12910 15808
rect 12974 15744 12982 15808
rect 12662 14720 12982 15744
rect 12662 14656 12670 14720
rect 12734 14656 12750 14720
rect 12814 14656 12830 14720
rect 12894 14656 12910 14720
rect 12974 14656 12982 14720
rect 12662 13632 12982 14656
rect 12662 13568 12670 13632
rect 12734 13568 12750 13632
rect 12814 13568 12830 13632
rect 12894 13568 12910 13632
rect 12974 13568 12982 13632
rect 12662 12544 12982 13568
rect 12662 12480 12670 12544
rect 12734 12480 12750 12544
rect 12814 12480 12830 12544
rect 12894 12480 12910 12544
rect 12974 12480 12982 12544
rect 12662 11456 12982 12480
rect 12662 11392 12670 11456
rect 12734 11392 12750 11456
rect 12814 11392 12830 11456
rect 12894 11392 12910 11456
rect 12974 11392 12982 11456
rect 12662 10368 12982 11392
rect 12662 10304 12670 10368
rect 12734 10304 12750 10368
rect 12814 10304 12830 10368
rect 12894 10304 12910 10368
rect 12974 10304 12982 10368
rect 12662 9280 12982 10304
rect 12662 9216 12670 9280
rect 12734 9216 12750 9280
rect 12814 9216 12830 9280
rect 12894 9216 12910 9280
rect 12974 9216 12982 9280
rect 12662 8192 12982 9216
rect 12662 8128 12670 8192
rect 12734 8128 12750 8192
rect 12814 8128 12830 8192
rect 12894 8128 12910 8192
rect 12974 8128 12982 8192
rect 12662 7104 12982 8128
rect 12662 7040 12670 7104
rect 12734 7040 12750 7104
rect 12814 7040 12830 7104
rect 12894 7040 12910 7104
rect 12974 7040 12982 7104
rect 12662 6016 12982 7040
rect 12662 5952 12670 6016
rect 12734 5952 12750 6016
rect 12814 5952 12830 6016
rect 12894 5952 12910 6016
rect 12974 5952 12982 6016
rect 12662 4928 12982 5952
rect 12662 4864 12670 4928
rect 12734 4864 12750 4928
rect 12814 4864 12830 4928
rect 12894 4864 12910 4928
rect 12974 4864 12982 4928
rect 12662 3840 12982 4864
rect 12662 3776 12670 3840
rect 12734 3776 12750 3840
rect 12814 3776 12830 3840
rect 12894 3776 12910 3840
rect 12974 3776 12982 3840
rect 12662 2752 12982 3776
rect 12662 2688 12670 2752
rect 12734 2688 12750 2752
rect 12814 2688 12830 2752
rect 12894 2688 12910 2752
rect 12974 2688 12982 2752
rect 12662 2128 12982 2688
rect 24380 17440 24700 17456
rect 24380 17376 24388 17440
rect 24452 17376 24468 17440
rect 24532 17376 24548 17440
rect 24612 17376 24628 17440
rect 24692 17376 24700 17440
rect 24380 16352 24700 17376
rect 24380 16288 24388 16352
rect 24452 16288 24468 16352
rect 24532 16288 24548 16352
rect 24612 16288 24628 16352
rect 24692 16288 24700 16352
rect 24380 15264 24700 16288
rect 24380 15200 24388 15264
rect 24452 15200 24468 15264
rect 24532 15200 24548 15264
rect 24612 15200 24628 15264
rect 24692 15200 24700 15264
rect 24380 14176 24700 15200
rect 24380 14112 24388 14176
rect 24452 14112 24468 14176
rect 24532 14112 24548 14176
rect 24612 14112 24628 14176
rect 24692 14112 24700 14176
rect 24380 13088 24700 14112
rect 24380 13024 24388 13088
rect 24452 13024 24468 13088
rect 24532 13024 24548 13088
rect 24612 13024 24628 13088
rect 24692 13024 24700 13088
rect 24380 12000 24700 13024
rect 24380 11936 24388 12000
rect 24452 11936 24468 12000
rect 24532 11936 24548 12000
rect 24612 11936 24628 12000
rect 24692 11936 24700 12000
rect 24380 10912 24700 11936
rect 24380 10848 24388 10912
rect 24452 10848 24468 10912
rect 24532 10848 24548 10912
rect 24612 10848 24628 10912
rect 24692 10848 24700 10912
rect 24380 9824 24700 10848
rect 24380 9760 24388 9824
rect 24452 9760 24468 9824
rect 24532 9760 24548 9824
rect 24612 9760 24628 9824
rect 24692 9760 24700 9824
rect 24380 8736 24700 9760
rect 24380 8672 24388 8736
rect 24452 8672 24468 8736
rect 24532 8672 24548 8736
rect 24612 8672 24628 8736
rect 24692 8672 24700 8736
rect 24380 7648 24700 8672
rect 24380 7584 24388 7648
rect 24452 7584 24468 7648
rect 24532 7584 24548 7648
rect 24612 7584 24628 7648
rect 24692 7584 24700 7648
rect 24380 6560 24700 7584
rect 24380 6496 24388 6560
rect 24452 6496 24468 6560
rect 24532 6496 24548 6560
rect 24612 6496 24628 6560
rect 24692 6496 24700 6560
rect 24380 5472 24700 6496
rect 24380 5408 24388 5472
rect 24452 5408 24468 5472
rect 24532 5408 24548 5472
rect 24612 5408 24628 5472
rect 24692 5408 24700 5472
rect 24380 4384 24700 5408
rect 24380 4320 24388 4384
rect 24452 4320 24468 4384
rect 24532 4320 24548 4384
rect 24612 4320 24628 4384
rect 24692 4320 24700 4384
rect 24380 3296 24700 4320
rect 24380 3232 24388 3296
rect 24452 3232 24468 3296
rect 24532 3232 24548 3296
rect 24612 3232 24628 3296
rect 24692 3232 24700 3296
rect 24380 2208 24700 3232
rect 24380 2144 24388 2208
rect 24452 2144 24468 2208
rect 24532 2144 24548 2208
rect 24612 2144 24628 2208
rect 24692 2144 24700 2208
rect 24380 2128 24700 2144
rect 36099 16896 36419 17456
rect 36099 16832 36107 16896
rect 36171 16832 36187 16896
rect 36251 16832 36267 16896
rect 36331 16832 36347 16896
rect 36411 16832 36419 16896
rect 36099 15808 36419 16832
rect 36099 15744 36107 15808
rect 36171 15744 36187 15808
rect 36251 15744 36267 15808
rect 36331 15744 36347 15808
rect 36411 15744 36419 15808
rect 36099 14720 36419 15744
rect 36099 14656 36107 14720
rect 36171 14656 36187 14720
rect 36251 14656 36267 14720
rect 36331 14656 36347 14720
rect 36411 14656 36419 14720
rect 36099 13632 36419 14656
rect 36099 13568 36107 13632
rect 36171 13568 36187 13632
rect 36251 13568 36267 13632
rect 36331 13568 36347 13632
rect 36411 13568 36419 13632
rect 36099 12544 36419 13568
rect 36099 12480 36107 12544
rect 36171 12480 36187 12544
rect 36251 12480 36267 12544
rect 36331 12480 36347 12544
rect 36411 12480 36419 12544
rect 36099 11456 36419 12480
rect 36099 11392 36107 11456
rect 36171 11392 36187 11456
rect 36251 11392 36267 11456
rect 36331 11392 36347 11456
rect 36411 11392 36419 11456
rect 36099 10368 36419 11392
rect 36099 10304 36107 10368
rect 36171 10304 36187 10368
rect 36251 10304 36267 10368
rect 36331 10304 36347 10368
rect 36411 10304 36419 10368
rect 36099 9280 36419 10304
rect 36099 9216 36107 9280
rect 36171 9216 36187 9280
rect 36251 9216 36267 9280
rect 36331 9216 36347 9280
rect 36411 9216 36419 9280
rect 36099 8192 36419 9216
rect 36099 8128 36107 8192
rect 36171 8128 36187 8192
rect 36251 8128 36267 8192
rect 36331 8128 36347 8192
rect 36411 8128 36419 8192
rect 36099 7104 36419 8128
rect 36099 7040 36107 7104
rect 36171 7040 36187 7104
rect 36251 7040 36267 7104
rect 36331 7040 36347 7104
rect 36411 7040 36419 7104
rect 36099 6016 36419 7040
rect 36099 5952 36107 6016
rect 36171 5952 36187 6016
rect 36251 5952 36267 6016
rect 36331 5952 36347 6016
rect 36411 5952 36419 6016
rect 36099 4928 36419 5952
rect 36099 4864 36107 4928
rect 36171 4864 36187 4928
rect 36251 4864 36267 4928
rect 36331 4864 36347 4928
rect 36411 4864 36419 4928
rect 36099 3840 36419 4864
rect 36099 3776 36107 3840
rect 36171 3776 36187 3840
rect 36251 3776 36267 3840
rect 36331 3776 36347 3840
rect 36411 3776 36419 3840
rect 36099 2752 36419 3776
rect 36099 2688 36107 2752
rect 36171 2688 36187 2752
rect 36251 2688 36267 2752
rect 36331 2688 36347 2752
rect 36411 2688 36419 2752
rect 36099 2128 36419 2688
rect 47817 17440 48137 17456
rect 47817 17376 47825 17440
rect 47889 17376 47905 17440
rect 47969 17376 47985 17440
rect 48049 17376 48065 17440
rect 48129 17376 48137 17440
rect 47817 16352 48137 17376
rect 47817 16288 47825 16352
rect 47889 16288 47905 16352
rect 47969 16288 47985 16352
rect 48049 16288 48065 16352
rect 48129 16288 48137 16352
rect 47817 15264 48137 16288
rect 47817 15200 47825 15264
rect 47889 15200 47905 15264
rect 47969 15200 47985 15264
rect 48049 15200 48065 15264
rect 48129 15200 48137 15264
rect 47817 14176 48137 15200
rect 47817 14112 47825 14176
rect 47889 14112 47905 14176
rect 47969 14112 47985 14176
rect 48049 14112 48065 14176
rect 48129 14112 48137 14176
rect 47817 13088 48137 14112
rect 47817 13024 47825 13088
rect 47889 13024 47905 13088
rect 47969 13024 47985 13088
rect 48049 13024 48065 13088
rect 48129 13024 48137 13088
rect 47817 12000 48137 13024
rect 47817 11936 47825 12000
rect 47889 11936 47905 12000
rect 47969 11936 47985 12000
rect 48049 11936 48065 12000
rect 48129 11936 48137 12000
rect 47817 10912 48137 11936
rect 59536 16896 59856 17456
rect 59536 16832 59544 16896
rect 59608 16832 59624 16896
rect 59688 16832 59704 16896
rect 59768 16832 59784 16896
rect 59848 16832 59856 16896
rect 59536 15808 59856 16832
rect 59536 15744 59544 15808
rect 59608 15744 59624 15808
rect 59688 15744 59704 15808
rect 59768 15744 59784 15808
rect 59848 15744 59856 15808
rect 59536 14720 59856 15744
rect 59536 14656 59544 14720
rect 59608 14656 59624 14720
rect 59688 14656 59704 14720
rect 59768 14656 59784 14720
rect 59848 14656 59856 14720
rect 59536 13632 59856 14656
rect 59536 13568 59544 13632
rect 59608 13568 59624 13632
rect 59688 13568 59704 13632
rect 59768 13568 59784 13632
rect 59848 13568 59856 13632
rect 59536 12544 59856 13568
rect 71254 17440 71574 17456
rect 71254 17376 71262 17440
rect 71326 17376 71342 17440
rect 71406 17376 71422 17440
rect 71486 17376 71502 17440
rect 71566 17376 71574 17440
rect 71254 16352 71574 17376
rect 71254 16288 71262 16352
rect 71326 16288 71342 16352
rect 71406 16288 71422 16352
rect 71486 16288 71502 16352
rect 71566 16288 71574 16352
rect 71254 15264 71574 16288
rect 71254 15200 71262 15264
rect 71326 15200 71342 15264
rect 71406 15200 71422 15264
rect 71486 15200 71502 15264
rect 71566 15200 71574 15264
rect 71254 14176 71574 15200
rect 71254 14112 71262 14176
rect 71326 14112 71342 14176
rect 71406 14112 71422 14176
rect 71486 14112 71502 14176
rect 71566 14112 71574 14176
rect 60227 13156 60293 13157
rect 60227 13092 60228 13156
rect 60292 13092 60293 13156
rect 60227 13091 60293 13092
rect 60230 12749 60290 13091
rect 71254 13088 71574 14112
rect 71254 13024 71262 13088
rect 71326 13024 71342 13088
rect 71406 13024 71422 13088
rect 71486 13024 71502 13088
rect 71566 13024 71574 13088
rect 60227 12748 60293 12749
rect 60227 12684 60228 12748
rect 60292 12684 60293 12748
rect 60227 12683 60293 12684
rect 59536 12480 59544 12544
rect 59608 12480 59624 12544
rect 59688 12480 59704 12544
rect 59768 12480 59784 12544
rect 59848 12480 59856 12544
rect 59536 11456 59856 12480
rect 59536 11392 59544 11456
rect 59608 11392 59624 11456
rect 59688 11392 59704 11456
rect 59768 11392 59784 11456
rect 59848 11392 59856 11456
rect 59307 11116 59373 11117
rect 59307 11052 59308 11116
rect 59372 11052 59373 11116
rect 59307 11051 59373 11052
rect 47817 10848 47825 10912
rect 47889 10848 47905 10912
rect 47969 10848 47985 10912
rect 48049 10848 48065 10912
rect 48129 10848 48137 10912
rect 47817 9824 48137 10848
rect 47817 9760 47825 9824
rect 47889 9760 47905 9824
rect 47969 9760 47985 9824
rect 48049 9760 48065 9824
rect 48129 9760 48137 9824
rect 47817 8736 48137 9760
rect 59310 8805 59370 11051
rect 59536 10368 59856 11392
rect 59536 10304 59544 10368
rect 59608 10304 59624 10368
rect 59688 10304 59704 10368
rect 59768 10304 59784 10368
rect 59848 10304 59856 10368
rect 59536 9280 59856 10304
rect 59536 9216 59544 9280
rect 59608 9216 59624 9280
rect 59688 9216 59704 9280
rect 59768 9216 59784 9280
rect 59848 9216 59856 9280
rect 59307 8804 59373 8805
rect 59307 8740 59308 8804
rect 59372 8740 59373 8804
rect 59307 8739 59373 8740
rect 47817 8672 47825 8736
rect 47889 8672 47905 8736
rect 47969 8672 47985 8736
rect 48049 8672 48065 8736
rect 48129 8672 48137 8736
rect 47817 7648 48137 8672
rect 47817 7584 47825 7648
rect 47889 7584 47905 7648
rect 47969 7584 47985 7648
rect 48049 7584 48065 7648
rect 48129 7584 48137 7648
rect 47817 6560 48137 7584
rect 47817 6496 47825 6560
rect 47889 6496 47905 6560
rect 47969 6496 47985 6560
rect 48049 6496 48065 6560
rect 48129 6496 48137 6560
rect 47817 5472 48137 6496
rect 47817 5408 47825 5472
rect 47889 5408 47905 5472
rect 47969 5408 47985 5472
rect 48049 5408 48065 5472
rect 48129 5408 48137 5472
rect 47817 4384 48137 5408
rect 47817 4320 47825 4384
rect 47889 4320 47905 4384
rect 47969 4320 47985 4384
rect 48049 4320 48065 4384
rect 48129 4320 48137 4384
rect 47817 3296 48137 4320
rect 47817 3232 47825 3296
rect 47889 3232 47905 3296
rect 47969 3232 47985 3296
rect 48049 3232 48065 3296
rect 48129 3232 48137 3296
rect 47817 2208 48137 3232
rect 47817 2144 47825 2208
rect 47889 2144 47905 2208
rect 47969 2144 47985 2208
rect 48049 2144 48065 2208
rect 48129 2144 48137 2208
rect 47817 2128 48137 2144
rect 59536 8192 59856 9216
rect 71254 12000 71574 13024
rect 71254 11936 71262 12000
rect 71326 11936 71342 12000
rect 71406 11936 71422 12000
rect 71486 11936 71502 12000
rect 71566 11936 71574 12000
rect 71254 10912 71574 11936
rect 71254 10848 71262 10912
rect 71326 10848 71342 10912
rect 71406 10848 71422 10912
rect 71486 10848 71502 10912
rect 71566 10848 71574 10912
rect 71254 9824 71574 10848
rect 71254 9760 71262 9824
rect 71326 9760 71342 9824
rect 71406 9760 71422 9824
rect 71486 9760 71502 9824
rect 71566 9760 71574 9824
rect 71254 8736 71574 9760
rect 71254 8672 71262 8736
rect 71326 8672 71342 8736
rect 71406 8672 71422 8736
rect 71486 8672 71502 8736
rect 71566 8672 71574 8736
rect 63539 8532 63605 8533
rect 63539 8468 63540 8532
rect 63604 8468 63605 8532
rect 63539 8467 63605 8468
rect 59536 8128 59544 8192
rect 59608 8128 59624 8192
rect 59688 8128 59704 8192
rect 59768 8128 59784 8192
rect 59848 8128 59856 8192
rect 59536 7104 59856 8128
rect 59536 7040 59544 7104
rect 59608 7040 59624 7104
rect 59688 7040 59704 7104
rect 59768 7040 59784 7104
rect 59848 7040 59856 7104
rect 59536 6016 59856 7040
rect 59536 5952 59544 6016
rect 59608 5952 59624 6016
rect 59688 5952 59704 6016
rect 59768 5952 59784 6016
rect 59848 5952 59856 6016
rect 59536 4928 59856 5952
rect 59536 4864 59544 4928
rect 59608 4864 59624 4928
rect 59688 4864 59704 4928
rect 59768 4864 59784 4928
rect 59848 4864 59856 4928
rect 59536 3840 59856 4864
rect 63542 4861 63602 8467
rect 71254 7648 71574 8672
rect 71254 7584 71262 7648
rect 71326 7584 71342 7648
rect 71406 7584 71422 7648
rect 71486 7584 71502 7648
rect 71566 7584 71574 7648
rect 71254 6560 71574 7584
rect 71254 6496 71262 6560
rect 71326 6496 71342 6560
rect 71406 6496 71422 6560
rect 71486 6496 71502 6560
rect 71566 6496 71574 6560
rect 71254 5472 71574 6496
rect 71254 5408 71262 5472
rect 71326 5408 71342 5472
rect 71406 5408 71422 5472
rect 71486 5408 71502 5472
rect 71566 5408 71574 5472
rect 63539 4860 63605 4861
rect 63539 4796 63540 4860
rect 63604 4796 63605 4860
rect 63539 4795 63605 4796
rect 59536 3776 59544 3840
rect 59608 3776 59624 3840
rect 59688 3776 59704 3840
rect 59768 3776 59784 3840
rect 59848 3776 59856 3840
rect 59536 2752 59856 3776
rect 59536 2688 59544 2752
rect 59608 2688 59624 2752
rect 59688 2688 59704 2752
rect 59768 2688 59784 2752
rect 59848 2688 59856 2752
rect 59536 2128 59856 2688
rect 71254 4384 71574 5408
rect 71254 4320 71262 4384
rect 71326 4320 71342 4384
rect 71406 4320 71422 4384
rect 71486 4320 71502 4384
rect 71566 4320 71574 4384
rect 71254 3296 71574 4320
rect 71254 3232 71262 3296
rect 71326 3232 71342 3296
rect 71406 3232 71422 3296
rect 71486 3232 71502 3296
rect 71566 3232 71574 3296
rect 71254 2208 71574 3232
rect 71254 2144 71262 2208
rect 71326 2144 71342 2208
rect 71406 2144 71422 2208
rect 71486 2144 71502 2208
rect 71566 2144 71574 2208
rect 71254 2128 71574 2144
rect 82973 16896 83293 17456
rect 82973 16832 82981 16896
rect 83045 16832 83061 16896
rect 83125 16832 83141 16896
rect 83205 16832 83221 16896
rect 83285 16832 83293 16896
rect 82973 15808 83293 16832
rect 82973 15744 82981 15808
rect 83045 15744 83061 15808
rect 83125 15744 83141 15808
rect 83205 15744 83221 15808
rect 83285 15744 83293 15808
rect 82973 14720 83293 15744
rect 82973 14656 82981 14720
rect 83045 14656 83061 14720
rect 83125 14656 83141 14720
rect 83205 14656 83221 14720
rect 83285 14656 83293 14720
rect 82973 13632 83293 14656
rect 82973 13568 82981 13632
rect 83045 13568 83061 13632
rect 83125 13568 83141 13632
rect 83205 13568 83221 13632
rect 83285 13568 83293 13632
rect 82973 12544 83293 13568
rect 82973 12480 82981 12544
rect 83045 12480 83061 12544
rect 83125 12480 83141 12544
rect 83205 12480 83221 12544
rect 83285 12480 83293 12544
rect 82973 11456 83293 12480
rect 82973 11392 82981 11456
rect 83045 11392 83061 11456
rect 83125 11392 83141 11456
rect 83205 11392 83221 11456
rect 83285 11392 83293 11456
rect 82973 10368 83293 11392
rect 82973 10304 82981 10368
rect 83045 10304 83061 10368
rect 83125 10304 83141 10368
rect 83205 10304 83221 10368
rect 83285 10304 83293 10368
rect 82973 9280 83293 10304
rect 82973 9216 82981 9280
rect 83045 9216 83061 9280
rect 83125 9216 83141 9280
rect 83205 9216 83221 9280
rect 83285 9216 83293 9280
rect 82973 8192 83293 9216
rect 82973 8128 82981 8192
rect 83045 8128 83061 8192
rect 83125 8128 83141 8192
rect 83205 8128 83221 8192
rect 83285 8128 83293 8192
rect 82973 7104 83293 8128
rect 82973 7040 82981 7104
rect 83045 7040 83061 7104
rect 83125 7040 83141 7104
rect 83205 7040 83221 7104
rect 83285 7040 83293 7104
rect 82973 6016 83293 7040
rect 82973 5952 82981 6016
rect 83045 5952 83061 6016
rect 83125 5952 83141 6016
rect 83205 5952 83221 6016
rect 83285 5952 83293 6016
rect 82973 4928 83293 5952
rect 82973 4864 82981 4928
rect 83045 4864 83061 4928
rect 83125 4864 83141 4928
rect 83205 4864 83221 4928
rect 83285 4864 83293 4928
rect 82973 3840 83293 4864
rect 82973 3776 82981 3840
rect 83045 3776 83061 3840
rect 83125 3776 83141 3840
rect 83205 3776 83221 3840
rect 83285 3776 83293 3840
rect 82973 2752 83293 3776
rect 82973 2688 82981 2752
rect 83045 2688 83061 2752
rect 83125 2688 83141 2752
rect 83205 2688 83221 2752
rect 83285 2688 83293 2752
rect 82973 2128 83293 2688
rect 94691 17440 95011 17456
rect 94691 17376 94699 17440
rect 94763 17376 94779 17440
rect 94843 17376 94859 17440
rect 94923 17376 94939 17440
rect 95003 17376 95011 17440
rect 94691 16352 95011 17376
rect 94691 16288 94699 16352
rect 94763 16288 94779 16352
rect 94843 16288 94859 16352
rect 94923 16288 94939 16352
rect 95003 16288 95011 16352
rect 94691 15264 95011 16288
rect 94691 15200 94699 15264
rect 94763 15200 94779 15264
rect 94843 15200 94859 15264
rect 94923 15200 94939 15264
rect 95003 15200 95011 15264
rect 94691 14176 95011 15200
rect 94691 14112 94699 14176
rect 94763 14112 94779 14176
rect 94843 14112 94859 14176
rect 94923 14112 94939 14176
rect 95003 14112 95011 14176
rect 94691 13088 95011 14112
rect 94691 13024 94699 13088
rect 94763 13024 94779 13088
rect 94843 13024 94859 13088
rect 94923 13024 94939 13088
rect 95003 13024 95011 13088
rect 94691 12000 95011 13024
rect 94691 11936 94699 12000
rect 94763 11936 94779 12000
rect 94843 11936 94859 12000
rect 94923 11936 94939 12000
rect 95003 11936 95011 12000
rect 94691 10912 95011 11936
rect 94691 10848 94699 10912
rect 94763 10848 94779 10912
rect 94843 10848 94859 10912
rect 94923 10848 94939 10912
rect 95003 10848 95011 10912
rect 94691 9824 95011 10848
rect 94691 9760 94699 9824
rect 94763 9760 94779 9824
rect 94843 9760 94859 9824
rect 94923 9760 94939 9824
rect 95003 9760 95011 9824
rect 94691 8736 95011 9760
rect 94691 8672 94699 8736
rect 94763 8672 94779 8736
rect 94843 8672 94859 8736
rect 94923 8672 94939 8736
rect 95003 8672 95011 8736
rect 94691 7648 95011 8672
rect 94691 7584 94699 7648
rect 94763 7584 94779 7648
rect 94843 7584 94859 7648
rect 94923 7584 94939 7648
rect 95003 7584 95011 7648
rect 94691 6560 95011 7584
rect 94691 6496 94699 6560
rect 94763 6496 94779 6560
rect 94843 6496 94859 6560
rect 94923 6496 94939 6560
rect 95003 6496 95011 6560
rect 94691 5472 95011 6496
rect 94691 5408 94699 5472
rect 94763 5408 94779 5472
rect 94843 5408 94859 5472
rect 94923 5408 94939 5472
rect 95003 5408 95011 5472
rect 94691 4384 95011 5408
rect 94691 4320 94699 4384
rect 94763 4320 94779 4384
rect 94843 4320 94859 4384
rect 94923 4320 94939 4384
rect 95003 4320 95011 4384
rect 94691 3296 95011 4320
rect 94691 3232 94699 3296
rect 94763 3232 94779 3296
rect 94843 3232 94859 3296
rect 94923 3232 94939 3296
rect 95003 3232 95011 3296
rect 94691 2208 95011 3232
rect 94691 2144 94699 2208
rect 94763 2144 94779 2208
rect 94843 2144 94859 2208
rect 94923 2144 94939 2208
rect 95003 2144 95011 2208
rect 94691 2128 95011 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__0446__1_A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 32660 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0446__2_A
timestamp 1662439860
transform 1 0 34224 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0447__A
timestamp 1662439860
transform -1 0 25024 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0458__A
timestamp 1662439860
transform -1 0 67528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0468__A
timestamp 1662439860
transform -1 0 90160 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0469__A
timestamp 1662439860
transform 1 0 79212 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0470__A
timestamp 1662439860
transform 1 0 90344 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0471__A
timestamp 1662439860
transform 1 0 85744 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0472__A
timestamp 1662439860
transform 1 0 64676 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0473__A
timestamp 1662439860
transform -1 0 78200 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0474__A
timestamp 1662439860
transform 1 0 66700 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0475__A
timestamp 1662439860
transform -1 0 94300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0476__A
timestamp 1662439860
transform -1 0 94300 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0477__A
timestamp 1662439860
transform 1 0 76084 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0478__A
timestamp 1662439860
transform 1 0 59156 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0479__A
timestamp 1662439860
transform 1 0 88320 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0480__A
timestamp 1662439860
transform -1 0 84456 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0481__A
timestamp 1662439860
transform -1 0 74244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0482__A
timestamp 1662439860
transform 1 0 85100 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0483__A
timestamp 1662439860
transform 1 0 74152 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0484__A
timestamp 1662439860
transform 1 0 58512 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0485__A
timestamp 1662439860
transform 1 0 77832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__A
timestamp 1662439860
transform 1 0 85100 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0487__A
timestamp 1662439860
transform -1 0 89884 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0488__A
timestamp 1662439860
transform -1 0 85284 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0489__A
timestamp 1662439860
transform -1 0 59616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0491__A
timestamp 1662439860
transform -1 0 22264 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0497__A
timestamp 1662439860
transform 1 0 5796 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__B
timestamp 1662439860
transform -1 0 2944 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0501__A
timestamp 1662439860
transform -1 0 20976 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0501__B
timestamp 1662439860
transform -1 0 18124 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0507__A
timestamp 1662439860
transform 1 0 43792 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0508__A
timestamp 1662439860
transform -1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0508__B
timestamp 1662439860
transform -1 0 5152 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0513__A
timestamp 1662439860
transform -1 0 59524 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0513__B
timestamp 1662439860
transform -1 0 59524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0514__A
timestamp 1662439860
transform 1 0 81788 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0517__A
timestamp 1662439860
transform -1 0 38824 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0517__B
timestamp 1662439860
transform -1 0 39008 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0518__A
timestamp 1662439860
transform -1 0 80224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__A
timestamp 1662439860
transform -1 0 88872 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__B
timestamp 1662439860
transform -1 0 81420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__A
timestamp 1662439860
transform 1 0 32384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__B
timestamp 1662439860
transform -1 0 37352 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__C
timestamp 1662439860
transform 1 0 31648 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__D_N
timestamp 1662439860
transform 1 0 31096 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__A
timestamp 1662439860
transform -1 0 53636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__B
timestamp 1662439860
transform -1 0 56580 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0528__A
timestamp 1662439860
transform 1 0 82064 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0531__B
timestamp 1662439860
transform 1 0 42964 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__A
timestamp 1662439860
transform -1 0 77924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0533__A
timestamp 1662439860
transform 1 0 64032 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0533__B
timestamp 1662439860
transform 1 0 59984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0536__A
timestamp 1662439860
transform 1 0 50508 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0536__B
timestamp 1662439860
transform 1 0 50876 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__A
timestamp 1662439860
transform -1 0 59340 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__B
timestamp 1662439860
transform -1 0 65780 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__D
timestamp 1662439860
transform -1 0 58236 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0538__A1
timestamp 1662439860
transform 1 0 11040 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0538__A2
timestamp 1662439860
transform 1 0 10488 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0539__A2
timestamp 1662439860
transform 1 0 11040 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__A
timestamp 1662439860
transform 1 0 10672 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__B
timestamp 1662439860
transform 1 0 11224 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__C_N
timestamp 1662439860
transform 1 0 10120 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0543__A
timestamp 1662439860
transform 1 0 6716 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__A
timestamp 1662439860
transform 1 0 9200 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__A
timestamp 1662439860
transform 1 0 65136 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__B
timestamp 1662439860
transform -1 0 58788 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__A
timestamp 1662439860
transform 1 0 54188 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__B
timestamp 1662439860
transform 1 0 54556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0548__B
timestamp 1662439860
transform 1 0 13432 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0548__C
timestamp 1662439860
transform 1 0 12512 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0549__A0
timestamp 1662439860
transform -1 0 38180 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0549__S
timestamp 1662439860
transform -1 0 38456 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0550__A
timestamp 1662439860
transform -1 0 24932 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__A
timestamp 1662439860
transform -1 0 32108 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__A
timestamp 1662439860
transform -1 0 68540 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__B
timestamp 1662439860
transform -1 0 69276 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0553__A
timestamp 1662439860
transform 1 0 61548 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0553__B
timestamp 1662439860
transform 1 0 62100 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0554__A
timestamp 1662439860
transform -1 0 58236 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0555__A1
timestamp 1662439860
transform 1 0 64216 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0555__S
timestamp 1662439860
transform 1 0 63664 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__A
timestamp 1662439860
transform -1 0 24380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__B
timestamp 1662439860
transform -1 0 25484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0557__A
timestamp 1662439860
transform 1 0 27140 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0557__B
timestamp 1662439860
transform -1 0 29900 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__A
timestamp 1662439860
transform -1 0 54740 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__B
timestamp 1662439860
transform 1 0 57224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__A
timestamp 1662439860
transform 1 0 61732 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__B
timestamp 1662439860
transform -1 0 56948 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__A1
timestamp 1662439860
transform 1 0 54280 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0563__A
timestamp 1662439860
transform 1 0 43608 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__A
timestamp 1662439860
transform -1 0 79488 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__B
timestamp 1662439860
transform 1 0 56672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__C
timestamp 1662439860
transform 1 0 54464 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0566__A
timestamp 1662439860
transform -1 0 41584 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__A
timestamp 1662439860
transform -1 0 43332 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__C
timestamp 1662439860
transform 1 0 49680 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__A
timestamp 1662439860
transform -1 0 5888 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__B
timestamp 1662439860
transform -1 0 7636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__A
timestamp 1662439860
transform 1 0 29992 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__B
timestamp 1662439860
transform -1 0 30728 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__A
timestamp 1662439860
transform -1 0 87308 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__B
timestamp 1662439860
transform 1 0 84364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__A
timestamp 1662439860
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__B
timestamp 1662439860
transform 1 0 5888 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__A
timestamp 1662439860
transform -1 0 7820 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__A
timestamp 1662439860
transform 1 0 9108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__A
timestamp 1662439860
transform 1 0 87400 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__B
timestamp 1662439860
transform -1 0 86572 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__B
timestamp 1662439860
transform -1 0 85376 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__A
timestamp 1662439860
transform 1 0 58052 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__B
timestamp 1662439860
transform -1 0 59432 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__A
timestamp 1662439860
transform 1 0 13340 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__B
timestamp 1662439860
transform -1 0 12328 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__A
timestamp 1662439860
transform -1 0 42964 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__B
timestamp 1662439860
transform -1 0 42412 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__A
timestamp 1662439860
transform -1 0 88780 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__B
timestamp 1662439860
transform 1 0 81236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__B
timestamp 1662439860
transform -1 0 89424 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__C
timestamp 1662439860
transform 1 0 85652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__A
timestamp 1662439860
transform 1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__B
timestamp 1662439860
transform -1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__A
timestamp 1662439860
transform -1 0 41952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__B
timestamp 1662439860
transform -1 0 42504 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__A
timestamp 1662439860
transform -1 0 59340 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__A
timestamp 1662439860
transform -1 0 37720 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__A
timestamp 1662439860
transform -1 0 23736 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0598__A
timestamp 1662439860
transform -1 0 38824 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__A
timestamp 1662439860
transform 1 0 12604 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__A
timestamp 1662439860
transform -1 0 69092 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__B
timestamp 1662439860
transform -1 0 22172 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__A
timestamp 1662439860
transform 1 0 46552 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__C
timestamp 1662439860
transform 1 0 83812 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__D
timestamp 1662439860
transform 1 0 83168 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__B
timestamp 1662439860
transform -1 0 21620 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__A
timestamp 1662439860
transform -1 0 74428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__B
timestamp 1662439860
transform 1 0 74704 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__B
timestamp 1662439860
transform -1 0 59524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__A0
timestamp 1662439860
transform -1 0 67528 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__A1
timestamp 1662439860
transform -1 0 65320 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__A
timestamp 1662439860
transform -1 0 71208 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__A
timestamp 1662439860
transform 1 0 63112 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__A
timestamp 1662439860
transform -1 0 62376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__A
timestamp 1662439860
transform -1 0 70380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A
timestamp 1662439860
transform 1 0 65136 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A
timestamp 1662439860
transform 1 0 40112 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A
timestamp 1662439860
transform -1 0 32384 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__A
timestamp 1662439860
transform 1 0 44252 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A
timestamp 1662439860
transform 1 0 29440 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A
timestamp 1662439860
transform -1 0 46644 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A
timestamp 1662439860
transform 1 0 36708 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__A
timestamp 1662439860
transform -1 0 35420 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__A
timestamp 1662439860
transform -1 0 43700 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A
timestamp 1662439860
transform 1 0 32568 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A
timestamp 1662439860
transform -1 0 53728 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__A
timestamp 1662439860
transform 1 0 36156 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A
timestamp 1662439860
transform -1 0 49496 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A
timestamp 1662439860
transform -1 0 46000 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A
timestamp 1662439860
transform -1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__B
timestamp 1662439860
transform 1 0 31648 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A
timestamp 1662439860
transform -1 0 41584 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__B
timestamp 1662439860
transform -1 0 42136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__B
timestamp 1662439860
transform -1 0 70564 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__C
timestamp 1662439860
transform 1 0 50324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A
timestamp 1662439860
transform 1 0 68632 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__C
timestamp 1662439860
transform -1 0 65228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__B
timestamp 1662439860
transform 1 0 70380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A
timestamp 1662439860
transform 1 0 61180 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__B
timestamp 1662439860
transform 1 0 62836 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__A
timestamp 1662439860
transform 1 0 64308 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__C
timestamp 1662439860
transform -1 0 63940 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A
timestamp 1662439860
transform 1 0 20884 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A
timestamp 1662439860
transform -1 0 64676 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__B1
timestamp 1662439860
transform 1 0 69184 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__A
timestamp 1662439860
transform 1 0 65412 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A
timestamp 1662439860
transform 1 0 19412 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__B1
timestamp 1662439860
transform 1 0 59708 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A
timestamp 1662439860
transform 1 0 63204 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A
timestamp 1662439860
transform 1 0 68080 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__B1
timestamp 1662439860
transform 1 0 66884 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A
timestamp 1662439860
transform -1 0 64676 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__B1
timestamp 1662439860
transform -1 0 63940 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A
timestamp 1662439860
transform -1 0 68816 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A
timestamp 1662439860
transform 1 0 35328 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A1
timestamp 1662439860
transform -1 0 61640 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A2
timestamp 1662439860
transform 1 0 64860 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A
timestamp 1662439860
transform 1 0 60628 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A
timestamp 1662439860
transform -1 0 59340 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B1
timestamp 1662439860
transform 1 0 61732 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__A
timestamp 1662439860
transform 1 0 67344 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B1
timestamp 1662439860
transform -1 0 51520 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A
timestamp 1662439860
transform 1 0 52164 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__A
timestamp 1662439860
transform 1 0 46000 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__B1
timestamp 1662439860
transform 1 0 50876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__B1
timestamp 1662439860
transform 1 0 49680 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A
timestamp 1662439860
transform 1 0 44252 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A
timestamp 1662439860
transform -1 0 43424 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__B1
timestamp 1662439860
transform 1 0 46920 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B1
timestamp 1662439860
transform -1 0 57316 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__B1
timestamp 1662439860
transform 1 0 57868 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__C1
timestamp 1662439860
transform 1 0 69736 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__B
timestamp 1662439860
transform 1 0 65044 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A
timestamp 1662439860
transform 1 0 84732 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__C
timestamp 1662439860
transform 1 0 76084 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A
timestamp 1662439860
transform -1 0 85376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A
timestamp 1662439860
transform 1 0 76820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B1
timestamp 1662439860
transform -1 0 84732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B1
timestamp 1662439860
transform -1 0 81052 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__B1
timestamp 1662439860
transform 1 0 81788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__B1
timestamp 1662439860
transform 1 0 75072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A1
timestamp 1662439860
transform 1 0 75900 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A
timestamp 1662439860
transform 1 0 73324 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__A
timestamp 1662439860
transform -1 0 76452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B1
timestamp 1662439860
transform 1 0 74244 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__B1
timestamp 1662439860
transform -1 0 77556 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A
timestamp 1662439860
transform 1 0 81420 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A
timestamp 1662439860
transform 1 0 73968 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__B1
timestamp 1662439860
transform 1 0 69184 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__B1
timestamp 1662439860
transform 1 0 71392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A
timestamp 1662439860
transform -1 0 78844 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__B1
timestamp 1662439860
transform -1 0 78108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A
timestamp 1662439860
transform -1 0 89976 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A
timestamp 1662439860
transform -1 0 90896 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__A
timestamp 1662439860
transform 1 0 65412 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__B1
timestamp 1662439860
transform 1 0 90344 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A
timestamp 1662439860
transform -1 0 86112 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__B1
timestamp 1662439860
transform -1 0 86940 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A
timestamp 1662439860
transform 1 0 86572 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__C1
timestamp 1662439860
transform -1 0 85192 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A
timestamp 1662439860
transform -1 0 80224 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1662439860
transform -1 0 94208 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A
timestamp 1662439860
transform -1 0 79764 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__B
timestamp 1662439860
transform -1 0 81696 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A1
timestamp 1662439860
transform 1 0 81880 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A2
timestamp 1662439860
transform 1 0 80132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__B1
timestamp 1662439860
transform -1 0 76636 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A1
timestamp 1662439860
transform 1 0 79580 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A2
timestamp 1662439860
transform 1 0 75440 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__B
timestamp 1662439860
transform 1 0 59892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A
timestamp 1662439860
transform 1 0 59248 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A1
timestamp 1662439860
transform -1 0 58788 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__C1
timestamp 1662439860
transform 1 0 62284 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__B
timestamp 1662439860
transform 1 0 78660 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A1
timestamp 1662439860
transform 1 0 71944 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__B1
timestamp 1662439860
transform -1 0 74888 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__B2
timestamp 1662439860
transform 1 0 73600 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A
timestamp 1662439860
transform -1 0 71116 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__B
timestamp 1662439860
transform 1 0 74152 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A2
timestamp 1662439860
transform -1 0 85928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__B1
timestamp 1662439860
transform -1 0 85468 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A
timestamp 1662439860
transform 1 0 76084 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__B
timestamp 1662439860
transform 1 0 75808 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A_N
timestamp 1662439860
transform -1 0 76544 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__B_N
timestamp 1662439860
transform -1 0 78200 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__D
timestamp 1662439860
transform -1 0 76084 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A1
timestamp 1662439860
transform 1 0 79304 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A3
timestamp 1662439860
transform -1 0 81972 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__B1
timestamp 1662439860
transform 1 0 81236 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A1
timestamp 1662439860
transform -1 0 85376 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A2
timestamp 1662439860
transform -1 0 79028 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A1
timestamp 1662439860
transform 1 0 80592 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A1
timestamp 1662439860
transform -1 0 81420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A2
timestamp 1662439860
transform -1 0 81144 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__A
timestamp 1662439860
transform 1 0 22908 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__B
timestamp 1662439860
transform -1 0 22540 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__C
timestamp 1662439860
transform 1 0 24104 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__B
timestamp 1662439860
transform 1 0 37720 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__D
timestamp 1662439860
transform -1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__A
timestamp 1662439860
transform 1 0 47104 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__B
timestamp 1662439860
transform 1 0 46276 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__C
timestamp 1662439860
transform 1 0 45632 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A
timestamp 1662439860
transform 1 0 45448 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__B
timestamp 1662439860
transform 1 0 47748 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A
timestamp 1662439860
transform 1 0 21988 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__B
timestamp 1662439860
transform 1 0 22264 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__A
timestamp 1662439860
transform 1 0 41400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__C
timestamp 1662439860
transform -1 0 42780 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__B
timestamp 1662439860
transform 1 0 38272 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__C
timestamp 1662439860
transform 1 0 41952 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A
timestamp 1662439860
transform 1 0 48392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__B
timestamp 1662439860
transform 1 0 46000 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__C
timestamp 1662439860
transform 1 0 46552 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__B1
timestamp 1662439860
transform 1 0 46828 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__A
timestamp 1662439860
transform 1 0 43976 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A
timestamp 1662439860
transform 1 0 51612 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__B
timestamp 1662439860
transform 1 0 52164 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A
timestamp 1662439860
transform -1 0 53912 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B1
timestamp 1662439860
transform 1 0 57408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A
timestamp 1662439860
transform 1 0 58052 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A
timestamp 1662439860
transform -1 0 52072 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__B1
timestamp 1662439860
transform 1 0 51980 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A
timestamp 1662439860
transform 1 0 47840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A
timestamp 1662439860
transform 1 0 46000 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A_N
timestamp 1662439860
transform 1 0 44528 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__B1
timestamp 1662439860
transform 1 0 44896 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A
timestamp 1662439860
transform 1 0 45172 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A2
timestamp 1662439860
transform 1 0 40112 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__A
timestamp 1662439860
transform 1 0 37996 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A
timestamp 1662439860
transform 1 0 34224 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__B1
timestamp 1662439860
transform 1 0 38180 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__A
timestamp 1662439860
transform -1 0 41032 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B
timestamp 1662439860
transform -1 0 39192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__A_N
timestamp 1662439860
transform 1 0 39560 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__B1
timestamp 1662439860
transform -1 0 40848 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A1
timestamp 1662439860
transform 1 0 39376 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A
timestamp 1662439860
transform -1 0 40940 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A
timestamp 1662439860
transform 1 0 40112 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1662439860
transform -1 0 39100 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A2
timestamp 1662439860
transform -1 0 38640 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__B1
timestamp 1662439860
transform 1 0 38824 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A2
timestamp 1662439860
transform -1 0 46736 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__B1
timestamp 1662439860
transform 1 0 45172 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A
timestamp 1662439860
transform -1 0 46460 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A
timestamp 1662439860
transform 1 0 20976 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__B1
timestamp 1662439860
transform 1 0 17848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A
timestamp 1662439860
transform -1 0 23000 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__B
timestamp 1662439860
transform 1 0 22908 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A
timestamp 1662439860
transform -1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__B
timestamp 1662439860
transform 1 0 23368 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__B1
timestamp 1662439860
transform -1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A
timestamp 1662439860
transform 1 0 24748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__B
timestamp 1662439860
transform 1 0 24104 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__B1
timestamp 1662439860
transform 1 0 25392 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1662439860
transform 1 0 41860 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__B
timestamp 1662439860
transform -1 0 43240 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__C1
timestamp 1662439860
transform 1 0 44528 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A
timestamp 1662439860
transform -1 0 32476 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__B
timestamp 1662439860
transform 1 0 33764 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__A
timestamp 1662439860
transform 1 0 58696 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A
timestamp 1662439860
transform 1 0 51428 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__B
timestamp 1662439860
transform 1 0 51612 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__B
timestamp 1662439860
transform -1 0 63480 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A
timestamp 1662439860
transform 1 0 39560 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__B
timestamp 1662439860
transform 1 0 27968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A
timestamp 1662439860
transform 1 0 22540 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A
timestamp 1662439860
transform -1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__B
timestamp 1662439860
transform -1 0 37996 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__D
timestamp 1662439860
transform -1 0 38548 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A
timestamp 1662439860
transform 1 0 44068 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__B
timestamp 1662439860
transform 1 0 30636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__B
timestamp 1662439860
transform -1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__B
timestamp 1662439860
transform 1 0 19412 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__C
timestamp 1662439860
transform -1 0 15456 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__B
timestamp 1662439860
transform -1 0 44068 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__D
timestamp 1662439860
transform -1 0 43792 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__B1
timestamp 1662439860
transform -1 0 39560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__B
timestamp 1662439860
transform 1 0 37720 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__C
timestamp 1662439860
transform 1 0 39192 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A
timestamp 1662439860
transform 1 0 39376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__B1
timestamp 1662439860
transform 1 0 37628 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__B
timestamp 1662439860
transform 1 0 45080 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__B1
timestamp 1662439860
transform 1 0 43056 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A
timestamp 1662439860
transform 1 0 46184 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A
timestamp 1662439860
transform 1 0 23000 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__B
timestamp 1662439860
transform -1 0 17664 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A_N
timestamp 1662439860
transform 1 0 37628 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__B
timestamp 1662439860
transform -1 0 37352 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A1
timestamp 1662439860
transform 1 0 36800 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__B1
timestamp 1662439860
transform 1 0 35880 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A2
timestamp 1662439860
transform 1 0 23092 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__B1
timestamp 1662439860
transform -1 0 17112 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A
timestamp 1662439860
transform -1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1662439860
transform 1 0 21988 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A2
timestamp 1662439860
transform 1 0 16836 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__B1
timestamp 1662439860
transform -1 0 15732 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 1662439860
transform -1 0 14628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A
timestamp 1662439860
transform -1 0 17572 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__B1
timestamp 1662439860
transform 1 0 16560 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A2
timestamp 1662439860
transform 1 0 17664 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A
timestamp 1662439860
transform 1 0 15272 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__B1
timestamp 1662439860
transform 1 0 23736 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A
timestamp 1662439860
transform 1 0 23000 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__B1
timestamp 1662439860
transform 1 0 22816 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A
timestamp 1662439860
transform 1 0 18216 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__B1
timestamp 1662439860
transform 1 0 16836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__B
timestamp 1662439860
transform -1 0 34592 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__B
timestamp 1662439860
transform 1 0 35328 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__B1
timestamp 1662439860
transform 1 0 31004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__B
timestamp 1662439860
transform 1 0 33028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__B1
timestamp 1662439860
transform 1 0 35880 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__C1
timestamp 1662439860
transform 1 0 39744 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A
timestamp 1662439860
transform 1 0 37444 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__B
timestamp 1662439860
transform -1 0 38824 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A
timestamp 1662439860
transform 1 0 34132 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__B
timestamp 1662439860
transform 1 0 35788 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A
timestamp 1662439860
transform 1 0 30084 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__B
timestamp 1662439860
transform -1 0 31188 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A
timestamp 1662439860
transform -1 0 34868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__B
timestamp 1662439860
transform -1 0 33028 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A
timestamp 1662439860
transform -1 0 48392 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__B
timestamp 1662439860
transform -1 0 47196 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A
timestamp 1662439860
transform -1 0 47932 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__B
timestamp 1662439860
transform 1 0 42872 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__A
timestamp 1662439860
transform 1 0 43332 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__B
timestamp 1662439860
transform -1 0 72680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A_N
timestamp 1662439860
transform 1 0 71944 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__B
timestamp 1662439860
transform -1 0 35696 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A
timestamp 1662439860
transform -1 0 61180 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__B
timestamp 1662439860
transform 1 0 64768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__C
timestamp 1662439860
transform -1 0 57224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__A1
timestamp 1662439860
transform -1 0 49312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__B1
timestamp 1662439860
transform -1 0 47288 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A1
timestamp 1662439860
transform -1 0 53912 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__B2
timestamp 1662439860
transform 1 0 50324 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A1
timestamp 1662439860
transform -1 0 54648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A2
timestamp 1662439860
transform -1 0 53544 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__C1
timestamp 1662439860
transform -1 0 57592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A2
timestamp 1662439860
transform 1 0 53728 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A3
timestamp 1662439860
transform -1 0 54096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__C1
timestamp 1662439860
transform 1 0 58236 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__B
timestamp 1662439860
transform -1 0 9936 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A
timestamp 1662439860
transform 1 0 49956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__B
timestamp 1662439860
transform 1 0 50324 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__B1
timestamp 1662439860
transform 1 0 50876 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__A1
timestamp 1662439860
transform -1 0 47288 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A
timestamp 1662439860
transform 1 0 7360 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__B
timestamp 1662439860
transform -1 0 6992 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A
timestamp 1662439860
transform -1 0 42136 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A
timestamp 1662439860
transform 1 0 53084 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A
timestamp 1662439860
transform 1 0 85192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A
timestamp 1662439860
transform -1 0 90252 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A
timestamp 1662439860
transform -1 0 89148 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A
timestamp 1662439860
transform 1 0 73600 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A
timestamp 1662439860
transform -1 0 54832 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1662439860
transform 1 0 63204 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A
timestamp 1662439860
transform 1 0 88320 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A
timestamp 1662439860
transform 1 0 78016 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A
timestamp 1662439860
transform -1 0 89700 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__B
timestamp 1662439860
transform 1 0 23552 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A
timestamp 1662439860
transform 1 0 63204 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A
timestamp 1662439860
transform 1 0 70288 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A
timestamp 1662439860
transform -1 0 64124 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__B
timestamp 1662439860
transform -1 0 63572 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__A
timestamp 1662439860
transform -1 0 90896 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__A
timestamp 1662439860
transform 1 0 88228 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__B
timestamp 1662439860
transform 1 0 86296 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__A
timestamp 1662439860
transform -1 0 94300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A
timestamp 1662439860
transform -1 0 83260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__B
timestamp 1662439860
transform 1 0 82892 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__A
timestamp 1662439860
transform 1 0 59892 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__B
timestamp 1662439860
transform 1 0 60444 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__A
timestamp 1662439860
transform 1 0 66792 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__A
timestamp 1662439860
transform -1 0 39284 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__B
timestamp 1662439860
transform -1 0 36432 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__A
timestamp 1662439860
transform 1 0 82340 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__B
timestamp 1662439860
transform -1 0 37628 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A
timestamp 1662439860
transform 1 0 74152 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__A
timestamp 1662439860
transform 1 0 48024 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__B
timestamp 1662439860
transform 1 0 45540 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A
timestamp 1662439860
transform 1 0 79396 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__A
timestamp 1662439860
transform -1 0 86572 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__A
timestamp 1662439860
transform 1 0 41952 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__B
timestamp 1662439860
transform 1 0 39376 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__A
timestamp 1662439860
transform -1 0 94300 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__A
timestamp 1662439860
transform 1 0 54924 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__B
timestamp 1662439860
transform 1 0 54832 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A
timestamp 1662439860
transform -1 0 90712 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__A
timestamp 1662439860
transform 1 0 64952 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A
timestamp 1662439860
transform -1 0 4784 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__A
timestamp 1662439860
transform 1 0 4968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A
timestamp 1662439860
transform -1 0 15088 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__A
timestamp 1662439860
transform 1 0 82340 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__B
timestamp 1662439860
transform -1 0 81420 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A
timestamp 1662439860
transform 1 0 87952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__B
timestamp 1662439860
transform 1 0 87952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__A
timestamp 1662439860
transform -1 0 80592 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__B
timestamp 1662439860
transform -1 0 80040 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A
timestamp 1662439860
transform -1 0 83812 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__B
timestamp 1662439860
transform -1 0 88780 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A
timestamp 1662439860
transform -1 0 52164 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__B
timestamp 1662439860
transform -1 0 52348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__B
timestamp 1662439860
transform -1 0 36800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__A
timestamp 1662439860
transform -1 0 50508 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__B
timestamp 1662439860
transform -1 0 50508 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A
timestamp 1662439860
transform 1 0 42412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__B
timestamp 1662439860
transform 1 0 40940 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__A
timestamp 1662439860
transform -1 0 58788 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__A
timestamp 1662439860
transform -1 0 56212 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__B
timestamp 1662439860
transform -1 0 55660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__A
timestamp 1662439860
transform -1 0 31464 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__B
timestamp 1662439860
transform 1 0 28520 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A
timestamp 1662439860
transform -1 0 13340 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__B
timestamp 1662439860
transform 1 0 14536 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__A
timestamp 1662439860
transform 1 0 12972 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__B
timestamp 1662439860
transform 1 0 11040 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__A
timestamp 1662439860
transform 1 0 8556 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__B
timestamp 1662439860
transform 1 0 7268 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A
timestamp 1662439860
transform -1 0 30728 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__B
timestamp 1662439860
transform -1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__B
timestamp 1662439860
transform 1 0 32568 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A
timestamp 1662439860
transform -1 0 26772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__B
timestamp 1662439860
transform -1 0 24748 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__A
timestamp 1662439860
transform 1 0 28520 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__B
timestamp 1662439860
transform 1 0 29072 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__3_A
timestamp 1662439860
transform -1 0 30820 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__A
timestamp 1662439860
transform 1 0 16100 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__B
timestamp 1662439860
transform 1 0 14536 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__4_A
timestamp 1662439860
transform 1 0 35972 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__5_A
timestamp 1662439860
transform 1 0 62192 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__RESET_B
timestamp 1662439860
transform -1 0 46276 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__D
timestamp 1662439860
transform -1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__RESET_B
timestamp 1662439860
transform 1 0 44528 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__RESET_B
timestamp 1662439860
transform 1 0 49680 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__D
timestamp 1662439860
transform -1 0 45356 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__RESET_B
timestamp 1662439860
transform 1 0 44804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__RESET_B
timestamp 1662439860
transform 1 0 11960 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__RESET_B
timestamp 1662439860
transform 1 0 51060 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__RESET_B
timestamp 1662439860
transform 1 0 36800 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__CLK
timestamp 1662439860
transform 1 0 37168 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__CLK
timestamp 1662439860
transform 1 0 13156 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__D
timestamp 1662439860
transform -1 0 17020 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__CLK
timestamp 1662439860
transform 1 0 37720 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__CLK
timestamp 1662439860
transform -1 0 41216 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__CLK
timestamp 1662439860
transform -1 0 41860 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__D
timestamp 1662439860
transform -1 0 42780 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__CLK
timestamp 1662439860
transform -1 0 69736 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__CLK
timestamp 1662439860
transform 1 0 62284 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__CLK
timestamp 1662439860
transform -1 0 69920 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__CLK
timestamp 1662439860
transform 1 0 65412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__CLK
timestamp 1662439860
transform 1 0 58052 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__RESET_B
timestamp 1662439860
transform -1 0 54464 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__CLK
timestamp 1662439860
transform 1 0 43148 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__RESET_B
timestamp 1662439860
transform 1 0 41308 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__CLK
timestamp 1662439860
transform 1 0 46828 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__RESET_B
timestamp 1662439860
transform 1 0 43792 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__CLK
timestamp 1662439860
transform -1 0 56396 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__RESET_B
timestamp 1662439860
transform -1 0 55016 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__CLK
timestamp 1662439860
transform 1 0 36800 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__RESET_B
timestamp 1662439860
transform -1 0 36984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__CLK
timestamp 1662439860
transform 1 0 50968 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__RESET_B
timestamp 1662439860
transform -1 0 51336 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__CLK
timestamp 1662439860
transform -1 0 61364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__CLK
timestamp 1662439860
transform 1 0 64308 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__CLK
timestamp 1662439860
transform -1 0 54280 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__CLK
timestamp 1662439860
transform -1 0 84180 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__CLK
timestamp 1662439860
transform -1 0 88964 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__CLK
timestamp 1662439860
transform 1 0 87676 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__CLK
timestamp 1662439860
transform 1 0 73508 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__CLK
timestamp 1662439860
transform -1 0 53360 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__CLK
timestamp 1662439860
transform -1 0 52624 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__CLK
timestamp 1662439860
transform 1 0 73416 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__CLK
timestamp 1662439860
transform 1 0 65780 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__CLK
timestamp 1662439860
transform -1 0 85744 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__CLK
timestamp 1662439860
transform -1 0 85836 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__CLK
timestamp 1662439860
transform 1 0 70288 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__CLK
timestamp 1662439860
transform 1 0 70932 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__CLK
timestamp 1662439860
transform 1 0 86848 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__CLK
timestamp 1662439860
transform -1 0 82800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__CLK
timestamp 1662439860
transform 1 0 90896 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__CLK
timestamp 1662439860
transform 1 0 84824 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__CLK
timestamp 1662439860
transform 1 0 93380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__CLK
timestamp 1662439860
transform 1 0 74980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__RESET_B
timestamp 1662439860
transform 1 0 68356 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__RESET_B
timestamp 1662439860
transform -1 0 66148 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__CLK
timestamp 1662439860
transform 1 0 82064 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__RESET_B
timestamp 1662439860
transform -1 0 68540 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__CLK
timestamp 1662439860
transform 1 0 72772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__CLK
timestamp 1662439860
transform 1 0 80592 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__CLK
timestamp 1662439860
transform -1 0 80684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__CLK
timestamp 1662439860
transform 1 0 94116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__CLK
timestamp 1662439860
transform -1 0 91080 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__CLK
timestamp 1662439860
transform -1 0 94392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__CLK
timestamp 1662439860
transform 1 0 83352 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__CLK
timestamp 1662439860
transform -1 0 58788 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__CLK
timestamp 1662439860
transform -1 0 69368 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__CLK
timestamp 1662439860
transform -1 0 91448 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__CLK
timestamp 1662439860
transform -1 0 90804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__CLK
timestamp 1662439860
transform -1 0 62652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__CLK
timestamp 1662439860
transform -1 0 78476 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__CLK
timestamp 1662439860
transform -1 0 80500 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__CLK
timestamp 1662439860
transform -1 0 66516 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__CLK
timestamp 1662439860
transform -1 0 89332 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__CLK
timestamp 1662439860
transform -1 0 78844 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__CLK
timestamp 1662439860
transform -1 0 85928 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__CLK
timestamp 1662439860
transform -1 0 92000 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__CLK
timestamp 1662439860
transform -1 0 92276 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__RESET_B
timestamp 1662439860
transform 1 0 93196 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__CLK
timestamp 1662439860
transform 1 0 64308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__D
timestamp 1662439860
transform 1 0 65780 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__CLK
timestamp 1662439860
transform 1 0 53728 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__RESET_B
timestamp 1662439860
transform -1 0 51888 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__CLK
timestamp 1662439860
transform -1 0 58604 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__RESET_B
timestamp 1662439860
transform -1 0 55660 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__CLK
timestamp 1662439860
transform 1 0 65412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__CLK
timestamp 1662439860
transform -1 0 86572 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__RESET_B
timestamp 1662439860
transform 1 0 83168 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__CLK
timestamp 1662439860
transform 1 0 67620 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__D
timestamp 1662439860
transform 1 0 68540 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__RESET_B
timestamp 1662439860
transform 1 0 65780 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__CLK
timestamp 1662439860
transform 1 0 63756 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__RESET_B
timestamp 1662439860
transform 1 0 63204 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__CLK
timestamp 1662439860
transform 1 0 64860 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__RESET_B
timestamp 1662439860
transform 1 0 64308 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__RESET_B
timestamp 1662439860
transform 1 0 91540 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__RESET_B
timestamp 1662439860
transform 1 0 79580 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__D
timestamp 1662439860
transform -1 0 22632 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__RESET_B
timestamp 1662439860
transform 1 0 68540 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__CLK
timestamp 1662439860
transform 1 0 10304 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__CLK
timestamp 1662439860
transform 1 0 6256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__CLK
timestamp 1662439860
transform 1 0 6532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__CLK
timestamp 1662439860
transform 1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__D
timestamp 1662439860
transform -1 0 36984 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__CLK
timestamp 1662439860
transform 1 0 66884 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__CLK
timestamp 1662439860
transform 1 0 69184 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__CLK
timestamp 1662439860
transform 1 0 67068 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__CLK
timestamp 1662439860
transform 1 0 74704 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__CLK
timestamp 1662439860
transform 1 0 67436 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__CLK
timestamp 1662439860
transform -1 0 77740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__CLK
timestamp 1662439860
transform 1 0 66516 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__CLK
timestamp 1662439860
transform -1 0 80316 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__CLK
timestamp 1662439860
transform -1 0 73232 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__CLK
timestamp 1662439860
transform 1 0 74888 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__CLK
timestamp 1662439860
transform -1 0 68172 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__CLK
timestamp 1662439860
transform -1 0 63388 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__CLK
timestamp 1662439860
transform -1 0 54464 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__D
timestamp 1662439860
transform -1 0 20424 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__RESET_B
timestamp 1662439860
transform 1 0 29072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__D
timestamp 1662439860
transform -1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__RESET_B
timestamp 1662439860
transform 1 0 32292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__RESET_B
timestamp 1662439860
transform 1 0 25208 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__RESET_B
timestamp 1662439860
transform 1 0 29348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__SET_B
timestamp 1662439860
transform 1 0 30452 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__RESET_B
timestamp 1662439860
transform 1 0 29900 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__CLK
timestamp 1662439860
transform 1 0 63756 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__D
timestamp 1662439860
transform -1 0 59432 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__CLK
timestamp 1662439860
transform 1 0 64308 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__CLK
timestamp 1662439860
transform -1 0 55016 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__CLK
timestamp 1662439860
transform -1 0 53268 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__CLK
timestamp 1662439860
transform -1 0 54280 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__CLK
timestamp 1662439860
transform -1 0 57500 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__CLK
timestamp 1662439860
transform 1 0 63756 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__CLK
timestamp 1662439860
transform 1 0 55476 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__CLK
timestamp 1662439860
transform -1 0 31740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__CLK
timestamp 1662439860
transform 1 0 36800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__CLK
timestamp 1662439860
transform 1 0 29808 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__RESET_B
timestamp 1662439860
transform 1 0 40020 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__D
timestamp 1662439860
transform -1 0 39928 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__RESET_B
timestamp 1662439860
transform -1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__RESET_B
timestamp 1662439860
transform 1 0 39652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__RESET_B
timestamp 1662439860
transform 1 0 40204 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__CLK
timestamp 1662439860
transform 1 0 37444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__RESET_B
timestamp 1662439860
transform 1 0 34224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__CLK
timestamp 1662439860
transform 1 0 49496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__D
timestamp 1662439860
transform 1 0 48760 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__RESET_B
timestamp 1662439860
transform 1 0 50600 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__CLK
timestamp 1662439860
transform 1 0 55936 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__D
timestamp 1662439860
transform -1 0 56672 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__RESET_B
timestamp 1662439860
transform 1 0 57040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__CLK
timestamp 1662439860
transform -1 0 61916 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__RESET_B
timestamp 1662439860
transform 1 0 64308 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__RESET_B
timestamp 1662439860
transform 1 0 63204 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1357__A
timestamp 1662439860
transform -1 0 77188 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__A
timestamp 1662439860
transform -1 0 69828 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__A
timestamp 1662439860
transform 1 0 68540 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__A
timestamp 1662439860
transform -1 0 52624 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__A
timestamp 1662439860
transform -1 0 93380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__A
timestamp 1662439860
transform 1 0 92644 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__A
timestamp 1662439860
transform -1 0 93288 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__A
timestamp 1662439860
transform -1 0 92644 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0__0306__A
timestamp 1662439860
transform -1 0 42872 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_master_A
timestamp 1662439860
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout31_A
timestamp 1662439860
transform 1 0 64860 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout32_A
timestamp 1662439860
transform 1 0 76452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout33_A
timestamp 1662439860
transform -1 0 94024 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout37_A
timestamp 1662439860
transform -1 0 82524 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout39_A
timestamp 1662439860
transform 1 0 86204 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout40_A
timestamp 1662439860
transform -1 0 89332 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout42_A
timestamp 1662439860
transform 1 0 2024 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout43_A
timestamp 1662439860
transform 1 0 5520 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout45_A
timestamp 1662439860
transform -1 0 17572 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout47_A
timestamp 1662439860
transform -1 0 24840 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout48_A
timestamp 1662439860
transform 1 0 32476 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout49_A
timestamp 1662439860
transform 1 0 27692 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout50_A
timestamp 1662439860
transform -1 0 36432 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout51_A
timestamp 1662439860
transform 1 0 4968 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout52_A
timestamp 1662439860
transform -1 0 62100 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout53_A
timestamp 1662439860
transform -1 0 62468 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout54_A
timestamp 1662439860
transform 1 0 50324 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout55_A
timestamp 1662439860
transform 1 0 76912 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout58_A
timestamp 1662439860
transform -1 0 83352 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout59_A
timestamp 1662439860
transform -1 0 75440 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1662439860
transform -1 0 43700 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1662439860
transform -1 0 92368 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1662439860
transform -1 0 43700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1662439860
transform -1 0 93012 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1662439860
transform -1 0 35788 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1662439860
transform -1 0 83260 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1662439860
transform -1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1662439860
transform -1 0 83352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1662439860
transform -1 0 1748 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1662439860
transform -1 0 1748 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output22_A
timestamp 1662439860
transform -1 0 58880 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output24_A
timestamp 1662439860
transform 1 0 61364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 8280 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 9108 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 9936 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
timestamp 1662439860
transform -1 0 7820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_A
timestamp 1662439860
transform 1 0 44344 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 4232 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 5428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_A
timestamp 1662439860
transform -1 0 33764 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
timestamp 1662439860
transform -1 0 1840 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_A
timestamp 1662439860
transform -1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
timestamp 1662439860
transform -1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
timestamp 1662439860
transform -1 0 1840 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 1748 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_A
timestamp 1662439860
transform -1 0 31832 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 9752 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
timestamp 1662439860
transform -1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf_A
timestamp 1662439860
transform -1 0 54188 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf_TE_B
timestamp 1662439860
transform -1 0 52992 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 11132 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_A
timestamp 1662439860
transform -1 0 60076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 6624 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_A
timestamp 1662439860
transform -1 0 58144 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_TE_B
timestamp 1662439860
transform -1 0 58972 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 10764 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_A
timestamp 1662439860
transform -1 0 60812 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 9476 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_A
timestamp 1662439860
transform -1 0 58512 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_A
timestamp 1662439860
transform -1 0 59064 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_TE_B
timestamp 1662439860
transform -1 0 60168 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 11684 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_TE_B
timestamp 1662439860
transform -1 0 48852 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 15916 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_A
timestamp 1662439860
transform 1 0 49680 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 13340 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.ro_block_I.ro_pol.tribuf.t_buf_TE_B
timestamp 1662439860
transform -1 0 77096 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.ro_block_I.ro_pol_eve.tribuf.t_buf_TE_B
timestamp 1662439860
transform -1 0 83996 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 88964 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
timestamp 1662439860
transform -1 0 94300 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 91264 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 88964 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 91172 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 93656 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
timestamp 1662439860
transform -1 0 88596 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 89516 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_GATE_N
timestamp 1662439860
transform -1 0 90804 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_A
timestamp 1662439860
transform -1 0 94116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 85376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_GATE_N
timestamp 1662439860
transform 1 0 90068 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
timestamp 1662439860
transform -1 0 92736 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
timestamp 1662439860
transform -1 0 86756 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
timestamp 1662439860
transform -1 0 87308 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 90068 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_A
timestamp 1662439860
transform -1 0 83076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 87860 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 85284 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_A
timestamp 1662439860
transform 1 0 58512 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
timestamp 1662439860
transform -1 0 92092 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 82616 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_GATE_N
timestamp 1662439860
transform -1 0 82708 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_A
timestamp 1662439860
transform -1 0 91080 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
timestamp 1662439860
transform -1 0 81696 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_GATE_N
timestamp 1662439860
transform -1 0 83260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_A
timestamp 1662439860
transform -1 0 75532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_TE_B
timestamp 1662439860
transform -1 0 77372 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 83904 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_GATE_N
timestamp 1662439860
transform -1 0 84824 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_TE_B
timestamp 1662439860
transform -1 0 47380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
timestamp 1662439860
transform 1 0 83444 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_GATE_N
timestamp 1662439860
transform 1 0 82984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.ro_block_I.ro_pol.tribuf.t_buf_TE_B
timestamp 1662439860
transform -1 0 65228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.ro_block_Q.ro_pol.tribuf.t_buf_TE_B
timestamp 1662439860
transform -1 0 53084 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf_TE_B
timestamp 1662439860
transform -1 0 54556 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1662439860
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1662439860
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1662439860
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1662439860
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1662439860
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1662439860
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1662439860
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1662439860
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1662439860
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_121 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 12236 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_127 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 12788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1662439860
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1662439860
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1662439860
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1662439860
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1662439860
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1662439860
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1662439860
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1662439860
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_210
timestamp 1662439860
transform 1 0 20424 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1662439860
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1662439860
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1662439860
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1662439860
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1662439860
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1662439860
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1662439860
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1662439860
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1662439860
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_293
timestamp 1662439860
transform 1 0 28060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_298
timestamp 1662439860
transform 1 0 28520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1662439860
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1662439860
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1662439860
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1662439860
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1662439860
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1662439860
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1662439860
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1662439860
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1662439860
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_384
timestamp 1662439860
transform 1 0 36432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1662439860
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1662439860
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_405
timestamp 1662439860
transform 1 0 38364 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_413
timestamp 1662439860
transform 1 0 39100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1662439860
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1662439860
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1662439860
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1662439860
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1662439860
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_463
timestamp 1662439860
transform 1 0 43700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_470
timestamp 1662439860
transform 1 0 44344 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1662439860
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1662439860
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1662439860
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1662439860
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_517
timestamp 1662439860
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1662439860
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1662439860
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_545
timestamp 1662439860
transform 1 0 51244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1662439860
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_561
timestamp 1662439860
transform 1 0 52716 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_567
timestamp 1662439860
transform 1 0 53268 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_571
timestamp 1662439860
transform 1 0 53636 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_581
timestamp 1662439860
transform 1 0 54556 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_587
timestamp 1662439860
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1662439860
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_601
timestamp 1662439860
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1662439860
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_617
timestamp 1662439860
transform 1 0 57868 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_629
timestamp 1662439860
transform 1 0 58972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 1662439860
transform 1 0 60076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_645
timestamp 1662439860
transform 1 0 60444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_651
timestamp 1662439860
transform 1 0 60996 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_657
timestamp 1662439860
transform 1 0 61548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1662439860
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_673
timestamp 1662439860
transform 1 0 63020 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_685
timestamp 1662439860
transform 1 0 64124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_689
timestamp 1662439860
transform 1 0 64492 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1662439860
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1662439860
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_713
timestamp 1662439860
transform 1 0 66700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1662439860
transform 1 0 67804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_729
timestamp 1662439860
transform 1 0 68172 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_735
timestamp 1662439860
transform 1 0 68724 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_747
timestamp 1662439860
transform 1 0 69828 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_755
timestamp 1662439860
transform 1 0 70564 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_757
timestamp 1662439860
transform 1 0 70748 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_769
timestamp 1662439860
transform 1 0 71852 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 1662439860
transform 1 0 72956 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_785
timestamp 1662439860
transform 1 0 73324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_797
timestamp 1662439860
transform 1 0 74428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_808
timestamp 1662439860
transform 1 0 75440 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_813
timestamp 1662439860
transform 1 0 75900 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_819
timestamp 1662439860
transform 1 0 76452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_831
timestamp 1662439860
transform 1 0 77556 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_839
timestamp 1662439860
transform 1 0 78292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_841
timestamp 1662439860
transform 1 0 78476 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_845
timestamp 1662439860
transform 1 0 78844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_857
timestamp 1662439860
transform 1 0 79948 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_865
timestamp 1662439860
transform 1 0 80684 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_869
timestamp 1662439860
transform 1 0 81052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_881
timestamp 1662439860
transform 1 0 82156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_889
timestamp 1662439860
transform 1 0 82892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_894
timestamp 1662439860
transform 1 0 83352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_897
timestamp 1662439860
transform 1 0 83628 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_903
timestamp 1662439860
transform 1 0 84180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_915
timestamp 1662439860
transform 1 0 85284 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_923
timestamp 1662439860
transform 1 0 86020 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_925
timestamp 1662439860
transform 1 0 86204 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_933
timestamp 1662439860
transform 1 0 86940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_945
timestamp 1662439860
transform 1 0 88044 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_951
timestamp 1662439860
transform 1 0 88596 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_953
timestamp 1662439860
transform 1 0 88780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_965
timestamp 1662439860
transform 1 0 89884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_973
timestamp 1662439860
transform 1 0 90620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_978
timestamp 1662439860
transform 1 0 91080 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_981
timestamp 1662439860
transform 1 0 91356 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_993
timestamp 1662439860
transform 1 0 92460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_999
timestamp 1662439860
transform 1 0 93012 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1007
timestamp 1662439860
transform 1 0 93748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1009
timestamp 1662439860
transform 1 0 93932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1015
timestamp 1662439860
transform 1 0 94484 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1662439860
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1662439860
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1662439860
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1662439860
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1662439860
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1662439860
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1662439860
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1662439860
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1662439860
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1662439860
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1662439860
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1662439860
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1662439860
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1662439860
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1662439860
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1662439860
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1662439860
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1662439860
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1662439860
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1662439860
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1662439860
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1662439860
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1662439860
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1662439860
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1662439860
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1662439860
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1662439860
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1662439860
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1662439860
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1662439860
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1662439860
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1662439860
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1662439860
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1662439860
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1662439860
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1662439860
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1662439860
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1662439860
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1662439860
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1662439860
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1662439860
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1662439860
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_393
timestamp 1662439860
transform 1 0 37260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_416
timestamp 1662439860
transform 1 0 39376 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_422
timestamp 1662439860
transform 1 0 39928 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_434
timestamp 1662439860
transform 1 0 41032 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1662439860
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1662439860
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1662439860
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1662439860
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1662439860
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1662439860
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1662439860
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1662439860
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1662439860
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1662439860
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_541
timestamp 1662439860
transform 1 0 50876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_546
timestamp 1662439860
transform 1 0 51336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_552
timestamp 1662439860
transform 1 0 51888 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1662439860
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_565
timestamp 1662439860
transform 1 0 53084 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_571
timestamp 1662439860
transform 1 0 53636 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_574
timestamp 1662439860
transform 1 0 53912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_580
timestamp 1662439860
transform 1 0 54464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_586
timestamp 1662439860
transform 1 0 55016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_590
timestamp 1662439860
transform 1 0 55384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_593
timestamp 1662439860
transform 1 0 55660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_601
timestamp 1662439860
transform 1 0 56396 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_611
timestamp 1662439860
transform 1 0 57316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1662439860
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1662439860
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1662439860
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1662439860
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_655
timestamp 1662439860
transform 1 0 61364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_667
timestamp 1662439860
transform 1 0 62468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1662439860
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_673
timestamp 1662439860
transform 1 0 63020 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_695
timestamp 1662439860
transform 1 0 65044 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_701
timestamp 1662439860
transform 1 0 65596 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_713
timestamp 1662439860
transform 1 0 66700 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_725
timestamp 1662439860
transform 1 0 67804 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1662439860
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1662439860
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1662439860
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1662439860
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 1662439860
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1662439860
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1662439860
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1662439860
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_809
timestamp 1662439860
transform 1 0 75532 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_819
timestamp 1662439860
transform 1 0 76452 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_827
timestamp 1662439860
transform 1 0 77188 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_831
timestamp 1662439860
transform 1 0 77556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_837
timestamp 1662439860
transform 1 0 78108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_841
timestamp 1662439860
transform 1 0 78476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_850
timestamp 1662439860
transform 1 0 79304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_857
timestamp 1662439860
transform 1 0 79948 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_865
timestamp 1662439860
transform 1 0 80684 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_873
timestamp 1662439860
transform 1 0 81420 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_876
timestamp 1662439860
transform 1 0 81696 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_884
timestamp 1662439860
transform 1 0 82432 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_887
timestamp 1662439860
transform 1 0 82708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_893
timestamp 1662439860
transform 1 0 83260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_897
timestamp 1662439860
transform 1 0 83628 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_905
timestamp 1662439860
transform 1 0 84364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_910
timestamp 1662439860
transform 1 0 84824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_916
timestamp 1662439860
transform 1 0 85376 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_924
timestamp 1662439860
transform 1 0 86112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_928
timestamp 1662439860
transform 1 0 86480 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_931
timestamp 1662439860
transform 1 0 86756 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_937
timestamp 1662439860
transform 1 0 87308 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_949
timestamp 1662439860
transform 1 0 88412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_953
timestamp 1662439860
transform 1 0 88780 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_961
timestamp 1662439860
transform 1 0 89516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_966
timestamp 1662439860
transform 1 0 89976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_972
timestamp 1662439860
transform 1 0 90528 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_978
timestamp 1662439860
transform 1 0 91080 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_986
timestamp 1662439860
transform 1 0 91816 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_989
timestamp 1662439860
transform 1 0 92092 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_995
timestamp 1662439860
transform 1 0 92644 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1662439860
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1009
timestamp 1662439860
transform 1 0 93932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1015
timestamp 1662439860
transform 1 0 94484 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1662439860
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1662439860
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1662439860
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1662439860
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1662439860
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1662439860
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1662439860
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1662439860
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1662439860
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1662439860
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1662439860
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1662439860
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1662439860
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1662439860
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1662439860
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1662439860
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_157
timestamp 1662439860
transform 1 0 15548 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_163
timestamp 1662439860
transform 1 0 16100 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_175
timestamp 1662439860
transform 1 0 17204 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1662439860
transform 1 0 18308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1662439860
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1662439860
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1662439860
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1662439860
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1662439860
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1662439860
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1662439860
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1662439860
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1662439860
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1662439860
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1662439860
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1662439860
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1662439860
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1662439860
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1662439860
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1662439860
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1662439860
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1662439860
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1662439860
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1662439860
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1662439860
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_389
timestamp 1662439860
transform 1 0 36892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_395
timestamp 1662439860
transform 1 0 37444 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_417
timestamp 1662439860
transform 1 0 39468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1662439860
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_425
timestamp 1662439860
transform 1 0 40204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_437
timestamp 1662439860
transform 1 0 41308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_449
timestamp 1662439860
transform 1 0 42412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_461
timestamp 1662439860
transform 1 0 43516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_473
timestamp 1662439860
transform 1 0 44620 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1662439860
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1662439860
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1662439860
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1662439860
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1662439860
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1662439860
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_533
timestamp 1662439860
transform 1 0 50140 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_541
timestamp 1662439860
transform 1 0 50876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_544
timestamp 1662439860
transform 1 0 51152 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_572
timestamp 1662439860
transform 1 0 53728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_578
timestamp 1662439860
transform 1 0 54280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_584
timestamp 1662439860
transform 1 0 54832 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_589
timestamp 1662439860
transform 1 0 55292 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_613
timestamp 1662439860
transform 1 0 57500 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_619
timestamp 1662439860
transform 1 0 58052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_625
timestamp 1662439860
transform 1 0 58604 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_633
timestamp 1662439860
transform 1 0 59340 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_641
timestamp 1662439860
transform 1 0 60076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_645
timestamp 1662439860
transform 1 0 60444 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_649
timestamp 1662439860
transform 1 0 60812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_655
timestamp 1662439860
transform 1 0 61364 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_658
timestamp 1662439860
transform 1 0 61640 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_685
timestamp 1662439860
transform 1 0 64124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_691
timestamp 1662439860
transform 1 0 64676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_697
timestamp 1662439860
transform 1 0 65228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_701
timestamp 1662439860
transform 1 0 65596 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_705
timestamp 1662439860
transform 1 0 65964 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_717
timestamp 1662439860
transform 1 0 67068 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_725
timestamp 1662439860
transform 1 0 67804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_729
timestamp 1662439860
transform 1 0 68172 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_735
timestamp 1662439860
transform 1 0 68724 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_747
timestamp 1662439860
transform 1 0 69828 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1662439860
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_757
timestamp 1662439860
transform 1 0 70748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_763
timestamp 1662439860
transform 1 0 71300 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_766
timestamp 1662439860
transform 1 0 71576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_774
timestamp 1662439860
transform 1 0 72312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_778
timestamp 1662439860
transform 1 0 72680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_781
timestamp 1662439860
transform 1 0 72956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_787
timestamp 1662439860
transform 1 0 73508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_791
timestamp 1662439860
transform 1 0 73876 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_794
timestamp 1662439860
transform 1 0 74152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_806
timestamp 1662439860
transform 1 0 75256 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_813
timestamp 1662439860
transform 1 0 75900 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_817
timestamp 1662439860
transform 1 0 76268 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_825
timestamp 1662439860
transform 1 0 77004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_833
timestamp 1662439860
transform 1 0 77740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_854
timestamp 1662439860
transform 1 0 79672 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_860
timestamp 1662439860
transform 1 0 80224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_866
timestamp 1662439860
transform 1 0 80776 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_869
timestamp 1662439860
transform 1 0 81052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_875
timestamp 1662439860
transform 1 0 81604 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_890
timestamp 1662439860
transform 1 0 82984 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_896
timestamp 1662439860
transform 1 0 83536 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_902
timestamp 1662439860
transform 1 0 84088 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_908
timestamp 1662439860
transform 1 0 84640 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_911
timestamp 1662439860
transform 1 0 84916 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 1662439860
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1662439860
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_925
timestamp 1662439860
transform 1 0 86204 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_929
timestamp 1662439860
transform 1 0 86572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_939
timestamp 1662439860
transform 1 0 87492 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_945
timestamp 1662439860
transform 1 0 88044 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_951
timestamp 1662439860
transform 1 0 88596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_955
timestamp 1662439860
transform 1 0 88964 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_976
timestamp 1662439860
transform 1 0 90896 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_981
timestamp 1662439860
transform 1 0 91356 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_990
timestamp 1662439860
transform 1 0 92184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_996
timestamp 1662439860
transform 1 0 92736 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1002
timestamp 1662439860
transform 1 0 93288 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1014
timestamp 1662439860
transform 1 0 94392 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1662439860
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1662439860
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1662439860
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1662439860
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1662439860
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1662439860
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1662439860
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1662439860
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_81
timestamp 1662439860
transform 1 0 8556 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_89
timestamp 1662439860
transform 1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1662439860
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1662439860
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_117
timestamp 1662439860
transform 1 0 11868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_129
timestamp 1662439860
transform 1 0 12972 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_150
timestamp 1662439860
transform 1 0 14904 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 1662439860
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1662439860
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1662439860
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1662439860
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1662439860
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1662439860
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1662439860
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1662439860
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_239
timestamp 1662439860
transform 1 0 23092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_251
timestamp 1662439860
transform 1 0 24196 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_263
timestamp 1662439860
transform 1 0 25300 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_266
timestamp 1662439860
transform 1 0 25576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_275
timestamp 1662439860
transform 1 0 26404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1662439860
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1662439860
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1662439860
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1662439860
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1662439860
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1662439860
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1662439860
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1662439860
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_354
timestamp 1662439860
transform 1 0 33672 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_365
timestamp 1662439860
transform 1 0 34684 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_377
timestamp 1662439860
transform 1 0 35788 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_385
timestamp 1662439860
transform 1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_390
timestamp 1662439860
transform 1 0 36984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1662439860
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_415
timestamp 1662439860
transform 1 0 39284 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_421
timestamp 1662439860
transform 1 0 39836 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_427
timestamp 1662439860
transform 1 0 40388 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_433
timestamp 1662439860
transform 1 0 40940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_439
timestamp 1662439860
transform 1 0 41492 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1662439860
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_449
timestamp 1662439860
transform 1 0 42412 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_459
timestamp 1662439860
transform 1 0 43332 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_463
timestamp 1662439860
transform 1 0 43700 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_466
timestamp 1662439860
transform 1 0 43976 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_478
timestamp 1662439860
transform 1 0 45080 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_490
timestamp 1662439860
transform 1 0 46184 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1662439860
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1662439860
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_517
timestamp 1662439860
transform 1 0 48668 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_521
timestamp 1662439860
transform 1 0 49036 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_542
timestamp 1662439860
transform 1 0 50968 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_548
timestamp 1662439860
transform 1 0 51520 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_554
timestamp 1662439860
transform 1 0 52072 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_557
timestamp 1662439860
transform 1 0 52348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_561
timestamp 1662439860
transform 1 0 52716 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_567
timestamp 1662439860
transform 1 0 53268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_571
timestamp 1662439860
transform 1 0 53636 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_574
timestamp 1662439860
transform 1 0 53912 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_580
timestamp 1662439860
transform 1 0 54464 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_594
timestamp 1662439860
transform 1 0 55752 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_604
timestamp 1662439860
transform 1 0 56672 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_614
timestamp 1662439860
transform 1 0 57592 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_617
timestamp 1662439860
transform 1 0 57868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_621
timestamp 1662439860
transform 1 0 58236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_627
timestamp 1662439860
transform 1 0 58788 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_653
timestamp 1662439860
transform 1 0 61180 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_663
timestamp 1662439860
transform 1 0 62100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_669
timestamp 1662439860
transform 1 0 62652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_673
timestamp 1662439860
transform 1 0 63020 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_677
timestamp 1662439860
transform 1 0 63388 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_683
timestamp 1662439860
transform 1 0 63940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_689
timestamp 1662439860
transform 1 0 64492 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_695
timestamp 1662439860
transform 1 0 65044 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_701
timestamp 1662439860
transform 1 0 65596 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_707
timestamp 1662439860
transform 1 0 66148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_719
timestamp 1662439860
transform 1 0 67252 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1662439860
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_729
timestamp 1662439860
transform 1 0 68172 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_733
timestamp 1662439860
transform 1 0 68540 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_745
timestamp 1662439860
transform 1 0 69644 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_757
timestamp 1662439860
transform 1 0 70748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_761
timestamp 1662439860
transform 1 0 71116 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_782
timestamp 1662439860
transform 1 0 73048 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_785
timestamp 1662439860
transform 1 0 73324 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_791
timestamp 1662439860
transform 1 0 73876 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_797
timestamp 1662439860
transform 1 0 74428 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_803
timestamp 1662439860
transform 1 0 74980 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_806
timestamp 1662439860
transform 1 0 75256 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_812
timestamp 1662439860
transform 1 0 75808 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_815
timestamp 1662439860
transform 1 0 76084 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_821
timestamp 1662439860
transform 1 0 76636 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_832
timestamp 1662439860
transform 1 0 77648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_838
timestamp 1662439860
transform 1 0 78200 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_841
timestamp 1662439860
transform 1 0 78476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_863
timestamp 1662439860
transform 1 0 80500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_869
timestamp 1662439860
transform 1 0 81052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_875
timestamp 1662439860
transform 1 0 81604 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_879
timestamp 1662439860
transform 1 0 81972 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_882
timestamp 1662439860
transform 1 0 82248 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_888
timestamp 1662439860
transform 1 0 82800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_894
timestamp 1662439860
transform 1 0 83352 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_897
timestamp 1662439860
transform 1 0 83628 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_906
timestamp 1662439860
transform 1 0 84456 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_912
timestamp 1662439860
transform 1 0 85008 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_918
timestamp 1662439860
transform 1 0 85560 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_924
timestamp 1662439860
transform 1 0 86112 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_927
timestamp 1662439860
transform 1 0 86388 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 1662439860
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1662439860
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_953
timestamp 1662439860
transform 1 0 88780 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_957
timestamp 1662439860
transform 1 0 89148 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_965
timestamp 1662439860
transform 1 0 89884 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_970
timestamp 1662439860
transform 1 0 90344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_976
timestamp 1662439860
transform 1 0 90896 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_984
timestamp 1662439860
transform 1 0 91632 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1005
timestamp 1662439860
transform 1 0 93564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1009
timestamp 1662439860
transform 1 0 93932 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1013
timestamp 1662439860
transform 1 0 94300 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1662439860
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1662439860
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1662439860
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1662439860
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1662439860
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_53
timestamp 1662439860
transform 1 0 5980 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1662439860
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1662439860
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_101
timestamp 1662439860
transform 1 0 10396 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_107
timestamp 1662439860
transform 1 0 10948 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_119
timestamp 1662439860
transform 1 0 12052 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_131
timestamp 1662439860
transform 1 0 13156 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1662439860
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1662439860
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_156
timestamp 1662439860
transform 1 0 15456 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_168
timestamp 1662439860
transform 1 0 16560 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_180
timestamp 1662439860
transform 1 0 17664 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1662439860
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1662439860
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1662439860
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_221
timestamp 1662439860
transform 1 0 21436 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_229
timestamp 1662439860
transform 1 0 22172 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_232
timestamp 1662439860
transform 1 0 22448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_238
timestamp 1662439860
transform 1 0 23000 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_244
timestamp 1662439860
transform 1 0 23552 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1662439860
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_253
timestamp 1662439860
transform 1 0 24380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_259
timestamp 1662439860
transform 1 0 24932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_266
timestamp 1662439860
transform 1 0 25576 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_270
timestamp 1662439860
transform 1 0 25944 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_291
timestamp 1662439860
transform 1 0 27876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_303
timestamp 1662439860
transform 1 0 28980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1662439860
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1662439860
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_314
timestamp 1662439860
transform 1 0 29992 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_326
timestamp 1662439860
transform 1 0 31096 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_340
timestamp 1662439860
transform 1 0 32384 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_358
timestamp 1662439860
transform 1 0 34040 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_365
timestamp 1662439860
transform 1 0 34684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_373
timestamp 1662439860
transform 1 0 35420 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_381
timestamp 1662439860
transform 1 0 36156 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_403
timestamp 1662439860
transform 1 0 38180 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1662439860
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1662439860
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_421
timestamp 1662439860
transform 1 0 39836 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_447
timestamp 1662439860
transform 1 0 42228 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_453
timestamp 1662439860
transform 1 0 42780 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_457
timestamp 1662439860
transform 1 0 43148 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_460
timestamp 1662439860
transform 1 0 43424 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_468
timestamp 1662439860
transform 1 0 44160 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_471
timestamp 1662439860
transform 1 0 44436 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1662439860
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_477
timestamp 1662439860
transform 1 0 44988 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_481
timestamp 1662439860
transform 1 0 45356 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_485
timestamp 1662439860
transform 1 0 45724 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_493
timestamp 1662439860
transform 1 0 46460 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_497
timestamp 1662439860
transform 1 0 46828 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_500
timestamp 1662439860
transform 1 0 47104 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_508
timestamp 1662439860
transform 1 0 47840 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_520
timestamp 1662439860
transform 1 0 48944 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_524
timestamp 1662439860
transform 1 0 49312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_530
timestamp 1662439860
transform 1 0 49864 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_533
timestamp 1662439860
transform 1 0 50140 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_537
timestamp 1662439860
transform 1 0 50508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_543
timestamp 1662439860
transform 1 0 51060 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_551
timestamp 1662439860
transform 1 0 51796 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_554
timestamp 1662439860
transform 1 0 52072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_560
timestamp 1662439860
transform 1 0 52624 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_574
timestamp 1662439860
transform 1 0 53912 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_582
timestamp 1662439860
transform 1 0 54648 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_586
timestamp 1662439860
transform 1 0 55016 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_589
timestamp 1662439860
transform 1 0 55292 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_602
timestamp 1662439860
transform 1 0 56488 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_611
timestamp 1662439860
transform 1 0 57316 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_620
timestamp 1662439860
transform 1 0 58144 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_627
timestamp 1662439860
transform 1 0 58788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_633
timestamp 1662439860
transform 1 0 59340 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_639
timestamp 1662439860
transform 1 0 59892 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1662439860
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_645
timestamp 1662439860
transform 1 0 60444 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_649
timestamp 1662439860
transform 1 0 60812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_655
timestamp 1662439860
transform 1 0 61364 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_661
timestamp 1662439860
transform 1 0 61916 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_667
timestamp 1662439860
transform 1 0 62468 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_673
timestamp 1662439860
transform 1 0 63020 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_679
timestamp 1662439860
transform 1 0 63572 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_685
timestamp 1662439860
transform 1 0 64124 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_691
timestamp 1662439860
transform 1 0 64676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_697
timestamp 1662439860
transform 1 0 65228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_701
timestamp 1662439860
transform 1 0 65596 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_724
timestamp 1662439860
transform 1 0 67712 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1662439860
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1662439860
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_757
timestamp 1662439860
transform 1 0 70748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_761
timestamp 1662439860
transform 1 0 71116 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_769
timestamp 1662439860
transform 1 0 71852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_780
timestamp 1662439860
transform 1 0 72864 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_790
timestamp 1662439860
transform 1 0 73784 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_799
timestamp 1662439860
transform 1 0 74612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1662439860
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1662439860
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_813
timestamp 1662439860
transform 1 0 75900 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_817
timestamp 1662439860
transform 1 0 76268 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_821
timestamp 1662439860
transform 1 0 76636 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_829
timestamp 1662439860
transform 1 0 77372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_837
timestamp 1662439860
transform 1 0 78108 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_844
timestamp 1662439860
transform 1 0 78752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_857
timestamp 1662439860
transform 1 0 79948 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_863
timestamp 1662439860
transform 1 0 80500 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1662439860
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_869
timestamp 1662439860
transform 1 0 81052 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_885
timestamp 1662439860
transform 1 0 82524 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_893
timestamp 1662439860
transform 1 0 83260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_908
timestamp 1662439860
transform 1 0 84640 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_914
timestamp 1662439860
transform 1 0 85192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_918
timestamp 1662439860
transform 1 0 85560 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_922
timestamp 1662439860
transform 1 0 85928 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_925
timestamp 1662439860
transform 1 0 86204 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_945
timestamp 1662439860
transform 1 0 88044 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_956
timestamp 1662439860
transform 1 0 89056 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_965
timestamp 1662439860
transform 1 0 89884 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_971
timestamp 1662439860
transform 1 0 90436 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_978
timestamp 1662439860
transform 1 0 91080 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_981
timestamp 1662439860
transform 1 0 91356 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_985
timestamp 1662439860
transform 1 0 91724 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_993
timestamp 1662439860
transform 1 0 92460 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1002
timestamp 1662439860
transform 1 0 93288 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1008
timestamp 1662439860
transform 1 0 93840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1014
timestamp 1662439860
transform 1 0 94392 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1662439860
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1662439860
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_27
timestamp 1662439860
transform 1 0 3588 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_36
timestamp 1662439860
transform 1 0 4416 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_48
timestamp 1662439860
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1662439860
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_65
timestamp 1662439860
transform 1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1662439860
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1662439860
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1662439860
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1662439860
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_125
timestamp 1662439860
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1662439860
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1662439860
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1662439860
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1662439860
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1662439860
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1662439860
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1662439860
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1662439860
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1662439860
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1662439860
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_229
timestamp 1662439860
transform 1 0 22172 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp 1662439860
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_246
timestamp 1662439860
transform 1 0 23736 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_252
timestamp 1662439860
transform 1 0 24288 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1662439860
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1662439860
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_296
timestamp 1662439860
transform 1 0 28336 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_304
timestamp 1662439860
transform 1 0 29072 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_312
timestamp 1662439860
transform 1 0 29808 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1662439860
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1662439860
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_346
timestamp 1662439860
transform 1 0 32936 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_354
timestamp 1662439860
transform 1 0 33672 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_357
timestamp 1662439860
transform 1 0 33948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_361
timestamp 1662439860
transform 1 0 34316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_364
timestamp 1662439860
transform 1 0 34592 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_376
timestamp 1662439860
transform 1 0 35696 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_384
timestamp 1662439860
transform 1 0 36432 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_390
timestamp 1662439860
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_393
timestamp 1662439860
transform 1 0 37260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_402
timestamp 1662439860
transform 1 0 38088 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_408
timestamp 1662439860
transform 1 0 38640 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_414
timestamp 1662439860
transform 1 0 39192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_420
timestamp 1662439860
transform 1 0 39744 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_426
timestamp 1662439860
transform 1 0 40296 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_434
timestamp 1662439860
transform 1 0 41032 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_440
timestamp 1662439860
transform 1 0 41584 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_446
timestamp 1662439860
transform 1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_449
timestamp 1662439860
transform 1 0 42412 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_458
timestamp 1662439860
transform 1 0 43240 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_487
timestamp 1662439860
transform 1 0 45908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_493
timestamp 1662439860
transform 1 0 46460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_499
timestamp 1662439860
transform 1 0 47012 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1662439860
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_505
timestamp 1662439860
transform 1 0 47564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_516
timestamp 1662439860
transform 1 0 48576 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_522
timestamp 1662439860
transform 1 0 49128 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_528
timestamp 1662439860
transform 1 0 49680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_536
timestamp 1662439860
transform 1 0 50416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_540
timestamp 1662439860
transform 1 0 50784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_545
timestamp 1662439860
transform 1 0 51244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_551
timestamp 1662439860
transform 1 0 51796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_557
timestamp 1662439860
transform 1 0 52348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_561
timestamp 1662439860
transform 1 0 52716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_565
timestamp 1662439860
transform 1 0 53084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_573
timestamp 1662439860
transform 1 0 53820 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_599
timestamp 1662439860
transform 1 0 56212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1662439860
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1662439860
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_617
timestamp 1662439860
transform 1 0 57868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_623
timestamp 1662439860
transform 1 0 58420 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_629
timestamp 1662439860
transform 1 0 58972 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_635
timestamp 1662439860
transform 1 0 59524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_641
timestamp 1662439860
transform 1 0 60076 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_649
timestamp 1662439860
transform 1 0 60812 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_670
timestamp 1662439860
transform 1 0 62744 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_673
timestamp 1662439860
transform 1 0 63020 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_677
timestamp 1662439860
transform 1 0 63388 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_683
timestamp 1662439860
transform 1 0 63940 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_689
timestamp 1662439860
transform 1 0 64492 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_695
timestamp 1662439860
transform 1 0 65044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_701
timestamp 1662439860
transform 1 0 65596 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_711
timestamp 1662439860
transform 1 0 66516 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_717
timestamp 1662439860
transform 1 0 67068 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_725
timestamp 1662439860
transform 1 0 67804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_729
timestamp 1662439860
transform 1 0 68172 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_733
timestamp 1662439860
transform 1 0 68540 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_739
timestamp 1662439860
transform 1 0 69092 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_742
timestamp 1662439860
transform 1 0 69368 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_767
timestamp 1662439860
transform 1 0 71668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_778
timestamp 1662439860
transform 1 0 72680 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_785
timestamp 1662439860
transform 1 0 73324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_790
timestamp 1662439860
transform 1 0 73784 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_797
timestamp 1662439860
transform 1 0 74428 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_810
timestamp 1662439860
transform 1 0 75624 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_817
timestamp 1662439860
transform 1 0 76268 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_824
timestamp 1662439860
transform 1 0 76912 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_830
timestamp 1662439860
transform 1 0 77464 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_835
timestamp 1662439860
transform 1 0 77924 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1662439860
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_841
timestamp 1662439860
transform 1 0 78476 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_854
timestamp 1662439860
transform 1 0 79672 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_860
timestamp 1662439860
transform 1 0 80224 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_864
timestamp 1662439860
transform 1 0 80592 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_886
timestamp 1662439860
transform 1 0 82616 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_892
timestamp 1662439860
transform 1 0 83168 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_897
timestamp 1662439860
transform 1 0 83628 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_901
timestamp 1662439860
transform 1 0 83996 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_909
timestamp 1662439860
transform 1 0 84732 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_927
timestamp 1662439860
transform 1 0 86388 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1662439860
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1662439860
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_953
timestamp 1662439860
transform 1 0 88780 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_957
timestamp 1662439860
transform 1 0 89148 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_963
timestamp 1662439860
transform 1 0 89700 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_969
timestamp 1662439860
transform 1 0 90252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_975
timestamp 1662439860
transform 1 0 90804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_981
timestamp 1662439860
transform 1 0 91356 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1003
timestamp 1662439860
transform 1 0 93380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1662439860
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1009
timestamp 1662439860
transform 1 0 93932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1013
timestamp 1662439860
transform 1 0 94300 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1662439860
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1662439860
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1662439860
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1662439860
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_52
timestamp 1662439860
transform 1 0 5888 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1662439860
transform 1 0 6440 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1662439860
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1662439860
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_90
timestamp 1662439860
transform 1 0 9384 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_96
timestamp 1662439860
transform 1 0 9936 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_102
timestamp 1662439860
transform 1 0 10488 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_108
timestamp 1662439860
transform 1 0 11040 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_111
timestamp 1662439860
transform 1 0 11316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_123
timestamp 1662439860
transform 1 0 12420 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1662439860
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1662439860
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1662439860
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_147
timestamp 1662439860
transform 1 0 14628 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_166
timestamp 1662439860
transform 1 0 16376 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_178
timestamp 1662439860
transform 1 0 17480 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_190
timestamp 1662439860
transform 1 0 18584 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1662439860
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_206
timestamp 1662439860
transform 1 0 20056 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_213
timestamp 1662439860
transform 1 0 20700 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_221
timestamp 1662439860
transform 1 0 21436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_230
timestamp 1662439860
transform 1 0 22264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_240
timestamp 1662439860
transform 1 0 23184 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1662439860
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_253
timestamp 1662439860
transform 1 0 24380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_260
timestamp 1662439860
transform 1 0 25024 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_270
timestamp 1662439860
transform 1 0 25944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_298
timestamp 1662439860
transform 1 0 28520 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1662439860
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_309
timestamp 1662439860
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_337
timestamp 1662439860
transform 1 0 32108 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1662439860
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_365
timestamp 1662439860
transform 1 0 34684 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_371
timestamp 1662439860
transform 1 0 35236 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_374
timestamp 1662439860
transform 1 0 35512 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_380
timestamp 1662439860
transform 1 0 36064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_390
timestamp 1662439860
transform 1 0 36984 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_394
timestamp 1662439860
transform 1 0 37352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_397
timestamp 1662439860
transform 1 0 37628 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_403
timestamp 1662439860
transform 1 0 38180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_409
timestamp 1662439860
transform 1 0 38732 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_412
timestamp 1662439860
transform 1 0 39008 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_418
timestamp 1662439860
transform 1 0 39560 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_421
timestamp 1662439860
transform 1 0 39836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_426
timestamp 1662439860
transform 1 0 40296 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_432
timestamp 1662439860
transform 1 0 40848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_457
timestamp 1662439860
transform 1 0 43148 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_467
timestamp 1662439860
transform 1 0 44068 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_474
timestamp 1662439860
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_477
timestamp 1662439860
transform 1 0 44988 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_481
timestamp 1662439860
transform 1 0 45356 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_487
timestamp 1662439860
transform 1 0 45908 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_490
timestamp 1662439860
transform 1 0 46184 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_496
timestamp 1662439860
transform 1 0 46736 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_500
timestamp 1662439860
transform 1 0 47104 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_503
timestamp 1662439860
transform 1 0 47380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_509
timestamp 1662439860
transform 1 0 47932 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_520
timestamp 1662439860
transform 1 0 48944 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_530
timestamp 1662439860
transform 1 0 49864 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_533
timestamp 1662439860
transform 1 0 50140 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_541
timestamp 1662439860
transform 1 0 50876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_549
timestamp 1662439860
transform 1 0 51612 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_555
timestamp 1662439860
transform 1 0 52164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_561
timestamp 1662439860
transform 1 0 52716 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_564
timestamp 1662439860
transform 1 0 52992 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_570
timestamp 1662439860
transform 1 0 53544 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_576
timestamp 1662439860
transform 1 0 54096 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_582
timestamp 1662439860
transform 1 0 54648 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_589
timestamp 1662439860
transform 1 0 55292 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_598
timestamp 1662439860
transform 1 0 56120 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_602
timestamp 1662439860
transform 1 0 56488 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_609
timestamp 1662439860
transform 1 0 57132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_618
timestamp 1662439860
transform 1 0 57960 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_624
timestamp 1662439860
transform 1 0 58512 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_630
timestamp 1662439860
transform 1 0 59064 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_636
timestamp 1662439860
transform 1 0 59616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_642
timestamp 1662439860
transform 1 0 60168 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_645
timestamp 1662439860
transform 1 0 60444 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_654
timestamp 1662439860
transform 1 0 61272 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_683
timestamp 1662439860
transform 1 0 63940 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_696
timestamp 1662439860
transform 1 0 65136 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_701
timestamp 1662439860
transform 1 0 65596 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_724
timestamp 1662439860
transform 1 0 67712 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_730
timestamp 1662439860
transform 1 0 68264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_736
timestamp 1662439860
transform 1 0 68816 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_742
timestamp 1662439860
transform 1 0 69368 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_748
timestamp 1662439860
transform 1 0 69920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_754
timestamp 1662439860
transform 1 0 70472 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_757
timestamp 1662439860
transform 1 0 70748 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_761
timestamp 1662439860
transform 1 0 71116 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_767
timestamp 1662439860
transform 1 0 71668 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_789
timestamp 1662439860
transform 1 0 73692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_795
timestamp 1662439860
transform 1 0 74244 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_803
timestamp 1662439860
transform 1 0 74980 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_810
timestamp 1662439860
transform 1 0 75624 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_813
timestamp 1662439860
transform 1 0 75900 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_822
timestamp 1662439860
transform 1 0 76728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_832
timestamp 1662439860
transform 1 0 77648 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_840
timestamp 1662439860
transform 1 0 78384 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_848
timestamp 1662439860
transform 1 0 79120 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_866
timestamp 1662439860
transform 1 0 80776 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_869
timestamp 1662439860
transform 1 0 81052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_873
timestamp 1662439860
transform 1 0 81420 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_879
timestamp 1662439860
transform 1 0 81972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_885
timestamp 1662439860
transform 1 0 82524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_891
timestamp 1662439860
transform 1 0 83076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_897
timestamp 1662439860
transform 1 0 83628 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_903
timestamp 1662439860
transform 1 0 84180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_909
timestamp 1662439860
transform 1 0 84732 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_915
timestamp 1662439860
transform 1 0 85284 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_919
timestamp 1662439860
transform 1 0 85652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_922
timestamp 1662439860
transform 1 0 85928 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_925
timestamp 1662439860
transform 1 0 86204 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_945
timestamp 1662439860
transform 1 0 88044 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_963
timestamp 1662439860
transform 1 0 89700 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_969
timestamp 1662439860
transform 1 0 90252 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_975
timestamp 1662439860
transform 1 0 90804 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1662439860
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_981
timestamp 1662439860
transform 1 0 91356 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_997
timestamp 1662439860
transform 1 0 92828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1004
timestamp 1662439860
transform 1 0 93472 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1010
timestamp 1662439860
transform 1 0 94024 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1662439860
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1662439860
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_27
timestamp 1662439860
transform 1 0 3588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_35
timestamp 1662439860
transform 1 0 4324 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_40
timestamp 1662439860
transform 1 0 4784 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1662439860
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1662439860
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_73
timestamp 1662439860
transform 1 0 7820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_91
timestamp 1662439860
transform 1 0 9476 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1662439860
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1662439860
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_117
timestamp 1662439860
transform 1 0 11868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_129
timestamp 1662439860
transform 1 0 12972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_141
timestamp 1662439860
transform 1 0 14076 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_146
timestamp 1662439860
transform 1 0 14536 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_152
timestamp 1662439860
transform 1 0 15088 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1662439860
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1662439860
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_181
timestamp 1662439860
transform 1 0 17756 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_184
timestamp 1662439860
transform 1 0 18032 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_192
timestamp 1662439860
transform 1 0 18768 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_205
timestamp 1662439860
transform 1 0 19964 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_212
timestamp 1662439860
transform 1 0 20608 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_218
timestamp 1662439860
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_225
timestamp 1662439860
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_233
timestamp 1662439860
transform 1 0 22540 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_239
timestamp 1662439860
transform 1 0 23092 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_250
timestamp 1662439860
transform 1 0 24104 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1662439860
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1662439860
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_290
timestamp 1662439860
transform 1 0 27784 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_316
timestamp 1662439860
transform 1 0 30176 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_328
timestamp 1662439860
transform 1 0 31280 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1662439860
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_341
timestamp 1662439860
transform 1 0 32476 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_368
timestamp 1662439860
transform 1 0 34960 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_374
timestamp 1662439860
transform 1 0 35512 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_378
timestamp 1662439860
transform 1 0 35880 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1662439860
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1662439860
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_393
timestamp 1662439860
transform 1 0 37260 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_404
timestamp 1662439860
transform 1 0 38272 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_412
timestamp 1662439860
transform 1 0 39008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_416
timestamp 1662439860
transform 1 0 39376 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_427
timestamp 1662439860
transform 1 0 40388 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_438
timestamp 1662439860
transform 1 0 41400 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_446
timestamp 1662439860
transform 1 0 42136 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_449
timestamp 1662439860
transform 1 0 42412 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_455
timestamp 1662439860
transform 1 0 42964 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_458
timestamp 1662439860
transform 1 0 43240 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_464
timestamp 1662439860
transform 1 0 43792 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_475
timestamp 1662439860
transform 1 0 44804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_486
timestamp 1662439860
transform 1 0 45816 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_493
timestamp 1662439860
transform 1 0 46460 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_499
timestamp 1662439860
transform 1 0 47012 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1662439860
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_505
timestamp 1662439860
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_516
timestamp 1662439860
transform 1 0 48576 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_523
timestamp 1662439860
transform 1 0 49220 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_534
timestamp 1662439860
transform 1 0 50232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_544
timestamp 1662439860
transform 1 0 51152 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_555
timestamp 1662439860
transform 1 0 52164 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1662439860
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_561
timestamp 1662439860
transform 1 0 52716 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_576
timestamp 1662439860
transform 1 0 54096 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_603
timestamp 1662439860
transform 1 0 56580 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_610
timestamp 1662439860
transform 1 0 57224 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_617
timestamp 1662439860
transform 1 0 57868 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_621
timestamp 1662439860
transform 1 0 58236 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_627
timestamp 1662439860
transform 1 0 58788 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_636
timestamp 1662439860
transform 1 0 59616 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_642
timestamp 1662439860
transform 1 0 60168 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_649
timestamp 1662439860
transform 1 0 60812 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_657
timestamp 1662439860
transform 1 0 61548 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1662439860
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1662439860
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_673
timestamp 1662439860
transform 1 0 63020 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_677
timestamp 1662439860
transform 1 0 63388 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_685
timestamp 1662439860
transform 1 0 64124 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_692
timestamp 1662439860
transform 1 0 64768 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_699
timestamp 1662439860
transform 1 0 65412 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_705
timestamp 1662439860
transform 1 0 65964 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_716
timestamp 1662439860
transform 1 0 66976 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_722
timestamp 1662439860
transform 1 0 67528 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_729
timestamp 1662439860
transform 1 0 68172 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_753
timestamp 1662439860
transform 1 0 70380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_761
timestamp 1662439860
transform 1 0 71116 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_768
timestamp 1662439860
transform 1 0 71760 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_779
timestamp 1662439860
transform 1 0 72772 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1662439860
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_785
timestamp 1662439860
transform 1 0 73324 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_790
timestamp 1662439860
transform 1 0 73784 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_802
timestamp 1662439860
transform 1 0 74888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_813
timestamp 1662439860
transform 1 0 75900 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_823
timestamp 1662439860
transform 1 0 76820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_830
timestamp 1662439860
transform 1 0 77464 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_836
timestamp 1662439860
transform 1 0 78016 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_841
timestamp 1662439860
transform 1 0 78476 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_845
timestamp 1662439860
transform 1 0 78844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_851
timestamp 1662439860
transform 1 0 79396 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_880
timestamp 1662439860
transform 1 0 82064 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_886
timestamp 1662439860
transform 1 0 82616 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_894
timestamp 1662439860
transform 1 0 83352 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_897
timestamp 1662439860
transform 1 0 83628 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_903
timestamp 1662439860
transform 1 0 84180 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_923
timestamp 1662439860
transform 1 0 86020 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_941
timestamp 1662439860
transform 1 0 87676 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_949
timestamp 1662439860
transform 1 0 88412 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_953
timestamp 1662439860
transform 1 0 88780 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_976
timestamp 1662439860
transform 1 0 90896 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_982
timestamp 1662439860
transform 1 0 91448 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_988
timestamp 1662439860
transform 1 0 92000 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1003
timestamp 1662439860
transform 1 0 93380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1662439860
transform 1 0 93748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1009
timestamp 1662439860
transform 1 0 93932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_1013
timestamp 1662439860
transform 1 0 94300 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1662439860
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_15
timestamp 1662439860
transform 1 0 2484 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1662439860
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1662439860
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_38
timestamp 1662439860
transform 1 0 4600 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_44
timestamp 1662439860
transform 1 0 5152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_56
timestamp 1662439860
transform 1 0 6256 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_62
timestamp 1662439860
transform 1 0 6808 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1662439860
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1662439860
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_93
timestamp 1662439860
transform 1 0 9660 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_111
timestamp 1662439860
transform 1 0 11316 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_129
timestamp 1662439860
transform 1 0 12972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1662439860
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1662439860
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1662439860
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_150
timestamp 1662439860
transform 1 0 14904 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_156
timestamp 1662439860
transform 1 0 15456 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_170
timestamp 1662439860
transform 1 0 16744 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_182
timestamp 1662439860
transform 1 0 17848 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_188
timestamp 1662439860
transform 1 0 18400 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1662439860
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1662439860
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_201
timestamp 1662439860
transform 1 0 19596 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_211
timestamp 1662439860
transform 1 0 20516 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_217
timestamp 1662439860
transform 1 0 21068 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_223
timestamp 1662439860
transform 1 0 21620 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_229
timestamp 1662439860
transform 1 0 22172 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_239
timestamp 1662439860
transform 1 0 23092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1662439860
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_253
timestamp 1662439860
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_259
timestamp 1662439860
transform 1 0 24932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_286
timestamp 1662439860
transform 1 0 27416 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_294
timestamp 1662439860
transform 1 0 28152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_303
timestamp 1662439860
transform 1 0 28980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1662439860
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_309
timestamp 1662439860
transform 1 0 29532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_315
timestamp 1662439860
transform 1 0 30084 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_342
timestamp 1662439860
transform 1 0 32568 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_353
timestamp 1662439860
transform 1 0 33580 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_357
timestamp 1662439860
transform 1 0 33948 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp 1662439860
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1662439860
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_388
timestamp 1662439860
transform 1 0 36800 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_394
timestamp 1662439860
transform 1 0 37352 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_398
timestamp 1662439860
transform 1 0 37720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_401
timestamp 1662439860
transform 1 0 37996 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_407
timestamp 1662439860
transform 1 0 38548 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_417
timestamp 1662439860
transform 1 0 39468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_421
timestamp 1662439860
transform 1 0 39836 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_429
timestamp 1662439860
transform 1 0 40572 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_436
timestamp 1662439860
transform 1 0 41216 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_442
timestamp 1662439860
transform 1 0 41768 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_445
timestamp 1662439860
transform 1 0 42044 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_456
timestamp 1662439860
transform 1 0 43056 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_466
timestamp 1662439860
transform 1 0 43976 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_474
timestamp 1662439860
transform 1 0 44712 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_477
timestamp 1662439860
transform 1 0 44988 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_483
timestamp 1662439860
transform 1 0 45540 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_487
timestamp 1662439860
transform 1 0 45908 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_509
timestamp 1662439860
transform 1 0 47932 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_519
timestamp 1662439860
transform 1 0 48852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_530
timestamp 1662439860
transform 1 0 49864 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_533
timestamp 1662439860
transform 1 0 50140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_555
timestamp 1662439860
transform 1 0 52164 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_562
timestamp 1662439860
transform 1 0 52808 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_568
timestamp 1662439860
transform 1 0 53360 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_574
timestamp 1662439860
transform 1 0 53912 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_578
timestamp 1662439860
transform 1 0 54280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_583
timestamp 1662439860
transform 1 0 54740 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1662439860
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_589
timestamp 1662439860
transform 1 0 55292 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_608
timestamp 1662439860
transform 1 0 57040 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_614
timestamp 1662439860
transform 1 0 57592 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_620
timestamp 1662439860
transform 1 0 58144 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_626
timestamp 1662439860
transform 1 0 58696 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_634
timestamp 1662439860
transform 1 0 59432 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_641
timestamp 1662439860
transform 1 0 60076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_645
timestamp 1662439860
transform 1 0 60444 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_654
timestamp 1662439860
transform 1 0 61272 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_665
timestamp 1662439860
transform 1 0 62284 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_673
timestamp 1662439860
transform 1 0 63020 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_677
timestamp 1662439860
transform 1 0 63388 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_698
timestamp 1662439860
transform 1 0 65320 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_701
timestamp 1662439860
transform 1 0 65596 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_730
timestamp 1662439860
transform 1 0 68264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_736
timestamp 1662439860
transform 1 0 68816 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_742
timestamp 1662439860
transform 1 0 69368 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_748
timestamp 1662439860
transform 1 0 69920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_754
timestamp 1662439860
transform 1 0 70472 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_757
timestamp 1662439860
transform 1 0 70748 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_784
timestamp 1662439860
transform 1 0 73232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_790
timestamp 1662439860
transform 1 0 73784 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_801
timestamp 1662439860
transform 1 0 74796 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_805
timestamp 1662439860
transform 1 0 75164 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_810
timestamp 1662439860
transform 1 0 75624 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_813
timestamp 1662439860
transform 1 0 75900 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_823
timestamp 1662439860
transform 1 0 76820 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_829
timestamp 1662439860
transform 1 0 77372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_835
timestamp 1662439860
transform 1 0 77924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_841
timestamp 1662439860
transform 1 0 78476 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_847
timestamp 1662439860
transform 1 0 79028 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_853
timestamp 1662439860
transform 1 0 79580 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_866
timestamp 1662439860
transform 1 0 80776 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_869
timestamp 1662439860
transform 1 0 81052 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_876
timestamp 1662439860
transform 1 0 81696 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_880
timestamp 1662439860
transform 1 0 82064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_901
timestamp 1662439860
transform 1 0 83996 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_910
timestamp 1662439860
transform 1 0 84824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_916
timestamp 1662439860
transform 1 0 85376 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_922
timestamp 1662439860
transform 1 0 85928 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_925
timestamp 1662439860
transform 1 0 86204 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_935
timestamp 1662439860
transform 1 0 87124 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_943
timestamp 1662439860
transform 1 0 87860 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_948
timestamp 1662439860
transform 1 0 88320 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_966
timestamp 1662439860
transform 1 0 89976 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_972
timestamp 1662439860
transform 1 0 90528 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_978
timestamp 1662439860
transform 1 0 91080 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_981
timestamp 1662439860
transform 1 0 91356 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_985
timestamp 1662439860
transform 1 0 91724 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_999
timestamp 1662439860
transform 1 0 93012 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1005
timestamp 1662439860
transform 1 0 93564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1011
timestamp 1662439860
transform 1 0 94116 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1015
timestamp 1662439860
transform 1 0 94484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1662439860
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_29
timestamp 1662439860
transform 1 0 3772 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1662439860
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1662439860
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_61
timestamp 1662439860
transform 1 0 6716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_67
timestamp 1662439860
transform 1 0 7268 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_93
timestamp 1662439860
transform 1 0 9660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_101
timestamp 1662439860
transform 1 0 10396 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_107
timestamp 1662439860
transform 1 0 10948 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1662439860
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1662439860
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_117
timestamp 1662439860
transform 1 0 11868 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_138
timestamp 1662439860
transform 1 0 13800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1662439860
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1662439860
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_173
timestamp 1662439860
transform 1 0 17020 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_179
timestamp 1662439860
transform 1 0 17572 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_182
timestamp 1662439860
transform 1 0 17848 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_189
timestamp 1662439860
transform 1 0 18492 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_196
timestamp 1662439860
transform 1 0 19136 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1662439860
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1662439860
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_240
timestamp 1662439860
transform 1 0 23184 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_246
timestamp 1662439860
transform 1 0 23736 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_252
timestamp 1662439860
transform 1 0 24288 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1662439860
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_281
timestamp 1662439860
transform 1 0 26956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_285
timestamp 1662439860
transform 1 0 27324 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_293
timestamp 1662439860
transform 1 0 28060 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_317
timestamp 1662439860
transform 1 0 30268 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_323
timestamp 1662439860
transform 1 0 30820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1662439860
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1662439860
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_341
timestamp 1662439860
transform 1 0 32476 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_368
timestamp 1662439860
transform 1 0 34960 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_372
timestamp 1662439860
transform 1 0 35328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_380
timestamp 1662439860
transform 1 0 36064 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1662439860
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_393
timestamp 1662439860
transform 1 0 37260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_399
timestamp 1662439860
transform 1 0 37812 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_405
timestamp 1662439860
transform 1 0 38364 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_416
timestamp 1662439860
transform 1 0 39376 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_427
timestamp 1662439860
transform 1 0 40388 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_438
timestamp 1662439860
transform 1 0 41400 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_446
timestamp 1662439860
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_449
timestamp 1662439860
transform 1 0 42412 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_458
timestamp 1662439860
transform 1 0 43240 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_466
timestamp 1662439860
transform 1 0 43976 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_469
timestamp 1662439860
transform 1 0 44252 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_475
timestamp 1662439860
transform 1 0 44804 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_478
timestamp 1662439860
transform 1 0 45080 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_484
timestamp 1662439860
transform 1 0 45632 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_490
timestamp 1662439860
transform 1 0 46184 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_496
timestamp 1662439860
transform 1 0 46736 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_502
timestamp 1662439860
transform 1 0 47288 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_505
timestamp 1662439860
transform 1 0 47564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_510
timestamp 1662439860
transform 1 0 48024 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_516
timestamp 1662439860
transform 1 0 48576 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_525
timestamp 1662439860
transform 1 0 49404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_550
timestamp 1662439860
transform 1 0 51704 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_557
timestamp 1662439860
transform 1 0 52348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_561
timestamp 1662439860
transform 1 0 52716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_576
timestamp 1662439860
transform 1 0 54096 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_580
timestamp 1662439860
transform 1 0 54464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_601
timestamp 1662439860
transform 1 0 56396 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_609
timestamp 1662439860
transform 1 0 57132 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_614
timestamp 1662439860
transform 1 0 57592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_617
timestamp 1662439860
transform 1 0 57868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_639
timestamp 1662439860
transform 1 0 59892 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_645
timestamp 1662439860
transform 1 0 60444 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_653
timestamp 1662439860
transform 1 0 61180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_663
timestamp 1662439860
transform 1 0 62100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_670
timestamp 1662439860
transform 1 0 62744 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_673
timestamp 1662439860
transform 1 0 63020 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_683
timestamp 1662439860
transform 1 0 63940 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_693
timestamp 1662439860
transform 1 0 64860 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_699
timestamp 1662439860
transform 1 0 65412 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_706
timestamp 1662439860
transform 1 0 66056 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_715
timestamp 1662439860
transform 1 0 66884 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_726
timestamp 1662439860
transform 1 0 67896 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_729
timestamp 1662439860
transform 1 0 68172 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_738
timestamp 1662439860
transform 1 0 69000 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_749
timestamp 1662439860
transform 1 0 70012 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_755
timestamp 1662439860
transform 1 0 70564 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_782
timestamp 1662439860
transform 1 0 73048 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_785
timestamp 1662439860
transform 1 0 73324 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_789
timestamp 1662439860
transform 1 0 73692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_797
timestamp 1662439860
transform 1 0 74428 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_805
timestamp 1662439860
transform 1 0 75164 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_813
timestamp 1662439860
transform 1 0 75900 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_820
timestamp 1662439860
transform 1 0 76544 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_826
timestamp 1662439860
transform 1 0 77096 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_838
timestamp 1662439860
transform 1 0 78200 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_841
timestamp 1662439860
transform 1 0 78476 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_846
timestamp 1662439860
transform 1 0 78936 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_859
timestamp 1662439860
transform 1 0 80132 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_884
timestamp 1662439860
transform 1 0 82432 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_894
timestamp 1662439860
transform 1 0 83352 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_897
timestamp 1662439860
transform 1 0 83628 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_910
timestamp 1662439860
transform 1 0 84824 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_916
timestamp 1662439860
transform 1 0 85376 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_925
timestamp 1662439860
transform 1 0 86204 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_931
timestamp 1662439860
transform 1 0 86756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_935
timestamp 1662439860
transform 1 0 87124 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_950
timestamp 1662439860
transform 1 0 88504 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_953
timestamp 1662439860
transform 1 0 88780 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_976
timestamp 1662439860
transform 1 0 90896 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_994
timestamp 1662439860
transform 1 0 92552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1002
timestamp 1662439860
transform 1 0 93288 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1009
timestamp 1662439860
transform 1 0 93932 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1013
timestamp 1662439860
transform 1 0 94300 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1662439860
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_15
timestamp 1662439860
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_20
timestamp 1662439860
transform 1 0 2944 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1662439860
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1662439860
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_35
timestamp 1662439860
transform 1 0 4324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_41
timestamp 1662439860
transform 1 0 4876 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_65
timestamp 1662439860
transform 1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_73
timestamp 1662439860
transform 1 0 7820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1662439860
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1662439860
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_101
timestamp 1662439860
transform 1 0 10396 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_109
timestamp 1662439860
transform 1 0 11132 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_132
timestamp 1662439860
transform 1 0 13248 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1662439860
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1662439860
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_163
timestamp 1662439860
transform 1 0 16100 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_173
timestamp 1662439860
transform 1 0 17020 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_179
timestamp 1662439860
transform 1 0 17572 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_185
timestamp 1662439860
transform 1 0 18124 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1662439860
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1662439860
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_208
timestamp 1662439860
transform 1 0 20240 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_219
timestamp 1662439860
transform 1 0 21252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_228
timestamp 1662439860
transform 1 0 22080 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_238
timestamp 1662439860
transform 1 0 23000 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1662439860
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_253
timestamp 1662439860
transform 1 0 24380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_261
timestamp 1662439860
transform 1 0 25116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_284
timestamp 1662439860
transform 1 0 27232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_288
timestamp 1662439860
transform 1 0 27600 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_291
timestamp 1662439860
transform 1 0 27876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_297
timestamp 1662439860
transform 1 0 28428 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_305
timestamp 1662439860
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_309
timestamp 1662439860
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_332
timestamp 1662439860
transform 1 0 31648 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_356
timestamp 1662439860
transform 1 0 33856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1662439860
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_365
timestamp 1662439860
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_388
timestamp 1662439860
transform 1 0 36800 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_394
timestamp 1662439860
transform 1 0 37352 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_400
timestamp 1662439860
transform 1 0 37904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_406
timestamp 1662439860
transform 1 0 38456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_412
timestamp 1662439860
transform 1 0 39008 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_418
timestamp 1662439860
transform 1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_421
timestamp 1662439860
transform 1 0 39836 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_425
timestamp 1662439860
transform 1 0 40204 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_433
timestamp 1662439860
transform 1 0 40940 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_443
timestamp 1662439860
transform 1 0 41860 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_451
timestamp 1662439860
transform 1 0 42596 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_458
timestamp 1662439860
transform 1 0 43240 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_468
timestamp 1662439860
transform 1 0 44160 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_474
timestamp 1662439860
transform 1 0 44712 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_477
timestamp 1662439860
transform 1 0 44988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_487
timestamp 1662439860
transform 1 0 45908 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_493
timestamp 1662439860
transform 1 0 46460 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_501
timestamp 1662439860
transform 1 0 47196 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_514
timestamp 1662439860
transform 1 0 48392 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_524
timestamp 1662439860
transform 1 0 49312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_530
timestamp 1662439860
transform 1 0 49864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_533
timestamp 1662439860
transform 1 0 50140 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_537
timestamp 1662439860
transform 1 0 50508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_541
timestamp 1662439860
transform 1 0 50876 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_548
timestamp 1662439860
transform 1 0 51520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_552
timestamp 1662439860
transform 1 0 51888 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_558
timestamp 1662439860
transform 1 0 52440 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_565
timestamp 1662439860
transform 1 0 53084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_571
timestamp 1662439860
transform 1 0 53636 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_577
timestamp 1662439860
transform 1 0 54188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_586
timestamp 1662439860
transform 1 0 55016 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_589
timestamp 1662439860
transform 1 0 55292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_596
timestamp 1662439860
transform 1 0 55936 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_620
timestamp 1662439860
transform 1 0 58144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_626
timestamp 1662439860
transform 1 0 58696 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_632
timestamp 1662439860
transform 1 0 59248 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_640
timestamp 1662439860
transform 1 0 59984 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_645
timestamp 1662439860
transform 1 0 60444 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_667
timestamp 1662439860
transform 1 0 62468 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_675
timestamp 1662439860
transform 1 0 63204 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_697
timestamp 1662439860
transform 1 0 65228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_701
timestamp 1662439860
transform 1 0 65596 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_710
timestamp 1662439860
transform 1 0 66424 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_716
timestamp 1662439860
transform 1 0 66976 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_740
timestamp 1662439860
transform 1 0 69184 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_747
timestamp 1662439860
transform 1 0 69828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_754
timestamp 1662439860
transform 1 0 70472 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_757
timestamp 1662439860
transform 1 0 70748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_767
timestamp 1662439860
transform 1 0 71668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_778
timestamp 1662439860
transform 1 0 72680 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_803
timestamp 1662439860
transform 1 0 74980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_809
timestamp 1662439860
transform 1 0 75532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_813
timestamp 1662439860
transform 1 0 75900 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_837
timestamp 1662439860
transform 1 0 78108 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_850
timestamp 1662439860
transform 1 0 79304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_854
timestamp 1662439860
transform 1 0 79672 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_858
timestamp 1662439860
transform 1 0 80040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_866
timestamp 1662439860
transform 1 0 80776 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_869
timestamp 1662439860
transform 1 0 81052 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_893
timestamp 1662439860
transform 1 0 83260 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_918
timestamp 1662439860
transform 1 0 85560 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_925
timestamp 1662439860
transform 1 0 86204 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_931
timestamp 1662439860
transform 1 0 86756 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_956
timestamp 1662439860
transform 1 0 89056 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_974
timestamp 1662439860
transform 1 0 90712 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_981
timestamp 1662439860
transform 1 0 91356 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1006
timestamp 1662439860
transform 1 0 93656 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1014
timestamp 1662439860
transform 1 0 94392 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1662439860
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_9
timestamp 1662439860
transform 1 0 1932 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_12
timestamp 1662439860
transform 1 0 2208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_23
timestamp 1662439860
transform 1 0 3220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_29
timestamp 1662439860
transform 1 0 3772 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_40
timestamp 1662439860
transform 1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_47
timestamp 1662439860
transform 1 0 5428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1662439860
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp 1662439860
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_74
timestamp 1662439860
transform 1 0 7912 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_78
timestamp 1662439860
transform 1 0 8280 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_82
timestamp 1662439860
transform 1 0 8648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1662439860
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1662439860
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_138
timestamp 1662439860
transform 1 0 13800 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_153
timestamp 1662439860
transform 1 0 15180 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_159
timestamp 1662439860
transform 1 0 15732 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1662439860
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp 1662439860
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_174
timestamp 1662439860
transform 1 0 17112 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_185
timestamp 1662439860
transform 1 0 18124 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_193
timestamp 1662439860
transform 1 0 18860 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_201
timestamp 1662439860
transform 1 0 19596 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_213
timestamp 1662439860
transform 1 0 20700 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1662439860
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1662439860
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_234
timestamp 1662439860
transform 1 0 22632 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_242
timestamp 1662439860
transform 1 0 23368 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_248
timestamp 1662439860
transform 1 0 23920 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_256
timestamp 1662439860
transform 1 0 24656 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp 1662439860
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1662439860
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_303
timestamp 1662439860
transform 1 0 28980 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_309
timestamp 1662439860
transform 1 0 29532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1662439860
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_337
timestamp 1662439860
transform 1 0 32108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_343
timestamp 1662439860
transform 1 0 32660 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_349
timestamp 1662439860
transform 1 0 33212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_376
timestamp 1662439860
transform 1 0 35696 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_386
timestamp 1662439860
transform 1 0 36616 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1662439860
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_400
timestamp 1662439860
transform 1 0 37904 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_410
timestamp 1662439860
transform 1 0 38824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_416
timestamp 1662439860
transform 1 0 39376 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_422
timestamp 1662439860
transform 1 0 39928 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_433
timestamp 1662439860
transform 1 0 40940 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_446
timestamp 1662439860
transform 1 0 42136 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_449
timestamp 1662439860
transform 1 0 42412 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_458
timestamp 1662439860
transform 1 0 43240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_462
timestamp 1662439860
transform 1 0 43608 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_470
timestamp 1662439860
transform 1 0 44344 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_480
timestamp 1662439860
transform 1 0 45264 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_486
timestamp 1662439860
transform 1 0 45816 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_492
timestamp 1662439860
transform 1 0 46368 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_502
timestamp 1662439860
transform 1 0 47288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_505
timestamp 1662439860
transform 1 0 47564 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_510
timestamp 1662439860
transform 1 0 48024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_514
timestamp 1662439860
transform 1 0 48392 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_521
timestamp 1662439860
transform 1 0 49036 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_525
timestamp 1662439860
transform 1 0 49404 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_533
timestamp 1662439860
transform 1 0 50140 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_537
timestamp 1662439860
transform 1 0 50508 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_558
timestamp 1662439860
transform 1 0 52440 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_561
timestamp 1662439860
transform 1 0 52716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_565
timestamp 1662439860
transform 1 0 53084 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_570
timestamp 1662439860
transform 1 0 53544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_577
timestamp 1662439860
transform 1 0 54188 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_583
timestamp 1662439860
transform 1 0 54740 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_587
timestamp 1662439860
transform 1 0 55108 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_608
timestamp 1662439860
transform 1 0 57040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_614
timestamp 1662439860
transform 1 0 57592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_617
timestamp 1662439860
transform 1 0 57868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_622
timestamp 1662439860
transform 1 0 58328 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_634
timestamp 1662439860
transform 1 0 59432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_659
timestamp 1662439860
transform 1 0 61732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_669
timestamp 1662439860
transform 1 0 62652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_673
timestamp 1662439860
transform 1 0 63020 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_677
timestamp 1662439860
transform 1 0 63388 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_685
timestamp 1662439860
transform 1 0 64124 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_695
timestamp 1662439860
transform 1 0 65044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_701
timestamp 1662439860
transform 1 0 65596 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_705
timestamp 1662439860
transform 1 0 65964 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_726
timestamp 1662439860
transform 1 0 67896 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_729
timestamp 1662439860
transform 1 0 68172 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_735
timestamp 1662439860
transform 1 0 68724 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_757
timestamp 1662439860
transform 1 0 70748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_782
timestamp 1662439860
transform 1 0 73048 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_785
timestamp 1662439860
transform 1 0 73324 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_800
timestamp 1662439860
transform 1 0 74704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_807
timestamp 1662439860
transform 1 0 75348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_832
timestamp 1662439860
transform 1 0 77648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_838
timestamp 1662439860
transform 1 0 78200 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_841
timestamp 1662439860
transform 1 0 78476 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_864
timestamp 1662439860
transform 1 0 80592 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_868
timestamp 1662439860
transform 1 0 80960 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_873
timestamp 1662439860
transform 1 0 81420 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_879
timestamp 1662439860
transform 1 0 81972 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_883
timestamp 1662439860
transform 1 0 82340 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_894
timestamp 1662439860
transform 1 0 83352 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_897
timestamp 1662439860
transform 1 0 83628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_901
timestamp 1662439860
transform 1 0 83996 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_905
timestamp 1662439860
transform 1 0 84364 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_934
timestamp 1662439860
transform 1 0 87032 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_947
timestamp 1662439860
transform 1 0 88228 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_951
timestamp 1662439860
transform 1 0 88596 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_953
timestamp 1662439860
transform 1 0 88780 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_969
timestamp 1662439860
transform 1 0 90252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_980
timestamp 1662439860
transform 1 0 91264 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_984
timestamp 1662439860
transform 1 0 91632 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1006
timestamp 1662439860
transform 1 0 93656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1009
timestamp 1662439860
transform 1 0 93932 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_1013
timestamp 1662439860
transform 1 0 94300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1662439860
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_8
timestamp 1662439860
transform 1 0 1840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1662439860
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1662439860
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_44
timestamp 1662439860
transform 1 0 5152 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_52
timestamp 1662439860
transform 1 0 5888 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_74
timestamp 1662439860
transform 1 0 7912 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1662439860
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1662439860
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_94
timestamp 1662439860
transform 1 0 9752 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_122
timestamp 1662439860
transform 1 0 12328 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_132
timestamp 1662439860
transform 1 0 13248 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1662439860
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1662439860
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 1662439860
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_149
timestamp 1662439860
transform 1 0 14812 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_159
timestamp 1662439860
transform 1 0 15732 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_166
timestamp 1662439860
transform 1 0 16376 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_174
timestamp 1662439860
transform 1 0 17112 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_181
timestamp 1662439860
transform 1 0 17756 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1662439860
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1662439860
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_206
timestamp 1662439860
transform 1 0 20056 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_217
timestamp 1662439860
transform 1 0 21068 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_227
timestamp 1662439860
transform 1 0 21988 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_234
timestamp 1662439860
transform 1 0 22632 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_240
timestamp 1662439860
transform 1 0 23184 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_253
timestamp 1662439860
transform 1 0 24380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_258
timestamp 1662439860
transform 1 0 24840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_264
timestamp 1662439860
transform 1 0 25392 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_291
timestamp 1662439860
transform 1 0 27876 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_302
timestamp 1662439860
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1662439860
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_313
timestamp 1662439860
transform 1 0 29900 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_321
timestamp 1662439860
transform 1 0 30636 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_327
timestamp 1662439860
transform 1 0 31188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_352
timestamp 1662439860
transform 1 0 33488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1662439860
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1662439860
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_388
timestamp 1662439860
transform 1 0 36800 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_399
timestamp 1662439860
transform 1 0 37812 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_406
timestamp 1662439860
transform 1 0 38456 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_417
timestamp 1662439860
transform 1 0 39468 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_421
timestamp 1662439860
transform 1 0 39836 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_427
timestamp 1662439860
transform 1 0 40388 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_431
timestamp 1662439860
transform 1 0 40756 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_437
timestamp 1662439860
transform 1 0 41308 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_440
timestamp 1662439860
transform 1 0 41584 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_465
timestamp 1662439860
transform 1 0 43884 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_474
timestamp 1662439860
transform 1 0 44712 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_477
timestamp 1662439860
transform 1 0 44988 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_486
timestamp 1662439860
transform 1 0 45816 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_496
timestamp 1662439860
transform 1 0 46736 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_502
timestamp 1662439860
transform 1 0 47288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_524
timestamp 1662439860
transform 1 0 49312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_530
timestamp 1662439860
transform 1 0 49864 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_533
timestamp 1662439860
transform 1 0 50140 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_550
timestamp 1662439860
transform 1 0 51704 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_575
timestamp 1662439860
transform 1 0 54004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_582
timestamp 1662439860
transform 1 0 54648 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_589
timestamp 1662439860
transform 1 0 55292 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_595
timestamp 1662439860
transform 1 0 55844 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_617
timestamp 1662439860
transform 1 0 57868 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_623
timestamp 1662439860
transform 1 0 58420 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_627
timestamp 1662439860
transform 1 0 58788 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_631
timestamp 1662439860
transform 1 0 59156 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_642
timestamp 1662439860
transform 1 0 60168 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_645
timestamp 1662439860
transform 1 0 60444 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_668
timestamp 1662439860
transform 1 0 62560 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_687
timestamp 1662439860
transform 1 0 64308 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1662439860
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1662439860
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_701
timestamp 1662439860
transform 1 0 65596 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_726
timestamp 1662439860
transform 1 0 67896 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_751
timestamp 1662439860
transform 1 0 70196 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_755
timestamp 1662439860
transform 1 0 70564 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_757
timestamp 1662439860
transform 1 0 70748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_762
timestamp 1662439860
transform 1 0 71208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_769
timestamp 1662439860
transform 1 0 71852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_786
timestamp 1662439860
transform 1 0 73416 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_810
timestamp 1662439860
transform 1 0 75624 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_813
timestamp 1662439860
transform 1 0 75900 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_819
timestamp 1662439860
transform 1 0 76452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_823
timestamp 1662439860
transform 1 0 76820 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_827
timestamp 1662439860
transform 1 0 77188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_851
timestamp 1662439860
transform 1 0 79396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_858
timestamp 1662439860
transform 1 0 80040 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_862
timestamp 1662439860
transform 1 0 80408 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_866
timestamp 1662439860
transform 1 0 80776 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_869
timestamp 1662439860
transform 1 0 81052 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_892
timestamp 1662439860
transform 1 0 83168 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_900
timestamp 1662439860
transform 1 0 83904 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_922
timestamp 1662439860
transform 1 0 85928 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_925
timestamp 1662439860
transform 1 0 86204 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_940
timestamp 1662439860
transform 1 0 87584 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_965
timestamp 1662439860
transform 1 0 89884 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_971
timestamp 1662439860
transform 1 0 90436 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_978
timestamp 1662439860
transform 1 0 91080 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_981
timestamp 1662439860
transform 1 0 91356 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1004
timestamp 1662439860
transform 1 0 93472 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1011
timestamp 1662439860
transform 1 0 94116 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1015
timestamp 1662439860
transform 1 0 94484 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1662439860
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1662439860
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_12
timestamp 1662439860
transform 1 0 2208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_30
timestamp 1662439860
transform 1 0 3864 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_36
timestamp 1662439860
transform 1 0 4416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1662439860
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1662439860
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_74
timestamp 1662439860
transform 1 0 7912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_92
timestamp 1662439860
transform 1 0 9568 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_98
timestamp 1662439860
transform 1 0 10120 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_104
timestamp 1662439860
transform 1 0 10672 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1662439860
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1662439860
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_119
timestamp 1662439860
transform 1 0 12052 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_129
timestamp 1662439860
transform 1 0 12972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_133
timestamp 1662439860
transform 1 0 13340 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_136
timestamp 1662439860
transform 1 0 13616 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_147
timestamp 1662439860
transform 1 0 14628 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_153
timestamp 1662439860
transform 1 0 15180 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_156
timestamp 1662439860
transform 1 0 15456 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1662439860
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1662439860
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_175
timestamp 1662439860
transform 1 0 17204 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_183
timestamp 1662439860
transform 1 0 17940 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_191
timestamp 1662439860
transform 1 0 18676 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_199
timestamp 1662439860
transform 1 0 19412 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_207
timestamp 1662439860
transform 1 0 20148 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_218
timestamp 1662439860
transform 1 0 21160 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1662439860
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_229
timestamp 1662439860
transform 1 0 22172 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_235
timestamp 1662439860
transform 1 0 22724 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_241
timestamp 1662439860
transform 1 0 23276 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_253
timestamp 1662439860
transform 1 0 24380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1662439860
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1662439860
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_304
timestamp 1662439860
transform 1 0 29072 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_312
timestamp 1662439860
transform 1 0 29808 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1662439860
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_337
timestamp 1662439860
transform 1 0 32108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_342
timestamp 1662439860
transform 1 0 32568 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_367
timestamp 1662439860
transform 1 0 34868 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_371
timestamp 1662439860
transform 1 0 35236 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_377
timestamp 1662439860
transform 1 0 35788 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_384
timestamp 1662439860
transform 1 0 36432 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1662439860
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_393
timestamp 1662439860
transform 1 0 37260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_397
timestamp 1662439860
transform 1 0 37628 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_400
timestamp 1662439860
transform 1 0 37904 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_406
timestamp 1662439860
transform 1 0 38456 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_416
timestamp 1662439860
transform 1 0 39376 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_420
timestamp 1662439860
transform 1 0 39744 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_427
timestamp 1662439860
transform 1 0 40388 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_438
timestamp 1662439860
transform 1 0 41400 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_446
timestamp 1662439860
transform 1 0 42136 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_449
timestamp 1662439860
transform 1 0 42412 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_455
timestamp 1662439860
transform 1 0 42964 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_458
timestamp 1662439860
transform 1 0 43240 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_469
timestamp 1662439860
transform 1 0 44252 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_484
timestamp 1662439860
transform 1 0 45632 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_490
timestamp 1662439860
transform 1 0 46184 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_496
timestamp 1662439860
transform 1 0 46736 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_502
timestamp 1662439860
transform 1 0 47288 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_505
timestamp 1662439860
transform 1 0 47564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_516
timestamp 1662439860
transform 1 0 48576 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_525
timestamp 1662439860
transform 1 0 49404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_550
timestamp 1662439860
transform 1 0 51704 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_558
timestamp 1662439860
transform 1 0 52440 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_561
timestamp 1662439860
transform 1 0 52716 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_568
timestamp 1662439860
transform 1 0 53360 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_574
timestamp 1662439860
transform 1 0 53912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_578
timestamp 1662439860
transform 1 0 54280 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_600
timestamp 1662439860
transform 1 0 56304 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_612
timestamp 1662439860
transform 1 0 57408 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_617
timestamp 1662439860
transform 1 0 57868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_622
timestamp 1662439860
transform 1 0 58328 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_629
timestamp 1662439860
transform 1 0 58972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_633
timestamp 1662439860
transform 1 0 59340 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_655
timestamp 1662439860
transform 1 0 61364 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_662
timestamp 1662439860
transform 1 0 62008 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_669
timestamp 1662439860
transform 1 0 62652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_673
timestamp 1662439860
transform 1 0 63020 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_680
timestamp 1662439860
transform 1 0 63664 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_688
timestamp 1662439860
transform 1 0 64400 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_709
timestamp 1662439860
transform 1 0 66332 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_715
timestamp 1662439860
transform 1 0 66884 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_719
timestamp 1662439860
transform 1 0 67252 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_726
timestamp 1662439860
transform 1 0 67896 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_729
timestamp 1662439860
transform 1 0 68172 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_735
timestamp 1662439860
transform 1 0 68724 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_756
timestamp 1662439860
transform 1 0 70656 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_762
timestamp 1662439860
transform 1 0 71208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_771
timestamp 1662439860
transform 1 0 72036 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_777
timestamp 1662439860
transform 1 0 72588 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_782
timestamp 1662439860
transform 1 0 73048 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_785
timestamp 1662439860
transform 1 0 73324 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_795
timestamp 1662439860
transform 1 0 74244 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_802
timestamp 1662439860
transform 1 0 74888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_809
timestamp 1662439860
transform 1 0 75532 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_816
timestamp 1662439860
transform 1 0 76176 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_820
timestamp 1662439860
transform 1 0 76544 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_827
timestamp 1662439860
transform 1 0 77188 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_833
timestamp 1662439860
transform 1 0 77740 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_838
timestamp 1662439860
transform 1 0 78200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_841
timestamp 1662439860
transform 1 0 78476 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_845
timestamp 1662439860
transform 1 0 78844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_862
timestamp 1662439860
transform 1 0 80408 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_887
timestamp 1662439860
transform 1 0 82708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_894
timestamp 1662439860
transform 1 0 83352 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_897
timestamp 1662439860
transform 1 0 83628 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_912
timestamp 1662439860
transform 1 0 85008 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_916
timestamp 1662439860
transform 1 0 85376 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_937
timestamp 1662439860
transform 1 0 87308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_944
timestamp 1662439860
transform 1 0 87952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_950
timestamp 1662439860
transform 1 0 88504 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_953
timestamp 1662439860
transform 1 0 88780 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_958
timestamp 1662439860
transform 1 0 89240 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_964
timestamp 1662439860
transform 1 0 89792 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_969
timestamp 1662439860
transform 1 0 90252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_993
timestamp 1662439860
transform 1 0 92460 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1003
timestamp 1662439860
transform 1 0 93380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1007
timestamp 1662439860
transform 1 0 93748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1009
timestamp 1662439860
transform 1 0 93932 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1014
timestamp 1662439860
transform 1 0 94392 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1662439860
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_8
timestamp 1662439860
transform 1 0 1840 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1662439860
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1662439860
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_34
timestamp 1662439860
transform 1 0 4232 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_61
timestamp 1662439860
transform 1 0 6716 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1662439860
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1662439860
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1662439860
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_89
timestamp 1662439860
transform 1 0 9292 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1662439860
transform 1 0 9660 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_96
timestamp 1662439860
transform 1 0 9936 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_109
timestamp 1662439860
transform 1 0 11132 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_115
timestamp 1662439860
transform 1 0 11684 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1662439860
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_141
timestamp 1662439860
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_154
timestamp 1662439860
transform 1 0 15272 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_178
timestamp 1662439860
transform 1 0 17480 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1662439860
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1662439860
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_201
timestamp 1662439860
transform 1 0 19596 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_228
timestamp 1662439860
transform 1 0 22080 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_234
timestamp 1662439860
transform 1 0 22632 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_240
timestamp 1662439860
transform 1 0 23184 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1662439860
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_253
timestamp 1662439860
transform 1 0 24380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_260
timestamp 1662439860
transform 1 0 25024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_287
timestamp 1662439860
transform 1 0 27508 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_297
timestamp 1662439860
transform 1 0 28428 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_303
timestamp 1662439860
transform 1 0 28980 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1662439860
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_309
timestamp 1662439860
transform 1 0 29532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_315
timestamp 1662439860
transform 1 0 30084 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_337
timestamp 1662439860
transform 1 0 32108 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 1662439860
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1662439860
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_373
timestamp 1662439860
transform 1 0 35420 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_377
timestamp 1662439860
transform 1 0 35788 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_380
timestamp 1662439860
transform 1 0 36064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_391
timestamp 1662439860
transform 1 0 37076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_399
timestamp 1662439860
transform 1 0 37812 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_410
timestamp 1662439860
transform 1 0 38824 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_418
timestamp 1662439860
transform 1 0 39560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_421
timestamp 1662439860
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_427
timestamp 1662439860
transform 1 0 40388 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_438
timestamp 1662439860
transform 1 0 41400 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_447
timestamp 1662439860
transform 1 0 42228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_455
timestamp 1662439860
transform 1 0 42964 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_465
timestamp 1662439860
transform 1 0 43884 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_474
timestamp 1662439860
transform 1 0 44712 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_477
timestamp 1662439860
transform 1 0 44988 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_487
timestamp 1662439860
transform 1 0 45908 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_494
timestamp 1662439860
transform 1 0 46552 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_505
timestamp 1662439860
transform 1 0 47564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_509
timestamp 1662439860
transform 1 0 47932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1662439860
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_522
timestamp 1662439860
transform 1 0 49128 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_530
timestamp 1662439860
transform 1 0 49864 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_533
timestamp 1662439860
transform 1 0 50140 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_537
timestamp 1662439860
transform 1 0 50508 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_562
timestamp 1662439860
transform 1 0 52808 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_574
timestamp 1662439860
transform 1 0 53912 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1662439860
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1662439860
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_589
timestamp 1662439860
transform 1 0 55292 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_598
timestamp 1662439860
transform 1 0 56120 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_604
timestamp 1662439860
transform 1 0 56672 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_626
timestamp 1662439860
transform 1 0 58696 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1662439860
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1662439860
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_645
timestamp 1662439860
transform 1 0 60444 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_660
timestamp 1662439860
transform 1 0 61824 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_671
timestamp 1662439860
transform 1 0 62836 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_679
timestamp 1662439860
transform 1 0 63572 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_687
timestamp 1662439860
transform 1 0 64308 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_692
timestamp 1662439860
transform 1 0 64768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_698
timestamp 1662439860
transform 1 0 65320 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_701
timestamp 1662439860
transform 1 0 65596 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_716
timestamp 1662439860
transform 1 0 66976 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_722
timestamp 1662439860
transform 1 0 67528 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_730
timestamp 1662439860
transform 1 0 68264 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_754
timestamp 1662439860
transform 1 0 70472 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_757
timestamp 1662439860
transform 1 0 70748 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_779
timestamp 1662439860
transform 1 0 72772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_803
timestamp 1662439860
transform 1 0 74980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_810
timestamp 1662439860
transform 1 0 75624 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_813
timestamp 1662439860
transform 1 0 75900 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_835
timestamp 1662439860
transform 1 0 77924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_842
timestamp 1662439860
transform 1 0 78568 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_849
timestamp 1662439860
transform 1 0 79212 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_853
timestamp 1662439860
transform 1 0 79580 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_861
timestamp 1662439860
transform 1 0 80316 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_867
timestamp 1662439860
transform 1 0 80868 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_869
timestamp 1662439860
transform 1 0 81052 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_874
timestamp 1662439860
transform 1 0 81512 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_880
timestamp 1662439860
transform 1 0 82064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_904
timestamp 1662439860
transform 1 0 84272 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_911
timestamp 1662439860
transform 1 0 84916 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_917
timestamp 1662439860
transform 1 0 85468 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_922
timestamp 1662439860
transform 1 0 85928 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_925
timestamp 1662439860
transform 1 0 86204 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_947
timestamp 1662439860
transform 1 0 88228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_953
timestamp 1662439860
transform 1 0 88780 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_959
timestamp 1662439860
transform 1 0 89332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_963
timestamp 1662439860
transform 1 0 89700 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_967
timestamp 1662439860
transform 1 0 90068 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_975
timestamp 1662439860
transform 1 0 90804 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_979
timestamp 1662439860
transform 1 0 91172 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_981
timestamp 1662439860
transform 1 0 91356 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1003
timestamp 1662439860
transform 1 0 93380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1010
timestamp 1662439860
transform 1 0 94024 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1662439860
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_9
timestamp 1662439860
transform 1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_33
timestamp 1662439860
transform 1 0 4140 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_43
timestamp 1662439860
transform 1 0 5060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1662439860
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1662439860
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1662439860
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_62
timestamp 1662439860
transform 1 0 6808 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_68
timestamp 1662439860
transform 1 0 7360 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_89
timestamp 1662439860
transform 1 0 9292 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_102
timestamp 1662439860
transform 1 0 10488 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1662439860
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1662439860
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_117
timestamp 1662439860
transform 1 0 11868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_122
timestamp 1662439860
transform 1 0 12328 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_146
timestamp 1662439860
transform 1 0 14536 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_150
timestamp 1662439860
transform 1 0 14904 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_156
timestamp 1662439860
transform 1 0 15456 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1662439860
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1662439860
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_178
timestamp 1662439860
transform 1 0 17480 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_187
timestamp 1662439860
transform 1 0 18308 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1662439860
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1662439860
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1662439860
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_247
timestamp 1662439860
transform 1 0 23828 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1662439860
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1662439860
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_285
timestamp 1662439860
transform 1 0 27324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_312
timestamp 1662439860
transform 1 0 29808 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_322
timestamp 1662439860
transform 1 0 30728 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_328
timestamp 1662439860
transform 1 0 31280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1662439860
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_337
timestamp 1662439860
transform 1 0 32108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_347
timestamp 1662439860
transform 1 0 33028 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_353
timestamp 1662439860
transform 1 0 33580 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_375
timestamp 1662439860
transform 1 0 35604 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_381
timestamp 1662439860
transform 1 0 36156 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1662439860
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1662439860
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_397
timestamp 1662439860
transform 1 0 37628 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_403
timestamp 1662439860
transform 1 0 38180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_414
timestamp 1662439860
transform 1 0 39192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_418
timestamp 1662439860
transform 1 0 39560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_440
timestamp 1662439860
transform 1 0 41584 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_446
timestamp 1662439860
transform 1 0 42136 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_449
timestamp 1662439860
transform 1 0 42412 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_458
timestamp 1662439860
transform 1 0 43240 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_469
timestamp 1662439860
transform 1 0 44252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_473
timestamp 1662439860
transform 1 0 44620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_495
timestamp 1662439860
transform 1 0 46644 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_499
timestamp 1662439860
transform 1 0 47012 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_502
timestamp 1662439860
transform 1 0 47288 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_505
timestamp 1662439860
transform 1 0 47564 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_511
timestamp 1662439860
transform 1 0 48116 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_520
timestamp 1662439860
transform 1 0 48944 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_531
timestamp 1662439860
transform 1 0 49956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_535
timestamp 1662439860
transform 1 0 50324 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_556
timestamp 1662439860
transform 1 0 52256 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_561
timestamp 1662439860
transform 1 0 52716 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_572
timestamp 1662439860
transform 1 0 53728 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_579
timestamp 1662439860
transform 1 0 54372 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_590
timestamp 1662439860
transform 1 0 55384 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_597
timestamp 1662439860
transform 1 0 56028 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_603
timestamp 1662439860
transform 1 0 56580 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_614
timestamp 1662439860
transform 1 0 57592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_617
timestamp 1662439860
transform 1 0 57868 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_639
timestamp 1662439860
transform 1 0 59892 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_645
timestamp 1662439860
transform 1 0 60444 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_649
timestamp 1662439860
transform 1 0 60812 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_670
timestamp 1662439860
transform 1 0 62744 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_673
timestamp 1662439860
transform 1 0 63020 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_695
timestamp 1662439860
transform 1 0 65044 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_719
timestamp 1662439860
transform 1 0 67252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_726
timestamp 1662439860
transform 1 0 67896 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_729
timestamp 1662439860
transform 1 0 68172 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_751
timestamp 1662439860
transform 1 0 70196 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_775
timestamp 1662439860
transform 1 0 72404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_782
timestamp 1662439860
transform 1 0 73048 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_785
timestamp 1662439860
transform 1 0 73324 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_790
timestamp 1662439860
transform 1 0 73784 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_796
timestamp 1662439860
transform 1 0 74336 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_804
timestamp 1662439860
transform 1 0 75072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_825
timestamp 1662439860
transform 1 0 77004 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_838
timestamp 1662439860
transform 1 0 78200 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_841
timestamp 1662439860
transform 1 0 78476 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_846
timestamp 1662439860
transform 1 0 78936 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_870
timestamp 1662439860
transform 1 0 81144 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_887
timestamp 1662439860
transform 1 0 82708 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_894
timestamp 1662439860
transform 1 0 83352 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_897
timestamp 1662439860
transform 1 0 83628 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_904
timestamp 1662439860
transform 1 0 84272 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_911
timestamp 1662439860
transform 1 0 84916 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_917
timestamp 1662439860
transform 1 0 85468 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_926
timestamp 1662439860
transform 1 0 86296 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_950
timestamp 1662439860
transform 1 0 88504 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_953
timestamp 1662439860
transform 1 0 88780 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_958
timestamp 1662439860
transform 1 0 89240 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_964
timestamp 1662439860
transform 1 0 89792 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_985
timestamp 1662439860
transform 1 0 91724 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1002
timestamp 1662439860
transform 1 0 93288 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1009
timestamp 1662439860
transform 1 0 93932 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1014
timestamp 1662439860
transform 1 0 94392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1662439860
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_8
timestamp 1662439860
transform 1 0 1840 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1662439860
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1662439860
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_45
timestamp 1662439860
transform 1 0 5244 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_49
timestamp 1662439860
transform 1 0 5612 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_52
timestamp 1662439860
transform 1 0 5888 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_65
timestamp 1662439860
transform 1 0 7084 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_71
timestamp 1662439860
transform 1 0 7636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1662439860
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1662439860
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_94
timestamp 1662439860
transform 1 0 9752 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_100
timestamp 1662439860
transform 1 0 10304 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_106
timestamp 1662439860
transform 1 0 10856 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_112
timestamp 1662439860
transform 1 0 11408 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_120
timestamp 1662439860
transform 1 0 12144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_126
timestamp 1662439860
transform 1 0 12696 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1662439860
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1662439860
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_147
timestamp 1662439860
transform 1 0 14628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_157
timestamp 1662439860
transform 1 0 15548 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_183
timestamp 1662439860
transform 1 0 17940 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_191
timestamp 1662439860
transform 1 0 18676 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1662439860
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1662439860
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_202
timestamp 1662439860
transform 1 0 19688 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1662439860
transform 1 0 20424 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_216
timestamp 1662439860
transform 1 0 20976 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_240
timestamp 1662439860
transform 1 0 23184 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1662439860
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_253
timestamp 1662439860
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_265
timestamp 1662439860
transform 1 0 25484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_269
timestamp 1662439860
transform 1 0 25852 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_291
timestamp 1662439860
transform 1 0 27876 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_297
timestamp 1662439860
transform 1 0 28428 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_300
timestamp 1662439860
transform 1 0 28704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1662439860
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_309
timestamp 1662439860
transform 1 0 29532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_313
timestamp 1662439860
transform 1 0 29900 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_316
timestamp 1662439860
transform 1 0 30176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_322
timestamp 1662439860
transform 1 0 30728 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_332
timestamp 1662439860
transform 1 0 31648 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_340
timestamp 1662439860
transform 1 0 32384 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1662439860
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_365
timestamp 1662439860
transform 1 0 34684 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_371
timestamp 1662439860
transform 1 0 35236 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_393
timestamp 1662439860
transform 1 0 37260 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_408
timestamp 1662439860
transform 1 0 38640 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_418
timestamp 1662439860
transform 1 0 39560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_421
timestamp 1662439860
transform 1 0 39836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_445
timestamp 1662439860
transform 1 0 42044 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_451
timestamp 1662439860
transform 1 0 42596 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_457
timestamp 1662439860
transform 1 0 43148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_474
timestamp 1662439860
transform 1 0 44712 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_477
timestamp 1662439860
transform 1 0 44988 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_485
timestamp 1662439860
transform 1 0 45724 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_511
timestamp 1662439860
transform 1 0 48116 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_519
timestamp 1662439860
transform 1 0 48852 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_529
timestamp 1662439860
transform 1 0 49772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_533
timestamp 1662439860
transform 1 0 50140 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_541
timestamp 1662439860
transform 1 0 50876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_548
timestamp 1662439860
transform 1 0 51520 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_574
timestamp 1662439860
transform 1 0 53912 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_583
timestamp 1662439860
transform 1 0 54740 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1662439860
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_589
timestamp 1662439860
transform 1 0 55292 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_601
timestamp 1662439860
transform 1 0 56396 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_612
timestamp 1662439860
transform 1 0 57408 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_620
timestamp 1662439860
transform 1 0 58144 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_630
timestamp 1662439860
transform 1 0 59064 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1662439860
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1662439860
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_645
timestamp 1662439860
transform 1 0 60444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_656
timestamp 1662439860
transform 1 0 61456 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_681
timestamp 1662439860
transform 1 0 63756 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_688
timestamp 1662439860
transform 1 0 64400 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_694
timestamp 1662439860
transform 1 0 64952 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_701
timestamp 1662439860
transform 1 0 65596 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_710
timestamp 1662439860
transform 1 0 66424 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_716
timestamp 1662439860
transform 1 0 66976 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_739
timestamp 1662439860
transform 1 0 69092 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_750
timestamp 1662439860
transform 1 0 70104 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_16_757
timestamp 1662439860
transform 1 0 70748 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_765
timestamp 1662439860
transform 1 0 71484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_782
timestamp 1662439860
transform 1 0 73048 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_788
timestamp 1662439860
transform 1 0 73600 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_792
timestamp 1662439860
transform 1 0 73968 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_800
timestamp 1662439860
transform 1 0 74704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_810
timestamp 1662439860
transform 1 0 75624 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_813
timestamp 1662439860
transform 1 0 75900 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_825
timestamp 1662439860
transform 1 0 77004 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_836
timestamp 1662439860
transform 1 0 78016 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_846
timestamp 1662439860
transform 1 0 78936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_850
timestamp 1662439860
transform 1 0 79304 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_854
timestamp 1662439860
transform 1 0 79672 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_860
timestamp 1662439860
transform 1 0 80224 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_864
timestamp 1662439860
transform 1 0 80592 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_869
timestamp 1662439860
transform 1 0 81052 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_897
timestamp 1662439860
transform 1 0 83628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_910
timestamp 1662439860
transform 1 0 84824 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_916
timestamp 1662439860
transform 1 0 85376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_922
timestamp 1662439860
transform 1 0 85928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_925
timestamp 1662439860
transform 1 0 86204 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_940
timestamp 1662439860
transform 1 0 87584 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_948
timestamp 1662439860
transform 1 0 88320 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_954
timestamp 1662439860
transform 1 0 88872 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_960
timestamp 1662439860
transform 1 0 89424 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_967
timestamp 1662439860
transform 1 0 90068 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_974
timestamp 1662439860
transform 1 0 90712 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_981
timestamp 1662439860
transform 1 0 91356 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1003
timestamp 1662439860
transform 1 0 93380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1010
timestamp 1662439860
transform 1 0 94024 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1662439860
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_7
timestamp 1662439860
transform 1 0 1748 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_15
timestamp 1662439860
transform 1 0 2484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_38
timestamp 1662439860
transform 1 0 4600 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_44
timestamp 1662439860
transform 1 0 5152 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_50
timestamp 1662439860
transform 1 0 5704 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1662439860
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_66
timestamp 1662439860
transform 1 0 7176 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_94
timestamp 1662439860
transform 1 0 9752 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_104
timestamp 1662439860
transform 1 0 10672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1662439860
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_119
timestamp 1662439860
transform 1 0 12052 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_122
timestamp 1662439860
transform 1 0 12328 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_133
timestamp 1662439860
transform 1 0 13340 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_142
timestamp 1662439860
transform 1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1662439860
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1662439860
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_176
timestamp 1662439860
transform 1 0 17296 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_203
timestamp 1662439860
transform 1 0 19780 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_213
timestamp 1662439860
transform 1 0 20700 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_219
timestamp 1662439860
transform 1 0 21252 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1662439860
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1662439860
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_247
timestamp 1662439860
transform 1 0 23828 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_253
timestamp 1662439860
transform 1 0 24380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1662439860
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1662439860
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_290
timestamp 1662439860
transform 1 0 27784 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_300
timestamp 1662439860
transform 1 0 28704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_311
timestamp 1662439860
transform 1 0 29716 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_317
timestamp 1662439860
transform 1 0 30268 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_324
timestamp 1662439860
transform 1 0 30912 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1662439860
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_337
timestamp 1662439860
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_341
timestamp 1662439860
transform 1 0 32476 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_344
timestamp 1662439860
transform 1 0 32752 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_361
timestamp 1662439860
transform 1 0 34316 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_365
timestamp 1662439860
transform 1 0 34684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_379
timestamp 1662439860
transform 1 0 35972 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_383
timestamp 1662439860
transform 1 0 36340 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_387
timestamp 1662439860
transform 1 0 36708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1662439860
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_393
timestamp 1662439860
transform 1 0 37260 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_399
timestamp 1662439860
transform 1 0 37812 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_413
timestamp 1662439860
transform 1 0 39100 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_430
timestamp 1662439860
transform 1 0 40664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_443
timestamp 1662439860
transform 1 0 41860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1662439860
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_449
timestamp 1662439860
transform 1 0 42412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_458
timestamp 1662439860
transform 1 0 43240 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_466
timestamp 1662439860
transform 1 0 43976 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_472
timestamp 1662439860
transform 1 0 44528 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1662439860
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1662439860
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_505
timestamp 1662439860
transform 1 0 47564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_511
timestamp 1662439860
transform 1 0 48116 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_525
timestamp 1662439860
transform 1 0 49404 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_546
timestamp 1662439860
transform 1 0 51336 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_558
timestamp 1662439860
transform 1 0 52440 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_561
timestamp 1662439860
transform 1 0 52716 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_566
timestamp 1662439860
transform 1 0 53176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_592
timestamp 1662439860
transform 1 0 55568 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_605
timestamp 1662439860
transform 1 0 56764 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_614
timestamp 1662439860
transform 1 0 57592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_617
timestamp 1662439860
transform 1 0 57868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_629
timestamp 1662439860
transform 1 0 58972 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_635
timestamp 1662439860
transform 1 0 59524 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_641
timestamp 1662439860
transform 1 0 60076 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_647
timestamp 1662439860
transform 1 0 60628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_653
timestamp 1662439860
transform 1 0 61180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_670
timestamp 1662439860
transform 1 0 62744 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_673
timestamp 1662439860
transform 1 0 63020 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_697
timestamp 1662439860
transform 1 0 65228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_703
timestamp 1662439860
transform 1 0 65780 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_724
timestamp 1662439860
transform 1 0 67712 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_729
timestamp 1662439860
transform 1 0 68172 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_751
timestamp 1662439860
transform 1 0 70196 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_768
timestamp 1662439860
transform 1 0 71760 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_781
timestamp 1662439860
transform 1 0 72956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_785
timestamp 1662439860
transform 1 0 73324 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_790
timestamp 1662439860
transform 1 0 73784 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_796
timestamp 1662439860
transform 1 0 74336 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_802
timestamp 1662439860
transform 1 0 74888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_806
timestamp 1662439860
transform 1 0 75256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_810
timestamp 1662439860
transform 1 0 75624 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_818
timestamp 1662439860
transform 1 0 76360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_830
timestamp 1662439860
transform 1 0 77464 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_837
timestamp 1662439860
transform 1 0 78108 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_841
timestamp 1662439860
transform 1 0 78476 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_849
timestamp 1662439860
transform 1 0 79212 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_855
timestamp 1662439860
transform 1 0 79764 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_868
timestamp 1662439860
transform 1 0 80960 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_894
timestamp 1662439860
transform 1 0 83352 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_897
timestamp 1662439860
transform 1 0 83628 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_906
timestamp 1662439860
transform 1 0 84456 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_916
timestamp 1662439860
transform 1 0 85376 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_924
timestamp 1662439860
transform 1 0 86112 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_945
timestamp 1662439860
transform 1 0 88044 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_951
timestamp 1662439860
transform 1 0 88596 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_953
timestamp 1662439860
transform 1 0 88780 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_958
timestamp 1662439860
transform 1 0 89240 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_984
timestamp 1662439860
transform 1 0 91632 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1001
timestamp 1662439860
transform 1 0 93196 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1007
timestamp 1662439860
transform 1 0 93748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1009
timestamp 1662439860
transform 1 0 93932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1014
timestamp 1662439860
transform 1 0 94392 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1662439860
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1662439860
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1662439860
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_29
timestamp 1662439860
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_46
timestamp 1662439860
transform 1 0 5336 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_56
timestamp 1662439860
transform 1 0 6256 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_60
timestamp 1662439860
transform 1 0 6624 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_63
timestamp 1662439860
transform 1 0 6900 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_69
timestamp 1662439860
transform 1 0 7452 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1662439860
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1662439860
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1662439860
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_109
timestamp 1662439860
transform 1 0 11132 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_117
timestamp 1662439860
transform 1 0 11868 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1662439860
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1662439860
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_164
timestamp 1662439860
transform 1 0 16192 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_190
timestamp 1662439860
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1662439860
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_219
timestamp 1662439860
transform 1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_226
timestamp 1662439860
transform 1 0 21896 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1662439860
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_253
timestamp 1662439860
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_259
timestamp 1662439860
transform 1 0 24932 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_265
timestamp 1662439860
transform 1 0 25484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_276
timestamp 1662439860
transform 1 0 26496 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_288
timestamp 1662439860
transform 1 0 27600 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_298
timestamp 1662439860
transform 1 0 28520 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1662439860
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_309
timestamp 1662439860
transform 1 0 29532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_319
timestamp 1662439860
transform 1 0 30452 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_330
timestamp 1662439860
transform 1 0 31464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_347
timestamp 1662439860
transform 1 0 33028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_358
timestamp 1662439860
transform 1 0 34040 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1662439860
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_370
timestamp 1662439860
transform 1 0 35144 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_394
timestamp 1662439860
transform 1 0 37352 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_418
timestamp 1662439860
transform 1 0 39560 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_421
timestamp 1662439860
transform 1 0 39836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_425
timestamp 1662439860
transform 1 0 40204 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_446
timestamp 1662439860
transform 1 0 42136 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_453
timestamp 1662439860
transform 1 0 42780 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_459
timestamp 1662439860
transform 1 0 43332 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_473
timestamp 1662439860
transform 1 0 44620 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_477
timestamp 1662439860
transform 1 0 44988 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_484
timestamp 1662439860
transform 1 0 45632 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_509
timestamp 1662439860
transform 1 0 47932 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_521
timestamp 1662439860
transform 1 0 49036 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_530
timestamp 1662439860
transform 1 0 49864 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_533
timestamp 1662439860
transform 1 0 50140 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_559
timestamp 1662439860
transform 1 0 52532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_567
timestamp 1662439860
transform 1 0 53268 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_577
timestamp 1662439860
transform 1 0 54188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_583
timestamp 1662439860
transform 1 0 54740 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1662439860
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_589
timestamp 1662439860
transform 1 0 55292 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_605
timestamp 1662439860
transform 1 0 56764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_612
timestamp 1662439860
transform 1 0 57408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_619
timestamp 1662439860
transform 1 0 58052 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_625
timestamp 1662439860
transform 1 0 58604 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_629
timestamp 1662439860
transform 1 0 58972 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_635
timestamp 1662439860
transform 1 0 59524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_641
timestamp 1662439860
transform 1 0 60076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_645
timestamp 1662439860
transform 1 0 60444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_650
timestamp 1662439860
transform 1 0 60904 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_665
timestamp 1662439860
transform 1 0 62284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_692
timestamp 1662439860
transform 1 0 64768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_698
timestamp 1662439860
transform 1 0 65320 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_701
timestamp 1662439860
transform 1 0 65596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_706
timestamp 1662439860
transform 1 0 66056 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_713
timestamp 1662439860
transform 1 0 66700 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_722
timestamp 1662439860
transform 1 0 67528 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_747
timestamp 1662439860
transform 1 0 69828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_754
timestamp 1662439860
transform 1 0 70472 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_757
timestamp 1662439860
transform 1 0 70748 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_783
timestamp 1662439860
transform 1 0 73140 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_810
timestamp 1662439860
transform 1 0 75624 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_813
timestamp 1662439860
transform 1 0 75900 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_820
timestamp 1662439860
transform 1 0 76544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_831
timestamp 1662439860
transform 1 0 77556 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_842
timestamp 1662439860
transform 1 0 78568 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_849
timestamp 1662439860
transform 1 0 79212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_855
timestamp 1662439860
transform 1 0 79764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_861
timestamp 1662439860
transform 1 0 80316 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_867
timestamp 1662439860
transform 1 0 80868 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_869
timestamp 1662439860
transform 1 0 81052 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_878
timestamp 1662439860
transform 1 0 81880 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_885
timestamp 1662439860
transform 1 0 82524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_898
timestamp 1662439860
transform 1 0 83720 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_922
timestamp 1662439860
transform 1 0 85928 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_925
timestamp 1662439860
transform 1 0 86204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_930
timestamp 1662439860
transform 1 0 86664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_947
timestamp 1662439860
transform 1 0 88228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_953
timestamp 1662439860
transform 1 0 88780 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_959
timestamp 1662439860
transform 1 0 89332 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_965
timestamp 1662439860
transform 1 0 89884 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_969
timestamp 1662439860
transform 1 0 90252 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_974
timestamp 1662439860
transform 1 0 90712 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_981
timestamp 1662439860
transform 1 0 91356 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1003
timestamp 1662439860
transform 1 0 93380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1009
timestamp 1662439860
transform 1 0 93932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_1014
timestamp 1662439860
transform 1 0 94392 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1662439860
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_15
timestamp 1662439860
transform 1 0 2484 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_23
timestamp 1662439860
transform 1 0 3220 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_37
timestamp 1662439860
transform 1 0 4508 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_47
timestamp 1662439860
transform 1 0 5428 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_51
timestamp 1662439860
transform 1 0 5796 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1662439860
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1662439860
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_66
timestamp 1662439860
transform 1 0 7176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_77
timestamp 1662439860
transform 1 0 8188 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_83
timestamp 1662439860
transform 1 0 8740 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_89
timestamp 1662439860
transform 1 0 9292 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_97
timestamp 1662439860
transform 1 0 10028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1662439860
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1662439860
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_118
timestamp 1662439860
transform 1 0 11960 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_130
timestamp 1662439860
transform 1 0 13064 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_133
timestamp 1662439860
transform 1 0 13340 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_140
timestamp 1662439860
transform 1 0 13984 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_144
timestamp 1662439860
transform 1 0 14352 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1662439860
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1662439860
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_177
timestamp 1662439860
transform 1 0 17388 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_184
timestamp 1662439860
transform 1 0 18032 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_188
timestamp 1662439860
transform 1 0 18400 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_192
timestamp 1662439860
transform 1 0 18768 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1662439860
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_225
timestamp 1662439860
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_234
timestamp 1662439860
transform 1 0 22632 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_258
timestamp 1662439860
transform 1 0 24840 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_265
timestamp 1662439860
transform 1 0 25484 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1662439860
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1662439860
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_285
timestamp 1662439860
transform 1 0 27324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_307
timestamp 1662439860
transform 1 0 29348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_311
timestamp 1662439860
transform 1 0 29716 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_314
timestamp 1662439860
transform 1 0 29992 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_321
timestamp 1662439860
transform 1 0 30636 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1662439860
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_337
timestamp 1662439860
transform 1 0 32108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_341
timestamp 1662439860
transform 1 0 32476 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_362
timestamp 1662439860
transform 1 0 34408 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_366
timestamp 1662439860
transform 1 0 34776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_372
timestamp 1662439860
transform 1 0 35328 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_382
timestamp 1662439860
transform 1 0 36248 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_390
timestamp 1662439860
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_393
timestamp 1662439860
transform 1 0 37260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_397
timestamp 1662439860
transform 1 0 37628 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_401
timestamp 1662439860
transform 1 0 37996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_426
timestamp 1662439860
transform 1 0 40296 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_432
timestamp 1662439860
transform 1 0 40848 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_435
timestamp 1662439860
transform 1 0 41124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_446
timestamp 1662439860
transform 1 0 42136 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_449
timestamp 1662439860
transform 1 0 42412 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_458
timestamp 1662439860
transform 1 0 43240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_464
timestamp 1662439860
transform 1 0 43792 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_488
timestamp 1662439860
transform 1 0 46000 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_502
timestamp 1662439860
transform 1 0 47288 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_505
timestamp 1662439860
transform 1 0 47564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_514
timestamp 1662439860
transform 1 0 48392 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_518
timestamp 1662439860
transform 1 0 48760 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_528
timestamp 1662439860
transform 1 0 49680 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_545
timestamp 1662439860
transform 1 0 51244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_556
timestamp 1662439860
transform 1 0 52256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_561
timestamp 1662439860
transform 1 0 52716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_583
timestamp 1662439860
transform 1 0 54740 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_600
timestamp 1662439860
transform 1 0 56304 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_606
timestamp 1662439860
transform 1 0 56856 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_612
timestamp 1662439860
transform 1 0 57408 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_617
timestamp 1662439860
transform 1 0 57868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_622
timestamp 1662439860
transform 1 0 58328 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_653
timestamp 1662439860
transform 1 0 61180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_659
timestamp 1662439860
transform 1 0 61732 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1662439860
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1662439860
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_673
timestamp 1662439860
transform 1 0 63020 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_696
timestamp 1662439860
transform 1 0 65136 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_703
timestamp 1662439860
transform 1 0 65780 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_709
timestamp 1662439860
transform 1 0 66332 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_713
timestamp 1662439860
transform 1 0 66700 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_721
timestamp 1662439860
transform 1 0 67436 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_725
timestamp 1662439860
transform 1 0 67804 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_729
timestamp 1662439860
transform 1 0 68172 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_736
timestamp 1662439860
transform 1 0 68816 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_742
timestamp 1662439860
transform 1 0 69368 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_750
timestamp 1662439860
transform 1 0 70104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_777
timestamp 1662439860
transform 1 0 72588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_783
timestamp 1662439860
transform 1 0 73140 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_785
timestamp 1662439860
transform 1 0 73324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_791
timestamp 1662439860
transform 1 0 73876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_797
timestamp 1662439860
transform 1 0 74428 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_801
timestamp 1662439860
transform 1 0 74796 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_806
timestamp 1662439860
transform 1 0 75256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_813
timestamp 1662439860
transform 1 0 75900 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_821
timestamp 1662439860
transform 1 0 76636 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_826
timestamp 1662439860
transform 1 0 77096 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_836
timestamp 1662439860
transform 1 0 78016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_841
timestamp 1662439860
transform 1 0 78476 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_863
timestamp 1662439860
transform 1 0 80500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_871
timestamp 1662439860
transform 1 0 81236 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_894
timestamp 1662439860
transform 1 0 83352 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_897
timestamp 1662439860
transform 1 0 83628 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_903
timestamp 1662439860
transform 1 0 84180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_910
timestamp 1662439860
transform 1 0 84824 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_914
timestamp 1662439860
transform 1 0 85192 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_918
timestamp 1662439860
transform 1 0 85560 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_922
timestamp 1662439860
transform 1 0 85928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_926
timestamp 1662439860
transform 1 0 86296 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_937
timestamp 1662439860
transform 1 0 87308 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_944
timestamp 1662439860
transform 1 0 87952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_950
timestamp 1662439860
transform 1 0 88504 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_953
timestamp 1662439860
transform 1 0 88780 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_962
timestamp 1662439860
transform 1 0 89608 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_990
timestamp 1662439860
transform 1 0 92184 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_997
timestamp 1662439860
transform 1 0 92828 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1004
timestamp 1662439860
transform 1 0 93472 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1009
timestamp 1662439860
transform 1 0 93932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1014
timestamp 1662439860
transform 1 0 94392 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1662439860
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_15
timestamp 1662439860
transform 1 0 2484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1662439860
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1662439860
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_38
timestamp 1662439860
transform 1 0 4600 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_44
timestamp 1662439860
transform 1 0 5152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_48
timestamp 1662439860
transform 1 0 5520 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_54
timestamp 1662439860
transform 1 0 6072 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_64
timestamp 1662439860
transform 1 0 6992 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_70
timestamp 1662439860
transform 1 0 7544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_74
timestamp 1662439860
transform 1 0 7912 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1662439860
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1662439860
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1662439860
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_114
timestamp 1662439860
transform 1 0 11592 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_127
timestamp 1662439860
transform 1 0 12788 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1662439860
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1662439860
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1662439860
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_166
timestamp 1662439860
transform 1 0 16376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_174
timestamp 1662439860
transform 1 0 17112 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1662439860
transform 1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1662439860
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1662439860
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1662439860
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_220
timestamp 1662439860
transform 1 0 21344 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_228
timestamp 1662439860
transform 1 0 22080 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1662439860
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1662439860
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_257
timestamp 1662439860
transform 1 0 24748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_267
timestamp 1662439860
transform 1 0 25668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_291
timestamp 1662439860
transform 1 0 27876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_299
timestamp 1662439860
transform 1 0 28612 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_303
timestamp 1662439860
transform 1 0 28980 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1662439860
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1662439860
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_331
timestamp 1662439860
transform 1 0 31556 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_337
timestamp 1662439860
transform 1 0 32108 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1662439860
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_365
timestamp 1662439860
transform 1 0 34684 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_374
timestamp 1662439860
transform 1 0 35512 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_381
timestamp 1662439860
transform 1 0 36156 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_385
timestamp 1662439860
transform 1 0 36524 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_388
timestamp 1662439860
transform 1 0 36800 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_394
timestamp 1662439860
transform 1 0 37352 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_418
timestamp 1662439860
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_421
timestamp 1662439860
transform 1 0 39836 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_426
timestamp 1662439860
transform 1 0 40296 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_450
timestamp 1662439860
transform 1 0 42504 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_474
timestamp 1662439860
transform 1 0 44712 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_477
timestamp 1662439860
transform 1 0 44988 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_499
timestamp 1662439860
transform 1 0 47012 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_523
timestamp 1662439860
transform 1 0 49220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_530
timestamp 1662439860
transform 1 0 49864 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_533
timestamp 1662439860
transform 1 0 50140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_537
timestamp 1662439860
transform 1 0 50508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_543
timestamp 1662439860
transform 1 0 51060 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_557
timestamp 1662439860
transform 1 0 52348 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_582
timestamp 1662439860
transform 1 0 54648 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_589
timestamp 1662439860
transform 1 0 55292 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_606
timestamp 1662439860
transform 1 0 56856 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_630
timestamp 1662439860
transform 1 0 59064 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1662439860
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1662439860
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_645
timestamp 1662439860
transform 1 0 60444 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_650
timestamp 1662439860
transform 1 0 60904 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_656
timestamp 1662439860
transform 1 0 61456 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_660
timestamp 1662439860
transform 1 0 61824 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_685
timestamp 1662439860
transform 1 0 64124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_692
timestamp 1662439860
transform 1 0 64768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_698
timestamp 1662439860
transform 1 0 65320 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_701
timestamp 1662439860
transform 1 0 65596 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_706
timestamp 1662439860
transform 1 0 66056 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_713
timestamp 1662439860
transform 1 0 66700 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_719
timestamp 1662439860
transform 1 0 67252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_743
timestamp 1662439860
transform 1 0 69460 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_750
timestamp 1662439860
transform 1 0 70104 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_757
timestamp 1662439860
transform 1 0 70748 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_762
timestamp 1662439860
transform 1 0 71208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_786
timestamp 1662439860
transform 1 0 73416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_810
timestamp 1662439860
transform 1 0 75624 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_813
timestamp 1662439860
transform 1 0 75900 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_818
timestamp 1662439860
transform 1 0 76360 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_824
timestamp 1662439860
transform 1 0 76912 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_846
timestamp 1662439860
transform 1 0 78936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_853
timestamp 1662439860
transform 1 0 79580 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_860
timestamp 1662439860
transform 1 0 80224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_866
timestamp 1662439860
transform 1 0 80776 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_869
timestamp 1662439860
transform 1 0 81052 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_873
timestamp 1662439860
transform 1 0 81420 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_879
timestamp 1662439860
transform 1 0 81972 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_885
timestamp 1662439860
transform 1 0 82524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_909
timestamp 1662439860
transform 1 0 84732 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_915
timestamp 1662439860
transform 1 0 85284 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_921
timestamp 1662439860
transform 1 0 85836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_925
timestamp 1662439860
transform 1 0 86204 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_929
timestamp 1662439860
transform 1 0 86572 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_934
timestamp 1662439860
transform 1 0 87032 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_959
timestamp 1662439860
transform 1 0 89332 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_966
timestamp 1662439860
transform 1 0 89976 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_973
timestamp 1662439860
transform 1 0 90620 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_979
timestamp 1662439860
transform 1 0 91172 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_981
timestamp 1662439860
transform 1 0 91356 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_985
timestamp 1662439860
transform 1 0 91724 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1006
timestamp 1662439860
transform 1 0 93656 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1012
timestamp 1662439860
transform 1 0 94208 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1662439860
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_15
timestamp 1662439860
transform 1 0 2484 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_41
timestamp 1662439860
transform 1 0 4876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1662439860
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1662439860
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_61
timestamp 1662439860
transform 1 0 6716 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1662439860
transform 1 0 7452 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_73
timestamp 1662439860
transform 1 0 7820 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_84
timestamp 1662439860
transform 1 0 8832 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_90
timestamp 1662439860
transform 1 0 9384 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_102
timestamp 1662439860
transform 1 0 10488 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1662439860
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1662439860
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_122
timestamp 1662439860
transform 1 0 12328 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_130
timestamp 1662439860
transform 1 0 13064 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_133
timestamp 1662439860
transform 1 0 13340 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_144
timestamp 1662439860
transform 1 0 14352 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_155
timestamp 1662439860
transform 1 0 15364 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_162
timestamp 1662439860
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1662439860
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_173
timestamp 1662439860
transform 1 0 17020 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_179
timestamp 1662439860
transform 1 0 17572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_191
timestamp 1662439860
transform 1 0 18676 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_213
timestamp 1662439860
transform 1 0 20700 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1662439860
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1662439860
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_247
timestamp 1662439860
transform 1 0 23828 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1662439860
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_281
timestamp 1662439860
transform 1 0 26956 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_287
timestamp 1662439860
transform 1 0 27508 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_291
timestamp 1662439860
transform 1 0 27876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_295
timestamp 1662439860
transform 1 0 28244 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_316
timestamp 1662439860
transform 1 0 30176 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_320
timestamp 1662439860
transform 1 0 30544 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_324
timestamp 1662439860
transform 1 0 30912 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1662439860
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1662439860
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_342
timestamp 1662439860
transform 1 0 32568 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_351
timestamp 1662439860
transform 1 0 33396 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_376
timestamp 1662439860
transform 1 0 35696 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_384
timestamp 1662439860
transform 1 0 36432 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1662439860
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_393
timestamp 1662439860
transform 1 0 37260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_397
timestamp 1662439860
transform 1 0 37628 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_400
timestamp 1662439860
transform 1 0 37904 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_407
timestamp 1662439860
transform 1 0 38548 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_434
timestamp 1662439860
transform 1 0 41032 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_445
timestamp 1662439860
transform 1 0 42044 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_449
timestamp 1662439860
transform 1 0 42412 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_464
timestamp 1662439860
transform 1 0 43792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_478
timestamp 1662439860
transform 1 0 45080 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_502
timestamp 1662439860
transform 1 0 47288 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_505
timestamp 1662439860
transform 1 0 47564 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_527
timestamp 1662439860
transform 1 0 49588 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_533
timestamp 1662439860
transform 1 0 50140 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_539
timestamp 1662439860
transform 1 0 50692 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_545
timestamp 1662439860
transform 1 0 51244 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_551
timestamp 1662439860
transform 1 0 51796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_557
timestamp 1662439860
transform 1 0 52348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_561
timestamp 1662439860
transform 1 0 52716 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_566
timestamp 1662439860
transform 1 0 53176 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_573
timestamp 1662439860
transform 1 0 53820 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_579
timestamp 1662439860
transform 1 0 54372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_585
timestamp 1662439860
transform 1 0 54924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1662439860
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1662439860
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_617
timestamp 1662439860
transform 1 0 57868 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_622
timestamp 1662439860
transform 1 0 58328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_628
timestamp 1662439860
transform 1 0 58880 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_655
timestamp 1662439860
transform 1 0 61364 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_661
timestamp 1662439860
transform 1 0 61916 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_667
timestamp 1662439860
transform 1 0 62468 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1662439860
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_673
timestamp 1662439860
transform 1 0 63020 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_680
timestamp 1662439860
transform 1 0 63664 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_686
timestamp 1662439860
transform 1 0 64216 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_711
timestamp 1662439860
transform 1 0 66516 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_717
timestamp 1662439860
transform 1 0 67068 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_723
timestamp 1662439860
transform 1 0 67620 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 1662439860
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_729
timestamp 1662439860
transform 1 0 68172 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_753
timestamp 1662439860
transform 1 0 70380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_778
timestamp 1662439860
transform 1 0 72680 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_785
timestamp 1662439860
transform 1 0 73324 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_790
timestamp 1662439860
transform 1 0 73784 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_796
timestamp 1662439860
transform 1 0 74336 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_802
timestamp 1662439860
transform 1 0 74888 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_811
timestamp 1662439860
transform 1 0 75716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_818
timestamp 1662439860
transform 1 0 76360 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_825
timestamp 1662439860
transform 1 0 77004 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_832
timestamp 1662439860
transform 1 0 77648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_838
timestamp 1662439860
transform 1 0 78200 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_841
timestamp 1662439860
transform 1 0 78476 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_864
timestamp 1662439860
transform 1 0 80592 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_870
timestamp 1662439860
transform 1 0 81144 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_876
timestamp 1662439860
transform 1 0 81696 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_882
timestamp 1662439860
transform 1 0 82248 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_888
timestamp 1662439860
transform 1 0 82800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_894
timestamp 1662439860
transform 1 0 83352 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_897
timestamp 1662439860
transform 1 0 83628 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_901
timestamp 1662439860
transform 1 0 83996 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_931
timestamp 1662439860
transform 1 0 86756 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_937
timestamp 1662439860
transform 1 0 87308 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_943
timestamp 1662439860
transform 1 0 87860 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_949
timestamp 1662439860
transform 1 0 88412 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_953
timestamp 1662439860
transform 1 0 88780 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_976
timestamp 1662439860
transform 1 0 90896 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_982
timestamp 1662439860
transform 1 0 91448 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_988
timestamp 1662439860
transform 1 0 92000 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_997
timestamp 1662439860
transform 1 0 92828 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_1003
timestamp 1662439860
transform 1 0 93380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1007
timestamp 1662439860
transform 1 0 93748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_1009
timestamp 1662439860
transform 1 0 93932 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_1013
timestamp 1662439860
transform 1 0 94300 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1662439860
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1662439860
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1662439860
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1662439860
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1662439860
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_53
timestamp 1662439860
transform 1 0 5980 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_59
timestamp 1662439860
transform 1 0 6532 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1662439860
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1662439860
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_89
timestamp 1662439860
transform 1 0 9292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_101
timestamp 1662439860
transform 1 0 10396 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_109
timestamp 1662439860
transform 1 0 11132 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_117
timestamp 1662439860
transform 1 0 11868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_121
timestamp 1662439860
transform 1 0 12236 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_125
timestamp 1662439860
transform 1 0 12604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_131
timestamp 1662439860
transform 1 0 13156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1662439860
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1662439860
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_145
timestamp 1662439860
transform 1 0 14444 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_148
timestamp 1662439860
transform 1 0 14720 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_159
timestamp 1662439860
transform 1 0 15732 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1662439860
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1662439860
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1662439860
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1662439860
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1662439860
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_222
timestamp 1662439860
transform 1 0 21528 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_247
timestamp 1662439860
transform 1 0 23828 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1662439860
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1662439860
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_258
timestamp 1662439860
transform 1 0 24840 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_264
timestamp 1662439860
transform 1 0 25392 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_268
timestamp 1662439860
transform 1 0 25760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1662439860
transform 1 0 26496 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_279
timestamp 1662439860
transform 1 0 26772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1662439860
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_309
timestamp 1662439860
transform 1 0 29532 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_315
timestamp 1662439860
transform 1 0 30084 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_322
timestamp 1662439860
transform 1 0 30728 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_330
timestamp 1662439860
transform 1 0 31464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_355
timestamp 1662439860
transform 1 0 33764 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_359
timestamp 1662439860
transform 1 0 34132 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1662439860
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_365
timestamp 1662439860
transform 1 0 34684 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_371
timestamp 1662439860
transform 1 0 35236 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_381
timestamp 1662439860
transform 1 0 36156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_398
timestamp 1662439860
transform 1 0 37720 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_405
timestamp 1662439860
transform 1 0 38364 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_409
timestamp 1662439860
transform 1 0 38732 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_414
timestamp 1662439860
transform 1 0 39192 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_421
timestamp 1662439860
transform 1 0 39836 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_425
timestamp 1662439860
transform 1 0 40204 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_447
timestamp 1662439860
transform 1 0 42228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_454
timestamp 1662439860
transform 1 0 42872 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_460
timestamp 1662439860
transform 1 0 43424 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_474
timestamp 1662439860
transform 1 0 44712 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_477
timestamp 1662439860
transform 1 0 44988 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_483
timestamp 1662439860
transform 1 0 45540 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_489
timestamp 1662439860
transform 1 0 46092 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_493
timestamp 1662439860
transform 1 0 46460 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_517
timestamp 1662439860
transform 1 0 48668 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_524
timestamp 1662439860
transform 1 0 49312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_530
timestamp 1662439860
transform 1 0 49864 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_533
timestamp 1662439860
transform 1 0 50140 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_537
timestamp 1662439860
transform 1 0 50508 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_543
timestamp 1662439860
transform 1 0 51060 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_547
timestamp 1662439860
transform 1 0 51428 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_569
timestamp 1662439860
transform 1 0 53452 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_576
timestamp 1662439860
transform 1 0 54096 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_582
timestamp 1662439860
transform 1 0 54648 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_589
timestamp 1662439860
transform 1 0 55292 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_593
timestamp 1662439860
transform 1 0 55660 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_601
timestamp 1662439860
transform 1 0 56396 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_607
timestamp 1662439860
transform 1 0 56948 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_628
timestamp 1662439860
transform 1 0 58880 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_634
timestamp 1662439860
transform 1 0 59432 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_638
timestamp 1662439860
transform 1 0 59800 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_642
timestamp 1662439860
transform 1 0 60168 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_645
timestamp 1662439860
transform 1 0 60444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_670
timestamp 1662439860
transform 1 0 62744 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_676
timestamp 1662439860
transform 1 0 63296 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_682
timestamp 1662439860
transform 1 0 63848 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_688
timestamp 1662439860
transform 1 0 64400 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_694
timestamp 1662439860
transform 1 0 64952 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_698
timestamp 1662439860
transform 1 0 65320 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_701
timestamp 1662439860
transform 1 0 65596 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_707
timestamp 1662439860
transform 1 0 66148 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_713
timestamp 1662439860
transform 1 0 66700 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_721
timestamp 1662439860
transform 1 0 67436 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_725
timestamp 1662439860
transform 1 0 67804 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_749
timestamp 1662439860
transform 1 0 70012 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_755
timestamp 1662439860
transform 1 0 70564 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_757
timestamp 1662439860
transform 1 0 70748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_766
timestamp 1662439860
transform 1 0 71576 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_773
timestamp 1662439860
transform 1 0 72220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_777
timestamp 1662439860
transform 1 0 72588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_798
timestamp 1662439860
transform 1 0 74520 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_804
timestamp 1662439860
transform 1 0 75072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_810
timestamp 1662439860
transform 1 0 75624 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_813
timestamp 1662439860
transform 1 0 75900 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_817
timestamp 1662439860
transform 1 0 76268 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_823
timestamp 1662439860
transform 1 0 76820 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_847
timestamp 1662439860
transform 1 0 79028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_854
timestamp 1662439860
transform 1 0 79672 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_861
timestamp 1662439860
transform 1 0 80316 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_867
timestamp 1662439860
transform 1 0 80868 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_869
timestamp 1662439860
transform 1 0 81052 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_873
timestamp 1662439860
transform 1 0 81420 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_879
timestamp 1662439860
transform 1 0 81972 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_885
timestamp 1662439860
transform 1 0 82524 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_900
timestamp 1662439860
transform 1 0 83904 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_906
timestamp 1662439860
transform 1 0 84456 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_910
timestamp 1662439860
transform 1 0 84824 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_914
timestamp 1662439860
transform 1 0 85192 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_920
timestamp 1662439860
transform 1 0 85744 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_925
timestamp 1662439860
transform 1 0 86204 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_940
timestamp 1662439860
transform 1 0 87584 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_953
timestamp 1662439860
transform 1 0 88780 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_957
timestamp 1662439860
transform 1 0 89148 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_962
timestamp 1662439860
transform 1 0 89608 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_968
timestamp 1662439860
transform 1 0 90160 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_974
timestamp 1662439860
transform 1 0 90712 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_981
timestamp 1662439860
transform 1 0 91356 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_985
timestamp 1662439860
transform 1 0 91724 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_991
timestamp 1662439860
transform 1 0 92276 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_997
timestamp 1662439860
transform 1 0 92828 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1009
timestamp 1662439860
transform 1 0 93932 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1015
timestamp 1662439860
transform 1 0 94484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1662439860
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1662439860
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1662439860
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1662439860
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1662439860
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1662439860
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1662439860
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1662439860
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1662439860
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1662439860
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1662439860
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1662439860
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1662439860
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_127
timestamp 1662439860
transform 1 0 12788 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_139
timestamp 1662439860
transform 1 0 13892 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_145
timestamp 1662439860
transform 1 0 14444 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_148
timestamp 1662439860
transform 1 0 14720 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_160
timestamp 1662439860
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1662439860
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1662439860
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_193
timestamp 1662439860
transform 1 0 18860 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1662439860
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 1662439860
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_230
timestamp 1662439860
transform 1 0 22264 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_237
timestamp 1662439860
transform 1 0 22908 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_244
timestamp 1662439860
transform 1 0 23552 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_272
timestamp 1662439860
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1662439860
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_314
timestamp 1662439860
transform 1 0 29992 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_331
timestamp 1662439860
transform 1 0 31556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1662439860
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_337
timestamp 1662439860
transform 1 0 32108 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_343
timestamp 1662439860
transform 1 0 32660 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_357
timestamp 1662439860
transform 1 0 33948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_374
timestamp 1662439860
transform 1 0 35512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_381
timestamp 1662439860
transform 1 0 36156 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_390
timestamp 1662439860
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1662439860
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_408
timestamp 1662439860
transform 1 0 38640 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_417
timestamp 1662439860
transform 1 0 39468 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_423
timestamp 1662439860
transform 1 0 40020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_427
timestamp 1662439860
transform 1 0 40388 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_431
timestamp 1662439860
transform 1 0 40756 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_435
timestamp 1662439860
transform 1 0 41124 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_442
timestamp 1662439860
transform 1 0 41768 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_449
timestamp 1662439860
transform 1 0 42412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_453
timestamp 1662439860
transform 1 0 42780 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_456
timestamp 1662439860
transform 1 0 43056 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_480
timestamp 1662439860
transform 1 0 45264 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1662439860
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1662439860
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_505
timestamp 1662439860
transform 1 0 47564 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_518
timestamp 1662439860
transform 1 0 48760 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_542
timestamp 1662439860
transform 1 0 50968 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_546
timestamp 1662439860
transform 1 0 51336 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_549
timestamp 1662439860
transform 1 0 51612 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_555
timestamp 1662439860
transform 1 0 52164 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1662439860
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_561
timestamp 1662439860
transform 1 0 52716 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_584
timestamp 1662439860
transform 1 0 54832 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1662439860
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1662439860
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_617
timestamp 1662439860
transform 1 0 57868 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_621
timestamp 1662439860
transform 1 0 58236 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_629
timestamp 1662439860
transform 1 0 58972 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_653
timestamp 1662439860
transform 1 0 61180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_660
timestamp 1662439860
transform 1 0 61824 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_666
timestamp 1662439860
transform 1 0 62376 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_673
timestamp 1662439860
transform 1 0 63020 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_677
timestamp 1662439860
transform 1 0 63388 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_683
timestamp 1662439860
transform 1 0 63940 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_689
timestamp 1662439860
transform 1 0 64492 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_714
timestamp 1662439860
transform 1 0 66792 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 1662439860
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 1662439860
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_729
timestamp 1662439860
transform 1 0 68172 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_734
timestamp 1662439860
transform 1 0 68632 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_738
timestamp 1662439860
transform 1 0 69000 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_742
timestamp 1662439860
transform 1 0 69368 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_766
timestamp 1662439860
transform 1 0 71576 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_778
timestamp 1662439860
transform 1 0 72680 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_785
timestamp 1662439860
transform 1 0 73324 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_796
timestamp 1662439860
transform 1 0 74336 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_802
timestamp 1662439860
transform 1 0 74888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_808
timestamp 1662439860
transform 1 0 75440 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_814
timestamp 1662439860
transform 1 0 75992 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_820
timestamp 1662439860
transform 1 0 76544 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_835
timestamp 1662439860
transform 1 0 77924 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_839
timestamp 1662439860
transform 1 0 78292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_841
timestamp 1662439860
transform 1 0 78476 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_846
timestamp 1662439860
transform 1 0 78936 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_852
timestamp 1662439860
transform 1 0 79488 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_867
timestamp 1662439860
transform 1 0 80868 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_873
timestamp 1662439860
transform 1 0 81420 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_894
timestamp 1662439860
transform 1 0 83352 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_897
timestamp 1662439860
transform 1 0 83628 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_908
timestamp 1662439860
transform 1 0 84640 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_912
timestamp 1662439860
transform 1 0 85008 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_915
timestamp 1662439860
transform 1 0 85284 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_921
timestamp 1662439860
transform 1 0 85836 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_925
timestamp 1662439860
transform 1 0 86204 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_928
timestamp 1662439860
transform 1 0 86480 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_934
timestamp 1662439860
transform 1 0 87032 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_940
timestamp 1662439860
transform 1 0 87584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_946
timestamp 1662439860
transform 1 0 88136 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_953
timestamp 1662439860
transform 1 0 88780 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_957
timestamp 1662439860
transform 1 0 89148 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_963
timestamp 1662439860
transform 1 0 89700 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_969
timestamp 1662439860
transform 1 0 90252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_973
timestamp 1662439860
transform 1 0 90620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_976
timestamp 1662439860
transform 1 0 90896 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_988
timestamp 1662439860
transform 1 0 92000 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_1000
timestamp 1662439860
transform 1 0 93104 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1009
timestamp 1662439860
transform 1 0 93932 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1015
timestamp 1662439860
transform 1 0 94484 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1662439860
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1662439860
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1662439860
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1662439860
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1662439860
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1662439860
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1662439860
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1662439860
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1662439860
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1662439860
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1662439860
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1662439860
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1662439860
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1662439860
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1662439860
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1662439860
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1662439860
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1662439860
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1662439860
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1662439860
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1662439860
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_197
timestamp 1662439860
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_208
timestamp 1662439860
transform 1 0 20240 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_215
timestamp 1662439860
transform 1 0 20884 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_227
timestamp 1662439860
transform 1 0 21988 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_233
timestamp 1662439860
transform 1 0 22540 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_237
timestamp 1662439860
transform 1 0 22908 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_243
timestamp 1662439860
transform 1 0 23460 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1662439860
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_253
timestamp 1662439860
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_257
timestamp 1662439860
transform 1 0 24748 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_260
timestamp 1662439860
transform 1 0 25024 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_272
timestamp 1662439860
transform 1 0 26128 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_284
timestamp 1662439860
transform 1 0 27232 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_299
timestamp 1662439860
transform 1 0 28612 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1662439860
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_309
timestamp 1662439860
transform 1 0 29532 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_317
timestamp 1662439860
transform 1 0 30268 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_323
timestamp 1662439860
transform 1 0 30820 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_329
timestamp 1662439860
transform 1 0 31372 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_333
timestamp 1662439860
transform 1 0 31740 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_343
timestamp 1662439860
transform 1 0 32660 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_360
timestamp 1662439860
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1662439860
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_370
timestamp 1662439860
transform 1 0 35144 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_376
timestamp 1662439860
transform 1 0 35696 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_380
timestamp 1662439860
transform 1 0 36064 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_383
timestamp 1662439860
transform 1 0 36340 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_389
timestamp 1662439860
transform 1 0 36892 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_395
timestamp 1662439860
transform 1 0 37444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_398
timestamp 1662439860
transform 1 0 37720 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_407
timestamp 1662439860
transform 1 0 38548 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_415
timestamp 1662439860
transform 1 0 39284 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1662439860
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_421
timestamp 1662439860
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_436
timestamp 1662439860
transform 1 0 41216 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_444
timestamp 1662439860
transform 1 0 41952 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_450
timestamp 1662439860
transform 1 0 42504 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_456
timestamp 1662439860
transform 1 0 43056 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_459
timestamp 1662439860
transform 1 0 43332 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_466
timestamp 1662439860
transform 1 0 43976 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_474
timestamp 1662439860
transform 1 0 44712 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_477
timestamp 1662439860
transform 1 0 44988 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_486
timestamp 1662439860
transform 1 0 45816 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_494
timestamp 1662439860
transform 1 0 46552 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_515
timestamp 1662439860
transform 1 0 48484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_522
timestamp 1662439860
transform 1 0 49128 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_528
timestamp 1662439860
transform 1 0 49680 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_533
timestamp 1662439860
transform 1 0 50140 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_537
timestamp 1662439860
transform 1 0 50508 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_540
timestamp 1662439860
transform 1 0 50784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_565
timestamp 1662439860
transform 1 0 53084 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_574
timestamp 1662439860
transform 1 0 53912 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_580
timestamp 1662439860
transform 1 0 54464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_586
timestamp 1662439860
transform 1 0 55016 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_589
timestamp 1662439860
transform 1 0 55292 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_595
timestamp 1662439860
transform 1 0 55844 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_599
timestamp 1662439860
transform 1 0 56212 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_607
timestamp 1662439860
transform 1 0 56948 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_628
timestamp 1662439860
transform 1 0 58880 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_634
timestamp 1662439860
transform 1 0 59432 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_638
timestamp 1662439860
transform 1 0 59800 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_642
timestamp 1662439860
transform 1 0 60168 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_645
timestamp 1662439860
transform 1 0 60444 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_651
timestamp 1662439860
transform 1 0 60996 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_672
timestamp 1662439860
transform 1 0 62928 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_678
timestamp 1662439860
transform 1 0 63480 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_686
timestamp 1662439860
transform 1 0 64216 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_696
timestamp 1662439860
transform 1 0 65136 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_701
timestamp 1662439860
transform 1 0 65596 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_708
timestamp 1662439860
transform 1 0 66240 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_715
timestamp 1662439860
transform 1 0 66884 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_722
timestamp 1662439860
transform 1 0 67528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_729
timestamp 1662439860
transform 1 0 68172 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_735
timestamp 1662439860
transform 1 0 68724 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_741
timestamp 1662439860
transform 1 0 69276 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_747
timestamp 1662439860
transform 1 0 69828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_753
timestamp 1662439860
transform 1 0 70380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_757
timestamp 1662439860
transform 1 0 70748 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_761
timestamp 1662439860
transform 1 0 71116 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_768
timestamp 1662439860
transform 1 0 71760 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_778
timestamp 1662439860
transform 1 0 72680 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_784
timestamp 1662439860
transform 1 0 73232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_790
timestamp 1662439860
transform 1 0 73784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_797
timestamp 1662439860
transform 1 0 74428 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_803
timestamp 1662439860
transform 1 0 74980 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_809
timestamp 1662439860
transform 1 0 75532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_813
timestamp 1662439860
transform 1 0 75900 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_820
timestamp 1662439860
transform 1 0 76544 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_849
timestamp 1662439860
transform 1 0 79212 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_855
timestamp 1662439860
transform 1 0 79764 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_861
timestamp 1662439860
transform 1 0 80316 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_867
timestamp 1662439860
transform 1 0 80868 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_869
timestamp 1662439860
transform 1 0 81052 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_873
timestamp 1662439860
transform 1 0 81420 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_885
timestamp 1662439860
transform 1 0 82524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_891
timestamp 1662439860
transform 1 0 83076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_899
timestamp 1662439860
transform 1 0 83812 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_907
timestamp 1662439860
transform 1 0 84548 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_919
timestamp 1662439860
transform 1 0 85652 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_923
timestamp 1662439860
transform 1 0 86020 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_925
timestamp 1662439860
transform 1 0 86204 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_929
timestamp 1662439860
transform 1 0 86572 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_941
timestamp 1662439860
transform 1 0 87676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_946
timestamp 1662439860
transform 1 0 88136 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_952
timestamp 1662439860
transform 1 0 88688 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_955
timestamp 1662439860
transform 1 0 88964 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_967
timestamp 1662439860
transform 1 0 90068 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_979
timestamp 1662439860
transform 1 0 91172 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_981
timestamp 1662439860
transform 1 0 91356 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_993
timestamp 1662439860
transform 1 0 92460 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_1005
timestamp 1662439860
transform 1 0 93564 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_1013
timestamp 1662439860
transform 1 0 94300 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1662439860
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1662439860
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1662439860
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1662439860
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1662439860
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1662439860
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1662439860
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1662439860
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1662439860
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1662439860
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1662439860
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1662439860
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1662439860
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1662439860
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1662439860
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1662439860
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1662439860
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1662439860
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1662439860
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_181
timestamp 1662439860
transform 1 0 17756 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1662439860
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_215
timestamp 1662439860
transform 1 0 20884 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1662439860
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1662439860
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1662439860
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1662439860
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1662439860
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1662439860
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1662439860
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1662439860
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_293
timestamp 1662439860
transform 1 0 28060 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_304
timestamp 1662439860
transform 1 0 29072 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_310
timestamp 1662439860
transform 1 0 29624 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_322
timestamp 1662439860
transform 1 0 30728 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_327
timestamp 1662439860
transform 1 0 31188 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1662439860
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_337
timestamp 1662439860
transform 1 0 32108 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_341
timestamp 1662439860
transform 1 0 32476 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_344
timestamp 1662439860
transform 1 0 32752 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_352
timestamp 1662439860
transform 1 0 33488 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_355
timestamp 1662439860
transform 1 0 33764 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_361
timestamp 1662439860
transform 1 0 34316 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_367
timestamp 1662439860
transform 1 0 34868 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_373
timestamp 1662439860
transform 1 0 35420 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_379
timestamp 1662439860
transform 1 0 35972 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1662439860
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1662439860
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_405
timestamp 1662439860
transform 1 0 38364 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_410
timestamp 1662439860
transform 1 0 38824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_420
timestamp 1662439860
transform 1 0 39744 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_426
timestamp 1662439860
transform 1 0 40296 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_433
timestamp 1662439860
transform 1 0 40940 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_437
timestamp 1662439860
transform 1 0 41308 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_440
timestamp 1662439860
transform 1 0 41584 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_446
timestamp 1662439860
transform 1 0 42136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_449
timestamp 1662439860
transform 1 0 42412 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_454
timestamp 1662439860
transform 1 0 42872 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_458
timestamp 1662439860
transform 1 0 43240 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_461
timestamp 1662439860
transform 1 0 43516 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_471
timestamp 1662439860
transform 1 0 44436 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_477
timestamp 1662439860
transform 1 0 44988 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_484
timestamp 1662439860
transform 1 0 45632 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_491
timestamp 1662439860
transform 1 0 46276 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_498
timestamp 1662439860
transform 1 0 46920 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_505
timestamp 1662439860
transform 1 0 47564 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_509
timestamp 1662439860
transform 1 0 47932 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_517
timestamp 1662439860
transform 1 0 48668 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_520
timestamp 1662439860
transform 1 0 48944 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_526
timestamp 1662439860
transform 1 0 49496 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_534
timestamp 1662439860
transform 1 0 50232 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1662439860
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_553
timestamp 1662439860
transform 1 0 51980 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_558
timestamp 1662439860
transform 1 0 52440 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_561
timestamp 1662439860
transform 1 0 52716 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_566
timestamp 1662439860
transform 1 0 53176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_572
timestamp 1662439860
transform 1 0 53728 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_578
timestamp 1662439860
transform 1 0 54280 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_584
timestamp 1662439860
transform 1 0 54832 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_587
timestamp 1662439860
transform 1 0 55108 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_593
timestamp 1662439860
transform 1 0 55660 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_604
timestamp 1662439860
transform 1 0 56672 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_610
timestamp 1662439860
transform 1 0 57224 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_617
timestamp 1662439860
transform 1 0 57868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_621
timestamp 1662439860
transform 1 0 58236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_627
timestamp 1662439860
transform 1 0 58788 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_633
timestamp 1662439860
transform 1 0 59340 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_660
timestamp 1662439860
transform 1 0 61824 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_666
timestamp 1662439860
transform 1 0 62376 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_673
timestamp 1662439860
transform 1 0 63020 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_677
timestamp 1662439860
transform 1 0 63388 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_683
timestamp 1662439860
transform 1 0 63940 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_689
timestamp 1662439860
transform 1 0 64492 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_693
timestamp 1662439860
transform 1 0 64860 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_696
timestamp 1662439860
transform 1 0 65136 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_706
timestamp 1662439860
transform 1 0 66056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_716
timestamp 1662439860
transform 1 0 66976 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_722
timestamp 1662439860
transform 1 0 67528 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_729
timestamp 1662439860
transform 1 0 68172 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_733
timestamp 1662439860
transform 1 0 68540 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_739
timestamp 1662439860
transform 1 0 69092 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_743
timestamp 1662439860
transform 1 0 69460 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_746
timestamp 1662439860
transform 1 0 69736 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_752
timestamp 1662439860
transform 1 0 70288 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_755
timestamp 1662439860
transform 1 0 70564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_762
timestamp 1662439860
transform 1 0 71208 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_772
timestamp 1662439860
transform 1 0 72128 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_778
timestamp 1662439860
transform 1 0 72680 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_785
timestamp 1662439860
transform 1 0 73324 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_797
timestamp 1662439860
transform 1 0 74428 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_809
timestamp 1662439860
transform 1 0 75532 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_815
timestamp 1662439860
transform 1 0 76084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_821
timestamp 1662439860
transform 1 0 76636 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_827
timestamp 1662439860
transform 1 0 77188 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_833
timestamp 1662439860
transform 1 0 77740 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_839
timestamp 1662439860
transform 1 0 78292 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_841
timestamp 1662439860
transform 1 0 78476 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_846
timestamp 1662439860
transform 1 0 78936 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_852
timestamp 1662439860
transform 1 0 79488 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_858
timestamp 1662439860
transform 1 0 80040 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_864
timestamp 1662439860
transform 1 0 80592 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_876
timestamp 1662439860
transform 1 0 81696 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_888
timestamp 1662439860
transform 1 0 82800 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_893
timestamp 1662439860
transform 1 0 83260 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_897
timestamp 1662439860
transform 1 0 83628 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_901
timestamp 1662439860
transform 1 0 83996 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_913
timestamp 1662439860
transform 1 0 85100 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_925
timestamp 1662439860
transform 1 0 86204 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_937
timestamp 1662439860
transform 1 0 87308 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_949
timestamp 1662439860
transform 1 0 88412 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_953
timestamp 1662439860
transform 1 0 88780 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_965
timestamp 1662439860
transform 1 0 89884 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_977
timestamp 1662439860
transform 1 0 90988 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_989
timestamp 1662439860
transform 1 0 92092 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1001
timestamp 1662439860
transform 1 0 93196 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1007
timestamp 1662439860
transform 1 0 93748 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1009
timestamp 1662439860
transform 1 0 93932 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1015
timestamp 1662439860
transform 1 0 94484 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1662439860
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_7
timestamp 1662439860
transform 1 0 1748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1662439860
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1662439860
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1662439860
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1662439860
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1662439860
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1662439860
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1662439860
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1662439860
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1662439860
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1662439860
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1662439860
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1662439860
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1662439860
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1662439860
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1662439860
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1662439860
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1662439860
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1662439860
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1662439860
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1662439860
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_197
timestamp 1662439860
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_203
timestamp 1662439860
transform 1 0 19780 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_207
timestamp 1662439860
transform 1 0 20148 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_210
timestamp 1662439860
transform 1 0 20424 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_222
timestamp 1662439860
transform 1 0 21528 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_234
timestamp 1662439860
transform 1 0 22632 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_246
timestamp 1662439860
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1662439860
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1662439860
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1662439860
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1662439860
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1662439860
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1662439860
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1662439860
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_321
timestamp 1662439860
transform 1 0 30636 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_329
timestamp 1662439860
transform 1 0 31372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_334
timestamp 1662439860
transform 1 0 31832 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_340
timestamp 1662439860
transform 1 0 32384 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_344
timestamp 1662439860
transform 1 0 32752 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_347
timestamp 1662439860
transform 1 0 33028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1662439860
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1662439860
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_365
timestamp 1662439860
transform 1 0 34684 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_373
timestamp 1662439860
transform 1 0 35420 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_377
timestamp 1662439860
transform 1 0 35788 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_385
timestamp 1662439860
transform 1 0 36524 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_397
timestamp 1662439860
transform 1 0 37628 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_405
timestamp 1662439860
transform 1 0 38364 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_410
timestamp 1662439860
transform 1 0 38824 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1662439860
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1662439860
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_433
timestamp 1662439860
transform 1 0 40940 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_436
timestamp 1662439860
transform 1 0 41216 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_440
timestamp 1662439860
transform 1 0 41584 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_443
timestamp 1662439860
transform 1 0 41860 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_449
timestamp 1662439860
transform 1 0 42412 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_455
timestamp 1662439860
transform 1 0 42964 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_463
timestamp 1662439860
transform 1 0 43700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1662439860
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_477
timestamp 1662439860
transform 1 0 44988 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_481
timestamp 1662439860
transform 1 0 45356 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_491
timestamp 1662439860
transform 1 0 46276 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_508
timestamp 1662439860
transform 1 0 47840 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_514
timestamp 1662439860
transform 1 0 48392 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_526
timestamp 1662439860
transform 1 0 49496 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_533
timestamp 1662439860
transform 1 0 50140 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_537
timestamp 1662439860
transform 1 0 50508 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_549
timestamp 1662439860
transform 1 0 51612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_557
timestamp 1662439860
transform 1 0 52348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_560
timestamp 1662439860
transform 1 0 52624 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_564
timestamp 1662439860
transform 1 0 52992 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_567
timestamp 1662439860
transform 1 0 53268 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_575
timestamp 1662439860
transform 1 0 54004 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_580
timestamp 1662439860
transform 1 0 54464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_586
timestamp 1662439860
transform 1 0 55016 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_589
timestamp 1662439860
transform 1 0 55292 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_593
timestamp 1662439860
transform 1 0 55660 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_599
timestamp 1662439860
transform 1 0 56212 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_607
timestamp 1662439860
transform 1 0 56948 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_613
timestamp 1662439860
transform 1 0 57500 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_621
timestamp 1662439860
transform 1 0 58236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_627
timestamp 1662439860
transform 1 0 58788 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_633
timestamp 1662439860
transform 1 0 59340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_642
timestamp 1662439860
transform 1 0 60168 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_645
timestamp 1662439860
transform 1 0 60444 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_667
timestamp 1662439860
transform 1 0 62468 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_691
timestamp 1662439860
transform 1 0 64676 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_697
timestamp 1662439860
transform 1 0 65228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_701
timestamp 1662439860
transform 1 0 65596 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_723
timestamp 1662439860
transform 1 0 67620 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_729
timestamp 1662439860
transform 1 0 68172 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_735
timestamp 1662439860
transform 1 0 68724 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_747
timestamp 1662439860
transform 1 0 69828 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_755
timestamp 1662439860
transform 1 0 70564 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_757
timestamp 1662439860
transform 1 0 70748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_769
timestamp 1662439860
transform 1 0 71852 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_772
timestamp 1662439860
transform 1 0 72128 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_784
timestamp 1662439860
transform 1 0 73232 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_796
timestamp 1662439860
transform 1 0 74336 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_808
timestamp 1662439860
transform 1 0 75440 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_813
timestamp 1662439860
transform 1 0 75900 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_821
timestamp 1662439860
transform 1 0 76636 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_826
timestamp 1662439860
transform 1 0 77096 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_838
timestamp 1662439860
transform 1 0 78200 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_850
timestamp 1662439860
transform 1 0 79304 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_862
timestamp 1662439860
transform 1 0 80408 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_869
timestamp 1662439860
transform 1 0 81052 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_881
timestamp 1662439860
transform 1 0 82156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_889
timestamp 1662439860
transform 1 0 82892 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_893
timestamp 1662439860
transform 1 0 83260 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_901
timestamp 1662439860
transform 1 0 83996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_913
timestamp 1662439860
transform 1 0 85100 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_921
timestamp 1662439860
transform 1 0 85836 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_925
timestamp 1662439860
transform 1 0 86204 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_937
timestamp 1662439860
transform 1 0 87308 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_949
timestamp 1662439860
transform 1 0 88412 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_961
timestamp 1662439860
transform 1 0 89516 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_973
timestamp 1662439860
transform 1 0 90620 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_979
timestamp 1662439860
transform 1 0 91172 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_981
timestamp 1662439860
transform 1 0 91356 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_993
timestamp 1662439860
transform 1 0 92460 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_997
timestamp 1662439860
transform 1 0 92828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1003
timestamp 1662439860
transform 1 0 93380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1009
timestamp 1662439860
transform 1 0 93932 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_1014
timestamp 1662439860
transform 1 0 94392 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1662439860
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_11
timestamp 1662439860
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_23
timestamp 1662439860
transform 1 0 3220 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1662439860
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_29
timestamp 1662439860
transform 1 0 3772 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_41
timestamp 1662439860
transform 1 0 4876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_48
timestamp 1662439860
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1662439860
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1662439860
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_81
timestamp 1662439860
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_85
timestamp 1662439860
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_97
timestamp 1662439860
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1662439860
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1662439860
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_121
timestamp 1662439860
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_127
timestamp 1662439860
transform 1 0 12788 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_139
timestamp 1662439860
transform 1 0 13892 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_141
timestamp 1662439860
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_153
timestamp 1662439860
transform 1 0 15180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1662439860
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1662439860
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1662439860
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_193
timestamp 1662439860
transform 1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_197
timestamp 1662439860
transform 1 0 19228 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_212
timestamp 1662439860
transform 1 0 20608 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1662439860
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1662439860
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_249
timestamp 1662439860
transform 1 0 24012 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_253
timestamp 1662439860
transform 1 0 24380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_265
timestamp 1662439860
transform 1 0 25484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1662439860
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1662439860
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_293
timestamp 1662439860
transform 1 0 28060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_298
timestamp 1662439860
transform 1 0 28520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_306
timestamp 1662439860
transform 1 0 29256 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_309
timestamp 1662439860
transform 1 0 29532 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_321
timestamp 1662439860
transform 1 0 30636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_333
timestamp 1662439860
transform 1 0 31740 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1662439860
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_349
timestamp 1662439860
transform 1 0 33212 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_357
timestamp 1662439860
transform 1 0 33948 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_362
timestamp 1662439860
transform 1 0 34408 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_365
timestamp 1662439860
transform 1 0 34684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_390
timestamp 1662439860
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1662439860
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_397
timestamp 1662439860
transform 1 0 37628 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_409
timestamp 1662439860
transform 1 0 38732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_417
timestamp 1662439860
transform 1 0 39468 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_421
timestamp 1662439860
transform 1 0 39836 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_433
timestamp 1662439860
transform 1 0 40940 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_445
timestamp 1662439860
transform 1 0 42044 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_449
timestamp 1662439860
transform 1 0 42412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_453
timestamp 1662439860
transform 1 0 42780 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_463
timestamp 1662439860
transform 1 0 43700 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_470
timestamp 1662439860
transform 1 0 44344 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_477
timestamp 1662439860
transform 1 0 44988 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_485
timestamp 1662439860
transform 1 0 45724 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_488
timestamp 1662439860
transform 1 0 46000 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_492
timestamp 1662439860
transform 1 0 46368 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_495
timestamp 1662439860
transform 1 0 46644 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_501
timestamp 1662439860
transform 1 0 47196 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1662439860
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1662439860
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_529
timestamp 1662439860
transform 1 0 49772 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_533
timestamp 1662439860
transform 1 0 50140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_545
timestamp 1662439860
transform 1 0 51244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_557
timestamp 1662439860
transform 1 0 52348 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1662439860
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1662439860
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_585
timestamp 1662439860
transform 1 0 54924 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_589
timestamp 1662439860
transform 1 0 55292 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_595
timestamp 1662439860
transform 1 0 55844 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_598
timestamp 1662439860
transform 1 0 56120 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_604
timestamp 1662439860
transform 1 0 56672 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_610
timestamp 1662439860
transform 1 0 57224 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1662439860
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_625
timestamp 1662439860
transform 1 0 58604 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_628
timestamp 1662439860
transform 1 0 58880 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_634
timestamp 1662439860
transform 1 0 59432 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_642
timestamp 1662439860
transform 1 0 60168 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_645
timestamp 1662439860
transform 1 0 60444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_655
timestamp 1662439860
transform 1 0 61364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_661
timestamp 1662439860
transform 1 0 61916 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_667
timestamp 1662439860
transform 1 0 62468 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 1662439860
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_673
timestamp 1662439860
transform 1 0 63020 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_677
timestamp 1662439860
transform 1 0 63388 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_683
timestamp 1662439860
transform 1 0 63940 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_689
timestamp 1662439860
transform 1 0 64492 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_695
timestamp 1662439860
transform 1 0 65044 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_699
timestamp 1662439860
transform 1 0 65412 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_701
timestamp 1662439860
transform 1 0 65596 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_705
timestamp 1662439860
transform 1 0 65964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_717
timestamp 1662439860
transform 1 0 67068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_725
timestamp 1662439860
transform 1 0 67804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_729
timestamp 1662439860
transform 1 0 68172 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_735
timestamp 1662439860
transform 1 0 68724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_747
timestamp 1662439860
transform 1 0 69828 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_755
timestamp 1662439860
transform 1 0 70564 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_757
timestamp 1662439860
transform 1 0 70748 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_769
timestamp 1662439860
transform 1 0 71852 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_781
timestamp 1662439860
transform 1 0 72956 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_785
timestamp 1662439860
transform 1 0 73324 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_797
timestamp 1662439860
transform 1 0 74428 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_809
timestamp 1662439860
transform 1 0 75532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_813
timestamp 1662439860
transform 1 0 75900 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_819
timestamp 1662439860
transform 1 0 76452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_831
timestamp 1662439860
transform 1 0 77556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_839
timestamp 1662439860
transform 1 0 78292 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_841
timestamp 1662439860
transform 1 0 78476 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_853
timestamp 1662439860
transform 1 0 79580 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_865
timestamp 1662439860
transform 1 0 80684 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_869
timestamp 1662439860
transform 1 0 81052 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_881
timestamp 1662439860
transform 1 0 82156 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_889
timestamp 1662439860
transform 1 0 82892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_894
timestamp 1662439860
transform 1 0 83352 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_897
timestamp 1662439860
transform 1 0 83628 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_922
timestamp 1662439860
transform 1 0 85928 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_925
timestamp 1662439860
transform 1 0 86204 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_929
timestamp 1662439860
transform 1 0 86572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_941
timestamp 1662439860
transform 1 0 87676 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_949
timestamp 1662439860
transform 1 0 88412 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_953
timestamp 1662439860
transform 1 0 88780 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_965
timestamp 1662439860
transform 1 0 89884 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_977
timestamp 1662439860
transform 1 0 90988 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_981
timestamp 1662439860
transform 1 0 91356 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_986
timestamp 1662439860
transform 1 0 91816 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_992
timestamp 1662439860
transform 1 0 92368 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_1004
timestamp 1662439860
transform 1 0 93472 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1009
timestamp 1662439860
transform 1 0 93932 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1015
timestamp 1662439860
transform 1 0 94484 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1662439860
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1662439860
transform -1 0 94852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1662439860
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1662439860
transform -1 0 94852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1662439860
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1662439860
transform -1 0 94852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1662439860
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1662439860
transform -1 0 94852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1662439860
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1662439860
transform -1 0 94852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1662439860
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1662439860
transform -1 0 94852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1662439860
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1662439860
transform -1 0 94852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1662439860
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1662439860
transform -1 0 94852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1662439860
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1662439860
transform -1 0 94852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1662439860
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1662439860
transform -1 0 94852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1662439860
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1662439860
transform -1 0 94852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1662439860
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1662439860
transform -1 0 94852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1662439860
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1662439860
transform -1 0 94852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1662439860
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1662439860
transform -1 0 94852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1662439860
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1662439860
transform -1 0 94852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1662439860
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1662439860
transform -1 0 94852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1662439860
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1662439860
transform -1 0 94852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1662439860
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1662439860
transform -1 0 94852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1662439860
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1662439860
transform -1 0 94852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1662439860
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1662439860
transform -1 0 94852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1662439860
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1662439860
transform -1 0 94852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1662439860
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1662439860
transform -1 0 94852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1662439860
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1662439860
transform -1 0 94852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1662439860
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1662439860
transform -1 0 94852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1662439860
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1662439860
transform -1 0 94852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1662439860
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1662439860
transform -1 0 94852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1662439860
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1662439860
transform -1 0 94852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1662439860
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1662439860
transform -1 0 94852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1662439860
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1662439860
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1662439860
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1662439860
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1662439860
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1662439860
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1662439860
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1662439860
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1662439860
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1662439860
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1662439860
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1662439860
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1662439860
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1662439860
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1662439860
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1662439860
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1662439860
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1662439860
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1662439860
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1662439860
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1662439860
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1662439860
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1662439860
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1662439860
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1662439860
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1662439860
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1662439860
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1662439860
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1662439860
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1662439860
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1662439860
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1662439860
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1662439860
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1662439860
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1662439860
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1662439860
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1662439860
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1662439860
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1662439860
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1662439860
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1662439860
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1662439860
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1662439860
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1662439860
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1662439860
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1662439860
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1662439860
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1662439860
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1662439860
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1662439860
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1662439860
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1662439860
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1662439860
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1662439860
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1662439860
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1662439860
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1662439860
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1662439860
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1662439860
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1662439860
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1662439860
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1662439860
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1662439860
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1662439860
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1662439860
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1662439860
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1662439860
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1662439860
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1662439860
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1662439860
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1662439860
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1662439860
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1662439860
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1662439860
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1662439860
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1662439860
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1662439860
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1662439860
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1662439860
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1662439860
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1662439860
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1662439860
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1662439860
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1662439860
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1662439860
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1662439860
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1662439860
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1662439860
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1662439860
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1662439860
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1662439860
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1662439860
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1662439860
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1662439860
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1662439860
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1662439860
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1662439860
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1662439860
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1662439860
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1662439860
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1662439860
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1662439860
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1662439860
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1662439860
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1662439860
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1662439860
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1662439860
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1662439860
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1662439860
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1662439860
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1662439860
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1662439860
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1662439860
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1662439860
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1662439860
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1662439860
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1662439860
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1662439860
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1662439860
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1662439860
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1662439860
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1662439860
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1662439860
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1662439860
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1662439860
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1662439860
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1662439860
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1662439860
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1662439860
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1662439860
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1662439860
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1662439860
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1662439860
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1662439860
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1662439860
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1662439860
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1662439860
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1662439860
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1662439860
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1662439860
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1662439860
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1662439860
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1662439860
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1662439860
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1662439860
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1662439860
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1662439860
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1662439860
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1662439860
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1662439860
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1662439860
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1662439860
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1662439860
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1662439860
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1662439860
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1662439860
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1662439860
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1662439860
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1662439860
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1662439860
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1662439860
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1662439860
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1662439860
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1662439860
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1662439860
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1662439860
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1662439860
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1662439860
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1662439860
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1662439860
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1662439860
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1662439860
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1662439860
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1662439860
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1662439860
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1662439860
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1662439860
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1662439860
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1662439860
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1662439860
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1662439860
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1662439860
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1662439860
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1662439860
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1662439860
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1662439860
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1662439860
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1662439860
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1662439860
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1662439860
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1662439860
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1662439860
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1662439860
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1662439860
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1662439860
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1662439860
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1662439860
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1662439860
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1662439860
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1662439860
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1662439860
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1662439860
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1662439860
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1662439860
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1662439860
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1662439860
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1662439860
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1662439860
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1662439860
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1662439860
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1662439860
transform 1 0 70656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1662439860
transform 1 0 75808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1662439860
transform 1 0 80960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1662439860
transform 1 0 86112 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1662439860
transform 1 0 91264 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1662439860
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1662439860
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1662439860
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1662439860
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1662439860
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1662439860
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1662439860
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1662439860
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1662439860
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1662439860
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1662439860
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1662439860
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1662439860
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1662439860
transform 1 0 73232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1662439860
transform 1 0 78384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1662439860
transform 1 0 83536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1662439860
transform 1 0 88688 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1662439860
transform 1 0 93840 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1662439860
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1662439860
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1662439860
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1662439860
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1662439860
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1662439860
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1662439860
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1662439860
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1662439860
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1662439860
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1662439860
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1662439860
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1662439860
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1662439860
transform 1 0 70656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1662439860
transform 1 0 75808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1662439860
transform 1 0 80960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1662439860
transform 1 0 86112 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1662439860
transform 1 0 91264 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1662439860
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1662439860
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1662439860
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1662439860
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1662439860
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1662439860
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1662439860
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1662439860
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1662439860
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1662439860
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1662439860
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1662439860
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1662439860
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1662439860
transform 1 0 73232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1662439860
transform 1 0 78384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1662439860
transform 1 0 83536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1662439860
transform 1 0 88688 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1662439860
transform 1 0 93840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1662439860
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1662439860
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1662439860
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1662439860
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1662439860
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1662439860
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1662439860
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1662439860
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1662439860
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1662439860
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1662439860
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1662439860
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1662439860
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1662439860
transform 1 0 70656 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1662439860
transform 1 0 75808 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1662439860
transform 1 0 80960 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1662439860
transform 1 0 86112 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1662439860
transform 1 0 91264 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1662439860
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1662439860
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1662439860
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1662439860
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1662439860
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1662439860
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1662439860
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1662439860
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1662439860
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1662439860
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1662439860
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1662439860
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1662439860
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1662439860
transform 1 0 73232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1662439860
transform 1 0 78384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1662439860
transform 1 0 83536 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1662439860
transform 1 0 88688 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1662439860
transform 1 0 93840 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1662439860
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1662439860
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1662439860
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1662439860
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1662439860
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1662439860
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1662439860
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1662439860
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1662439860
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1662439860
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1662439860
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1662439860
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1662439860
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1662439860
transform 1 0 70656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1662439860
transform 1 0 75808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1662439860
transform 1 0 80960 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1662439860
transform 1 0 86112 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1662439860
transform 1 0 91264 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1662439860
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1662439860
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1662439860
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1662439860
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1662439860
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1662439860
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1662439860
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1662439860
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1662439860
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1662439860
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1662439860
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1662439860
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1662439860
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1662439860
transform 1 0 73232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1662439860
transform 1 0 78384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1662439860
transform 1 0 83536 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1662439860
transform 1 0 88688 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1662439860
transform 1 0 93840 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1662439860
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1662439860
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1662439860
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1662439860
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1662439860
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1662439860
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1662439860
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1662439860
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1662439860
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1662439860
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1662439860
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1662439860
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1662439860
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1662439860
transform 1 0 70656 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1662439860
transform 1 0 75808 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1662439860
transform 1 0 80960 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1662439860
transform 1 0 86112 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1662439860
transform 1 0 91264 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1662439860
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1662439860
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1662439860
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1662439860
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1662439860
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1662439860
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1662439860
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1662439860
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1662439860
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1662439860
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1662439860
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1662439860
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1662439860
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1662439860
transform 1 0 73232 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1662439860
transform 1 0 78384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1662439860
transform 1 0 83536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1662439860
transform 1 0 88688 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1662439860
transform 1 0 93840 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1662439860
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1662439860
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1662439860
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1662439860
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1662439860
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1662439860
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1662439860
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1662439860
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1662439860
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1662439860
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1662439860
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1662439860
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1662439860
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1662439860
transform 1 0 70656 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1662439860
transform 1 0 75808 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1662439860
transform 1 0 80960 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1662439860
transform 1 0 86112 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1662439860
transform 1 0 91264 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1662439860
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1662439860
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1662439860
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1662439860
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1662439860
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1662439860
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1662439860
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1662439860
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1662439860
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1662439860
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1662439860
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1662439860
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1662439860
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1662439860
transform 1 0 73232 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1662439860
transform 1 0 78384 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1662439860
transform 1 0 83536 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1662439860
transform 1 0 88688 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1662439860
transform 1 0 93840 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1662439860
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1662439860
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1662439860
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1662439860
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1662439860
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1662439860
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1662439860
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1662439860
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1662439860
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1662439860
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1662439860
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1662439860
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1662439860
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1662439860
transform 1 0 70656 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1662439860
transform 1 0 75808 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1662439860
transform 1 0 80960 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1662439860
transform 1 0 86112 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1662439860
transform 1 0 91264 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1662439860
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1662439860
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1662439860
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1662439860
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1662439860
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1662439860
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1662439860
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1662439860
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1662439860
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1662439860
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1662439860
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1662439860
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1662439860
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1662439860
transform 1 0 73232 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1662439860
transform 1 0 78384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1662439860
transform 1 0 83536 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1662439860
transform 1 0 88688 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1662439860
transform 1 0 93840 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1662439860
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1662439860
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1662439860
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1662439860
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1662439860
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1662439860
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1662439860
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1662439860
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1662439860
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1662439860
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1662439860
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1662439860
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1662439860
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1662439860
transform 1 0 70656 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1662439860
transform 1 0 75808 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1662439860
transform 1 0 80960 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1662439860
transform 1 0 86112 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1662439860
transform 1 0 91264 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1662439860
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1662439860
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1662439860
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1662439860
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1662439860
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1662439860
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1662439860
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1662439860
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1662439860
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1662439860
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1662439860
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1662439860
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1662439860
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1662439860
transform 1 0 73232 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1662439860
transform 1 0 78384 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1662439860
transform 1 0 83536 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1662439860
transform 1 0 88688 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1662439860
transform 1 0 93840 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1662439860
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1662439860
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1662439860
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1662439860
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1662439860
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1662439860
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1662439860
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1662439860
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1662439860
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1662439860
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1662439860
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1662439860
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1662439860
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1662439860
transform 1 0 70656 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1662439860
transform 1 0 75808 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1662439860
transform 1 0 80960 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1662439860
transform 1 0 86112 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1662439860
transform 1 0 91264 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1662439860
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1662439860
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1662439860
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1662439860
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1662439860
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1662439860
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1662439860
transform 1 0 19136 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1662439860
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1662439860
transform 1 0 24288 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1662439860
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1662439860
transform 1 0 29440 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1662439860
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1662439860
transform 1 0 34592 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1662439860
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1662439860
transform 1 0 39744 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1662439860
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1662439860
transform 1 0 44896 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1662439860
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1662439860
transform 1 0 50048 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1662439860
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1662439860
transform 1 0 55200 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1662439860
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1662439860
transform 1 0 60352 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1662439860
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1662439860
transform 1 0 65504 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1662439860
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1662439860
transform 1 0 70656 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1662439860
transform 1 0 73232 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1662439860
transform 1 0 75808 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1662439860
transform 1 0 78384 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1662439860
transform 1 0 80960 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1662439860
transform 1 0 83536 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1662439860
transform 1 0 86112 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1662439860
transform 1 0 88688 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1662439860
transform 1 0 91264 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1662439860
transform 1 0 93840 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0445_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 21620 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0446__1 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 33120 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0446__2
timestamp 1662439860
transform -1 0 35144 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0447_
timestamp 1662439860
transform -1 0 24840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0448__6
timestamp 1662439860
transform -1 0 20240 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0449__7
timestamp 1662439860
transform -1 0 29256 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0450__8
timestamp 1662439860
transform -1 0 28612 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0451__9
timestamp 1662439860
transform -1 0 25760 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0452__10
timestamp 1662439860
transform 1 0 30452 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0453__11
timestamp 1662439860
transform -1 0 18952 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0454__12
timestamp 1662439860
transform -1 0 20884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0455__13
timestamp 1662439860
transform -1 0 20884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0456__14
timestamp 1662439860
transform 1 0 22632 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0457__15
timestamp 1662439860
transform -1 0 19780 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0458_
timestamp 1662439860
transform 1 0 66424 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0459__16
timestamp 1662439860
transform -1 0 66884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0460__17
timestamp 1662439860
transform -1 0 71208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0461__18
timestamp 1662439860
transform 1 0 80040 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0462__19
timestamp 1662439860
transform 1 0 79948 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0463__20
timestamp 1662439860
transform -1 0 65320 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0464__21
timestamp 1662439860
transform -1 0 79672 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0465__22
timestamp 1662439860
transform -1 0 78936 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466__23
timestamp 1662439860
transform 1 0 71484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0467__24
timestamp 1662439860
transform -1 0 78936 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0468_
timestamp 1662439860
transform -1 0 89608 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0469_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 76636 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0470_
timestamp 1662439860
transform -1 0 87952 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0471_
timestamp 1662439860
transform -1 0 84916 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1662439860
transform 1 0 58052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0473_
timestamp 1662439860
transform 1 0 76912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0474_
timestamp 1662439860
transform -1 0 58972 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0475_
timestamp 1662439860
transform 1 0 94116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0476_
timestamp 1662439860
transform 1 0 94116 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0477_
timestamp 1662439860
transform -1 0 75348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1662439860
transform 1 0 58052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1662439860
transform -1 0 81512 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0480_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 82892 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0481_
timestamp 1662439860
transform -1 0 73784 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0482_
timestamp 1662439860
transform -1 0 85560 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0483_
timestamp 1662439860
transform -1 0 70472 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1662439860
transform -1 0 54556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1662439860
transform -1 0 75532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0486_
timestamp 1662439860
transform 1 0 82248 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0487_
timestamp 1662439860
transform 1 0 87676 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0488_
timestamp 1662439860
transform 1 0 84088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0489_
timestamp 1662439860
transform -1 0 55936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490__25
timestamp 1662439860
transform -1 0 71208 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0491_
timestamp 1662439860
transform -1 0 22908 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0492__26
timestamp 1662439860
transform -1 0 15732 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0493__27
timestamp 1662439860
transform -1 0 16008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0494__28
timestamp 1662439860
transform 1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0495_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 15548 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0496_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3956 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _0497_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3956 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0498_
timestamp 1662439860
transform 1 0 14260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0499_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 15916 0 1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_1  _0500_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 3220 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0501_
timestamp 1662439860
transform -1 0 19320 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _0502_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 16928 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1662439860
transform -1 0 6808 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0504_
timestamp 1662439860
transform -1 0 12788 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  _0505_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 4324 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__xnor2_4  _0506_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 11592 0 1 13056
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0507_
timestamp 1662439860
transform 1 0 45356 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0508_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 4232 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0509_
timestamp 1662439860
transform -1 0 3496 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0510_
timestamp 1662439860
transform 1 0 3956 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0511_
timestamp 1662439860
transform 1 0 25116 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0512_
timestamp 1662439860
transform 1 0 10120 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _0513_
timestamp 1662439860
transform -1 0 55568 0 -1 11968
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1662439860
transform -1 0 79672 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0515_
timestamp 1662439860
transform 1 0 27968 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0516_
timestamp 1662439860
transform 1 0 24932 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _0517_
timestamp 1662439860
transform 1 0 40020 0 1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0518_
timestamp 1662439860
transform 1 0 78292 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0519_
timestamp 1662439860
transform 1 0 48852 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _0520_
timestamp 1662439860
transform 1 0 6256 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_4  _0521_
timestamp 1662439860
transform 1 0 81604 0 1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_6  _0522_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 77556 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0523_
timestamp 1662439860
transform -1 0 11132 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_2  _0524_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 36248 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _0525_
timestamp 1662439860
transform 1 0 27048 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0526_
timestamp 1662439860
transform 1 0 20148 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_4  _0527_
timestamp 1662439860
transform 1 0 51888 0 1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1662439860
transform 1 0 78936 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0529_
timestamp 1662439860
transform 1 0 48484 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0530_
timestamp 1662439860
transform 1 0 31096 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_4  _0531_
timestamp 1662439860
transform 1 0 46092 0 1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1662439860
transform 1 0 75348 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0533_
timestamp 1662439860
transform -1 0 59708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0534_
timestamp 1662439860
transform 1 0 46736 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0535_
timestamp 1662439860
transform 1 0 30360 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_4  _0536_
timestamp 1662439860
transform 1 0 50508 0 1 11968
box -38 -48 2062 592
use sky130_fd_sc_hd__or4_4  _0537_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 59064 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0538_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 12972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0539_
timestamp 1662439860
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0540_
timestamp 1662439860
transform 1 0 9844 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0541_
timestamp 1662439860
transform 1 0 13064 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0542_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 9752 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0543_
timestamp 1662439860
transform 1 0 6532 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0544_
timestamp 1662439860
transform 1 0 8004 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0545_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 55752 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0546_
timestamp 1662439860
transform -1 0 51520 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0547_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 52900 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0548_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 14996 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0549_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 41032 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0550_
timestamp 1662439860
transform -1 0 26496 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0551_
timestamp 1662439860
transform -1 0 34040 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0552_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 68356 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0553_
timestamp 1662439860
transform -1 0 57408 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0554_
timestamp 1662439860
transform 1 0 57776 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0555_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 61456 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0556_
timestamp 1662439860
transform -1 0 27784 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0557_
timestamp 1662439860
transform -1 0 29716 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0558_
timestamp 1662439860
transform 1 0 52900 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0559_
timestamp 1662439860
transform 1 0 54096 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0560_
timestamp 1662439860
transform -1 0 57408 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0561_
timestamp 1662439860
transform 1 0 53360 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0562_
timestamp 1662439860
transform -1 0 39192 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0563_
timestamp 1662439860
transform -1 0 48392 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1662439860
transform 1 0 78660 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0565_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 52440 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0566_
timestamp 1662439860
transform -1 0 43240 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0567_
timestamp 1662439860
transform 1 0 42596 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0568_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 49772 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0569_
timestamp 1662439860
transform -1 0 8648 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0570_
timestamp 1662439860
transform 1 0 32384 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_6  _0571_
timestamp 1662439860
transform 1 0 47932 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _0572_
timestamp 1662439860
transform -1 0 8648 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _0573_
timestamp 1662439860
transform -1 0 86756 0 -1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1662439860
transform 1 0 84916 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0575_
timestamp 1662439860
transform -1 0 6072 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0576_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 8832 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _0577_
timestamp 1662439860
transform 1 0 6624 0 1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_4  _0578_
timestamp 1662439860
transform 1 0 51796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0579_
timestamp 1662439860
transform 1 0 15824 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0580_
timestamp 1662439860
transform -1 0 87584 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  _0581_
timestamp 1662439860
transform 1 0 86664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0582_
timestamp 1662439860
transform -1 0 84272 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _0583_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 56764 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0584_
timestamp 1662439860
transform -1 0 13340 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0585_
timestamp 1662439860
transform 1 0 41400 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0586_
timestamp 1662439860
transform 1 0 44528 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0587_
timestamp 1662439860
transform 1 0 12696 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0588_
timestamp 1662439860
transform 1 0 79672 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _0589_
timestamp 1662439860
transform 1 0 81052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0590_
timestamp 1662439860
transform -1 0 84824 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0591_
timestamp 1662439860
transform -1 0 15272 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0592_
timestamp 1662439860
transform 1 0 41492 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1662439860
transform 1 0 58052 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0594_
timestamp 1662439860
transform 1 0 37720 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1662439860
transform -1 0 36156 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1662439860
transform 1 0 27600 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0597_
timestamp 1662439860
transform -1 0 23552 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0598_
timestamp 1662439860
transform 1 0 38824 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0599_
timestamp 1662439860
transform -1 0 12604 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1662439860
transform -1 0 68632 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1662439860
transform 1 0 69092 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0602_
timestamp 1662439860
transform 1 0 54372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 1662439860
transform -1 0 52808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0604_
timestamp 1662439860
transform -1 0 82340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1662439860
transform 1 0 83076 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0606_
timestamp 1662439860
transform -1 0 89608 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1662439860
transform -1 0 90620 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0608_
timestamp 1662439860
transform 1 0 87952 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1662439860
transform -1 0 86664 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0610_
timestamp 1662439860
transform 1 0 72680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 1662439860
transform -1 0 74888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0612_
timestamp 1662439860
transform -1 0 49864 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0613_
timestamp 1662439860
transform 1 0 52072 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0614_
timestamp 1662439860
transform 1 0 67896 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0615_
timestamp 1662439860
transform -1 0 63572 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1662439860
transform -1 0 86296 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0617_
timestamp 1662439860
transform -1 0 84180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 1662439860
transform -1 0 71208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0619_
timestamp 1662439860
transform 1 0 69736 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1662439860
transform 1 0 86020 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1662439860
transform -1 0 80592 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0622_
timestamp 1662439860
transform 1 0 57224 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1662439860
transform -1 0 55016 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 1662439860
transform -1 0 69828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0625_
timestamp 1662439860
transform 1 0 73876 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1662439860
transform 1 0 94116 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1662439860
transform 1 0 93748 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1662439860
transform 1 0 93840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0629_
timestamp 1662439860
transform -1 0 90252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0630_
timestamp 1662439860
transform -1 0 57408 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1662439860
transform 1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1662439860
transform -1 0 79212 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0633_
timestamp 1662439860
transform -1 0 78200 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1662439860
transform -1 0 60812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0635_
timestamp 1662439860
transform 1 0 64400 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0636_
timestamp 1662439860
transform 1 0 84640 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1662439860
transform -1 0 83352 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1662439860
transform 1 0 88964 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0639_
timestamp 1662439860
transform 1 0 85560 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1662439860
transform -1 0 90068 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1662439860
transform 1 0 93196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0642_
timestamp 1662439860
transform 1 0 19504 0 -1 7616
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1662439860
transform 1 0 49128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _0644_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 80960 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0645_
timestamp 1662439860
transform -1 0 21252 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0646_
timestamp 1662439860
transform 1 0 69460 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0647_
timestamp 1662439860
transform -1 0 59708 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0648_
timestamp 1662439860
transform -1 0 61456 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0649_
timestamp 1662439860
transform -1 0 62744 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0650_
timestamp 1662439860
transform 1 0 65780 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1662439860
transform 1 0 94116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0652_
timestamp 1662439860
transform 1 0 14260 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0653_
timestamp 1662439860
transform -1 0 9384 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0654_
timestamp 1662439860
transform 1 0 6716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1662439860
transform -1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1662439860
transform -1 0 8648 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1662439860
transform -1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0658_
timestamp 1662439860
transform 1 0 11684 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1662439860
transform -1 0 5428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0660_
timestamp 1662439860
transform 1 0 60628 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1662439860
transform 1 0 67528 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0662_
timestamp 1662439860
transform 1 0 61548 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 1662439860
transform 1 0 69828 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1662439860
transform -1 0 66700 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1662439860
transform 1 0 76084 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1662439860
transform 1 0 77372 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1662439860
transform -1 0 77004 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1662439860
transform 1 0 66424 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1662439860
transform 1 0 60628 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0670_
timestamp 1662439860
transform 1 0 76728 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 1662439860
transform -1 0 58972 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1662439860
transform -1 0 79580 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1662439860
transform -1 0 75716 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1662439860
transform 1 0 76268 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1662439860
transform 1 0 75624 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1662439860
transform -1 0 67804 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0677_
timestamp 1662439860
transform -1 0 66148 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1662439860
transform 1 0 40848 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1662439860
transform -1 0 40940 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1662439860
transform 1 0 39192 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1662439860
transform -1 0 31740 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1662439860
transform 1 0 45356 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1662439860
transform -1 0 29072 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1662439860
transform 1 0 46644 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1662439860
transform -1 0 35144 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1662439860
transform -1 0 35236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1662439860
transform 1 0 43700 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1662439860
transform -1 0 36984 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1662439860
transform 1 0 38272 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1662439860
transform -1 0 32568 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1662439860
transform 1 0 52900 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1662439860
transform -1 0 36156 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1662439860
transform 1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1662439860
transform 1 0 46000 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1662439860
transform -1 0 38364 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1662439860
transform 1 0 29808 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1662439860
transform -1 0 30912 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0698_
timestamp 1662439860
transform 1 0 35880 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1662439860
transform -1 0 35512 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0700_
timestamp 1662439860
transform 1 0 34776 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0701_
timestamp 1662439860
transform 1 0 31832 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0702_
timestamp 1662439860
transform 1 0 42596 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0703_
timestamp 1662439860
transform 1 0 70932 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0704_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 53912 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0705_
timestamp 1662439860
transform -1 0 49864 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0706_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 49220 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0707_
timestamp 1662439860
transform 1 0 64308 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0708_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 66424 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0709_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 53820 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0710_
timestamp 1662439860
transform -1 0 49680 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0711_
timestamp 1662439860
transform 1 0 49588 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0712_
timestamp 1662439860
transform -1 0 61180 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0713_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 63204 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _0714_
timestamp 1662439860
transform 1 0 4508 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_4  _0715_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 21068 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0716_
timestamp 1662439860
transform 1 0 63388 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0717_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 67344 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0718_
timestamp 1662439860
transform 1 0 67252 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0719_
timestamp 1662439860
transform -1 0 60168 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0720_
timestamp 1662439860
transform -1 0 62652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0721_
timestamp 1662439860
transform 1 0 19964 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0722_
timestamp 1662439860
transform -1 0 59432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0723_
timestamp 1662439860
transform 1 0 59340 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0724_
timestamp 1662439860
transform 1 0 65136 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0725_
timestamp 1662439860
transform -1 0 66056 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0726_
timestamp 1662439860
transform 1 0 69368 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0727_
timestamp 1662439860
transform 1 0 64492 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0728_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 61548 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0729_
timestamp 1662439860
transform 1 0 62652 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0730_
timestamp 1662439860
transform -1 0 69000 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0731_
timestamp 1662439860
transform 1 0 35972 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0732_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 61640 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0733_
timestamp 1662439860
transform -1 0 60812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0734_
timestamp 1662439860
transform 1 0 60628 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0735_
timestamp 1662439860
transform 1 0 59340 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0736_
timestamp 1662439860
transform -1 0 60076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0737_
timestamp 1662439860
transform 1 0 61640 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0738_
timestamp 1662439860
transform -1 0 49220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0739_
timestamp 1662439860
transform 1 0 50600 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0740_
timestamp 1662439860
transform 1 0 51244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0741_
timestamp 1662439860
transform 1 0 51520 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0742_
timestamp 1662439860
transform 1 0 47932 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0743_
timestamp 1662439860
transform -1 0 46460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0744_
timestamp 1662439860
transform -1 0 44804 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0745_
timestamp 1662439860
transform 1 0 48668 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0746_
timestamp 1662439860
transform -1 0 50876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0747_
timestamp 1662439860
transform 1 0 40756 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0748_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 50048 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0749_
timestamp 1662439860
transform 1 0 50876 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0750_
timestamp 1662439860
transform 1 0 55476 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1662439860
transform -1 0 49312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0752_
timestamp 1662439860
transform 1 0 47748 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0753_
timestamp 1662439860
transform -1 0 44712 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0754_
timestamp 1662439860
transform -1 0 43240 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0755_
timestamp 1662439860
transform 1 0 43424 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0756_
timestamp 1662439860
transform -1 0 47840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0757_
timestamp 1662439860
transform 1 0 45816 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0758_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 58420 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0759_
timestamp 1662439860
transform -1 0 57960 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0760_
timestamp 1662439860
transform -1 0 57316 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0761_
timestamp 1662439860
transform 1 0 56580 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0762_
timestamp 1662439860
transform 1 0 55844 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0763_
timestamp 1662439860
transform -1 0 57224 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0764_
timestamp 1662439860
transform 1 0 56580 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0765_
timestamp 1662439860
transform 1 0 60628 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0766_
timestamp 1662439860
transform 1 0 65780 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0767_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 72680 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0768_
timestamp 1662439860
transform 1 0 74520 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0769_
timestamp 1662439860
transform 1 0 64492 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0770_
timestamp 1662439860
transform -1 0 54096 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _0771_
timestamp 1662439860
transform -1 0 83260 0 1 7616
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0772_
timestamp 1662439860
transform -1 0 92184 0 -1 13056
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _0773_
timestamp 1662439860
transform 1 0 86388 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0774_
timestamp 1662439860
transform -1 0 73416 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0775_
timestamp 1662439860
transform 1 0 50508 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0776_
timestamp 1662439860
transform -1 0 67712 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0777_
timestamp 1662439860
transform -1 0 88228 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0778_
timestamp 1662439860
transform 1 0 65780 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0779_
timestamp 1662439860
transform 1 0 81512 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__or4_2  _0780_
timestamp 1662439860
transform -1 0 84732 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0781_
timestamp 1662439860
transform -1 0 73784 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0782_
timestamp 1662439860
transform -1 0 75624 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0783_
timestamp 1662439860
transform 1 0 75992 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0784_
timestamp 1662439860
transform 1 0 84364 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0785_
timestamp 1662439860
transform -1 0 84456 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0786_
timestamp 1662439860
transform 1 0 74152 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0787_
timestamp 1662439860
transform 1 0 76084 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0788_
timestamp 1662439860
transform -1 0 76820 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0789_
timestamp 1662439860
transform 1 0 81236 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0790_
timestamp 1662439860
transform 1 0 82800 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0791_
timestamp 1662439860
transform 1 0 82708 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0792_
timestamp 1662439860
transform 1 0 79672 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0793_
timestamp 1662439860
transform -1 0 80040 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0794_
timestamp 1662439860
transform 1 0 80408 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0795_
timestamp 1662439860
transform 1 0 80132 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0796_
timestamp 1662439860
transform -1 0 78936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0797_
timestamp 1662439860
transform -1 0 78200 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0798_
timestamp 1662439860
transform 1 0 78660 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0799_
timestamp 1662439860
transform 1 0 77188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0800_
timestamp 1662439860
transform -1 0 76820 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0801_
timestamp 1662439860
transform -1 0 75624 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0802_
timestamp 1662439860
transform -1 0 74796 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0803_
timestamp 1662439860
transform 1 0 75256 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0804_
timestamp 1662439860
transform -1 0 73784 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0805_
timestamp 1662439860
transform -1 0 72772 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0806_
timestamp 1662439860
transform -1 0 76268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0807_
timestamp 1662439860
transform 1 0 74336 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0808_
timestamp 1662439860
transform -1 0 66976 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0809_
timestamp 1662439860
transform -1 0 76912 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0810_
timestamp 1662439860
transform 1 0 77096 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0811_
timestamp 1662439860
transform 1 0 77556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0812_
timestamp 1662439860
transform 1 0 79028 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0813_
timestamp 1662439860
transform 1 0 74980 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0814_
timestamp 1662439860
transform -1 0 74428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0815_
timestamp 1662439860
transform -1 0 72864 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0816_
timestamp 1662439860
transform -1 0 73784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0817_
timestamp 1662439860
transform 1 0 71208 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0818_
timestamp 1662439860
transform -1 0 72680 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0819_
timestamp 1662439860
transform -1 0 73876 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0820_
timestamp 1662439860
transform -1 0 72312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0821_
timestamp 1662439860
transform -1 0 71852 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1662439860
transform 1 0 77372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0823_
timestamp 1662439860
transform 1 0 79120 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0824_
timestamp 1662439860
transform -1 0 78752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0825_
timestamp 1662439860
transform 1 0 78660 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0826_
timestamp 1662439860
transform -1 0 78108 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0827_
timestamp 1662439860
transform 1 0 76728 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0828_
timestamp 1662439860
transform 1 0 89976 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0829_
timestamp 1662439860
transform -1 0 89884 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0830_
timestamp 1662439860
transform 1 0 92828 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _0831_
timestamp 1662439860
transform 1 0 64492 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0832_
timestamp 1662439860
transform -1 0 91080 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0833_
timestamp 1662439860
transform 1 0 91816 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0834_
timestamp 1662439860
transform 1 0 85652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0835_
timestamp 1662439860
transform -1 0 87492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0836_
timestamp 1662439860
transform 1 0 88412 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0837_
timestamp 1662439860
transform 1 0 82708 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0838_
timestamp 1662439860
transform -1 0 84824 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0839_
timestamp 1662439860
transform 1 0 90620 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0840_
timestamp 1662439860
transform 1 0 78476 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0841_
timestamp 1662439860
transform 1 0 55844 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0842_
timestamp 1662439860
transform 1 0 73508 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0843_
timestamp 1662439860
transform 1 0 92092 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0844_
timestamp 1662439860
transform -1 0 93012 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0845_
timestamp 1662439860
transform 1 0 60628 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0846_
timestamp 1662439860
transform 1 0 79212 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0847_
timestamp 1662439860
transform 1 0 63112 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0848_
timestamp 1662439860
transform -1 0 85008 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0849_
timestamp 1662439860
transform 1 0 86388 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0850_
timestamp 1662439860
transform 1 0 92000 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _0851_
timestamp 1662439860
transform 1 0 57040 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0852_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 58512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0853_
timestamp 1662439860
transform 1 0 56120 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0854_
timestamp 1662439860
transform 1 0 57684 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0855_
timestamp 1662439860
transform 1 0 54740 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0856_
timestamp 1662439860
transform 1 0 66424 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0857_
timestamp 1662439860
transform -1 0 68172 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0858_
timestamp 1662439860
transform 1 0 65504 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0859_
timestamp 1662439860
transform 1 0 65780 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0860_
timestamp 1662439860
transform 1 0 67252 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0861_
timestamp 1662439860
transform -1 0 92828 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0862_
timestamp 1662439860
transform -1 0 78108 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0863_
timestamp 1662439860
transform 1 0 75072 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0864_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 74060 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0865_
timestamp 1662439860
transform 1 0 54280 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0866_
timestamp 1662439860
transform -1 0 57592 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0867_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 58972 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0868_
timestamp 1662439860
transform 1 0 71576 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0869_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 72128 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0870_
timestamp 1662439860
transform -1 0 57592 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0871_
timestamp 1662439860
transform 1 0 71024 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0872_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 78936 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0873_
timestamp 1662439860
transform 1 0 75348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _0874_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 76084 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0875_
timestamp 1662439860
transform -1 0 77556 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0876_
timestamp 1662439860
transform 1 0 77372 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _0877_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 77464 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _0878_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 78568 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0879_
timestamp 1662439860
transform -1 0 83352 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0880_
timestamp 1662439860
transform 1 0 15180 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0881_
timestamp 1662439860
transform 1 0 14260 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _0882_
timestamp 1662439860
transform 1 0 9016 0 -1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0883_
timestamp 1662439860
transform 1 0 11224 0 1 7616
box -38 -48 2062 592
use sky130_fd_sc_hd__or4_1  _0884_
timestamp 1662439860
transform -1 0 23184 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0885_
timestamp 1662439860
transform 1 0 23460 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0886_
timestamp 1662439860
transform 1 0 42688 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0887_
timestamp 1662439860
transform 1 0 48484 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0888_
timestamp 1662439860
transform -1 0 48392 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0889_
timestamp 1662439860
transform -1 0 22264 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0890_
timestamp 1662439860
transform 1 0 28520 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0891_
timestamp 1662439860
transform -1 0 43240 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0892_
timestamp 1662439860
transform 1 0 42596 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0893_
timestamp 1662439860
transform -1 0 49404 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0894_
timestamp 1662439860
transform 1 0 46184 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0895_
timestamp 1662439860
transform -1 0 45632 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0896_
timestamp 1662439860
transform 1 0 51980 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0897_
timestamp 1662439860
transform 1 0 53912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0898_
timestamp 1662439860
transform 1 0 53176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0899_
timestamp 1662439860
transform -1 0 56120 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0900_
timestamp 1662439860
transform 1 0 52072 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0901_
timestamp 1662439860
transform 1 0 50968 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0902_
timestamp 1662439860
transform -1 0 50140 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0903_
timestamp 1662439860
transform 1 0 47748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0904_
timestamp 1662439860
transform -1 0 47288 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0905_
timestamp 1662439860
transform -1 0 47196 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0906_
timestamp 1662439860
transform -1 0 45908 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0907_
timestamp 1662439860
transform 1 0 40296 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0908_
timestamp 1662439860
transform -1 0 38456 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0909_
timestamp 1662439860
transform -1 0 37812 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0910_
timestamp 1662439860
transform 1 0 40480 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0911_
timestamp 1662439860
transform -1 0 41860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0912_
timestamp 1662439860
transform -1 0 43056 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0913_
timestamp 1662439860
transform -1 0 40388 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0914_
timestamp 1662439860
transform 1 0 40020 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0915_
timestamp 1662439860
transform -1 0 42136 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0916_
timestamp 1662439860
transform -1 0 40388 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0917_
timestamp 1662439860
transform -1 0 41400 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0918_
timestamp 1662439860
transform -1 0 41216 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0919_
timestamp 1662439860
transform -1 0 40940 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0920_
timestamp 1662439860
transform 1 0 39100 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0921_
timestamp 1662439860
transform 1 0 38916 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0922_
timestamp 1662439860
transform -1 0 39376 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0923_
timestamp 1662439860
transform -1 0 23092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0924_
timestamp 1662439860
transform 1 0 45172 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0925_
timestamp 1662439860
transform -1 0 45816 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1662439860
transform -1 0 20700 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0927_
timestamp 1662439860
transform -1 0 19964 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0928_
timestamp 1662439860
transform 1 0 20332 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0929_
timestamp 1662439860
transform 1 0 23460 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0930_
timestamp 1662439860
transform -1 0 18768 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0931_
timestamp 1662439860
transform 1 0 19412 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0932_
timestamp 1662439860
transform 1 0 22540 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0933_
timestamp 1662439860
transform 1 0 23276 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0934_
timestamp 1662439860
transform 1 0 25944 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0935_
timestamp 1662439860
transform -1 0 25944 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0936_
timestamp 1662439860
transform -1 0 27784 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0937_
timestamp 1662439860
transform 1 0 24748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0938_
timestamp 1662439860
transform -1 0 25576 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0939_
timestamp 1662439860
transform -1 0 32936 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0940_
timestamp 1662439860
transform 1 0 43700 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0941_
timestamp 1662439860
transform 1 0 45172 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0942_
timestamp 1662439860
transform -1 0 41400 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0943_
timestamp 1662439860
transform -1 0 33580 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0944_
timestamp 1662439860
transform -1 0 56764 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0945_
timestamp 1662439860
transform -1 0 51244 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _0946_
timestamp 1662439860
transform -1 0 69092 0 1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _0947_
timestamp 1662439860
transform -1 0 73048 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0948_
timestamp 1662439860
transform 1 0 55660 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0949_
timestamp 1662439860
transform -1 0 62744 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _0950_
timestamp 1662439860
transform -1 0 83352 0 -1 13056
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _0951_
timestamp 1662439860
transform -1 0 71760 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _0952_
timestamp 1662439860
transform -1 0 70380 0 -1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _0953_
timestamp 1662439860
transform 1 0 40020 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__or4_2  _0954_
timestamp 1662439860
transform -1 0 28060 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0955_
timestamp 1662439860
transform -1 0 21988 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0956_
timestamp 1662439860
transform 1 0 19412 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0957_
timestamp 1662439860
transform 1 0 38824 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0958_
timestamp 1662439860
transform -1 0 44712 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0959_
timestamp 1662439860
transform -1 0 29164 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0960_
timestamp 1662439860
transform -1 0 22080 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0961_
timestamp 1662439860
transform -1 0 18768 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _0962_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 18216 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_1  _0963_
timestamp 1662439860
transform -1 0 44712 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0964_
timestamp 1662439860
transform 1 0 43332 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0965_
timestamp 1662439860
transform -1 0 39468 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0966_
timestamp 1662439860
transform 1 0 41768 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0967_
timestamp 1662439860
transform -1 0 41400 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0968_
timestamp 1662439860
transform 1 0 42596 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0969_
timestamp 1662439860
transform -1 0 44252 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0970_
timestamp 1662439860
transform -1 0 46552 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0971_
timestamp 1662439860
transform -1 0 45908 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0972_
timestamp 1662439860
transform -1 0 47564 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0973_
timestamp 1662439860
transform -1 0 18308 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0974_
timestamp 1662439860
transform 1 0 39836 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0975_
timestamp 1662439860
transform -1 0 40388 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0976_
timestamp 1662439860
transform -1 0 38824 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0977_
timestamp 1662439860
transform -1 0 19412 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0978_
timestamp 1662439860
transform 1 0 19412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0979_
timestamp 1662439860
transform 1 0 20516 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0980_
timestamp 1662439860
transform -1 0 16376 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0981_
timestamp 1662439860
transform 1 0 15824 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0982_
timestamp 1662439860
transform 1 0 16836 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0983_
timestamp 1662439860
transform -1 0 17756 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0984_
timestamp 1662439860
transform 1 0 15824 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0985_
timestamp 1662439860
transform 1 0 16744 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0986_
timestamp 1662439860
transform 1 0 17296 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0987_
timestamp 1662439860
transform 1 0 17480 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0988_
timestamp 1662439860
transform -1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0989_
timestamp 1662439860
transform 1 0 13984 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0990_
timestamp 1662439860
transform -1 0 22632 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0991_
timestamp 1662439860
transform -1 0 20700 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0992_
timestamp 1662439860
transform 1 0 20424 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0993_
timestamp 1662439860
transform -1 0 20148 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0994_
timestamp 1662439860
transform 1 0 23000 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0995_
timestamp 1662439860
transform 1 0 21988 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1662439860
transform -1 0 19136 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0997_
timestamp 1662439860
transform 1 0 19412 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0998_
timestamp 1662439860
transform -1 0 18492 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0999_
timestamp 1662439860
transform 1 0 18952 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1000_
timestamp 1662439860
transform -1 0 18860 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1001_
timestamp 1662439860
transform 1 0 14536 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1002_
timestamp 1662439860
transform 1 0 34040 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1003_
timestamp 1662439860
transform 1 0 35328 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1004_
timestamp 1662439860
transform 1 0 37444 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1005_
timestamp 1662439860
transform 1 0 33856 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1006_
timestamp 1662439860
transform 1 0 28244 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1007_
timestamp 1662439860
transform 1 0 36156 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1008_
timestamp 1662439860
transform 1 0 36064 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1009_
timestamp 1662439860
transform -1 0 36064 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1010_
timestamp 1662439860
transform 1 0 41492 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1011_
timestamp 1662439860
transform 1 0 43608 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1012_
timestamp 1662439860
transform -1 0 37076 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1013_
timestamp 1662439860
transform -1 0 38272 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1014_
timestamp 1662439860
transform -1 0 38640 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1015_
timestamp 1662439860
transform -1 0 35512 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1016_
timestamp 1662439860
transform -1 0 31556 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1017_
timestamp 1662439860
transform -1 0 34224 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1018_
timestamp 1662439860
transform -1 0 37720 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1019_
timestamp 1662439860
transform -1 0 47840 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1020_
timestamp 1662439860
transform 1 0 45632 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1021_
timestamp 1662439860
transform 1 0 43516 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1022_
timestamp 1662439860
transform 1 0 32752 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1023_
timestamp 1662439860
transform -1 0 34316 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _1024_
timestamp 1662439860
transform -1 0 35420 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1662439860
transform 1 0 34408 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1026_
timestamp 1662439860
transform -1 0 34040 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1027_
timestamp 1662439860
transform -1 0 33672 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1662439860
transform 1 0 29716 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1029_
timestamp 1662439860
transform 1 0 72128 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1662439860
transform -1 0 74428 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1031_
timestamp 1662439860
transform 1 0 72128 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1032_
timestamp 1662439860
transform 1 0 75072 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1662439860
transform -1 0 76544 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1034_
timestamp 1662439860
transform 1 0 34868 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1035_
timestamp 1662439860
transform -1 0 56396 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1036_
timestamp 1662439860
transform 1 0 48576 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1037_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 49312 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _1038_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 53912 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1039_
timestamp 1662439860
transform 1 0 52992 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1040_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 48576 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1041_
timestamp 1662439860
transform -1 0 9752 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1042_
timestamp 1662439860
transform 1 0 49404 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1043_
timestamp 1662439860
transform -1 0 50876 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_2  _1044_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 48208 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1045_
timestamp 1662439860
transform -1 0 7176 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1046__29
timestamp 1662439860
transform 1 0 18492 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047__30
timestamp 1662439860
transform -1 0 18032 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048__31
timestamp 1662439860
transform -1 0 18308 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049__32
timestamp 1662439860
transform -1 0 13984 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1050__33
timestamp 1662439860
transform 1 0 21252 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051__34
timestamp 1662439860
transform 1 0 25208 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052__35
timestamp 1662439860
transform -1 0 22632 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1053_
timestamp 1662439860
transform 1 0 42504 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1054__36
timestamp 1662439860
transform 1 0 46184 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1055__37
timestamp 1662439860
transform -1 0 45540 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1056__38
timestamp 1662439860
transform 1 0 49588 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1057__39
timestamp 1662439860
transform -1 0 45816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1058__40
timestamp 1662439860
transform -1 0 49312 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1059__41
timestamp 1662439860
transform 1 0 42596 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1060__42
timestamp 1662439860
transform -1 0 38548 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1061__43
timestamp 1662439860
transform -1 0 40296 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1062_
timestamp 1662439860
transform 1 0 2852 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1063__44
timestamp 1662439860
transform -1 0 40388 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1064_
timestamp 1662439860
transform 1 0 9384 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1065__45
timestamp 1662439860
transform -1 0 41768 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _1066_
timestamp 1662439860
transform 1 0 2852 0 -1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_6  _1067_
timestamp 1662439860
transform 1 0 87400 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1662439860
transform -1 0 53084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1069_
timestamp 1662439860
transform 1 0 80500 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1070_
timestamp 1662439860
transform 1 0 89700 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1071_
timestamp 1662439860
transform -1 0 89240 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1662439860
transform -1 0 73048 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1073_
timestamp 1662439860
transform -1 0 54648 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1074_
timestamp 1662439860
transform 1 0 62560 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1075_
timestamp 1662439860
transform -1 0 84824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1662439860
transform -1 0 71852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1077_
timestamp 1662439860
transform -1 0 89240 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1078_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 21988 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_4  _1079_
timestamp 1662439860
transform -1 0 91080 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1662439860
transform -1 0 62744 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1662439860
transform -1 0 70472 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1082_
timestamp 1662439860
transform 1 0 63480 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1083_
timestamp 1662439860
transform 1 0 90436 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1084_
timestamp 1662439860
transform 1 0 86664 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1085_
timestamp 1662439860
transform -1 0 94024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1086_
timestamp 1662439860
transform 1 0 83260 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1087_
timestamp 1662439860
transform 1 0 54740 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1088_
timestamp 1662439860
transform -1 0 62008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1089_
timestamp 1662439860
transform 1 0 37904 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1662439860
transform -1 0 80040 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1091_
timestamp 1662439860
transform 1 0 42596 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1092_
timestamp 1662439860
transform -1 0 67896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1093_
timestamp 1662439860
transform 1 0 48208 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1662439860
transform 1 0 75900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1095_
timestamp 1662439860
transform 1 0 85928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1096_
timestamp 1662439860
transform 1 0 43516 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 1662439860
transform 1 0 89792 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1098_
timestamp 1662439860
transform 1 0 55108 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  _1099_
timestamp 1662439860
transform 1 0 90344 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1100_
timestamp 1662439860
transform 1 0 65504 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1101__46
timestamp 1662439860
transform 1 0 73600 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1102__47
timestamp 1662439860
transform 1 0 67252 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1103_
timestamp 1662439860
transform 1 0 3956 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1104_
timestamp 1662439860
transform 1 0 4140 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1105_
timestamp 1662439860
transform -1 0 14904 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1106__48
timestamp 1662439860
transform -1 0 64400 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1107_
timestamp 1662439860
transform -1 0 81880 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1108__49
timestamp 1662439860
transform -1 0 66056 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1109_
timestamp 1662439860
transform -1 0 88780 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1110__50
timestamp 1662439860
transform -1 0 64768 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1111_
timestamp 1662439860
transform -1 0 80868 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1112_
timestamp 1662439860
transform -1 0 84456 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1113__51
timestamp 1662439860
transform 1 0 73508 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1114_
timestamp 1662439860
transform 1 0 51612 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1115__52
timestamp 1662439860
transform -1 0 66056 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1116_
timestamp 1662439860
transform 1 0 39468 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1117__53
timestamp 1662439860
transform -1 0 63664 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1118_
timestamp 1662439860
transform 1 0 50140 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1119__54
timestamp 1662439860
transform -1 0 72220 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1120__55
timestamp 1662439860
transform 1 0 73508 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1121_
timestamp 1662439860
transform 1 0 43424 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_1  _1122_
timestamp 1662439860
transform 1 0 58052 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1123__56
timestamp 1662439860
transform 1 0 61548 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1124_
timestamp 1662439860
transform 1 0 55752 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1125__57
timestamp 1662439860
transform 1 0 56396 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1126_
timestamp 1662439860
transform 1 0 11224 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1127__58
timestamp 1662439860
transform 1 0 59892 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1128_
timestamp 1662439860
transform -1 0 31832 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1129__59
timestamp 1662439860
transform -1 0 60168 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1130_
timestamp 1662439860
transform 1 0 13708 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1131__60
timestamp 1662439860
transform -1 0 53912 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1132_
timestamp 1662439860
transform 1 0 11684 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1133_
timestamp 1662439860
transform 1 0 7544 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1134__61
timestamp 1662439860
transform -1 0 53176 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1135_
timestamp 1662439860
transform -1 0 31464 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1136__62
timestamp 1662439860
transform -1 0 54096 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1137_
timestamp 1662439860
transform -1 0 38640 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1138__63
timestamp 1662439860
transform -1 0 56212 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1139_
timestamp 1662439860
transform 1 0 26036 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1140__64
timestamp 1662439860
transform 1 0 59892 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1141__65
timestamp 1662439860
transform -1 0 53820 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1142_
timestamp 1662439860
transform -1 0 30452 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1143__3
timestamp 1662439860
transform 1 0 30360 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1144_
timestamp 1662439860
transform 1 0 14720 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1145__4
timestamp 1662439860
transform -1 0 36708 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1146_
timestamp 1662439860
transform 1 0 3312 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1147__5
timestamp 1662439860
transform -1 0 59708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1148_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 1932 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1149_
timestamp 1662439860
transform -1 0 18584 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1150_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 17664 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1151_
timestamp 1662439860
transform 1 0 4600 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1152_
timestamp 1662439860
transform 1 0 2760 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1153_
timestamp 1662439860
transform 1 0 19412 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1154_
timestamp 1662439860
transform -1 0 13616 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1155_
timestamp 1662439860
transform -1 0 13800 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1156_
timestamp 1662439860
transform 1 0 7452 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1157_
timestamp 1662439860
transform 1 0 22172 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1158_
timestamp 1662439860
transform 1 0 21344 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1159_
timestamp 1662439860
transform -1 0 24840 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1160_
timestamp 1662439860
transform 1 0 14536 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1161_
timestamp 1662439860
transform 1 0 22264 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1162_
timestamp 1662439860
transform 1 0 21988 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1163_
timestamp 1662439860
transform 1 0 46644 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1164_
timestamp 1662439860
transform 1 0 21988 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1165_
timestamp 1662439860
transform 1 0 45172 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1166_
timestamp 1662439860
transform 1 0 2300 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1167_
timestamp 1662439860
transform 1 0 47380 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1168_
timestamp 1662439860
transform 1 0 7912 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1169_
timestamp 1662439860
transform 1 0 45448 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1170_
timestamp 1662439860
transform 1 0 12696 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1171_
timestamp 1662439860
transform 1 0 47748 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1172_
timestamp 1662439860
transform -1 0 12328 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1173_
timestamp 1662439860
transform -1 0 42136 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1174_
timestamp 1662439860
transform -1 0 39560 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1175_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 16192 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1176_
timestamp 1662439860
transform 1 0 38364 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1177_
timestamp 1662439860
transform 1 0 14444 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1178_
timestamp 1662439860
transform 1 0 38916 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1179_
timestamp 1662439860
transform 1 0 14260 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1180_
timestamp 1662439860
transform 1 0 40296 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1181_
timestamp 1662439860
transform 1 0 69736 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1182_
timestamp 1662439860
transform -1 0 67896 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1183_
timestamp 1662439860
transform 1 0 59800 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1184_
timestamp 1662439860
transform -1 0 73048 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1185_
timestamp 1662439860
transform -1 0 68264 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1186_
timestamp 1662439860
transform 1 0 63480 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1187_
timestamp 1662439860
transform 1 0 61824 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1188_
timestamp 1662439860
transform 1 0 54464 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1189_
timestamp 1662439860
transform 1 0 41216 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1190_
timestamp 1662439860
transform 1 0 43976 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1191_
timestamp 1662439860
transform -1 0 56212 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1192_
timestamp 1662439860
transform 1 0 36340 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1193_
timestamp 1662439860
transform 1 0 49128 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1194_
timestamp 1662439860
transform -1 0 61180 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1195_
timestamp 1662439860
transform -1 0 62744 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1196_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 75716 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1197_
timestamp 1662439860
transform -1 0 67712 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1198_
timestamp 1662439860
transform 1 0 54556 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1199_
timestamp 1662439860
transform 1 0 50324 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1200_
timestamp 1662439860
transform 1 0 81236 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1201_
timestamp 1662439860
transform 1 0 85100 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1202_
timestamp 1662439860
transform 1 0 88964 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1203_
timestamp 1662439860
transform 1 0 87400 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1204_
timestamp 1662439860
transform -1 0 88044 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1205_
timestamp 1662439860
transform 1 0 81512 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1206_
timestamp 1662439860
transform 1 0 73140 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1207_
timestamp 1662439860
transform 1 0 68816 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1208_
timestamp 1662439860
transform 1 0 50416 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1209_
timestamp 1662439860
transform -1 0 52440 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1210_
timestamp 1662439860
transform 1 0 68356 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1211_
timestamp 1662439860
transform 1 0 63204 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1212_
timestamp 1662439860
transform -1 0 85928 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1213_
timestamp 1662439860
transform 1 0 82892 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1214_
timestamp 1662439860
transform -1 0 70472 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1215_
timestamp 1662439860
transform 1 0 70932 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1216_
timestamp 1662439860
transform 1 0 86664 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1217_
timestamp 1662439860
transform 1 0 79304 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1218_
timestamp 1662439860
transform -1 0 90896 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1219_
timestamp 1662439860
transform 1 0 82156 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1220_
timestamp 1662439860
transform -1 0 89056 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1221_
timestamp 1662439860
transform 1 0 71300 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1222_
timestamp 1662439860
transform -1 0 70380 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1223_
timestamp 1662439860
transform 1 0 65780 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1224_
timestamp 1662439860
transform 1 0 79948 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1225_
timestamp 1662439860
transform 1 0 68080 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1226_
timestamp 1662439860
transform 1 0 69736 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1227_
timestamp 1662439860
transform 1 0 71208 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1228_
timestamp 1662439860
transform -1 0 79672 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1229_
timestamp 1662439860
transform 1 0 78660 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1230_
timestamp 1662439860
transform -1 0 93564 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1231_
timestamp 1662439860
transform 1 0 89056 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1232_
timestamp 1662439860
transform 1 0 91724 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1233_
timestamp 1662439860
transform 1 0 80684 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1234_
timestamp 1662439860
transform 1 0 58052 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1235_
timestamp 1662439860
transform 1 0 55200 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1236_
timestamp 1662439860
transform 1 0 67344 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1237_
timestamp 1662439860
transform 1 0 73784 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1238_
timestamp 1662439860
transform 1 0 89792 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1239_
timestamp 1662439860
transform 1 0 91540 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1240_
timestamp 1662439860
transform 1 0 90620 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1241_
timestamp 1662439860
transform 1 0 91540 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1242_
timestamp 1662439860
transform 1 0 56304 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1243_
timestamp 1662439860
transform 1 0 60628 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1244_
timestamp 1662439860
transform 1 0 76084 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1245_
timestamp 1662439860
transform 1 0 77556 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1246_
timestamp 1662439860
transform 1 0 58052 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1247_
timestamp 1662439860
transform 1 0 64492 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1248_
timestamp 1662439860
transform -1 0 84272 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1249_
timestamp 1662439860
transform 1 0 75164 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1250_
timestamp 1662439860
transform -1 0 87308 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1251_
timestamp 1662439860
transform 1 0 86388 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1252_
timestamp 1662439860
transform 1 0 89884 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1253_
timestamp 1662439860
transform -1 0 93656 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1254_
timestamp 1662439860
transform -1 0 64124 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1255_
timestamp 1662439860
transform -1 0 53728 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1256_
timestamp 1662439860
transform 1 0 55660 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1257_
timestamp 1662439860
transform -1 0 65044 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1258_
timestamp 1662439860
transform -1 0 85928 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1259_
timestamp 1662439860
transform -1 0 67620 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1260_
timestamp 1662439860
transform -1 0 62468 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1261_
timestamp 1662439860
transform 1 0 62836 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1262_
timestamp 1662439860
transform 1 0 91540 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1263_
timestamp 1662439860
transform 1 0 14168 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1264_
timestamp 1662439860
transform 1 0 73508 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1265_
timestamp 1662439860
transform 1 0 19964 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1266_
timestamp 1662439860
transform 1 0 67896 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1267_
timestamp 1662439860
transform -1 0 14904 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1268_
timestamp 1662439860
transform 1 0 6808 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1269_
timestamp 1662439860
transform 1 0 6716 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1270_
timestamp 1662439860
transform 1 0 3956 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1271_
timestamp 1662439860
transform 1 0 5980 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1272_
timestamp 1662439860
transform 1 0 4140 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1273_
timestamp 1662439860
transform -1 0 13800 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1274_
timestamp 1662439860
transform 1 0 4968 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1275_
timestamp 1662439860
transform 1 0 29900 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1276_
timestamp 1662439860
transform 1 0 34868 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1277_
timestamp 1662439860
transform 1 0 33580 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1278_
timestamp 1662439860
transform 1 0 32844 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1279_
timestamp 1662439860
transform 1 0 25760 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1280_
timestamp 1662439860
transform 1 0 25300 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1281_
timestamp 1662439860
transform 1 0 34868 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1282_
timestamp 1662439860
transform 1 0 29900 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1283_
timestamp 1662439860
transform 1 0 32476 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1284_
timestamp 1662439860
transform 1 0 34868 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1285_
timestamp 1662439860
transform 1 0 26680 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1286_
timestamp 1662439860
transform 1 0 24840 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1287_
timestamp 1662439860
transform -1 0 26496 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1288_
timestamp 1662439860
transform -1 0 31832 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1289_
timestamp 1662439860
transform 1 0 30176 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1290_
timestamp 1662439860
transform 1 0 32844 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1291_
timestamp 1662439860
transform 1 0 61824 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1292_
timestamp 1662439860
transform -1 0 79212 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1293_
timestamp 1662439860
transform 1 0 63296 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1294_
timestamp 1662439860
transform -1 0 72680 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1295_
timestamp 1662439860
transform 1 0 62652 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1296_
timestamp 1662439860
transform -1 0 79028 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1297_
timestamp 1662439860
transform -1 0 80500 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1298_
timestamp 1662439860
transform 1 0 71576 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1299_
timestamp 1662439860
transform -1 0 66516 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1300_
timestamp 1662439860
transform 1 0 63204 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1301_
timestamp 1662439860
transform 1 0 77004 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1302_
timestamp 1662439860
transform 1 0 62192 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1303_
timestamp 1662439860
transform 1 0 78660 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1304_
timestamp 1662439860
transform 1 0 70472 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1305_
timestamp 1662439860
transform -1 0 73140 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1306_
timestamp 1662439860
transform 1 0 68172 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1307_
timestamp 1662439860
transform -1 0 62744 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1308_
timestamp 1662439860
transform 1 0 64860 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1309_
timestamp 1662439860
transform 1 0 55200 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1310_
timestamp 1662439860
transform 1 0 18308 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1311_
timestamp 1662439860
transform 1 0 31556 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1312_
timestamp 1662439860
transform 1 0 32476 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1313_
timestamp 1662439860
transform 1 0 24564 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1314_
timestamp 1662439860
transform 1 0 32936 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1315_
timestamp 1662439860
transform 1 0 25392 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1316_
timestamp 1662439860
transform 1 0 27692 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1317_
timestamp 1662439860
transform 1 0 25944 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1318_
timestamp 1662439860
transform 1 0 27140 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1319_
timestamp 1662439860
transform 1 0 24564 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1320_
timestamp 1662439860
transform -1 0 26588 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1321_
timestamp 1662439860
transform -1 0 26496 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1322_
timestamp 1662439860
transform -1 0 27232 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1323_
timestamp 1662439860
transform -1 0 30268 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1324_
timestamp 1662439860
transform -1 0 30176 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1325_
timestamp 1662439860
transform -1 0 34408 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1326_
timestamp 1662439860
transform -1 0 32568 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1327_
timestamp 1662439860
transform -1 0 61824 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1328_
timestamp 1662439860
transform -1 0 23828 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1329_
timestamp 1662439860
transform -1 0 61180 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1330_
timestamp 1662439860
transform 1 0 19412 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1331_
timestamp 1662439860
transform -1 0 54832 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1332_
timestamp 1662439860
transform 1 0 19044 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1333_
timestamp 1662439860
transform 1 0 19412 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1334_
timestamp 1662439860
transform 1 0 51152 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1335_
timestamp 1662439860
transform -1 0 30176 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1336_
timestamp 1662439860
transform 1 0 51520 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1337_
timestamp 1662439860
transform -1 0 26680 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1338_
timestamp 1662439860
transform -1 0 57132 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1339_
timestamp 1662439860
transform 1 0 27140 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1340_
timestamp 1662439860
transform -1 0 61364 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1341_
timestamp 1662439860
transform -1 0 54648 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1342_
timestamp 1662439860
transform -1 0 29992 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1343_
timestamp 1662439860
transform 1 0 29716 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1344_
timestamp 1662439860
transform 1 0 18768 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1345_
timestamp 1662439860
transform -1 0 37352 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1346_
timestamp 1662439860
transform 1 0 32568 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1347_
timestamp 1662439860
transform -1 0 39468 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1348_
timestamp 1662439860
transform -1 0 39376 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1349_
timestamp 1662439860
transform 1 0 37444 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1350_
timestamp 1662439860
transform 1 0 40388 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1351_
timestamp 1662439860
transform -1 0 36984 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1352_
timestamp 1662439860
transform 1 0 49128 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1353_
timestamp 1662439860
transform 1 0 57040 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1354_
timestamp 1662439860
transform 1 0 61088 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1355_
timestamp 1662439860
transform 1 0 59064 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__buf_2  _1356_
timestamp 1662439860
transform 1 0 28244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1357_
timestamp 1662439860
transform 1 0 76084 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1358_
timestamp 1662439860
transform 1 0 28704 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1359_
timestamp 1662439860
transform -1 0 75440 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1360_
timestamp 1662439860
transform 1 0 20056 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1361_
timestamp 1662439860
transform -1 0 67436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1362_
timestamp 1662439860
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1363_
timestamp 1662439860
transform -1 0 68172 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1364_
timestamp 1662439860
transform 1 0 5244 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1365_
timestamp 1662439860
transform 1 0 52164 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1366_
timestamp 1662439860
transform -1 0 11960 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1367_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 90804 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1368_
timestamp 1662439860
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1369_
timestamp 1662439860
transform 1 0 79672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1370_
timestamp 1662439860
transform -1 0 92828 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1371_
timestamp 1662439860
transform -1 0 92828 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1372_
timestamp 1662439860
transform -1 0 93472 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1373_
timestamp 1662439860
transform -1 0 92184 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1374_
timestamp 1662439860
transform -1 0 3312 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1375_
timestamp 1662439860
transform 1 0 53360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0301_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 43424 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0304_
timestamp 1662439860
transform 1 0 68356 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0305_
timestamp 1662439860
transform -1 0 58880 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0306_
timestamp 1662439860
transform 1 0 42872 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0307_
timestamp 1662439860
transform 1 0 24288 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0308_
timestamp 1662439860
transform 1 0 72680 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0311_
timestamp 1662439860
transform -1 0 21160 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_master
timestamp 1662439860
transform 1 0 11960 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w0.cclk_I
timestamp 1662439860
transform -1 0 31648 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0301_
timestamp 1662439860
transform -1 0 39560 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0304_
timestamp 1662439860
transform -1 0 67252 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0305_
timestamp 1662439860
transform -1 0 54740 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0306_
timestamp 1662439860
transform -1 0 42504 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0307_
timestamp 1662439860
transform -1 0 23828 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0308_
timestamp 1662439860
transform -1 0 69460 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0311_
timestamp 1662439860
transform -1 0 17480 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0301_
timestamp 1662439860
transform 1 0 44160 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0304_
timestamp 1662439860
transform 1 0 70564 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0305_
timestamp 1662439860
transform 1 0 57224 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0306_
timestamp 1662439860
transform 1 0 46828 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0307_
timestamp 1662439860
transform 1 0 26036 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0308_
timestamp 1662439860
transform 1 0 73784 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0311_
timestamp 1662439860
transform 1 0 19688 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk_master
timestamp 1662439860
transform -1 0 9660 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_w0.cclk_I
timestamp 1662439860
transform -1 0 27876 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk_master
timestamp 1662439860
transform -1 0 9660 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_w0.cclk_I
timestamp 1662439860
transform -1 0 28980 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk_master
timestamp 1662439860
transform 1 0 12972 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_w0.cclk_I
timestamp 1662439860
transform 1 0 30268 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk_master
timestamp 1662439860
transform 1 0 14260 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_w0.cclk_I
timestamp 1662439860
transform 1 0 32016 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 1662439860
transform 1 0 63756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout32
timestamp 1662439860
transform -1 0 76452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout33
timestamp 1662439860
transform -1 0 93380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout34
timestamp 1662439860
transform 1 0 92920 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp 1662439860
transform 1 0 75992 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout36
timestamp 1662439860
transform -1 0 79212 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout37
timestamp 1662439860
transform 1 0 77464 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout38
timestamp 1662439860
transform 1 0 86756 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout39
timestamp 1662439860
transform 1 0 86388 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout40
timestamp 1662439860
transform 1 0 84824 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp 1662439860
transform 1 0 10028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout42
timestamp 1662439860
transform -1 0 2208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout43
timestamp 1662439860
transform -1 0 6256 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout44
timestamp 1662439860
transform 1 0 16836 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 1662439860
transform -1 0 17112 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout46
timestamp 1662439860
transform -1 0 24104 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout47
timestamp 1662439860
transform -1 0 25024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout48
timestamp 1662439860
transform -1 0 35420 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 1662439860
transform 1 0 27876 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout50
timestamp 1662439860
transform 1 0 37536 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout51
timestamp 1662439860
transform 1 0 4876 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout52
timestamp 1662439860
transform 1 0 62100 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout53
timestamp 1662439860
transform -1 0 61364 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout54
timestamp 1662439860
transform 1 0 50324 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout55
timestamp 1662439860
transform -1 0 71668 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout56
timestamp 1662439860
transform -1 0 88412 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout57
timestamp 1662439860
transform 1 0 87952 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout58
timestamp 1662439860
transform 1 0 83812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout59
timestamp 1662439860
transform -1 0 75256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1662439860
transform 1 0 44068 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1662439860
transform 1 0 91540 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1662439860
transform 1 0 44068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 91540 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1662439860
transform 1 0 36156 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1662439860
transform 1 0 83628 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1662439860
transform -1 0 36432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1662439860
transform -1 0 84180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input9
timestamp 1662439860
transform 1 0 1564 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1662439860
transform -1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output11
timestamp 1662439860
transform 1 0 28244 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1662439860
transform 1 0 76084 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output13
timestamp 1662439860
transform 1 0 28244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1662439860
transform 1 0 76084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output15
timestamp 1662439860
transform 1 0 20332 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1662439860
transform 1 0 68356 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output17
timestamp 1662439860
transform 1 0 20792 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1662439860
transform 1 0 68356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1662439860
transform -1 0 4876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1662439860
transform -1 0 52348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1662439860
transform 1 0 12420 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1662439860
transform -1 0 60168 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1662439860
transform -1 0 12788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1662439860
transform -1 0 60996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1662439860
transform 1 0 94024 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1662439860
transform 1 0 94024 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1662439860
transform 1 0 94024 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1662439860
transform 1 0 94024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1662439860
transform 1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1662439860
transform -1 0 52348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 6624 0 -1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 33672 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn
timestamp 1662439860
transform -1 0 8372 0 1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
timestamp 1662439860
transform 1 0 35328 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn
timestamp 1662439860
transform 1 0 8280 0 -1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
timestamp 1662439860
transform 1 0 44712 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn
timestamp 1662439860
transform -1 0 7912 0 -1 8704
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
timestamp 1662439860
transform 1 0 46000 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn
timestamp 1662439860
transform 1 0 4784 0 -1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
timestamp 1662439860
transform -1 0 46828 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn
timestamp 1662439860
transform 1 0 3956 0 1 10880
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
timestamp 1662439860
transform -1 0 35696 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn
timestamp 1662439860
transform 1 0 2208 0 1 10880
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
timestamp 1662439860
transform 1 0 32476 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn
timestamp 1662439860
transform 1 0 2576 0 -1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
timestamp 1662439860
transform 1 0 27416 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn
timestamp 1662439860
transform 1 0 2208 0 1 8704
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
timestamp 1662439860
transform -1 0 26680 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn
timestamp 1662439860
transform 1 0 2208 0 1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
timestamp 1662439860
transform 1 0 31832 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn
timestamp 1662439860
transform 1 0 8188 0 -1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
timestamp 1662439860
transform -1 0 41584 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn
timestamp 1662439860
transform 1 0 6532 0 -1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
timestamp 1662439860
transform -1 0 52808 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn
timestamp 1662439860
transform 1 0 9844 0 -1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
timestamp 1662439860
transform -1 0 61364 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn
timestamp 1662439860
transform 1 0 7176 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
timestamp 1662439860
transform -1 0 56304 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn
timestamp 1662439860
transform 1 0 9108 0 1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
timestamp 1662439860
transform -1 0 62560 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn
timestamp 1662439860
transform -1 0 10396 0 1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
timestamp 1662439860
transform 1 0 56764 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn
timestamp 1662439860
transform 1 0 9568 0 -1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
timestamp 1662439860
transform -1 0 57868 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn
timestamp 1662439860
transform 1 0 10028 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
timestamp 1662439860
transform 1 0 47380 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn
timestamp 1662439860
transform -1 0 15548 0 1 3264
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
timestamp 1662439860
transform 1 0 49772 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn
timestamp 1662439860
transform -1 0 12972 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
timestamp 1662439860
transform -1 0 43884 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_2  w0.ro_block_I.ro_pol.tribuf.t_buf dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 77096 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  w0.ro_block_I.ro_pol_eve.tribuf.t_buf
timestamp 1662439860
transform 1 0 83812 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  w0.ro_block_Q.ro_pol.tribuf.t_buf dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 27140 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  w0.ro_block_Q.ro_pol_eve.tribuf.t_buf
timestamp 1662439860
transform 1 0 31188 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn
timestamp 1662439860
transform 1 0 88688 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
timestamp 1662439860
transform -1 0 93656 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn
timestamp 1662439860
transform 1 0 89424 0 1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
timestamp 1662439860
transform 1 0 88964 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn
timestamp 1662439860
transform -1 0 90252 0 -1 8704
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
timestamp 1662439860
transform 1 0 83628 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn
timestamp 1662439860
transform 1 0 87216 0 -1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
timestamp 1662439860
transform 1 0 78660 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn
timestamp 1662439860
transform 1 0 91264 0 -1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
timestamp 1662439860
transform 1 0 80500 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn
timestamp 1662439860
transform 1 0 91540 0 1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
timestamp 1662439860
transform 1 0 68816 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn
timestamp 1662439860
transform -1 0 89700 0 1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
timestamp 1662439860
transform -1 0 78108 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn
timestamp 1662439860
transform 1 0 86388 0 -1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
timestamp 1662439860
transform -1 0 93472 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn
timestamp 1662439860
transform 1 0 84732 0 -1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
timestamp 1662439860
transform -1 0 74980 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn
timestamp 1662439860
transform 1 0 92092 0 -1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
timestamp 1662439860
transform 1 0 71760 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn
timestamp 1662439860
transform 1 0 86756 0 -1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
timestamp 1662439860
transform 1 0 83996 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn
timestamp 1662439860
transform 1 0 86756 0 1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
timestamp 1662439860
transform 1 0 68264 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn
timestamp 1662439860
transform -1 0 88044 0 1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
timestamp 1662439860
transform -1 0 82708 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn
timestamp 1662439860
transform -1 0 88044 0 -1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
timestamp 1662439860
transform 1 0 65964 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn
timestamp 1662439860
transform -1 0 86388 0 -1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
timestamp 1662439860
transform -1 0 54004 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn
timestamp 1662439860
transform 1 0 92092 0 -1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
timestamp 1662439860
transform -1 0 65228 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn
timestamp 1662439860
transform 1 0 81236 0 1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
timestamp 1662439860
transform 1 0 87952 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn
timestamp 1662439860
transform 1 0 81696 0 1 3264
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
timestamp 1662439860
transform -1 0 73048 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn
timestamp 1662439860
transform 1 0 83352 0 1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
timestamp 1662439860
transform 1 0 46000 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn
timestamp 1662439860
transform -1 0 80776 0 1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
timestamp 1662439860
transform 1 0 49772 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_2  wrapper_cell_loop\[0\].w1.ro_block_I.ro_pol.tribuf.t_buf
timestamp 1662439860
transform -1 0 65136 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  wrapper_cell_loop\[0\].w1.ro_block_I.ro_pol_eve.tribuf.t_buf
timestamp 1662439860
transform 1 0 73508 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  wrapper_cell_loop\[0\].w1.ro_block_Q.ro_pol.tribuf.t_buf
timestamp 1662439860
transform -1 0 54096 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  wrapper_cell_loop\[0\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf
timestamp 1662439860
transform -1 0 55752 0 -1 4352
box -38 -48 1234 592
<< labels >>
flabel metal2 s 28170 19200 28226 20000 0 FreeSans 224 90 0 0 cclk_I[0]
port 0 nsew signal tristate
flabel metal2 s 75642 19200 75698 20000 0 FreeSans 224 90 0 0 cclk_I[1]
port 1 nsew signal tristate
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 cclk_Q[0]
port 2 nsew signal tristate
flabel metal2 s 75642 0 75698 800 0 FreeSans 224 90 0 0 cclk_Q[1]
port 3 nsew signal tristate
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 clk_master
port 4 nsew signal input
flabel metal2 s 20258 19200 20314 20000 0 FreeSans 224 90 0 0 clkdiv2_I[0]
port 5 nsew signal tristate
flabel metal2 s 67730 19200 67786 20000 0 FreeSans 224 90 0 0 clkdiv2_I[1]
port 6 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 clkdiv2_Q[0]
port 7 nsew signal tristate
flabel metal2 s 67730 0 67786 800 0 FreeSans 224 90 0 0 clkdiv2_Q[1]
port 8 nsew signal tristate
flabel metal2 s 43994 19200 44050 20000 0 FreeSans 224 90 0 0 comp_high_I[0]
port 9 nsew signal input
flabel metal2 s 91466 19200 91522 20000 0 FreeSans 224 90 0 0 comp_high_I[1]
port 10 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 comp_high_Q[0]
port 11 nsew signal input
flabel metal2 s 91466 0 91522 800 0 FreeSans 224 90 0 0 comp_high_Q[1]
port 12 nsew signal input
flabel metal2 s 4434 19200 4490 20000 0 FreeSans 224 90 0 0 cos_out[0]
port 13 nsew signal tristate
flabel metal2 s 51906 19200 51962 20000 0 FreeSans 224 90 0 0 cos_out[1]
port 14 nsew signal tristate
flabel metal2 s 12346 19200 12402 20000 0 FreeSans 224 90 0 0 fb1_I[0]
port 15 nsew signal tristate
flabel metal2 s 59818 19200 59874 20000 0 FreeSans 224 90 0 0 fb1_I[1]
port 16 nsew signal tristate
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 fb1_Q[0]
port 17 nsew signal tristate
flabel metal2 s 59818 0 59874 800 0 FreeSans 224 90 0 0 fb1_Q[1]
port 18 nsew signal tristate
flabel metal2 s 36082 19200 36138 20000 0 FreeSans 224 90 0 0 phi1b_dig_I[0]
port 19 nsew signal input
flabel metal2 s 83554 19200 83610 20000 0 FreeSans 224 90 0 0 phi1b_dig_I[1]
port 20 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 phi1b_dig_Q[0]
port 21 nsew signal input
flabel metal2 s 83554 0 83610 800 0 FreeSans 224 90 0 0 phi1b_dig_Q[1]
port 22 nsew signal input
flabel metal3 s 95200 17280 96000 17400 0 FreeSans 480 0 0 0 read_out_I[0]
port 23 nsew signal tristate
flabel metal3 s 95200 12384 96000 12504 0 FreeSans 480 0 0 0 read_out_I[1]
port 24 nsew signal tristate
flabel metal3 s 95200 7488 96000 7608 0 FreeSans 480 0 0 0 read_out_Q[0]
port 25 nsew signal tristate
flabel metal3 s 95200 2592 96000 2712 0 FreeSans 480 0 0 0 read_out_Q[1]
port 26 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 rstb
port 27 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 sin_out[0]
port 28 nsew signal tristate
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 sin_out[1]
port 29 nsew signal tristate
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 ud_en
port 30 nsew signal input
flabel metal4 s 12662 2128 12982 17456 0 FreeSans 1920 90 0 0 vccd1
port 31 nsew power bidirectional
flabel metal4 s 36099 2128 36419 17456 0 FreeSans 1920 90 0 0 vccd1
port 31 nsew power bidirectional
flabel metal4 s 59536 2128 59856 17456 0 FreeSans 1920 90 0 0 vccd1
port 31 nsew power bidirectional
flabel metal4 s 82973 2128 83293 17456 0 FreeSans 1920 90 0 0 vccd1
port 31 nsew power bidirectional
flabel metal4 s 24380 2128 24700 17456 0 FreeSans 1920 90 0 0 vssd1
port 32 nsew ground bidirectional
flabel metal4 s 47817 2128 48137 17456 0 FreeSans 1920 90 0 0 vssd1
port 32 nsew ground bidirectional
flabel metal4 s 71254 2128 71574 17456 0 FreeSans 1920 90 0 0 vssd1
port 32 nsew ground bidirectional
flabel metal4 s 94691 2128 95011 17456 0 FreeSans 1920 90 0 0 vssd1
port 32 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 96000 20000
<< end >>
