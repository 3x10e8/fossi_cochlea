* NGSPICE file created from digital_unison.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlrtn_1 abstract view
.subckt sky130_fd_sc_hd__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

.subckt digital_unison cclk_I[0] cclk_I[1] cclk_I[2] cclk_I[3] cclk_I[4] cclk_I[5]
+ cclk_I[6] cclk_I[7] cclk_Q[0] cclk_Q[1] cclk_Q[2] cclk_Q[3] cclk_Q[4] cclk_Q[5]
+ cclk_Q[6] cclk_Q[7] clk_master clkdiv2_I[0] clkdiv2_I[1] clkdiv2_I[2] clkdiv2_I[3]
+ clkdiv2_I[4] clkdiv2_I[5] clkdiv2_I[6] clkdiv2_I[7] clkdiv2_Q[0] clkdiv2_Q[1] clkdiv2_Q[2]
+ clkdiv2_Q[3] clkdiv2_Q[4] clkdiv2_Q[5] clkdiv2_Q[6] clkdiv2_Q[7] comp_high_I[0]
+ comp_high_I[1] comp_high_I[2] comp_high_I[3] comp_high_I[4] comp_high_I[5] comp_high_I[6]
+ comp_high_I[7] comp_high_Q[0] comp_high_Q[1] comp_high_Q[2] comp_high_Q[3] comp_high_Q[4]
+ comp_high_Q[5] comp_high_Q[6] comp_high_Q[7] cos_out[0] cos_out[1] cos_out[2] cos_out[3]
+ cos_out[4] cos_out[5] cos_out[6] cos_out[7] fb1_I[0] fb1_I[1] fb1_I[2] fb1_I[3]
+ fb1_I[4] fb1_I[5] fb1_I[6] fb1_I[7] fb1_Q[0] fb1_Q[1] fb1_Q[2] fb1_Q[3] fb1_Q[4]
+ fb1_Q[5] fb1_Q[6] fb1_Q[7] phi1b_dig_I[0] phi1b_dig_I[1] phi1b_dig_I[2] phi1b_dig_I[3]
+ phi1b_dig_I[4] phi1b_dig_I[5] phi1b_dig_I[6] phi1b_dig_I[7] phi1b_dig_Q[0] phi1b_dig_Q[1]
+ phi1b_dig_Q[2] phi1b_dig_Q[3] phi1b_dig_Q[4] phi1b_dig_Q[5] phi1b_dig_Q[6] phi1b_dig_Q[7]
+ read_out_I[0] read_out_I[1] read_out_Q[0] read_out_Q[1] rstb sin_out[0] sin_out[1]
+ sin_out[2] sin_out[3] sin_out[4] sin_out[5] sin_out[6] sin_out[7] ud_en vccd1 vssd1
XFILLER_7_2570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3140__A1 _4064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3155_ _3777_/A vssd1 vssd1 vccd1 vccd1 _3155_/X sky130_fd_sc_hd__buf_1
X_2106_ _4463_/D _4464_/Q vssd1 vssd1 vccd1 vccd1 _2107_/B sky130_fd_sc_hd__and2b_1
X_3086_ _4990_/Q _3086_/B vssd1 vssd1 vccd1 vccd1 _3086_/X sky130_fd_sc_hd__and2b_1
XFILLER_23_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_2409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2037_ _4426_/Q vssd1 vssd1 vccd1 vccd1 _2049_/A sky130_fd_sc_hd__inv_2
XANTENNA__2455__A _3658_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout162_A _5013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4728__CLK _5013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3988_ _4451_/Q vssd1 vssd1 vccd1 vccd1 _4452_/D sky130_fd_sc_hd__inv_2
XFILLER_17_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2939_ _4931_/D _4905_/Q _4903_/Q vssd1 vssd1 vccd1 vccd1 _2939_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__4878__CLK _1765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3286__A _3895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4490__RESET_B fanout202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2190__A _4555_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4609_ _2470_/A1 _4609_/D _3340_/Y vssd1 vssd1 vccd1 vccd1 _4609_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_RESET_B
+ fanout239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4578__RESET_B fanout228/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1996__A2 _4397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_2998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_2119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3924__A _3924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_2710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_3383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_3269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_3121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4960_ _4962_/CLK _4960_/D fanout212/X vssd1 vssd1 vccd1 vccd1 _4960_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_3154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_3165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3911_ _3907_/Y _3914_/B _3914_/C vssd1 vssd1 vccd1 vccd1 _3913_/B sky130_fd_sc_hd__mux2_4
X_4891_ _4901_/CLK _4891_/D fanout236/X vssd1 vssd1 vccd1 vccd1 _4891_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_2453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4930__RESET_B fanout236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3842_ _4360_/Q vssd1 vssd1 vccd1 vccd1 _3848_/A sky130_fd_sc_hd__buf_4
XFILLER_11_3906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_2620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_2041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2724_ _4808_/Q _4807_/Q _4806_/Q _2760_/A vssd1 vssd1 vccd1 vccd1 _2747_/B sky130_fd_sc_hd__or4_1
XFILLER_9_4012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2655_ _4763_/Q _2659_/B _2661_/A vssd1 vssd1 vccd1 vccd1 _2704_/C sky130_fd_sc_hd__o21ai_1
XFILLER_31_1985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_4078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_3103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2586_ _4713_/Q _2550_/D _2579_/B vssd1 vssd1 vccd1 vccd1 _2587_/B sky130_fd_sc_hd__a21bo_1
XFILLER_5_3208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4400__CLK _4402_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4325_ _5040_/A _4325_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _4325_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_29_2582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout105 _3135_/Y vssd1 vssd1 vccd1 vccd1 _4997_/CLK sky130_fd_sc_hd__clkbuf_4
Xfanout116 _4811_/CLK vssd1 vssd1 vccd1 vccd1 _4812_/CLK sky130_fd_sc_hd__buf_2
Xfanout127 fanout128/X vssd1 vssd1 vccd1 vccd1 _3643_/A sky130_fd_sc_hd__buf_2
XFILLER_5_2518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout138 _4655_/Q vssd1 vssd1 vccd1 vccd1 _5060_/A sky130_fd_sc_hd__buf_6
XFILLER_29_1881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout149 _2114_/Y vssd1 vssd1 vccd1 vccd1 _5033_/A sky130_fd_sc_hd__buf_4
X_4256_ _4256_/A vssd1 vssd1 vccd1 vccd1 _4841_/D sky130_fd_sc_hd__clkinv_2
XFILLER_25_1767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4187_ _4248_/D vssd1 vssd1 vccd1 vccd1 _4187_/Y sky130_fd_sc_hd__inv_8
XFILLER_20_3781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4550__CLK _2470_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3138_ _2972_/X _3137_/X _3941_/B vssd1 vssd1 vccd1 vccd1 _3138_/X sky130_fd_sc_hd__a21o_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_2297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2185__A _4494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3069_ _4985_/Q _3069_/B vssd1 vssd1 vccd1 vccd1 _3069_/Y sky130_fd_sc_hd__nor2_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_3107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2913__A _2916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_4117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3744__A _3748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3463__B _3923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_2153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_3753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_2855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_4142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_4006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4423__CLK _1952_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2440_ _4638_/Q _4637_/Q vssd1 vssd1 vccd1 vccd1 _2440_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_26_2700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_3445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2371_ _4606_/Q _4605_/Q vssd1 vssd1 vccd1 vccd1 _2371_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_26_3489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4188__C _4248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4573__CLK _3855_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4110_ _4638_/Q vssd1 vssd1 vccd1 vccd1 _4637_/D sky130_fd_sc_hd__inv_2
XFILLER_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5090_ _5090_/A vssd1 vssd1 vccd1 vccd1 _5090_/X sky130_fd_sc_hd__buf_4
XFILLER_20_3022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4041_ _4537_/Q vssd1 vssd1 vccd1 vccd1 _4536_/D sky130_fd_sc_hd__inv_2
XFILLER_20_2321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_2595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
+ _4997_/Q _3124_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_20_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4429__RESET_B fanout194/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4943_ _4943_/CLK _4943_/D _3528__52/Y vssd1 vssd1 vccd1 vccd1 _4943_/Q sky130_fd_sc_hd__dfrtp_1
X_4874_ _4187_/Y _4874_/D _3484_/Y vssd1 vssd1 vccd1 vccd1 _4874_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_1402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3825_ _4339_/Q vssd1 vssd1 vccd1 vccd1 _4338_/D sky130_fd_sc_hd__inv_2
XFILLER_31_3173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout125_A _4709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3756_ _3948_/A vssd1 vssd1 vccd1 vccd1 _3756_/Y sky130_fd_sc_hd__inv_2
X_2707_ _4778_/Q _4777_/Q vssd1 vssd1 vccd1 vccd1 _2707_/Y sky130_fd_sc_hd__xnor2_2
X_3687_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3687_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4916__CLK _4916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2638_ _4131_/C _2456_/Y _2978_/B _3875_/D vssd1 vssd1 vccd1 vccd1 _2638_/X sky130_fd_sc_hd__a211o_1
XFILLER_27_2519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2569_ _4708_/Q _2569_/B vssd1 vssd1 vccd1 vccd1 _2569_/X sky130_fd_sc_hd__and2b_1
X_4308_ _3845_/Y _4308_/D _3162__62/Y vssd1 vssd1 vccd1 vccd1 _4308_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_3865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4239_ _4827_/Q vssd1 vssd1 vccd1 vccd1 _4828_/D sky130_fd_sc_hd__inv_2
XFILLER_21_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2908__A _4895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3654__84 _3654__84/A vssd1 vssd1 vccd1 vccd1 _3654__84/Y sky130_fd_sc_hd__inv_2
XFILLER_19_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_2924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3739__A _3748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_2968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2362__B _2362_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_2670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_2018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_2917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_2939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_4098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout157/X fanout203/X vssd1 vssd1 vccd1 vccd1 _5082_/A sky130_fd_sc_hd__dlrtn_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3649__A _4195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1940_ _3882_/A _1952_/A1 _3910_/A _1939_/X vssd1 vssd1 vccd1 vccd1 _1941_/C sky130_fd_sc_hd__a31o_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1871_ _1871_/A _1871_/B vssd1 vssd1 vccd1 vccd1 _4311_/D sky130_fd_sc_hd__xnor2_1
XFILLER_32_3493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3610_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3610_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4939__CLK _4943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4590_ _4590_/CLK _4590_/D fanout229/X vssd1 vssd1 vccd1 vccd1 _4590_/Q sky130_fd_sc_hd__dfrtp_2
X_3541_ _4127_/A _4129_/A vssd1 vssd1 vccd1 vccd1 _3541_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_10_3791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3384__A _3947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2119__A2 _3941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2423_ _4622_/Q _2423_/B vssd1 vssd1 vccd1 vccd1 _4622_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_2602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_3358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2354_ _4648_/D _4590_/Q _4588_/Q vssd1 vssd1 vccd1 vccd1 _2354_/Y sky130_fd_sc_hd__nor3_1
XFILLER_26_2574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2728__A _2996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5073_ _5073_/A vssd1 vssd1 vccd1 vccd1 _5073_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4319__CLK _4324_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2285_ _3684_/Y _3710_/Y vssd1 vssd1 vccd1 vccd1 _2285_/Y sky130_fd_sc_hd__nor2_4
XFILLER_6_1967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4024_ _4502_/Q vssd1 vssd1 vccd1 vccd1 _4503_/D sky130_fd_sc_hd__inv_2
XFILLER_6_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4469__CLK _3257_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3559__A _3571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_3809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_2501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4926_ input31/X _4926_/D fanout228/X vssd1 vssd1 vccd1 vccd1 _4927_/D sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout242_A fanout257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_2512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3278__B _3442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2182__B _4497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4857_ _4865_/CLK _4857_/D fanout228/X vssd1 vssd1 vccd1 vccd1 _4857_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_1833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_2589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3808_ _4304_/Q vssd1 vssd1 vccd1 vccd1 _4305_/D sky130_fd_sc_hd__inv_2
XFILLER_11_2821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4788_ _3438_/Y _4788_/D _3647_/Y vssd1 vssd1 vccd1 vccd1 _4788_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_2291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3739_ _3748_/A vssd1 vssd1 vccd1 vccd1 _3739_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3294__A _4004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_2305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_2112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_2972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3188__B _3886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_2765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1717__A _4946_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_4127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3932__A _3932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_2944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[5\].w1.ro_block_I.ro_pol_eve.tribuf.t_buf _2967_/A _2815_/Y vssd1
+ vssd1 vccd1 vccd1 _5089_/A sky130_fd_sc_hd__ebufn_8
XFILLER_7_2966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4774__RESET_B fanout253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2548__A _4745_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4703__RESET_B _3669_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2809__B1 _3914_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2070_ _4432_/Q _2070_/B vssd1 vssd1 vccd1 vccd1 _4432_/D sky130_fd_sc_hd__xnor2_1
X_3476__46 _3523__49/A vssd1 vssd1 vccd1 vccd1 _3476__46/Y sky130_fd_sc_hd__inv_2
XANTENNA__4611__CLK _4623_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_2587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3379__A _3393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_2821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2972_ _4003_/C _2978_/C _2978_/D vssd1 vssd1 vccd1 vccd1 _2972_/X sky130_fd_sc_hd__a21bo_1
X_4711_ _4712_/CLK _4711_/D fanout245/X vssd1 vssd1 vccd1 vccd1 _4711_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1923_ _4343_/Q _4342_/Q vssd1 vssd1 vccd1 vccd1 _1923_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_34_2865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf _4274_/Q _1853_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_12_3875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4642_ _3358_/Y _4642_/D _3687_/Y vssd1 vssd1 vccd1 vccd1 _4642_/Q sky130_fd_sc_hd__dfrtp_2
X_1854_ _4309_/Q _4308_/Q vssd1 vssd1 vccd1 vccd1 _1854_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_15_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_4027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4573_ _3855_/Y _4573_/D _3320__29/Y vssd1 vssd1 vccd1 vccd1 _4573_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2730__B _4799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1785_ _4279_/Q _4278_/Q _4277_/Q _1799_/B vssd1 vssd1 vccd1 vccd1 _1790_/B sky130_fd_sc_hd__or4_1
XFILLER_11_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3191__73_A _3193__75/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4003__A _4131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout120/X fanout249/X vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__dlrtn_1
X_3455_ _4065_/A _3543_/B vssd1 vssd1 vccd1 vccd1 _3455_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_26_3050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_3083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2406_ _2377_/D _2405_/X _2344_/X vssd1 vssd1 vccd1 vccd1 _2407_/B sky130_fd_sc_hd__o21ai_1
X_3386_ _3935_/A _3440_/B vssd1 vssd1 vccd1 vccd1 _3386_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_6_2432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_2202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_3971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2337_ _4584_/Q _4583_/Q _2304_/D _2334_/B vssd1 vssd1 vccd1 vccd1 _2338_/B sky130_fd_sc_hd__a31o_1
XFILLER_6_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2458__A _3908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_2476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout192_A fanout193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5056_ _5056_/A vssd1 vssd1 vccd1 vccd1 _5056_/X sky130_fd_sc_hd__buf_2
XFILLER_6_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2268_ _4541_/Q _4540_/Q vssd1 vssd1 vccd1 vccd1 _2268_/Y sky130_fd_sc_hd__xnor2_2
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
+ _4801_/Q _2781_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_35_4009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4291__CLK _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4007_ _3932_/B _3935_/B _4007_/S vssd1 vssd1 vccd1 vccd1 _4009_/B sky130_fd_sc_hd__mux2_1
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2199_ _4509_/Q _4508_/Q vssd1 vssd1 vccd1 vccd1 _2199_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_25_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_3753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3289__A _5058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2193__A _2608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_4031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_4042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4909_ _3504_/Y _4909_/D _3614_/Y vssd1 vssd1 vccd1 vccd1 _4909_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2921__A _4896_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_4086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_3385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2640__B _2640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3752__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_3553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_3492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_2841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input18_A phi1b_dig_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_2827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_2849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
+ _4859_/Q _2881_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_3624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2550__B _4712_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_4060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_4143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output86_A _5083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_TE_B _1921_/Y vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3662__A _3669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3947_/A _3438_/B vssd1 vssd1 vccd1 vccd1 _3240_/Y sky130_fd_sc_hd__xnor2_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _3925_/A _3442_/B vssd1 vssd1 vccd1 vccd1 _3171_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_7_2796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2122_ _4007_/S _2122_/B vssd1 vssd1 vccd1 vccd1 _5093_/A sky130_fd_sc_hd__xnor2_1
XFILLER_23_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2053_ _4430_/Q _2053_/B vssd1 vssd1 vccd1 vccd1 _2054_/B sky130_fd_sc_hd__nor2_1
XFILLER_1_2351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_2362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_4097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2955_ _4919_/Q _4918_/Q vssd1 vssd1 vccd1 vccd1 _2955_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_34_2673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_2504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout128/X fanout246/X vssd1 vssd1 vccd1 vccd1 _5077_/A sky130_fd_sc_hd__dlrtn_1
X_1906_ _1904_/X _1905_/Y _1823_/X vssd1 vssd1 vccd1 vccd1 _1907_/B sky130_fd_sc_hd__o21ai_1
X_2886_ _4887_/Q _4886_/Q vssd1 vssd1 vccd1 vccd1 _2886_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__3556__B _3556_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_3694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4625_ _5043_/A _4625_/D fanout222/X vssd1 vssd1 vccd1 vccd1 _4625_/Q sky130_fd_sc_hd__dfstp_1
X_1837_ _1909_/A _1837_/B vssd1 vssd1 vccd1 vccd1 _1838_/B sky130_fd_sc_hd__nand2_1
XFILLER_15_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_2993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_3206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4556_ input27/X _4556_/D fanout199/X vssd1 vssd1 vccd1 vccd1 _4557_/D sky130_fd_sc_hd__dfrtp_1
X_1768_ _5030_/Q _1768_/B vssd1 vssd1 vccd1 vccd1 _5031_/D sky130_fd_sc_hd__xnor2_1
XFILLER_28_3145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3507_ _3519_/A vssd1 vssd1 vccd1 vccd1 _3507_/Y sky130_fd_sc_hd__inv_2
X_4487_ _5042_/A _4487_/D fanout201/X vssd1 vssd1 vccd1 vccd1 _4487_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_3189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1699_ _3556_/A _3556_/B vssd1 vssd1 vccd1 vccd1 _1761_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__3572__A _3924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3438_ _3946_/A _3438_/B vssd1 vssd1 vccd1 vccd1 _3438_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2188__A _2327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5039_ _5047_/A vssd1 vssd1 vccd1 vccd1 _5039_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_2098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2916__A _2916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1820__A _1909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2635__B _2635_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_2415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_2437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_2893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3747__A _3748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2651__A _4834_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_2757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_3193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
+ _4589_/Q _2373_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__3482__A _3498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput42 _5039_/X vssd1 vssd1 vccd1 vccd1 cclk_I[7] sky130_fd_sc_hd__buf_2
Xoutput53 _5050_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_I[2] sky130_fd_sc_hd__buf_2
XFILLER_20_4108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput64 _5061_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_Q[5] sky130_fd_sc_hd__buf_2
XFILLER_8_3773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput75 _5072_/X vssd1 vssd1 vccd1 vccd1 fb1_I[0] sky130_fd_sc_hd__buf_2
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_2048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput86 _5083_/X vssd1 vssd1 vccd1 vccd1 fb1_Q[3] sky130_fd_sc_hd__buf_2
Xoutput97 _5094_/X vssd1 vssd1 vccd1 vccd1 sin_out[2] sky130_fd_sc_hd__buf_2
XFILLER_7_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_4051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_4073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_4095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_4037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_2646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_3525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_2960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2740_ _4800_/Q _2740_/B vssd1 vssd1 vccd1 vccd1 _4800_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__2561__A _4707_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2671_ _4765_/Q _2671_/B vssd1 vssd1 vccd1 vccd1 _4765_/D sky130_fd_sc_hd__xnor2_1
X_4410_ _3220_/Y _4410_/D _3756_/Y vssd1 vssd1 vccd1 vccd1 _4410_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3316__27_A _3366__32/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4341_ _3186_/Y _4341_/D _3765__105/Y vssd1 vssd1 vccd1 vccd1 _4341_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_3329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_3498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3392__A _3912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1905__A _4351_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4272_ _3151_/Y _4272_/D _5048_/A vssd1 vssd1 vccd1 vccd1 _4272_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3223_ _3233_/A vssd1 vssd1 vccd1 vccd1 _3223_/Y sky130_fd_sc_hd__inv_2
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3140__A2 _4188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2105_ _2105_/A vssd1 vssd1 vccd1 vccd1 _2107_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_2479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2736__A _4799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3085_ _4991_/Q _3085_/B vssd1 vssd1 vccd1 vccd1 _3086_/B sky130_fd_sc_hd__nor2_1
XFILLER_3_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2036_ _4431_/Q _4430_/Q _4429_/Q _2036_/D vssd1 vssd1 vccd1 vccd1 _2046_/C sky130_fd_sc_hd__and4_1
XANTENNA__2455__B _3684_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout155_A _4981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_2134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3987_ _4452_/Q vssd1 vssd1 vccd1 vccd1 _4451_/D sky130_fd_sc_hd__inv_2
XANTENNA__3567__A _3571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_2178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2938_ _4931_/D _4905_/Q _4903_/Q vssd1 vssd1 vccd1 vccd1 _2938_/X sky130_fd_sc_hd__and3_1
XFILLER_30_2312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_2323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_2334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3286__B _3372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2869_ _2867_/X _2868_/Y _2858_/X vssd1 vssd1 vccd1 vccd1 _2870_/B sky130_fd_sc_hd__o21ai_1
XFILLER_30_2367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4806__RESET_B fanout256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4608_ _3339_/Y _4608_/D _3697_/Y vssd1 vssd1 vccd1 vccd1 _4608_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_30_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4539_ _3296_/Y _4539_/D _3718_/Y vssd1 vssd1 vccd1 vccd1 _4539_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1815__A _3114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_2285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_2966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3477__A _3905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_2289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_2543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_3580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4972__CLK _3541_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_4041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3940__A _3940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_2755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2556__A _4712_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4352__CLK input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3419__38 _3425__41/A vssd1 vssd1 vccd1 vccd1 _3419__38/Y sky130_fd_sc_hd__inv_2
XANTENNA__2275__B _4556_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3910_ _3910_/A _3910_/B vssd1 vssd1 vccd1 vccd1 _3914_/C sky130_fd_sc_hd__nand2_1
X_4890_ _5046_/A _4890_/D fanout237/X vssd1 vssd1 vccd1 vccd1 _4890_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2633__A1 _3941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3841_ _4358_/Q vssd1 vssd1 vccd1 vccd1 _4358_/D sky130_fd_sc_hd__inv_2
XFILLER_18_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3387__A _3393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_2020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2723_ _4838_/D _4812_/Q _4810_/Q _4809_/Q vssd1 vssd1 vccd1 vccd1 _2760_/A sky130_fd_sc_hd__or4_1
XFILLER_9_4002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_3301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2654_ _4766_/Q _4765_/Q _4764_/Q _2665_/B vssd1 vssd1 vccd1 vccd1 _2659_/B sky130_fd_sc_hd__or4_2
XFILLER_9_3323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2585_ _4711_/Q _2585_/B vssd1 vssd1 vccd1 vccd1 _4711_/D sky130_fd_sc_hd__xnor2_1
XFILLER_25_3115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_3137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4324_ _4324_/CLK _4324_/D fanout194/X vssd1 vssd1 vccd1 vccd1 _4324_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_25_2403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout106 _3135_/Y vssd1 vssd1 vccd1 vccd1 _5047_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_2655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout117 _4803_/CLK vssd1 vssd1 vccd1 vccd1 _4811_/CLK sky130_fd_sc_hd__clkbuf_4
Xfanout128 _3632_/A vssd1 vssd1 vccd1 vccd1 fanout128/X sky130_fd_sc_hd__buf_2
X_4255_ _4844_/Q _4255_/B vssd1 vssd1 vccd1 vccd1 _4845_/D sky130_fd_sc_hd__xnor2_1
Xfanout139 _2285_/Y vssd1 vssd1 vccd1 vccd1 _5042_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4186_ _4189_/A _4190_/A vssd1 vssd1 vccd1 vccd1 _4248_/D sky130_fd_sc_hd__xnor2_4
XFILLER_28_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_2171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_2182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3137_ _2978_/B _3136_/X _4248_/A vssd1 vssd1 vccd1 vccd1 _3137_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_3865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3068_ _4986_/Q _4985_/Q _3068_/C vssd1 vssd1 vccd1 vccd1 _3068_/X sky130_fd_sc_hd__and3_1
XFILLER_19_2207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2185__B _2185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2019_ _4462_/D _4389_/Q vssd1 vssd1 vccd1 vccd1 _2020_/D sky130_fd_sc_hd__xnor2_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_4129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3297__A _3309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4995__CLK _5047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_TE_B
+ _2030_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_3721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_3765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4375__CLK _3598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_2867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2376__A _4620_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_2878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__0630_ clkbuf_0__0630_/X vssd1 vssd1 vccd1 vccd1 _3732__95/A sky130_fd_sc_hd__clkbuf_16
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4799__RESET_B fanout247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4741__D _4741_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_2097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3935__A _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_4103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4310__RESET_B fanout194/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
+ _4393_/Q _2027_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_26_3424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_2712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4718__CLK _4718_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2370_ _4604_/Q _4603_/Q vssd1 vssd1 vccd1 vccd1 _2370_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3670__A _5060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4040_ _4534_/Q vssd1 vssd1 vccd1 vccd1 _4535_/D sky130_fd_sc_hd__inv_2
XFILLER_4_3275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_2541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_3297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4868__CLK _4905_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout144/X fanout215/X vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_0_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4942_ _3527_/Y _4942_/D _3603__77/Y vssd1 vssd1 vccd1 vccd1 _4942_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_2705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4873_ _3483_/Y _4873_/D _3625_/Y vssd1 vssd1 vccd1 vccd1 _4873_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_3862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_3873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4469__RESET_B fanout201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3824_ _4336_/Q vssd1 vssd1 vccd1 vccd1 _4337_/D sky130_fd_sc_hd__inv_2
XFILLER_21_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3755_ _3948_/A vssd1 vssd1 vccd1 vccd1 _3755_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3845__A _3882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2706_ _3114_/A _4776_/Q vssd1 vssd1 vccd1 vccd1 _4776_/D sky130_fd_sc_hd__xor2_1
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_GATE_N
+ _3632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3686_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3686_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout118_A _5045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2637_ _4124_/B _4003_/C vssd1 vssd1 vccd1 vccd1 _2978_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4398__CLK _4402_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2568_ _4709_/Q _2568_/B vssd1 vssd1 vccd1 vccd1 _2569_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_2474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4307_ _3888_/A _4307_/D _3775__114/Y vssd1 vssd1 vccd1 vccd1 _4307_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_3905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3580__A _3587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2499_ _2490_/C _2498_/X _2344_/X vssd1 vssd1 vccd1 vccd1 _2500_/B sky130_fd_sc_hd__o21ai_1
XFILLER_21_2108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_2277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4238_ _4828_/Q vssd1 vssd1 vccd1 vccd1 _4827_/D sky130_fd_sc_hd__inv_2
XFILLER_22_3877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4169_ _4724_/Q vssd1 vssd1 vccd1 vccd1 _4725_/D sky130_fd_sc_hd__inv_2
XFILLER_3_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2924__A _3030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5023__CLK input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_4040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4892__RESET_B fanout236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_2936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_4084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_2237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3755__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_3711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_2907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3418__37_A _3469__42/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3490__A _3498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3089__A1 _4992_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_2725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1870_ _1868_/X _1869_/Y _1791_/X vssd1 vssd1 vccd1 vccd1 _1871_/B sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_1_0_0_w0.cclk_I_A clkbuf_0_w0.cclk_I/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_2771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3665__A _3669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3540_ _3550_/A vssd1 vssd1 vccd1 vccd1 _3540_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4540__CLK _4063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3384__B _3438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_TE_B
+ _2023_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2422_ _2375_/C _2418_/Y _2344_/X vssd1 vssd1 vccd1 vccd1 _2423_/B sky130_fd_sc_hd__o21ai_1
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4690__CLK _4916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_2542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2353_ _4648_/D _4590_/Q _4588_/Q vssd1 vssd1 vccd1 vccd1 _2353_/X sky130_fd_sc_hd__and3_1
XFILLER_26_2553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_2586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5072_ _5072_/A vssd1 vssd1 vccd1 vccd1 _5072_/X sky130_fd_sc_hd__clkbuf_1
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout158/X fanout205/X vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__dlrtn_1
X_2284_ _2284_/A vssd1 vssd1 vccd1 vccd1 _2284_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3258__18_A _3262__21/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4023_ _4503_/Q vssd1 vssd1 vccd1 vccd1 _4502_/D sky130_fd_sc_hd__inv_2
XFILLER_0_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_2196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4925_ _3520_/Y _4925_/D _3605_/Y vssd1 vssd1 vccd1 vccd1 _4925_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_3247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_3258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout235_A input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4856_ _4905_/CLK _4856_/D fanout226/X vssd1 vssd1 vccd1 vccd1 _4856_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_3692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3807_ _4305_/Q vssd1 vssd1 vccd1 vccd1 _4304_/D sky130_fd_sc_hd__inv_2
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4787_ _5013_/CLK _4787_/D _3437_/Y vssd1 vssd1 vccd1 vccd1 _4787_/Q sky130_fd_sc_hd__dfrtp_2
X_1999_ _4398_/Q _1962_/D _1992_/B vssd1 vssd1 vccd1 vccd1 _2000_/B sky130_fd_sc_hd__a21bo_1
XFILLER_11_2833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3738_ _3738_/A vssd1 vssd1 vccd1 vccd1 _3748_/A sky130_fd_sc_hd__buf_8
XFILLER_10_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3294__B _3491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3669_ _3669_/A vssd1 vssd1 vccd1 vccd1 _3669_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_3939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3576_/A fanout251/X vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_9_2282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1823__A _2922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5020__RESET_B fanout207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4556__D _4556_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_3779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_4113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4413__CLK _3931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_3445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4563__CLK _5030_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3485__A _4189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_3541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_2978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_2809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4466__D _4466_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2809__A1 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4743__RESET_B fanout212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4906__CLK _1700_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[2\].w1.ro_block_I.ro_pol_eve.tribuf.t_buf _2453_/A _2301_/Y vssd1
+ vssd1 vccd1 vccd1 _5089_/A sky130_fd_sc_hd__ebufn_8
X_2971_ _3929_/A _4063_/C _4123_/B vssd1 vssd1 vccd1 vccd1 _2978_/D sky130_fd_sc_hd__a21oi_1
X_4710_ _4712_/CLK _4710_/D fanout243/X vssd1 vssd1 vccd1 vccd1 _4710_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1922_ _4341_/Q _4340_/Q vssd1 vssd1 vccd1 vccd1 _1922_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_2877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_3843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1853_ _4307_/Q _4306_/Q vssd1 vssd1 vccd1 vccd1 _1853_/Y sky130_fd_sc_hd__xnor2_2
X_4641_ _4852_/CLK _4641_/D _3357_/Y vssd1 vssd1 vccd1 vccd1 _4641_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_2118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_2287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_3887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1908__A _4351_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4572_ _3319_/Y _4572_/D _3707__92/Y vssd1 vssd1 vccd1 vccd1 _4572_/Q sky130_fd_sc_hd__dfrtp_1
X_1784_ _4282_/Q _4281_/Q _4280_/Q _1810_/B vssd1 vssd1 vccd1 vccd1 _1799_/B sky130_fd_sc_hd__or4_1
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_A
+ _4614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4003__B _4131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3454_ _3466_/A vssd1 vssd1 vccd1 vccd1 _3454_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2405_ _4618_/Q _2405_/B vssd1 vssd1 vccd1 vccd1 _2405_/X sky130_fd_sc_hd__and2b_1
X_3385_ _3393_/A vssd1 vssd1 vccd1 vccd1 _3385_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_3095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2336_ _4581_/Q _2336_/B vssd1 vssd1 vccd1 vccd1 _4581_/D sky130_fd_sc_hd__xnor2_1
XFILLER_29_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2458__B _2807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4436__CLK _5041_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5055_ _5055_/A vssd1 vssd1 vccd1 vccd1 _5055_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2267_ _4539_/Q _4538_/Q vssd1 vssd1 vccd1 vccd1 _2267_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_6_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4006_ _4473_/Q _4472_/Q vssd1 vssd1 vccd1 vccd1 _4007_/S sky130_fd_sc_hd__xnor2_2
X_2198_ _4507_/Q _4506_/Q vssd1 vssd1 vccd1 vccd1 _2198_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_26_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_3721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4586__CLK _4623_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2193__B _4497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_2018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout119/X fanout248/X vssd1 vssd1 vccd1 vccd1 _5078_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_16_2029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_3629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4908_ _4247_/Y _4908_/D _3503_/Y vssd1 vssd1 vccd1 vccd1 _4908_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_2917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4839_ input22/X _4839_/D fanout227/X vssd1 vssd1 vccd1 vccd1 _4840_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_11_3353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1818__A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_2685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_3510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4929__CLK input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_3821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_2416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4309__CLK _3882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2550__C _4711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3943__A _4131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_2957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1950__A1 _3888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4459__CLK _1952_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output79_A _5076_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2559__A _2996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3760__100 _3759__99/A vssd1 vssd1 vccd1 vccd1 _3760__100/Y sky130_fd_sc_hd__inv_2
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4995__RESET_B fanout242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3170_ _3923_/A vssd1 vssd1 vccd1 vccd1 _3442_/B sky130_fd_sc_hd__buf_12
XANTENNA__2278__B _2278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3213__17_A _3264__22/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2121_ _2121_/A _2121_/B vssd1 vssd1 vccd1 vccd1 _2122_/B sky130_fd_sc_hd__or2_1
XFILLER_23_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_3042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_2589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2052_ _4427_/Q _2052_/B vssd1 vssd1 vccd1 vccd1 _4427_/D sky130_fd_sc_hd__xnor2_1
XFILLER_1_3097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_4010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_4032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_3331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_2349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_3949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2954_ _4917_/Q _4916_/Q vssd1 vssd1 vccd1 vccd1 _2954_/Y sky130_fd_sc_hd__xnor2_2
Xclkbuf_1_0__f__1628_ clkbuf_0__1628_/X vssd1 vssd1 vccd1 vccd1 _3169__65/A sky130_fd_sc_hd__clkbuf_16
XFILLER_34_2685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_2062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1905_ _4351_/D _4325_/Q _4323_/Q vssd1 vssd1 vccd1 vccd1 _1905_/Y sky130_fd_sc_hd__nor3_1
XFILLER_15_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2885_ _4885_/Q _4884_/Q vssd1 vssd1 vccd1 vccd1 _2885_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_30_2538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4624_ _4626_/CLK _4624_/D fanout236/X vssd1 vssd1 vccd1 vccd1 _4624_/Q sky130_fd_sc_hd__dfrtp_1
X_1836_ _4347_/D _4289_/Q vssd1 vssd1 vccd1 vccd1 _1837_/B sky130_fd_sc_hd__xnor2_1
XFILLER_11_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1767_ _5031_/Q _1768_/B vssd1 vssd1 vccd1 vccd1 _5030_/D sky130_fd_sc_hd__xnor2_1
X_4555_ input27/X _4555_/D fanout202/X vssd1 vssd1 vccd1 vccd1 _4556_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_28_3157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3506_ _4189_/A _4190_/A vssd1 vssd1 vccd1 vccd1 _3506_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_2423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1698_ _4936_/Q vssd1 vssd1 vccd1 vccd1 _3556_/B sky130_fd_sc_hd__clkbuf_4
X_4486_ _5042_/A _4486_/D fanout201/X vssd1 vssd1 vccd1 vccd1 _4486_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_28_2456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3572__B _3923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3437_ _3445_/A vssd1 vssd1 vccd1 vccd1 _3437_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_2478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_2489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_2230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _3470_/A vssd1 vssd1 vccd1 vccd1 _3368_/X sky130_fd_sc_hd__buf_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2319_ _4578_/Q _2315_/C _2316_/B vssd1 vssd1 vccd1 vccd1 _2320_/B sky130_fd_sc_hd__a21bo_1
XFILLER_22_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3299_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3299_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3160__60 _3169__65/A vssd1 vssd1 vccd1 vccd1 _3160__60/Y sky130_fd_sc_hd__inv_2
X_5038_ _5046_/A vssd1 vssd1 vccd1 vccd1 _5038_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4834__D _4834_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
+ _4990_/Q _3116_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_13_2725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4601__CLK _4981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput43 _5040_/X vssd1 vssd1 vccd1 vccd1 cclk_Q[0] sky130_fd_sc_hd__clkbuf_1
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput54 _5051_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_I[3] sky130_fd_sc_hd__buf_2
XFILLER_4_3605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_3533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput65 _5062_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_Q[6] sky130_fd_sc_hd__buf_2
Xoutput76 _5073_/X vssd1 vssd1 vccd1 vccd1 fb1_I[1] sky130_fd_sc_hd__buf_2
XFILLER_24_3555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput87 _5084_/X vssd1 vssd1 vccd1 vccd1 fb1_Q[4] sky130_fd_sc_hd__buf_2
XFILLER_1_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput98 _5095_/X vssd1 vssd1 vccd1 vccd1 sin_out[3] sky130_fd_sc_hd__buf_2
XANTENNA__4751__CLK _5030_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input30_A phi1b_dig_Q[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_4085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_3290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_2650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3003__A _3030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_2603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3938__A _3946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2842__A _2916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_2825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_4112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_2257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2670_ _2680_/A _2670_/B vssd1 vssd1 vccd1 vccd1 _2671_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_3411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4281__CLK _4281_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3673__A _4135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4340_ _2294_/B1 _4340_/D _3185__70/Y vssd1 vssd1 vccd1 vccd1 _4340_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_2743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3392__B _3446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_2776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4271_ _3846_/A _4271_/D _5048_/A vssd1 vssd1 vccd1 vccd1 _4271_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_3273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3222_ _3925_/A _3442_/B vssd1 vssd1 vccd1 vccd1 _3222_/Y sky130_fd_sc_hd__xnor2_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_GATE_N _4363_/CLK
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_2353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_2375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2104_ _4464_/Q _4463_/D vssd1 vssd1 vccd1 vccd1 _2105_/A sky130_fd_sc_hd__and2b_1
XFILLER_23_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3084_ _4988_/Q _3084_/B vssd1 vssd1 vccd1 vccd1 _4988_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__2736__B _2736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2580__A_N _4711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2035_ _4434_/Q _4433_/Q _4432_/Q _2035_/D vssd1 vssd1 vccd1 vccd1 _2036_/D sky130_fd_sc_hd__and4_1
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5056_/A fanout190/X vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_18_3871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3848__A _3848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_3893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_3757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3986_ _4449_/Q vssd1 vssd1 vccd1 vccd1 _4450_/D sky130_fd_sc_hd__inv_2
XANTENNA_fanout148_A _2114_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2937_ _4901_/Q _2937_/B vssd1 vssd1 vccd1 vccd1 _4901_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__4624__CLK _4626_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2868_ _4927_/D _4869_/Q _4867_/Q vssd1 vssd1 vccd1 vccd1 _2868_/Y sky130_fd_sc_hd__nor3_1
XFILLER_12_3492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3767__106 _3770__109/A vssd1 vssd1 vccd1 vccd1 _3767__106/Y sky130_fd_sc_hd__inv_2
X_4607_ _3861_/Y _4607_/D _3338_/Y vssd1 vssd1 vccd1 vccd1 _4607_/Q sky130_fd_sc_hd__dfrtp_1
X_1819_ _4283_/Q _1778_/D _1810_/B vssd1 vssd1 vccd1 vccd1 _1820_/B sky130_fd_sc_hd__a21bo_1
X_2799_ _3877_/A _2799_/B vssd1 vssd1 vccd1 vccd1 _2799_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3583__A _3587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
+ _4705_/Q _2616_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__4774__CLK _4812_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4538_ _4063_/C _4538_/D _3295_/Y vssd1 vssd1 vccd1 vccd1 _4538_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_2253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4469_ _3257_/Y _4469_/D fanout201/X vssd1 vssd1 vccd1 vccd1 _4469_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2927__A _3030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_TE_B
+ _2544_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_4093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3758__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3477__B _3913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_A
+ _4763_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3493__A _3946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_3628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_4086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_2892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2837__A _4859_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_2684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2556__B _4711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
+ _4763_/Q _2713_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_18_3101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_2491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4647__CLK input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2633__A2 _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3668__A _3669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2572__A _2922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3840_ _4357_/Q vssd1 vssd1 vccd1 vccd1 _4357_/D sky130_fd_sc_hd__inv_2
XFILLER_18_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_2600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2722_ _4800_/Q _4799_/Q _2730_/C _2733_/A vssd1 vssd1 vccd1 vccd1 _2774_/B sky130_fd_sc_hd__a31o_1
XANTENNA__4797__CLK _4811_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_2666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2653_ _4769_/Q _4768_/Q _4767_/Q _2675_/B vssd1 vssd1 vccd1 vccd1 _2665_/B sky130_fd_sc_hd__or4_1
XFILLER_29_3230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2149__A1 _4485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_2098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_4069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2584_ _2680_/A _2584_/B vssd1 vssd1 vccd1 vccd1 _2585_/B sky130_fd_sc_hd__nand2_1
XFILLER_12_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_3127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4323_ _4324_/CLK _4323_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _4323_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_3149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout107 _4905_/CLK vssd1 vssd1 vccd1 vccd1 _4865_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_9_2667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout118 _5045_/A vssd1 vssd1 vccd1 vccd1 _4803_/CLK sky130_fd_sc_hd__buf_2
Xfanout129 _5061_/A vssd1 vssd1 vccd1 vccd1 _3632_/A sky130_fd_sc_hd__buf_4
XFILLER_7_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4254_ _4845_/Q _4255_/B vssd1 vssd1 vccd1 vccd1 _4844_/D sky130_fd_sc_hd__xnor2_1
XFILLER_29_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3205_ _3600_/A vssd1 vssd1 vccd1 vccd1 _3205_/X sky130_fd_sc_hd__buf_1
XANTENNA__3197__5_A _3199__7/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4185_ _4750_/Q vssd1 vssd1 vccd1 vccd1 _4190_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_3_2233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_3761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout136/X fanout239/X vssd1 vssd1 vccd1 vccd1 _5084_/A sky130_fd_sc_hd__dlrtn_1
X_3136_ _4123_/A _4123_/B vssd1 vssd1 vccd1 vccd1 _3136_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3067_ _4983_/Q _3067_/B vssd1 vssd1 vccd1 vccd1 _4983_/D sky130_fd_sc_hd__xor2_1
XFILLER_23_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2018_ _4402_/Q _2018_/B vssd1 vssd1 vccd1 vccd1 _4402_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__2085__B1 _2003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_3109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3578__A _3587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3969_ _4418_/Q vssd1 vssd1 vccd1 vccd1 _4417_/D sky130_fd_sc_hd__inv_2
XFILLER_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3736__98 _3759__99/A vssd1 vssd1 vccd1 vccd1 _3736__98/Y sky130_fd_sc_hd__inv_2
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf _4282_/Q _1845_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XANTENNA__4559__D _4559_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_3788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5033__A _5033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2376__B _4619_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3267__23 _3365__31/A vssd1 vssd1 vccd1 vccd1 _3267__23/Y sky130_fd_sc_hd__inv_2
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3488__A _3498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2392__A _2412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_2606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2379__A1 _4614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_3097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3935__B _3935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4768__RESET_B fanout256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_4115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_2829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_2757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_3287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_2553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2286__B _2286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4941_ _4943_/CLK _4941_/D _3526__51/Y vssd1 vssd1 vccd1 vccd1 _4941_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_17_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4932__D _4932_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3398__A _3414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4872_ _4247_/Y _4872_/D _3482_/Y vssd1 vssd1 vccd1 vccd1 _4872_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3823_ _4337_/Q vssd1 vssd1 vccd1 vccd1 _4336_/D sky130_fd_sc_hd__inv_2
XFILLER_21_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_A
+ _4896_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3476__46_A _3523__49/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3754_ _3948_/A vssd1 vssd1 vccd1 vccd1 _3754_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_3197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_2474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2705_ _4775_/Q _2705_/B vssd1 vssd1 vccd1 vccd1 _4775_/D sky130_fd_sc_hd__xor2_1
X_3685_ _3696_/A vssd1 vssd1 vccd1 vccd1 _3695_/A sky130_fd_sc_hd__buf_6
XANTENNA__4438__RESET_B fanout198/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2636_ _2459_/B _2457_/Y _2632_/X vssd1 vssd1 vccd1 vccd1 _2636_/X sky130_fd_sc_hd__o21a_1
XFILLER_12_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2567_ _4706_/Q _2567_/B vssd1 vssd1 vccd1 vccd1 _4706_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__3861__A _3897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_2453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4306_ _1952_/A1 _4306_/D _3161__61/Y vssd1 vssd1 vccd1 vccd1 _4306_/Q sky130_fd_sc_hd__dfrtp_1
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout144/X fanout217/X vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_5_2317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_2245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2498_ _4672_/Q _2498_/B vssd1 vssd1 vccd1 vccd1 _2498_/X sky130_fd_sc_hd__and2b_1
XFILLER_2_3917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4812__CLK _4812_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4237_ _4825_/Q vssd1 vssd1 vccd1 vccd1 _4826_/D sky130_fd_sc_hd__inv_2
XANTENNA__2477__A _4741_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_2052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4168_ _4725_/Q vssd1 vssd1 vccd1 vccd1 _4724_/D sky130_fd_sc_hd__inv_2
XFILLER_20_3580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_2085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3119_ _5008_/Q _5007_/Q vssd1 vssd1 vccd1 vccd1 _3119_/Y sky130_fd_sc_hd__xnor2_2
X_4099_ _4609_/Q vssd1 vssd1 vccd1 vccd1 _4610_/D sky130_fd_sc_hd__clkinv_2
XFILLER_19_2005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4962__CLK _4962_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4342__CLK _1952_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
+ _4524_/Q _2267_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_30_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_4023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4492__CLK _5042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_4078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2387__A _4614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3089__A2 _4991_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2818__C _4861_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_2665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_4141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3011__A _4951_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4949__RESET_B fanout210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3946__A _3946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4531__RESET_B fanout212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3470_ _3470_/A vssd1 vssd1 vccd1 vccd1 _3470_/X sky130_fd_sc_hd__buf_1
XFILLER_6_3305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2421_ _4621_/Q _2421_/B vssd1 vssd1 vccd1 vccd1 _4621_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__4835__CLK input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_2615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2352_ _4586_/Q _2352_/B vssd1 vssd1 vccd1 vccd1 _4586_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__4927__D _4927_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5071_ _5071_/A vssd1 vssd1 vccd1 vccd1 _5071_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_3051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2297__A _3929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2283_ _2283_/A _2283_/B vssd1 vssd1 vccd1 vccd1 _2284_/A sky130_fd_sc_hd__or2_1
XFILLER_26_2598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4985__CLK _4997_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4022_ _4500_/Q vssd1 vssd1 vccd1 vccd1 _4501_/D sky130_fd_sc_hd__inv_2
XANTENNA__2288__B1 _3892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
+ _4582_/Q _2365_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_2203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4924_ _4943_/CLK _4924_/D _3519_/Y vssd1 vssd1 vccd1 vccd1 _4924_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4855_ _4905_/CLK _4855_/D fanout228/X vssd1 vssd1 vccd1 vccd1 _4855_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_2558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3806_ _4302_/Q vssd1 vssd1 vccd1 vccd1 _4303_/D sky130_fd_sc_hd__inv_2
XANTENNA__4365__CLK _4472_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout130_A _4748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4786_ _3436_/Y _4786_/D _3648_/Y vssd1 vssd1 vccd1 vccd1 _4786_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout228_A fanout230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1998_ _4396_/Q _1998_/B vssd1 vssd1 vccd1 vccd1 _4396_/D sky130_fd_sc_hd__xnor2_1
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3737_ _5057_/A vssd1 vssd1 vccd1 vccd1 _3737_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_2878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4272__RESET_B _5048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3668_ _3669_/A vssd1 vssd1 vccd1 vccd1 _3668_/Y sky130_fd_sc_hd__inv_2
X_2619_ _4743_/Q _4742_/D vssd1 vssd1 vccd1 vccd1 _2620_/A sky130_fd_sc_hd__and2b_1
XFILLER_27_2329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3591__A _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3182__69 _3189__72/A vssd1 vssd1 vccd1 vccd1 _3182__69/Y sky130_fd_sc_hd__inv_2
XFILLER_22_3642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_3675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2000__A _2061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4708__CLK _4712_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3766__A _3777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2670__A _2680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_2057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3485__B _4190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_2322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5055_/A fanout244/X vssd1 vssd1 vccd1 vccd1 _5079_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_14_2491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4858__CLK _4865_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3163__63_A _3169__65/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_2896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_3185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2845__A _2916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3199__7 _3199__7/A vssd1 vssd1 vccd1 vccd1 _4368_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2970_ _3929_/A _4248_/A vssd1 vssd1 vccd1 vccd1 _2978_/C sky130_fd_sc_hd__nand2_1
XFILLER_34_3557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1921_ _4339_/Q _4338_/Q vssd1 vssd1 vccd1 vccd1 _1921_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_19_2391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3676__A _4135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4640_ _3356_/Y _4640_/D _3688_/Y vssd1 vssd1 vccd1 vccd1 _4640_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4712__RESET_B fanout256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1852_ _4305_/Q _4304_/Q vssd1 vssd1 vccd1 vccd1 _1852_/Y sky130_fd_sc_hd__xnor2_2
X_4571_ _3855_/Y _4571_/D _3318__28/Y vssd1 vssd1 vccd1 vccd1 _4571_/Q sky130_fd_sc_hd__dfrtp_1
X_1783_ _4285_/Q _4284_/Q _4283_/Q _1826_/A vssd1 vssd1 vccd1 vccd1 _1810_/B sky130_fd_sc_hd__or4_4
XFILLER_28_3339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4003__C _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3453_ _4127_/A _4129_/A vssd1 vssd1 vccd1 vccd1 _3453_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_26_3030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5013__CLK _5013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2404_ _4619_/Q _2404_/B vssd1 vssd1 vccd1 vccd1 _2405_/B sky130_fd_sc_hd__nor2_1
X_3384_ _3947_/A _3438_/B vssd1 vssd1 vccd1 vccd1 _3384_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_6_3157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_3940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_2351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2335_ _2305_/D _2334_/X _2173_/X vssd1 vssd1 vccd1 vccd1 _2336_/B sky130_fd_sc_hd__o21ai_1
XFILLER_23_3962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5054_ _5062_/A vssd1 vssd1 vccd1 vccd1 _5054_/X sky130_fd_sc_hd__clkbuf_1
X_2266_ _4537_/Q _4536_/Q vssd1 vssd1 vccd1 vccd1 _2266_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_22_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4005_ _4005_/A _4005_/B vssd1 vssd1 vccd1 vccd1 _4471_/D sky130_fd_sc_hd__xnor2_1
X_2197_ _4505_/Q _4504_/Q vssd1 vssd1 vccd1 vccd1 _2197_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout178_A _3857_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_3744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_3012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4907_ _3502_/Y _4907_/D _3615_/Y vssd1 vssd1 vccd1 vccd1 _4907_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_2907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3586__A _3587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_4066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2490__A _4671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4838_ input22/X _4838_/D fanout231/X vssd1 vssd1 vccd1 vccd1 _4839_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_33_2377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4769_ _4812_/CLK _4769_/D fanout250/X vssd1 vssd1 vccd1 vccd1 _4769_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_28_3862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_2126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3159__59_A _3159__59/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_2771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4530__CLK _4532_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5041__A _5041_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_3221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4680__CLK _4719_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3496__A _3498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_2564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_2428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2727__A1 _4799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_4040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1950__A2 _3914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_2693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_2607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2120_ _3931_/A _2118_/X _2119_/X _3901_/A vssd1 vssd1 vccd1 vccd1 _2121_/B sky130_fd_sc_hd__o22a_1
XFILLER_3_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2051_ _2061_/A _2051_/B vssd1 vssd1 vccd1 vccd1 _2052_/B sky130_fd_sc_hd__nand2_1
XANTENNA__2575__A _4708_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_4044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_2317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2415__B1 _2344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2953_ _4915_/Q _4914_/Q vssd1 vssd1 vccd1 vccd1 _2953_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_34_3387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_2653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1904_ _4351_/D _4325_/Q _4323_/Q vssd1 vssd1 vccd1 vccd1 _1904_/X sky130_fd_sc_hd__and3_1
X_2884_ _4883_/Q _4882_/Q vssd1 vssd1 vccd1 vccd1 _2884_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_34_2697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_2528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4623_ _4623_/CLK _4623_/D fanout236/X vssd1 vssd1 vccd1 vccd1 _4623_/Q sky130_fd_sc_hd__dfrtp_1
X_1835_ _4286_/Q _1835_/B vssd1 vssd1 vccd1 vccd1 _4286_/D sky130_fd_sc_hd__xnor2_1
XFILLER_12_2951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout180/X fanout184/X vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__dlrtn_1
X_4554_ input27/X _4554_/D fanout207/X vssd1 vssd1 vccd1 vccd1 _4555_/D sky130_fd_sc_hd__dfrtp_4
X_1766_ _4250_/B _3144_/A _1765_/X vssd1 vssd1 vccd1 vccd1 _1768_/B sky130_fd_sc_hd__a21bo_1
X_3505_ _3519_/A vssd1 vssd1 vccd1 vccd1 _3505_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4403__CLK _4429_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4485_ _5042_/A _4485_/D fanout205/X vssd1 vssd1 vccd1 vccd1 _4485_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_2507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1697_ _4935_/Q vssd1 vssd1 vccd1 vccd1 _3556_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_8_2518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3436_ _4004_/A _3491_/B vssd1 vssd1 vccd1 vccd1 _3436_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__3143__A1 _4248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _3895_/A _3372_/B vssd1 vssd1 vccd1 vccd1 _3367_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_6_2242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ _2318_/A _2318_/B vssd1 vssd1 vccd1 vccd1 _4576_/D sky130_fd_sc_hd__xnor2_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3298_ _3935_/A _3440_/B vssd1 vssd1 vccd1 vccd1 _3298_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_26_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5037_ _5045_/A vssd1 vssd1 vccd1 vccd1 _5037_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2485__A _4676_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2249_ _2248_/Y _2206_/C _4529_/Q vssd1 vssd1 vccd1 vccd1 _2250_/B sky130_fd_sc_hd__mux2_1
XFILLER_19_3806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_w0.ro_block_Q.ro_pol.tribuf.t_buf_TE_B _1770_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2406__B1 _2344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_2737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_2185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_3785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5036__A _5044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_3501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_3681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput44 _5041_/X vssd1 vssd1 vccd1 vccd1 cclk_Q[1] sky130_fd_sc_hd__buf_2
Xoutput55 _5052_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_I[4] sky130_fd_sc_hd__buf_2
XFILLER_7_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput66 _5063_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_Q[7] sky130_fd_sc_hd__buf_2
Xoutput77 _5074_/X vssd1 vssd1 vccd1 vccd1 fb1_I[2] sky130_fd_sc_hd__buf_2
XFILLER_27_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput88 _5085_/X vssd1 vssd1 vccd1 vccd1 fb1_Q[5] sky130_fd_sc_hd__buf_2
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput99 _5096_/X vssd1 vssd1 vccd1 vccd1 sin_out[4] sky130_fd_sc_hd__buf_2
XFILLER_24_2844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input23_A phi1b_dig_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_4017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_2673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4375__RESET_B fanout214/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3938__B _3945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_3950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3070__B1 _2143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_2203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2561__C _2561_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4426__CLK _5033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output91_A _5088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4576__CLK _5043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4270_ _3150_/Y _4270_/D _4359_/CLK vssd1 vssd1 vccd1 vccd1 _4270_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_2608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_2788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3221_ _3233_/A vssd1 vssd1 vccd1 vccd1 _3221_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_3285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_3149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_2365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2103_ _4460_/Q _4459_/Q vssd1 vssd1 vccd1 vccd1 _2103_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_7_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3083_ _3109_/A _3083_/B vssd1 vssd1 vccd1 vccd1 _3084_/B sky130_fd_sc_hd__nand2_1
XFILLER_3_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2034_ _4436_/Q _4435_/Q _2034_/C vssd1 vssd1 vccd1 vccd1 _2035_/D sky130_fd_sc_hd__and3_1
XFILLER_1_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3848__B _3848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3985_ _4450_/Q vssd1 vssd1 vccd1 vccd1 _4449_/D sky130_fd_sc_hd__inv_2
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2936_ _2889_/C _2932_/Y _2858_/X vssd1 vssd1 vccd1 vccd1 _2937_/B sky130_fd_sc_hd__o21ai_1
XFILLER_17_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_2483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_0_0_clk_master clkbuf_3_1_0_clk_master/A vssd1 vssd1 vccd1 vccd1 _5056_/A
+ sky130_fd_sc_hd__clkbuf_8
X_2867_ _4927_/D _4869_/Q _4867_/Q vssd1 vssd1 vccd1 vccd1 _2867_/X sky130_fd_sc_hd__and3_1
XFILLER_30_2347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3864__A _3905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_2770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4606_ _3337_/Y _4606_/D _3698_/Y vssd1 vssd1 vccd1 vccd1 _4606_/Q sky130_fd_sc_hd__dfrtp_1
X_1818_ _3112_/A vssd1 vssd1 vccd1 vccd1 _1909_/A sky130_fd_sc_hd__buf_4
XFILLER_11_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2798_ _3929_/A _4123_/B _2462_/Y _2457_/Y _4003_/C vssd1 vssd1 vccd1 vccd1 _2799_/B
+ sky130_fd_sc_hd__a221oi_1
X_4537_ _3294_/Y _4537_/D _3719_/Y vssd1 vssd1 vccd1 vccd1 _4537_/Q sky130_fd_sc_hd__dfrtp_1
X_1749_ _5010_/Q vssd1 vssd1 vccd1 vccd1 _5009_/D sky130_fd_sc_hd__inv_2
XFILLER_28_2210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_3904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4468_ input18/X _4468_/D fanout197/X vssd1 vssd1 vccd1 vccd1 _4468_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_3865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4399_ _4402_/CLK _4399_/D fanout189/X vssd1 vssd1 vccd1 vccd1 _4399_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5048_/A fanout191/X vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__dlrtn_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3104__A _5024_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_3614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2943__A _3030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_2946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3643_/A fanout243/X vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__dlrtn_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4449__CLK _3931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2381__C _4620_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_3279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4599__CLK _4920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_2870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3493__B _3945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_4104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_2939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3200__8_A _3201__9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4556__RESET_B fanout199/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_2538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf _4324_/Q _1924_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_20_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3014__A _4952_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2556__C _4710_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2853__A _4861_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_2401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_4014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_2309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2721_ _4798_/Q vssd1 vssd1 vccd1 vccd1 _2733_/A sky130_fd_sc_hd__inv_2
XFILLER_12_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_2055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2652_ _4772_/Q _4771_/Q _4770_/Q _2690_/A vssd1 vssd1 vccd1 vccd1 _2675_/B sky130_fd_sc_hd__or4_1
XFILLER_9_4037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_3242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_3253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2583_ _4713_/Q _4712_/Q _2550_/D _2580_/B vssd1 vssd1 vccd1 vccd1 _2584_/B sky130_fd_sc_hd__a31o_1
XFILLER_9_2602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4322_ _4324_/CLK _4322_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _4322_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout108 _5046_/A vssd1 vssd1 vccd1 vccd1 _4905_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout119 _5062_/A vssd1 vssd1 vccd1 vccd1 fanout119/X sky130_fd_sc_hd__clkbuf_2
X_4253_ _4248_/C _4251_/Y _4252_/Y vssd1 vssd1 vccd1 vccd1 _4255_/B sky130_fd_sc_hd__o21ai_1
XFILLER_25_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4184_ _4749_/Q vssd1 vssd1 vccd1 vccd1 _4189_/A sky130_fd_sc_hd__buf_12
X_3135_ _3576_/Y _5027_/D vssd1 vssd1 vccd1 vccd1 _3135_/Y sky130_fd_sc_hd__nor2_8
XFILLER_0_3834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_2256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_2289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3066_ _3066_/A _3112_/B _3112_/C vssd1 vssd1 vccd1 vccd1 _3067_/B sky130_fd_sc_hd__and3_1
XFILLER_3_1555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2017_ _2061_/A _2017_/B vssd1 vssd1 vccd1 vccd1 _2018_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout160_A _4000_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_GATE_N _4359_/CLK
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_TE_B
+ _2201_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_2821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3968_ _4415_/Q vssd1 vssd1 vccd1 vccd1 _4416_/D sky130_fd_sc_hd__inv_2
XANTENNA__4741__CLK input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2919_ _4897_/Q _2919_/B vssd1 vssd1 vccd1 vccd1 _2919_/X sky130_fd_sc_hd__and2b_1
XFILLER_10_2707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3594__A _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3899_ _3899_/A _3914_/A vssd1 vssd1 vccd1 vccd1 _3900_/B sky130_fd_sc_hd__nand2_1
XFILLER_12_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_2729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_1_w0.cclk_I clkbuf_1_1_1_w0.cclk_I/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_w0.cclk_I/A
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__4891__CLK _4901_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2003__A _2922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_3745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2938__A _4931_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_2825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
+ _4894_/Q _2953_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3659_/A fanout240/X vssd1 vssd1 vccd1 vccd1 _5076_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__2376__C _4618_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4271__CLK _3846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2673__A _2680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2379__A2 _4613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_4091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_2976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_GATE_N
+ fanout128/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3879__A2 _3925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_4070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2839__B1 _2687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_3277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4614__CLK _4623_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4390__RESET_B fanout194/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2286__C _3931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3679__A _4135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4940_ _3525_/Y _4940_/D _3604__78/Y vssd1 vssd1 vccd1 vccd1 _4940_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4764__CLK _4811_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1814__A1 _4283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4871_ _1761_/B _4871_/D _3626_/Y vssd1 vssd1 vccd1 vccd1 _4871_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_2253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_2729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3822_ _4334_/Q vssd1 vssd1 vccd1 vccd1 _4335_/D sky130_fd_sc_hd__inv_2
XFILLER_20_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
+ _4952_/Q _3048_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_3753_ _3948_/A vssd1 vssd1 vccd1 vccd1 _3753_/Y sky130_fd_sc_hd__inv_2
Xwrapper_cell_loop\[1\].w1.ro_block_Q.ro_pol.tribuf.t_buf _2279_/X _2128_/Y vssd1
+ vssd1 vccd1 vccd1 _5090_/A sky130_fd_sc_hd__ebufn_8
X_2704_ _3112_/A _2704_/B _2704_/C _2704_/D vssd1 vssd1 vccd1 vccd1 _2705_/B sky130_fd_sc_hd__and4_1
X_3684_ _3684_/A vssd1 vssd1 vccd1 vccd1 _3684_/Y sky130_fd_sc_hd__clkinv_4
X_2635_ _4192_/S _2635_/B vssd1 vssd1 vccd1 vccd1 _5096_/A sky130_fd_sc_hd__xnor2_1
XFILLER_9_3122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_3072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2566_ _2566_/A _2566_/B vssd1 vssd1 vccd1 vccd1 _2567_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4305_ _3892_/B _4305_/D _3776__115/Y vssd1 vssd1 vccd1 vccd1 _4305_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2497_ _4673_/Q _2497_/B vssd1 vssd1 vccd1 vccd1 _2498_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_1742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_2487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4236_ _4826_/Q vssd1 vssd1 vccd1 vccd1 _4825_/D sky130_fd_sc_hd__inv_2
XANTENNA__4294__CLK _3932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4167_ _4722_/Q vssd1 vssd1 vccd1 vccd1 _4723_/D sky130_fd_sc_hd__inv_2
XFILLER_25_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_2064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3118_ _5006_/Q _5005_/Q vssd1 vssd1 vccd1 vccd1 _3118_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_20_3592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4098_ _4610_/Q vssd1 vssd1 vccd1 vccd1 _4609_/D sky130_fd_sc_hd__inv_2
XFILLER_20_2880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3589__A _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3049_ _4972_/Q _4971_/Q vssd1 vssd1 vccd1 vccd1 _3049_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_19_2017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3007__B1 _2858_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_3975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1837__A _1909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_3757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4637__CLK _3922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2668__A _4764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_3470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5044__A _5044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2387__B _4613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4787__CLK _5013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_2749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3499__A _3916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3011__B _3011_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_2448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_TE_B
+ _2194_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_2773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4989__RESET_B fanout235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_3201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2420_ _2566_/A _2420_/B vssd1 vssd1 vccd1 vccd1 _2421_/B sky130_fd_sc_hd__nand2_1
X_3176__67 _3189__72/A vssd1 vssd1 vccd1 vccd1 _3176__67/Y sky130_fd_sc_hd__inv_2
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
+ _4682_/Q _2547_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_26_3267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2351_ _2303_/C _2347_/Y _2344_/X vssd1 vssd1 vccd1 vccd1 _2352_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__2578__A _4709_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5070_ _5070_/A vssd1 vssd1 vccd1 vccd1 _5070_/X sky130_fd_sc_hd__clkbuf_2
X_2282_ _4560_/D _4561_/Q vssd1 vssd1 vccd1 vccd1 _2283_/B sky130_fd_sc_hd__and2b_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4021_ _4501_/Q vssd1 vssd1 vccd1 vccd1 _4500_/D sky130_fd_sc_hd__inv_2
XFILLER_20_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_3205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4923_ _3518_/Y _4923_/D _3607_/Y vssd1 vssd1 vccd1 vccd1 _4923_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_3249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4854_ _4865_/CLK _4854_/D fanout228/X vssd1 vssd1 vccd1 vccd1 _4854_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3805_ _4303_/Q vssd1 vssd1 vccd1 vccd1 _4302_/D sky130_fd_sc_hd__inv_2
X_4785_ _2809_/A1 _4785_/D _3435_/Y vssd1 vssd1 vccd1 vccd1 _4785_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_18_1393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1997_ _2061_/A _1997_/B vssd1 vssd1 vccd1 vccd1 _1998_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout123_A _4719_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3667_ _3669_/A vssd1 vssd1 vccd1 vccd1 _3667_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3872__A _3888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2618_ _4739_/Q _4738_/Q vssd1 vssd1 vccd1 vccd1 _2618_/Y sky130_fd_sc_hd__xnor2_4
X_3598_ _3598_/A vssd1 vssd1 vccd1 vccd1 _3598_/X sky130_fd_sc_hd__buf_1
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2488__A _2996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2549_ _4715_/Q _4714_/Q _2549_/C vssd1 vssd1 vccd1 vccd1 _2550_/D sky130_fd_sc_hd__and3_1
XFILLER_22_3610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_2021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4219_ _4791_/Q vssd1 vssd1 vccd1 vccd1 _4792_/D sky130_fd_sc_hd__inv_2
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_2986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3112__A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_3403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2654__C _4764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_2713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1983__A_N _4393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3189__72_A _3189__72/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5039__A _5047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_A
+ _4710_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_3565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_2936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_3361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_2739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_2441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_2474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1920_ _4337_/Q _4336_/Q vssd1 vssd1 vccd1 vccd1 _1920_/Y sky130_fd_sc_hd__xnor2_4
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1851_ _4303_/Q _4302_/Q vssd1 vssd1 vccd1 vccd1 _1851_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4570_ _3317_/Y _4570_/D _3708__93/Y vssd1 vssd1 vccd1 vccd1 _4570_/Q sky130_fd_sc_hd__dfrtp_1
X_1782_ _4347_/D _4289_/Q _4287_/Q _4286_/Q vssd1 vssd1 vccd1 vccd1 _1826_/A sky130_fd_sc_hd__or4_1
X_3521_ _5062_/A vssd1 vssd1 vccd1 vccd1 _3521_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_3_5_0_clk_master clkbuf_3_5_0_clk_master/A vssd1 vssd1 vccd1 vccd1 _3598_/A
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__4752__RESET_B fanout223/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3692__A _3695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1953__B1 _3845_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3452_ _3466_/A vssd1 vssd1 vccd1 vccd1 _3452_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4952__CLK _4962_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2403_ _4616_/Q _2403_/B vssd1 vssd1 vccd1 vccd1 _4616_/D sky130_fd_sc_hd__xnor2_1
XFILLER_26_2330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3383_ _3393_/A vssd1 vssd1 vccd1 vccd1 _3383_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_3169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_2424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2334_ _4582_/Q _2334_/B vssd1 vssd1 vccd1 vccd1 _2334_/X sky130_fd_sc_hd__and2b_1
XFILLER_6_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_2446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_2457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_3996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5053_ _5061_/A vssd1 vssd1 vccd1 vccd1 _5053_/X sky130_fd_sc_hd__clkbuf_1
X_2265_ _4535_/Q _4534_/Q vssd1 vssd1 vccd1 vccd1 _2265_/Y sky130_fd_sc_hd__xnor2_2
X_4004_ _4004_/A _4005_/B vssd1 vssd1 vccd1 vccd1 _4470_/D sky130_fd_sc_hd__xnor2_1
XFILLER_2_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2196_ _4503_/Q _4502_/Q vssd1 vssd1 vccd1 vccd1 _2196_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4332__CLK _3931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4906_ _1700_/Y _4906_/D _3501_/Y vssd1 vssd1 vccd1 vccd1 _4906_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_3057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4482__CLK _4533_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4837_ input22/X input6/X fanout233/X vssd1 vssd1 vccd1 vccd1 _4838_/D sky130_fd_sc_hd__dfrtp_4
XANTENNA__2490__B _4670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4768_ _4811_/CLK _4768_/D fanout256/X vssd1 vssd1 vccd1 vccd1 _4768_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_2665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3719_ _3721_/A vssd1 vssd1 vccd1 vccd1 _3719_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4493__RESET_B fanout208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4699_ _3390_/Y _4699_/D _3672_/Y vssd1 vssd1 vccd1 vccd1 _4699_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_3924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_2105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout157/X fanout203/X vssd1 vssd1 vccd1 vccd1 _5082_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_22_4141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_2070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_3681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2946__A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_2980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_3233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3777__A _3777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4825__CLK _4920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
+ _4428_/Q _2099_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_31_3709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_3889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_3277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4975__CLK _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_2131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_4113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_4074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_2514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_2683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_2536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_2619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4355__CLK _4359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_2321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2050_ _4428_/Q _2046_/C _2047_/B vssd1 vssd1 vccd1 vccd1 _2051_/B sky130_fd_sc_hd__a21bo_1
XFILLER_19_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3687__A _3695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2952_ _4913_/Q _4912_/Q vssd1 vssd1 vccd1 vccd1 _2952_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_30_3219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1903_ _4321_/Q _1903_/B vssd1 vssd1 vccd1 vccd1 _4321_/D sky130_fd_sc_hd__xnor2_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2883_ _4881_/Q _4880_/Q vssd1 vssd1 vccd1 vccd1 _2883_/Y sky130_fd_sc_hd__xnor2_2
X_1834_ _1832_/X _1833_/Y _1823_/X vssd1 vssd1 vccd1 vccd1 _1835_/B sky130_fd_sc_hd__o21ai_1
X_4622_ _4626_/CLK _4622_/D fanout233/X vssd1 vssd1 vccd1 vccd1 _4622_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4553_ _3310_/Y _4553_/D _3710_/Y vssd1 vssd1 vccd1 vccd1 _4553_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_3104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1765_ _1765_/A _4248_/B _4248_/C _3144_/A vssd1 vssd1 vccd1 vccd1 _1765_/X sky130_fd_sc_hd__or4_1
X_3504_ _4249_/A _4250_/A vssd1 vssd1 vccd1 vccd1 _3504_/Y sky130_fd_sc_hd__xnor2_2
X_4484_ _4533_/CLK _4484_/D fanout206/X vssd1 vssd1 vccd1 vccd1 _4484_/Q sky130_fd_sc_hd__dfrtp_4
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
+ _4486_/Q _2198_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_1696_ _4924_/Q vssd1 vssd1 vccd1 vccd1 _4925_/D sky130_fd_sc_hd__inv_2
XFILLER_28_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3435_ _3445_/A vssd1 vssd1 vccd1 vccd1 _3435_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_2210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3143__A2 _3138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2351__B1 _2344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_2182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ _2315_/X _2316_/Y _1975_/X vssd1 vssd1 vccd1 vccd1 _2318_/B sky130_fd_sc_hd__o21a_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout190_A fanout193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2766__A _4838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3297_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3297_/Y sky130_fd_sc_hd__inv_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_2068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5036_ _5044_/A vssd1 vssd1 vccd1 vccd1 _5036_/X sky130_fd_sc_hd__clkbuf_1
X_2248_ _2248_/A vssd1 vssd1 vccd1 vccd1 _2248_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2485__B _4675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4848__CLK _3865_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2179_ _4492_/Q _2179_/B vssd1 vssd1 vccd1 vccd1 _4492_/D sky130_fd_sc_hd__xnor2_1
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3749_/A fanout188/X vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_35_2407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_4118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3597__A _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4998__CLK _5047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4674__RESET_B fanout247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_2153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_2197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3783__124 _3784__125/A vssd1 vssd1 vccd1 vccd1 _3783__124/Y sky130_fd_sc_hd__inv_2
XFILLER_28_3660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2590__B1 _2518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput45 _5042_/X vssd1 vssd1 vccd1 vccd1 cclk_Q[2] sky130_fd_sc_hd__buf_2
XFILLER_28_3693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput56 _5053_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_I[5] sky130_fd_sc_hd__buf_2
Xoutput67 _5064_/X vssd1 vssd1 vccd1 vccd1 cos_out[0] sky130_fd_sc_hd__buf_2
XFILLER_27_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput78 _5075_/X vssd1 vssd1 vccd1 vccd1 fb1_I[3] sky130_fd_sc_hd__buf_2
XFILLER_8_3787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_4021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput89 _5086_/X vssd1 vssd1 vccd1 vccd1 fb1_Q[6] sky130_fd_sc_hd__buf_2
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5052__A _5060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_4029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input16_A comp_high_Q[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_2685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout120/X fanout249/X vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_2_1951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_3328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_2627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5003__CLK _4247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3300__A _3925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_2974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4131__A _4131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_2806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output84_A _5081_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2581__B1 _2518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3220_ _3935_/A _3440_/B vssd1 vssd1 vccd1 vccd1 _3220_/Y sky130_fd_sc_hd__xnor2_1
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3151_ _3838_/A _3839_/A vssd1 vssd1 vccd1 vccd1 _3151_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_7_1862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2102_ _4458_/Q _4457_/Q vssd1 vssd1 vccd1 vccd1 _2102_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_3_2449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3082_ _4989_/Q _3058_/D _3075_/B vssd1 vssd1 vccd1 vccd1 _3083_/B sky130_fd_sc_hd__a21bo_1
XFILLER_23_2388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2033_ _4466_/D _4440_/Q _4438_/Q _4437_/Q vssd1 vssd1 vccd1 vccd1 _2034_/C sky130_fd_sc_hd__and4_1
XFILLER_35_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_3163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3210__A _3848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3984_ _4447_/Q vssd1 vssd1 vccd1 vccd1 _4448_/D sky130_fd_sc_hd__inv_2
XFILLER_17_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2935_ _4900_/Q _2935_/B vssd1 vssd1 vccd1 vccd1 _4900_/D sky130_fd_sc_hd__xnor2_1
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_A
+ _4859_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2866_ _4865_/Q _2866_/B vssd1 vssd1 vccd1 vccd1 _4865_/D sky130_fd_sc_hd__xnor2_1
Xclkbuf_1_0_1_w0.cclk_I clkbuf_1_0_1_w0.cclk_I/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_w0.cclk_I/A
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__3864__B _3913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4605_ _4852_/CLK _4605_/D _3336_/Y vssd1 vssd1 vccd1 vccd1 _4605_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1817_ _1839_/A vssd1 vssd1 vccd1 vccd1 _3112_/A sky130_fd_sc_hd__buf_12
X_2797_ _3605_/Y _3631_/Y vssd1 vssd1 vccd1 vccd1 _5045_/A sky130_fd_sc_hd__nor2_4
XFILLER_30_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4536_ _2809_/A1 _4536_/D _3293_/Y vssd1 vssd1 vccd1 vccd1 _4536_/Q sky130_fd_sc_hd__dfrtp_1
X_1748_ _5007_/Q vssd1 vssd1 vccd1 vccd1 _5008_/D sky130_fd_sc_hd__inv_2
XANTENNA__4520__CLK _4532_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4467_ input18/X _4467_/D fanout197/X vssd1 vssd1 vccd1 vccd1 _4468_/D sky130_fd_sc_hd__dfrtp_1
X_1679_ _4909_/Q vssd1 vssd1 vccd1 vccd1 _4908_/D sky130_fd_sc_hd__inv_2
XFILLER_5_3916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4398_ _4402_/CLK _4398_/D fanout189/X vssd1 vssd1 vccd1 vccd1 _4398_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2324__B1 _2173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_TE_B
+ _2713_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input8_A comp_high_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4670__CLK _4718_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2496__A _4670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3349_ _3361_/A vssd1 vssd1 vccd1 vccd1 _3349_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_2062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5019_ input32/X _5019_/D fanout214/X vssd1 vssd1 vccd1 vccd1 _5020_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_27_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5026__CLK input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4855__RESET_B fanout228/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_2969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_3837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2381__D _2418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3203__11 _3201__9/A vssd1 vssd1 vccd1 vccd1 _4376_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5047__A _5047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_4022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2563__B1 _1975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_2918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_3218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_2883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout128/X fanout246/X vssd1 vssd1 vccd1 vccd1 _5077_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_2_3161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2556__D _2579_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2853__B _2853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4126__A _4126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_4037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3030__A _3030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_3347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_3358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2720_ _4803_/Q _4802_/Q _4801_/Q _2720_/D vssd1 vssd1 vccd1 vccd1 _2730_/C sky130_fd_sc_hd__and4_1
XFILLER_9_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2651_ _4834_/D _4776_/Q _4774_/Q _4773_/Q vssd1 vssd1 vccd1 vccd1 _2690_/A sky130_fd_sc_hd__or4_1
XFILLER_9_4049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2582_ _4710_/Q _2582_/B vssd1 vssd1 vccd1 vccd1 _4710_/D sky130_fd_sc_hd__xnor2_1
X_4321_ _4324_/CLK _4321_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _4321_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout109 _5046_/A vssd1 vssd1 vccd1 vccd1 _4901_/CLK sky130_fd_sc_hd__buf_2
X_4252_ _4126_/A _4248_/C _4251_/Y vssd1 vssd1 vccd1 vccd1 _4252_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_3061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4183_ _4738_/Q vssd1 vssd1 vccd1 vccd1 _4739_/D sky130_fd_sc_hd__inv_2
XFILLER_23_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3205__A _3600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3134_ _3134_/A vssd1 vssd1 vccd1 vccd1 _3134_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3065_ _4985_/Q _3069_/B _3071_/A vssd1 vssd1 vccd1 vccd1 _3112_/C sky130_fd_sc_hd__o21ai_1
XFILLER_3_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2016_ _4462_/D _4404_/Q vssd1 vssd1 vccd1 vccd1 _2017_/B sky130_fd_sc_hd__xnor2_1
X_3773__112 _3776__115/A vssd1 vssd1 vccd1 vccd1 _3773__112/Y sky130_fd_sc_hd__inv_2
XFILLER_23_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3681__88 _3683__90/A vssd1 vssd1 vccd1 vccd1 _3681__88/Y sky130_fd_sc_hd__inv_2
XANTENNA__4266__RESET_B _5056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout153_A _3930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_2991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3967_ _4416_/Q vssd1 vssd1 vccd1 vccd1 _4415_/D sky130_fd_sc_hd__inv_2
XANTENNA__3875__A _3899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_2281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2918_ _4898_/Q _2918_/B vssd1 vssd1 vccd1 vccd1 _2919_/B sky130_fd_sc_hd__nor2_1
X_3898_ _3909_/A _3898_/B vssd1 vssd1 vccd1 vccd1 _3900_/A sky130_fd_sc_hd__nand2_4
XFILLER_30_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2849_ _2819_/D _2848_/X _2687_/X vssd1 vssd1 vccd1 vccd1 _2850_/B sky130_fd_sc_hd__o21ai_1
XFILLER_30_2178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4519_ _4532_/CLK _4519_/D fanout211/X vssd1 vssd1 vccd1 vccd1 _4519_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_3641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2938__B _4905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_2490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_4117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_3245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_2325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4909__CLK _3504_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_2210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4870_ _1700_/Y _4870_/D _3481_/Y vssd1 vssd1 vccd1 vccd1 _4870_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_3854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_2265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_3865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3821_ _4335_/Q vssd1 vssd1 vccd1 vccd1 _4334_/D sky130_fd_sc_hd__inv_2
XFILLER_18_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3695__A _3695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3752_ _3948_/A vssd1 vssd1 vccd1 vccd1 _3752_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2703_ _4834_/D _4761_/Q vssd1 vssd1 vccd1 vccd1 _2704_/D sky130_fd_sc_hd__xnor2_1
XFILLER_31_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2634_ _4063_/C _2631_/X _2632_/X _2802_/A _3875_/D vssd1 vssd1 vccd1 vccd1 _2635_/B
+ sky130_fd_sc_hd__o32a_2
XFILLER_31_1786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2565_ _4707_/Q _2561_/C _2562_/B vssd1 vssd1 vccd1 vccd1 _2566_/B sky130_fd_sc_hd__a21bo_1
XFILLER_29_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4304_ _2294_/B1 _4304_/D _3160__60/Y vssd1 vssd1 vccd1 vccd1 _4304_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_2372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2496_ _4670_/Q _2496_/B vssd1 vssd1 vccd1 vccd1 _4670_/D sky130_fd_sc_hd__xnor2_1
XFILLER_22_3825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4439__CLK _5033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4235_ _4823_/Q vssd1 vssd1 vccd1 vccd1 _4824_/D sky130_fd_sc_hd__inv_2
XFILLER_25_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4166_ _4723_/Q vssd1 vssd1 vccd1 vccd1 _4722_/D sky130_fd_sc_hd__inv_2
XANTENNA_w0.ro_block_Q.ro_pol_eve.tribuf.t_buf_TE_B _1771_/Y vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3117_ _5004_/Q _5003_/Q vssd1 vssd1 vccd1 vccd1 _3117_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__2774__A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4097_ _4607_/Q vssd1 vssd1 vccd1 vccd1 _4608_/D sky130_fd_sc_hd__inv_2
XANTENNA__4589__CLK _5043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3048_ _4970_/Q _4969_/Q vssd1 vssd1 vccd1 vccd1 _3048_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__4439__SET_B fanout195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_2029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2586__B1_N _2579_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4999_ _3552_/X _4999_/D _3586_/Y vssd1 vssd1 vccd1 vccd1 _4999_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_2516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_4014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_4108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_3429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_2781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5060__A _5060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3499__B _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3774__113_A _3776__115/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_2173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2509__B1 _2344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1763__A _5029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2350_ _4585_/Q _2350_/B vssd1 vssd1 vccd1 vccd1 _4585_/D sky130_fd_sc_hd__xnor2_1
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2281_ _2281_/A vssd1 vssd1 vccd1 vccd1 _2283_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4020_ _4498_/Q vssd1 vssd1 vccd1 vccd1 _4499_/D sky130_fd_sc_hd__inv_2
XANTENNA__4731__CLK _3407_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2594__A _2680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4922_ _4981_/CLK _4922_/D _3517_/Y vssd1 vssd1 vccd1 vccd1 _4922_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_3217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4853_ _3479_/Y _4853_/D _3627__79/Y vssd1 vssd1 vccd1 vccd1 _4853_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3804_ _4300_/Q vssd1 vssd1 vccd1 vccd1 _4301_/D sky130_fd_sc_hd__inv_2
XFILLER_20_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4784_ _3434_/Y _4784_/D _3649_/Y vssd1 vssd1 vccd1 vccd1 _4784_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1996_ _4398_/Q _4397_/Q _1962_/D _1993_/B vssd1 vssd1 vccd1 vccd1 _1997_/B sky130_fd_sc_hd__a31o_1
XFILLER_14_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_2295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout116_A _4811_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3666_ _3669_/A vssd1 vssd1 vccd1 vccd1 _3666_/Y sky130_fd_sc_hd__inv_2
X_2617_ _4737_/Q _4736_/Q vssd1 vssd1 vccd1 vccd1 _2617_/Y sky130_fd_sc_hd__xnor2_4
X_3597_ _3597_/A vssd1 vssd1 vccd1 vccd1 _3597_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2548_ _4745_/D _4719_/Q _4717_/Q _4716_/Q vssd1 vssd1 vccd1 vccd1 _2549_/C sky130_fd_sc_hd__and4_1
XFILLER_6_3841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2920__B1 _2858_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_GATE_N
+ _5063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2479_ _4677_/Q _4676_/Q _4675_/Q _2479_/D vssd1 vssd1 vccd1 vccd1 _2480_/D sky130_fd_sc_hd__and4_2
XFILLER_2_3749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4218_ _4792_/Q vssd1 vssd1 vccd1 vccd1 _4791_/D sky130_fd_sc_hd__inv_2
XFILLER_5_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4281__RESET_B fanout201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4149_ _4688_/Q vssd1 vssd1 vccd1 vccd1 _4689_/D sky130_fd_sc_hd__inv_2
XFILLER_0_3473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3260__20 _3264__22/A vssd1 vssd1 vccd1 vccd1 _3260__20/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2739__B1 _2687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_3809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_2379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout144/X fanout215/X vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__dlrtn_1
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
+ _4798_/Q _2784_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_3577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_4074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3303__A _3309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_3548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__1642_ clkbuf_0__1642_/X vssd1 vssd1 vccd1 vccd1 _3365__31/A sky130_fd_sc_hd__clkbuf_16
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1850_ _4301_/Q _4300_/Q vssd1 vssd1 vccd1 vccd1 _1850_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_19_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_3868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4284__CLK _4288_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_2571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1781_ _4277_/Q _4276_/Q _1789_/C _1793_/A vssd1 vssd1 vccd1 vccd1 _1841_/B sky130_fd_sc_hd__a31o_1
XFILLER_30_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3520_ _3916_/A _3915_/A vssd1 vssd1 vccd1 vccd1 _3520_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_10_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3451_ _4189_/A _4190_/A vssd1 vssd1 vccd1 vccd1 _3451_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_26_3021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2402_ _2412_/A _2402_/B vssd1 vssd1 vccd1 vccd1 _2403_/B sky130_fd_sc_hd__nand2_1
X_3382_ _4004_/A _3491_/B vssd1 vssd1 vccd1 vccd1 _3382_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_1917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_2342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2333_ _4583_/Q _2333_/B vssd1 vssd1 vccd1 vccd1 _2334_/B sky130_fd_sc_hd__nor2_1
XFILLER_26_2375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_3986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5052_ _5060_/A vssd1 vssd1 vccd1 vccd1 _5052_/X sky130_fd_sc_hd__clkbuf_1
X_2264_ _2608_/A _4533_/Q vssd1 vssd1 vccd1 vccd1 _4533_/D sky130_fd_sc_hd__xor2_1
XFILLER_22_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4003_ _4131_/A _4131_/B _4003_/C _4131_/C vssd1 vssd1 vccd1 vccd1 _4005_/B sky130_fd_sc_hd__or4_2
XFILLER_22_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2195_ _4501_/Q _4500_/Q vssd1 vssd1 vccd1 vccd1 _2195_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_4_2193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
+ _4856_/Q _2884_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_20_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4905_ _4905_/CLK _4905_/D fanout231/X vssd1 vssd1 vccd1 vccd1 _4905_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_17_3779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4627__CLK _4248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf _4317_/Q _1916_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_33_3069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_3470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout233_A fanout234/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4836_ input30/X _4836_/D fanout238/X vssd1 vssd1 vccd1 vccd1 _4836_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2490__C _2490_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4767_ _4809_/CLK _4767_/D fanout252/X vssd1 vssd1 vccd1 vccd1 _4767_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__3883__A _3883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1979_ _4392_/Q _1973_/C _1974_/B vssd1 vssd1 vccd1 vccd1 _1980_/B sky130_fd_sc_hd__a21bo_1
XFILLER_11_2644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4777__CLK _4247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3718_ _3721_/A vssd1 vssd1 vccd1 vccd1 _3718_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_2677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4698_ _2807_/A _4698_/D _3389_/Y vssd1 vssd1 vccd1 vccd1 _4698_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_14_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3649_ _4195_/A vssd1 vssd1 vccd1 vccd1 _3649_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4809__RESET_B fanout255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3146__B1 _2468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4462__RESET_B fanout199/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3312__24 _3366__32/A vssd1 vssd1 vccd1 vccd1 _4564_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_3557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2962__A _2962_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_3289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout158/X fanout205/X vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_29_3606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_3628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_2154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_4031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_3639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_4064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_4086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3137__B1 _4248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_3205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_3001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_3067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4129__A _4129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2872__A _2916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_3345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2951_ _4911_/Q _4910_/Q vssd1 vssd1 vccd1 vccd1 _2951_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_17_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_3209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1902_ _1856_/C _1898_/Y _1823_/X vssd1 vssd1 vccd1 vccd1 _1903_/B sky130_fd_sc_hd__o21ai_1
XFILLER_31_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2882_ _4879_/Q _4878_/Q vssd1 vssd1 vccd1 vccd1 _2882_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_30_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_3080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4621_ _4626_/CLK _4621_/D fanout233/X vssd1 vssd1 vccd1 vccd1 _4621_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1833_ _4347_/D _4289_/Q _4287_/Q vssd1 vssd1 vccd1 vccd1 _1833_/Y sky130_fd_sc_hd__nor3_1
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_TE_B
+ _2780_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_4090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4552_ _2294_/B1 _4552_/D _3309_/Y vssd1 vssd1 vccd1 vccd1 _4552_/Q sky130_fd_sc_hd__dfrtp_1
X_1764_ _5031_/Q _5030_/Q vssd1 vssd1 vccd1 vccd1 _3144_/A sky130_fd_sc_hd__xnor2_4
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_A
+ _4524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3503_ _3519_/A vssd1 vssd1 vccd1 vccd1 _3503_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1935__B _3737_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4902__RESET_B fanout231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4483_ _5042_/A _4483_/D fanout202/X vssd1 vssd1 vccd1 vccd1 _4483_/Q sky130_fd_sc_hd__dfrtp_1
X_1695_ _4925_/Q vssd1 vssd1 vccd1 vccd1 _4924_/D sky130_fd_sc_hd__inv_2
XANTENNA__3208__A _3848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3434_ _4065_/A _3543_/B vssd1 vssd1 vccd1 vccd1 _3434_/Y sky130_fd_sc_hd__xnor2_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1951__A _3882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2316_ _4577_/Q _2316_/B vssd1 vssd1 vccd1 vccd1 _2316_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_3844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _3947_/A _3438_/B vssd1 vssd1 vccd1 vccd1 _3296_/Y sky130_fd_sc_hd__xnor2_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5035_ _5043_/A vssd1 vssd1 vccd1 vccd1 _5035_/X sky130_fd_sc_hd__clkbuf_1
X_2247_ _4527_/Q _2247_/B vssd1 vssd1 vccd1 vccd1 _4527_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2485__C _4674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2178_ _2178_/A _2178_/B vssd1 vssd1 vccd1 vccd1 _2179_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_3109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_2121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_GATE_N
+ _3375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4819_ _1765_/A _4819_/D _3454_/Y vssd1 vssd1 vccd1 vccd1 _4819_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2022__A _2608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput35 _5032_/X vssd1 vssd1 vccd1 vccd1 cclk_I[0] sky130_fd_sc_hd__clkbuf_1
XFILLER_7_2008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput46 _5043_/X vssd1 vssd1 vccd1 vccd1 cclk_Q[3] sky130_fd_sc_hd__buf_2
XFILLER_27_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput57 _5054_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_I[6] sky130_fd_sc_hd__buf_2
XFILLER_2_4000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput68 _5065_/X vssd1 vssd1 vccd1 vccd1 cos_out[1] sky130_fd_sc_hd__buf_2
Xoutput79 _5076_/X vssd1 vssd1 vccd1 vccd1 fb1_I[4] sky130_fd_sc_hd__buf_2
XFILLER_24_3569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1861__A _4351_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_2918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3203__11_A _3201__9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3300__B _3442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_3529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_3930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_2839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_3414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
+ _4617_/Q _2437_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__4131__B _4131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_2713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_2818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4322__CLK _4324_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout119/X fanout248/X vssd1 vssd1 vccd1 vccd1 _5078_/A sky130_fd_sc_hd__dlrtn_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2867__A _4927_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_3118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3150_ _3838_/A _3839_/A vssd1 vssd1 vccd1 vccd1 _3150_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_23_2334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_2597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4472__CLK _4472_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2101_ _4456_/Q _4455_/Q vssd1 vssd1 vccd1 vccd1 _2101_/Y sky130_fd_sc_hd__xnor2_4
X_3081_ _4987_/Q _3081_/B vssd1 vssd1 vccd1 vccd1 _4987_/D sky130_fd_sc_hd__xnor2_1
X_2032_ _4424_/Q _4423_/Q vssd1 vssd1 vccd1 vccd1 _2032_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_1_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3698__A _4071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2621__A_N _4742_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_3705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3364__30_A _3366__32/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3983_ _4448_/Q vssd1 vssd1 vccd1 vccd1 _4447_/D sky130_fd_sc_hd__inv_2
XFILLER_16_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_2430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3210__B _3847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2934_ _3030_/A _2934_/B vssd1 vssd1 vccd1 vccd1 _2935_/B sky130_fd_sc_hd__nand2_1
XFILLER_15_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2865_ _2817_/C _2861_/Y _2858_/X vssd1 vssd1 vccd1 vccd1 _2866_/B sky130_fd_sc_hd__o21ai_1
XFILLER_34_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4604_ _3335_/Y _4604_/D _3699_/Y vssd1 vssd1 vccd1 vccd1 _4604_/Q sky130_fd_sc_hd__dfrtp_1
X_1816_ _4281_/Q _1816_/B vssd1 vssd1 vccd1 vccd1 _4281_/D sky130_fd_sc_hd__xnor2_1
X_2796_ _2796_/A vssd1 vssd1 vccd1 vccd1 _2796_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_2783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4535_ _3292_/Y _4535_/D _3720_/Y vssd1 vssd1 vccd1 vccd1 _4535_/Q sky130_fd_sc_hd__dfrtp_1
X_1747_ _5008_/Q vssd1 vssd1 vccd1 vccd1 _5007_/D sky130_fd_sc_hd__inv_2
XFILLER_11_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_3801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_2306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4466_ input18/X _4466_/D fanout198/X vssd1 vssd1 vccd1 vccd1 _4467_/D sky130_fd_sc_hd__dfrtp_1
X_1678_ _4906_/Q vssd1 vssd1 vccd1 vccd1 _4907_/D sky130_fd_sc_hd__inv_2
XFILLER_28_2256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4815__CLK _4187_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4397_ _4402_/CLK _4397_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _4397_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_3878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3348_ _4004_/A _3491_/B vssd1 vssd1 vccd1 vccd1 _3348_/Y sky130_fd_sc_hd__xnor2_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
+ _4675_/Q _2539_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_3279_ _3287_/A vssd1 vssd1 vccd1 vccd1 _3279_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4965__CLK _1700_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5018_ _3572_/Y _5018_/D _3576_/Y vssd1 vssd1 vccd1 vccd1 _5018_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_6_1395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_4030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_3638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3401__A _4065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_3395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2017__A _2061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4895__RESET_B fanout234/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_2282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_4045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_4117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_3480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4495__CLK _4533_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2687__A _2858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5063__A _5063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_2704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_3399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_2748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_4141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3311__A _4469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_2414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4126__B _4248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_2447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2794__A_N _4839_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_4049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4565__RESET_B fanout212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_2035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2650_ _4764_/Q _4763_/Q _2658_/C _2661_/A vssd1 vssd1 vccd1 vccd1 _2704_/B sky130_fd_sc_hd__a31o_1
XFILLER_12_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_4028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4838__CLK input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2581_ _2551_/D _2580_/X _2518_/X vssd1 vssd1 vccd1 vccd1 _2582_/B sky130_fd_sc_hd__o21ai_1
XFILLER_9_3327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4320_ _4324_/CLK _4320_/D fanout189/X vssd1 vssd1 vccd1 vccd1 _4320_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_2626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_2407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4251_ _4845_/Q _4844_/Q vssd1 vssd1 vccd1 vccd1 _4251_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_25_2429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4988__CLK _4997_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4182_ _4739_/Q vssd1 vssd1 vccd1 vccd1 _4738_/D sky130_fd_sc_hd__inv_2
XFILLER_23_2153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3133_ _3133_/A _3133_/B vssd1 vssd1 vccd1 vccd1 _3134_/A sky130_fd_sc_hd__or2_1
XFILLER_7_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3064_ _4988_/Q _4987_/Q _4986_/Q _3075_/B vssd1 vssd1 vccd1 vccd1 _3069_/B sky130_fd_sc_hd__or4_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2015_ _4401_/Q _2015_/B vssd1 vssd1 vccd1 vccd1 _4401_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__3221__A _3233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
+ _4390_/Q _2030_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_17_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3966_ _4413_/Q vssd1 vssd1 vccd1 vccd1 _4414_/D sky130_fd_sc_hd__inv_2
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2917_ _4895_/Q _2917_/B vssd1 vssd1 vccd1 vccd1 _4895_/D sky130_fd_sc_hd__xnor2_1
XFILLER_17_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3897_ _3897_/A vssd1 vssd1 vccd1 vccd1 _3898_/B sky130_fd_sc_hd__buf_4
XFILLER_17_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2848_ _4861_/Q _2848_/B vssd1 vssd1 vccd1 vccd1 _2848_/X sky130_fd_sc_hd__and2b_1
XFILLER_30_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2779_ _4818_/Q _4817_/Q vssd1 vssd1 vccd1 vccd1 _2779_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__3891__A _3891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4518_ _4532_/CLK _4518_/D fanout219/X vssd1 vssd1 vccd1 vccd1 _4518_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_2_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_2042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_2053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4449_ _3931_/A _4449_/D _3245_/Y vssd1 vssd1 vccd1 vccd1 _4449_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_2147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_3697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_2963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_2849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3657__86 _3683__90/A vssd1 vssd1 vccd1 vccd1 _3657__86/Y sky130_fd_sc_hd__inv_2
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_2035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2970__A _3929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_2333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5058__A _5058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_4129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_3428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_GATE_N _5048_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3306__A _3903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_2589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4137__A _4660_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3041__A _5020_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4510__CLK _2286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1814__A3 _1778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3820_ _4332_/Q vssd1 vssd1 vccd1 vccd1 _4333_/D sky130_fd_sc_hd__inv_2
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3751_ _3948_/A vssd1 vssd1 vccd1 vccd1 _3751_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4660__CLK _2470_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_2444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2702_ _4774_/Q _2702_/B vssd1 vssd1 vccd1 vccd1 _4774_/D sky130_fd_sc_hd__xnor2_1
XFILLER_13_3590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2633_ _3941_/B _4003_/C _4131_/C _2456_/Y _3929_/A vssd1 vssd1 vccd1 vccd1 _2802_/A
+ sky130_fd_sc_hd__a221o_1
X_2564_ _2564_/A _2564_/B vssd1 vssd1 vccd1 vccd1 _4705_/D sky130_fd_sc_hd__xnor2_1
X_4303_ _3910_/A _4303_/D _3778__119/Y vssd1 vssd1 vccd1 vccd1 _4303_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_2215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2495_ _2566_/A _2495_/B vssd1 vssd1 vccd1 vccd1 _2496_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_3973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3216__A _3233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4234_ _4824_/Q vssd1 vssd1 vccd1 vccd1 _4823_/D sky130_fd_sc_hd__inv_2
XFILLER_22_3837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4165_ _4720_/Q vssd1 vssd1 vccd1 vccd1 _4721_/D sky130_fd_sc_hd__inv_2
XFILLER_25_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3116_ _5002_/Q _5001_/Q vssd1 vssd1 vccd1 vccd1 _3116_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_7_1490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4096_ _4608_/Q vssd1 vssd1 vccd1 vccd1 _4607_/D sky130_fd_sc_hd__inv_2
XFILLER_3_2088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3047_ _4968_/Q _4967_/Q vssd1 vssd1 vccd1 vccd1 _3047_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4487__RESET_B fanout201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3886__A _3886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2790__A _2790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4998_ _5047_/A _4998_/D fanout242/X vssd1 vssd1 vccd1 vccd1 _4998_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_3977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_3365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3949_ _4382_/Q vssd1 vssd1 vccd1 vccd1 _4381_/D sky130_fd_sc_hd__inv_2
XFILLER_14_1930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_3737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_3577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_3358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_2865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4533__CLK _4533_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_2668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4683__CLK _4717_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_2753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2205__A _4559_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_2797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout136/X fanout239/X vssd1 vssd1 vccd1 vccd1 _5084_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2509__A1 _2480_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1763__B _1763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2280_ _4561_/Q _4560_/D vssd1 vssd1 vccd1 vccd1 _2281_/A sky130_fd_sc_hd__and2b_1
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2875__A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4998__RESET_B fanout242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_2375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4927__RESET_B fanout214/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_2189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4921_ _3516_/Y _4921_/D _3608_/Y vssd1 vssd1 vccd1 vccd1 _4921_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_3229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4852_ _4852_/CLK _4852_/D _3478__47/Y vssd1 vssd1 vccd1 vccd1 _4852_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_3641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3803_ _4301_/Q vssd1 vssd1 vccd1 vccd1 _4300_/D sky130_fd_sc_hd__inv_2
XFILLER_18_2096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4783_ _1765_/A _4783_/D _3433_/Y vssd1 vssd1 vccd1 vccd1 _4783_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_18_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1995_ _4395_/Q _1995_/B vssd1 vssd1 vccd1 vccd1 _4395_/D sky130_fd_sc_hd__xnor2_1
XFILLER_33_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4406__CLK _4064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3665_ _3669_/A vssd1 vssd1 vccd1 vccd1 _3665_/Y sky130_fd_sc_hd__inv_2
X_2616_ _4735_/Q _4734_/Q vssd1 vssd1 vccd1 vccd1 _2616_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_31_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout109_A _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3596_ _3597_/A vssd1 vssd1 vccd1 vccd1 _3596_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_2220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2547_ _4703_/Q _4702_/Q vssd1 vssd1 vccd1 vccd1 _2547_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_6_3831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4556__CLK input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2478_ _4679_/Q _4678_/Q _2478_/C vssd1 vssd1 vccd1 vccd1 _2479_/D sky130_fd_sc_hd__and3_1
XFILLER_2_3717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_2297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_2067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4217_ _4789_/Q vssd1 vssd1 vccd1 vccd1 _4790_/D sky130_fd_sc_hd__inv_2
XFILLER_5_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4148_ _4689_/Q vssd1 vssd1 vccd1 vccd1 _4688_/D sky130_fd_sc_hd__inv_2
XFILLER_20_3380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4668__RESET_B fanout242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_4106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_4117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4079_ _4573_/Q vssd1 vssd1 vccd1 vccd1 _4574_/D sky130_fd_sc_hd__inv_2
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3158__58 _3159__59/A vssd1 vssd1 vccd1 vccd1 _3158__58/Y sky130_fd_sc_hd__inv_2
XFILLER_30_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_4020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_4086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5071__A _5071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_3249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_2515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3684_/A fanout216/X vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__dlrtn_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4429__CLK _4429_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1780_ _4275_/Q vssd1 vssd1 vccd1 vccd1 _1793_/A sky130_fd_sc_hd__inv_2
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_2583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1938__C1 _1952_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1774__A _1839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4579__CLK _4590_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3450_ _3466_/A vssd1 vssd1 vccd1 vccd1 _3450_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_2619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2401_ _4617_/Q _2377_/D _2394_/B vssd1 vssd1 vccd1 vccd1 _2402_/B sky130_fd_sc_hd__a21bo_1
XFILLER_26_3044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3381_ _3393_/A vssd1 vssd1 vccd1 vccd1 _3381_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_2404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_2415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2332_ _4580_/Q _2332_/B vssd1 vssd1 vccd1 vccd1 _4580_/D sky130_fd_sc_hd__xnor2_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_2218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5051_ _5059_/A vssd1 vssd1 vccd1 vccd1 _5051_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2263_ _4532_/Q _2263_/B vssd1 vssd1 vccd1 vccd1 _4532_/D sky130_fd_sc_hd__xor2_1
X_4002_ _4123_/A vssd1 vssd1 vccd1 vccd1 _4003_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_6_1769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2194_ _4499_/Q _4498_/Q vssd1 vssd1 vccd1 vccd1 _2194_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_4_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4904_ _5046_/A _4904_/D fanout236/X vssd1 vssd1 vccd1 vccd1 _4904_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_21_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4835_ input30/X _4835_/D fanout238/X vssd1 vssd1 vccd1 vccd1 _4836_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_15_2781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4766_ _4809_/CLK _4766_/D fanout255/X vssd1 vssd1 vccd1 vccd1 _4766_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout226_A fanout230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1978_ _3112_/A vssd1 vssd1 vccd1 vccd1 _2061_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3883__B _3883_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3717_ _3721_/A vssd1 vssd1 vccd1 vccd1 _3717_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4697_ _3388_/Y _4697_/D _3673_/Y vssd1 vssd1 vccd1 vccd1 _4697_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4060__A _4126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3648_ _4195_/A vssd1 vssd1 vccd1 vccd1 _3648_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_3854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3146__A1 _4064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3579_ _3587_/A vssd1 vssd1 vccd1 vccd1 _3579_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_3661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_3475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3404__A _3414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_2741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_3486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_2785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_3582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_2881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_2917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_4098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4871__CLK _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
+ _4987_/Q _3119_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_21_2251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_2345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_4003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_2295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_2309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[4\].w1.ro_block_I.ro_pol.tribuf.t_buf _2796_/X _2643_/Y vssd1
+ vssd1 vccd1 vccd1 _5088_/A sky130_fd_sc_hd__ebufn_8
XFILLER_16_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2950_ _4909_/Q _4908_/Q vssd1 vssd1 vccd1 vccd1 _2950_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_34_3357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_2000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1901_ _4320_/Q _1901_/B vssd1 vssd1 vccd1 vccd1 _4320_/D sky130_fd_sc_hd__xnor2_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2881_ _4877_/Q _4876_/Q vssd1 vssd1 vccd1 vccd1 _2881_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_31_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_2055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4620_ _4623_/CLK _4620_/D fanout234/X vssd1 vssd1 vccd1 vccd1 _4620_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_30_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1832_ _4347_/D _4289_/Q _4287_/Q vssd1 vssd1 vccd1 vccd1 _1832_/X sky130_fd_sc_hd__and3_1
XFILLER_12_3666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4551_ _3308_/Y _4551_/D _3712_/Y vssd1 vssd1 vccd1 vccd1 _4551_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_2965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1763_ _5029_/Q _1763_/B vssd1 vssd1 vccd1 vccd1 _5029_/D sky130_fd_sc_hd__xnor2_1
XFILLER_11_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_2987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3502_ _3556_/A _3556_/B vssd1 vssd1 vccd1 vccd1 _3502_/Y sky130_fd_sc_hd__xnor2_2
X_4482_ _4533_/CLK _4482_/D fanout208/X vssd1 vssd1 vccd1 vccd1 _4482_/Q sky130_fd_sc_hd__dfrtp_2
X_1694_ _4922_/Q vssd1 vssd1 vccd1 vccd1 _4923_/D sky130_fd_sc_hd__inv_2
XANTENNA__3208__B _3847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3433_ _3445_/A vssd1 vssd1 vccd1 vccd1 _3433_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_2449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2315_ _4578_/Q _4577_/Q _2315_/C vssd1 vssd1 vccd1 vccd1 _2315_/X sky130_fd_sc_hd__and3_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3295_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_2037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3224__A _3917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5034_/A vssd1 vssd1 vccd1 vccd1 _5034_/X sky130_fd_sc_hd__clkbuf_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ _2207_/D _2245_/Y _2173_/X vssd1 vssd1 vccd1 vccd1 _2247_/B sky130_fd_sc_hd__o21ai_1
XFILLER_22_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5055_/A fanout244/X vssd1 vssd1 vccd1 vccd1 _5079_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__2485__D _2507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_3809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2177_ _2176_/Y _2133_/C _4493_/Q vssd1 vssd1 vccd1 vccd1 _2178_/B sky130_fd_sc_hd__mux2_1
XANTENNA_fanout176_A _4060_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3878__B _4131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4744__CLK input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_3891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_3121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4818_ _3453_/Y _4818_/D _3639_/Y vssd1 vssd1 vccd1 vccd1 _4818_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_2177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_2420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_TE_B _1922_/Y vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4894__CLK _4901_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4749_ _5030_/CLK _4749_/D fanout224/X vssd1 vssd1 vccd1 vccd1 _4749_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_2475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput36 _5033_/X vssd1 vssd1 vccd1 vccd1 cclk_I[1] sky130_fd_sc_hd__buf_2
Xoutput47 _5044_/X vssd1 vssd1 vccd1 vccd1 cclk_Q[4] sky130_fd_sc_hd__buf_2
Xoutput58 _5055_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_I[7] sky130_fd_sc_hd__buf_2
Xoutput69 _5066_/X vssd1 vssd1 vccd1 vccd1 cos_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4683__RESET_B fanout255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4612__RESET_B fanout234/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_2869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4274__CLK _4281_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_4009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_3611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_3065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3309__A _3309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2213__A _4526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_2725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2869__B1 _2858_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4617__CLK _4626_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3044__A _3114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2100_ _4454_/Q _4453_/Q vssd1 vssd1 vccd1 vccd1 _2100_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_23_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3080_ _3109_/A _3080_/B vssd1 vssd1 vccd1 vccd1 _3081_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_3968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2031_ _4422_/Q _4421_/Q vssd1 vssd1 vccd1 vccd1 _2031_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_23_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_2153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_2197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3982_ _4445_/Q vssd1 vssd1 vccd1 vccd1 _4446_/D sky130_fd_sc_hd__inv_2
XFILLER_14_3717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_3897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_3165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2933_ _2932_/Y _2889_/C _4901_/Q vssd1 vssd1 vccd1 vccd1 _2934_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2864_ _4864_/Q _2864_/B vssd1 vssd1 vccd1 vccd1 _4864_/D sky130_fd_sc_hd__xnor2_1
XFILLER_30_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_2497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4603_ _4943_/CLK _4603_/D _3334_/Y vssd1 vssd1 vccd1 vccd1 _4603_/Q sky130_fd_sc_hd__dfrtp_1
X_1815_ _3114_/A _1815_/B vssd1 vssd1 vccd1 vccd1 _1816_/B sky130_fd_sc_hd__nand2_1
X_2795_ _2795_/A _2795_/B vssd1 vssd1 vccd1 vccd1 _2796_/A sky130_fd_sc_hd__or2_1
XFILLER_12_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3219__A _3233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4534_ _4248_/A _4534_/D _3290_/Y vssd1 vssd1 vccd1 vccd1 _4534_/Q sky130_fd_sc_hd__dfrtp_1
X_1746_ _5005_/Q vssd1 vssd1 vccd1 vccd1 _5006_/D sky130_fd_sc_hd__inv_2
XFILLER_29_3960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4465_ input18/X input2/X fanout197/X vssd1 vssd1 vccd1 vccd1 _4466_/D sky130_fd_sc_hd__dfrtp_4
X_1677_ _4907_/Q vssd1 vssd1 vccd1 vccd1 _4906_/D sky130_fd_sc_hd__inv_2
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
+ _4775_/Q _2716_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_8_2318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3416_ _5060_/A vssd1 vssd1 vccd1 vccd1 _3416_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_2329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4396_ _4402_/CLK _4396_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _4396_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__4297__CLK _3877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3347_ _3361_/A vssd1 vssd1 vccd1 vccd1 _3347_/Y sky130_fd_sc_hd__inv_2
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3278_ _3925_/A _3442_/B vssd1 vssd1 vccd1 vccd1 _3278_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_22_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3889__A _3889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5017_ _3922_/X _5017_/D _3571_/Y vssd1 vssd1 vccd1 vccd1 _5017_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_2891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2229_ _4524_/Q _4523_/Q _2208_/D _2226_/B vssd1 vssd1 vccd1 vccd1 _2230_/B sky130_fd_sc_hd__a31o_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3401__B _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_4086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_2651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3129__A _3129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2033__A _4466_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_2895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4864__RESET_B fanout228/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_4035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_4129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_2633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_2738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input21_A phi1b_dig_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout180/X fanout184/X vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_20_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2208__A _4524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_4017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_2459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf _4279_/Q _1848_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_31_2604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_2014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_2648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_2058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3039__A _3109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2580_ _4711_/Q _2580_/B vssd1 vssd1 vccd1 vccd1 _2580_/X sky130_fd_sc_hd__and2b_1
XFILLER_9_3317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_3339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_TE_B _1915_/Y vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1782__A _4347_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4250_ _4250_/A _4250_/B vssd1 vssd1 vccd1 vccd1 _4843_/D sky130_fd_sc_hd__xnor2_1
XFILLER_29_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4181_ _4736_/Q vssd1 vssd1 vccd1 vccd1 _4737_/D sky130_fd_sc_hd__inv_2
X_3132_ _5025_/D _5026_/Q vssd1 vssd1 vccd1 vccd1 _3133_/B sky130_fd_sc_hd__and2b_1
XFILLER_23_2165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3063_ _4991_/Q _4990_/Q _4989_/Q _3085_/B vssd1 vssd1 vccd1 vccd1 _3075_/B sky130_fd_sc_hd__or4_1
XFILLER_23_2198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3502__A _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2014_ _2012_/X _2013_/Y _2003_/X vssd1 vssd1 vccd1 vccd1 _2015_/B sky130_fd_sc_hd__o21ai_1
XFILLER_3_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_2971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3965_ _4414_/Q vssd1 vssd1 vccd1 vccd1 _4413_/D sky130_fd_sc_hd__inv_2
XFILLER_14_3569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3875__C _3901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2916_ _2916_/A _2916_/B vssd1 vssd1 vccd1 vccd1 _2917_/B sky130_fd_sc_hd__nand2_1
XANTENNA__2242__A1 _4527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3896_ _3896_/A vssd1 vssd1 vccd1 vccd1 _3903_/A sky130_fd_sc_hd__buf_12
XANTENNA_fanout139_A _2285_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_2125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2847_ _4862_/Q _2847_/B vssd1 vssd1 vccd1 vccd1 _2848_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2778_ _4816_/Q _4815_/Q vssd1 vssd1 vccd1 vccd1 _2778_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_30_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4517_ _3288_/Y _4517_/D _3721_/Y vssd1 vssd1 vccd1 vccd1 _4517_/Q sky130_fd_sc_hd__dfrtp_2
X_1729_ _4974_/Q vssd1 vssd1 vccd1 vccd1 _4973_/D sky130_fd_sc_hd__inv_2
XANTENNA__4275__RESET_B fanout199/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4932__CLK input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4448_ _3244_/Y _4448_/D _3744_/Y vssd1 vssd1 vccd1 vccd1 _4448_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_3665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_2098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4379_ _4472_/CLK _4379_/D fanout210/X vssd1 vssd1 vccd1 vccd1 _4379_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_3529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3412__A _3414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4312__CLK _5040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2970__B _4248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_2913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_4083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_3079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4462__CLK input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5074__A _5074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_3120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3306__B _3420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_2535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3322__A _3696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3041__B _4947_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
+ _4521_/Q _2270_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_11_3709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_3135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3750_ _3948_/A vssd1 vssd1 vccd1 vccd1 _3750_/Y sky130_fd_sc_hd__inv_2
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5048_/A fanout191/X vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2701_ _2771_/A _2701_/B vssd1 vssd1 vccd1 vccd1 _2702_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_2456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2632_ _3914_/B _2462_/Y _3898_/B vssd1 vssd1 vccd1 vccd1 _2632_/X sky130_fd_sc_hd__o21a_1
XFILLER_31_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2563_ _2561_/X _2562_/Y _1975_/X vssd1 vssd1 vccd1 vccd1 _2564_/B sky130_fd_sc_hd__o21a_1
XFILLER_9_2402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_3086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_2413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3643_/A fanout243/X vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__dlrtn_1
X_4302_ _3899_/A _4302_/D _3159__59/Y vssd1 vssd1 vccd1 vccd1 _4302_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_26_3941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_2363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_2446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2494_ _4671_/Q _2490_/C _2491_/B vssd1 vssd1 vccd1 vccd1 _2495_/B sky130_fd_sc_hd__a21bo_1
XFILLER_9_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_2457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_2385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4233_ _4821_/Q vssd1 vssd1 vccd1 vccd1 _4822_/D sky130_fd_sc_hd__inv_2
XFILLER_25_2238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4164_ _4721_/Q vssd1 vssd1 vccd1 vccd1 _4720_/D sky130_fd_sc_hd__inv_2
XFILLER_4_3781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3115_ _5000_/Q _4999_/Q vssd1 vssd1 vccd1 vccd1 _3115_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_23_1250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4095_ _4605_/Q vssd1 vssd1 vccd1 vccd1 _4606_/D sky130_fd_sc_hd__inv_2
XFILLER_0_2911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3232__A _3891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3046_ _4966_/Q _4965_/Q vssd1 vssd1 vccd1 vccd1 _3046_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_2977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2463__A1 _2631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout256_A fanout257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4485__CLK _5042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4997_ _4997_/CLK _4997_/D fanout232/X vssd1 vssd1 vccd1 vccd1 _4997_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4063__A _4131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3948_ _3948_/A vssd1 vssd1 vccd1 vccd1 _4354_/D sky130_fd_sc_hd__inv_2
XFILLER_14_2643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3879_ _3870_/Y _3925_/B _3878_/X vssd1 vssd1 vccd1 vccd1 _3881_/B sky130_fd_sc_hd__a21oi_1
XFILLER_30_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
+ _4579_/Q _2368_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__3407__A _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_4027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_3495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5069__A _5069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_3499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_2765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_2142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2205__B _4533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3681__88_A _3683__90/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2509__A2 _2508_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3317__A _3891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4358__CLK _4359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2891__A _4896_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4920_ _4920_/CLK _4920_/D _3515_/Y vssd1 vssd1 vccd1 vccd1 _4920_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_2020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4851_ _3477_/Y _4851_/D _3628__80/Y vssd1 vssd1 vccd1 vccd1 _4851_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_3631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_2518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_2075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3802_ _4298_/Q vssd1 vssd1 vccd1 vccd1 _4299_/D sky130_fd_sc_hd__inv_2
XFILLER_18_1352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4782_ _3432_/Y _4782_/D _3650_/Y vssd1 vssd1 vccd1 vccd1 _4782_/Q sky130_fd_sc_hd__dfrtp_4
X_1994_ _1963_/D _1993_/X _1823_/X vssd1 vssd1 vccd1 vccd1 _1995_/B sky130_fd_sc_hd__o21ai_1
XFILLER_15_3697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_2963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3733_ _3777_/A vssd1 vssd1 vccd1 vccd1 _3733_/X sky130_fd_sc_hd__buf_1
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_A
+ _4487_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3664_ _3669_/A vssd1 vssd1 vccd1 vccd1 _3664_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2615_ _4733_/Q _4732_/Q vssd1 vssd1 vccd1 vccd1 _2615_/Y sky130_fd_sc_hd__xnor2_4
X_3595_ _3597_/A vssd1 vssd1 vccd1 vccd1 _3595_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3227__A _3233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2546_ _4701_/Q _4700_/Q vssd1 vssd1 vccd1 vccd1 _2546_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_9_2232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_2276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2477_ _4741_/D _4683_/Q _4681_/Q _4680_/Q vssd1 vssd1 vccd1 vccd1 _2478_/C sky130_fd_sc_hd__and4_1
XFILLER_5_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_2912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_3898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4216_ _4790_/Q vssd1 vssd1 vccd1 vccd1 _4789_/D sky130_fd_sc_hd__inv_2
XFILLER_25_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_2923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_2945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4147_ _4686_/Q vssd1 vssd1 vccd1 vccd1 _4687_/D sky130_fd_sc_hd__inv_2
XFILLER_21_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3779__120 _3781__122/A vssd1 vssd1 vccd1 vccd1 _3779__120/Y sky130_fd_sc_hd__inv_2
XFILLER_25_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4078_ _4574_/Q vssd1 vssd1 vccd1 vccd1 _4573_/D sky130_fd_sc_hd__inv_2
XFILLER_23_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_4129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3897__A _3897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3029_ _3028_/Y _2986_/C _4958_/Q vssd1 vssd1 vccd1 vccd1 _3030_/B sky130_fd_sc_hd__mux2_1
X_3627__79 _3654__84/A vssd1 vssd1 vccd1 vccd1 _3627__79/Y sky130_fd_sc_hd__inv_2
XFILLER_16_3417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_2705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_GATE_N
+ fanout128/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_2304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_TE_B
+ _2024_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4500__CLK _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_2812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_4065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1880__A _1909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout250 fanout256/X vssd1 vssd1 vccd1 vccd1 fanout250/X sky130_fd_sc_hd__buf_2
XFILLER_1_3217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_2663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4650__CLK input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_2499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3600__A _3600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4378__RESET_B fanout219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2216__A _2996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_2237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1938__B1 _3845_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_2595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_2609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2400_ _4615_/Q _2400_/B vssd1 vssd1 vccd1 vccd1 _4615_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_3106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3380_ _4065_/A _3543_/B vssd1 vssd1 vccd1 vccd1 _3380_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_23_3911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2331_ _2412_/A _2331_/B vssd1 vssd1 vccd1 vccd1 _2332_/B sky130_fd_sc_hd__nand2_1
XFILLER_3_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_3089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5050_ _5058_/A vssd1 vssd1 vccd1 vccd1 _5050_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_3977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2262_ _3066_/A _2262_/B _2262_/C _2262_/D vssd1 vssd1 vccd1 vccd1 _2263_/B sky130_fd_sc_hd__and4_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4001_ _4001_/A vssd1 vssd1 vccd1 vccd1 _4004_/A sky130_fd_sc_hd__buf_12
XFILLER_23_3999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2193_ _2608_/A _4497_/Q vssd1 vssd1 vccd1 vccd1 _4497_/D sky130_fd_sc_hd__xor2_1
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3510__A _4065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4903_ _4905_/CLK _4903_/D fanout235/X vssd1 vssd1 vccd1 vccd1 _4903_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_4015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4834_ input30/X _4834_/D fanout237/X vssd1 vssd1 vccd1 vccd1 _4835_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_33_2337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4765_ _4811_/CLK _4765_/D fanout256/X vssd1 vssd1 vccd1 vccd1 _4765_/Q sky130_fd_sc_hd__dfrtp_2
X_1977_ _1977_/A _1977_/B vssd1 vssd1 vccd1 vccd1 _4390_/D sky130_fd_sc_hd__xnor2_1
XFILLER_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_2793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4523__CLK _4533_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3716_ _3721_/A vssd1 vssd1 vccd1 vccd1 _3716_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout219_A fanout220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4696_ _4981_/CLK _4696_/D _3387_/Y vssd1 vssd1 vccd1 vccd1 _4696_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3647_ _4195_/A vssd1 vssd1 vccd1 vccd1 _3647_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3146__A2 _4248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_3877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3578_ _3587_/A vssd1 vssd1 vccd1 vccd1 _3578_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4673__CLK _4718_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2529_ _2527_/X _2528_/Y _2518_/X vssd1 vssd1 vccd1 vccd1 _2530_/B sky130_fd_sc_hd__o21ai_1
XFILLER_9_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_2825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_2753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_2797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_3837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3420__A _3896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3082__A1 _4989_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4471__RESET_B fanout212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2036__A _4431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_2568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_2893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_2112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2345__B1 _2344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_3229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_2506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5082__A _5082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_2368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_4026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3330__A _3340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_4059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3472__44 _3528__52/A vssd1 vssd1 vccd1 vccd1 _3472__44/Y sky130_fd_sc_hd__inv_2
XFILLER_34_3369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1900_ _1909_/A _1900_/B vssd1 vssd1 vccd1 vccd1 _1901_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4546__CLK _4852_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2880_ _4875_/Q _4874_/Q vssd1 vssd1 vccd1 vccd1 _2880_/Y sky130_fd_sc_hd__xnor2_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1831_ _4285_/Q _1831_/B vssd1 vssd1 vccd1 vccd1 _4285_/D sky130_fd_sc_hd__xnor2_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1762_ _5028_/Q _1763_/B vssd1 vssd1 vccd1 vccd1 _5028_/D sky130_fd_sc_hd__xnor2_1
X_4550_ _2470_/A1 _4550_/D _3307_/Y vssd1 vssd1 vccd1 vccd1 _4550_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_1388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3501_ _3519_/A vssd1 vssd1 vccd1 vccd1 _3501_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4696__CLK _4981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1693_ _4923_/Q vssd1 vssd1 vccd1 vccd1 _4922_/D sky130_fd_sc_hd__inv_2
X_4481_ _3268_/Y _4481_/D _3732__95/Y vssd1 vssd1 vccd1 vccd1 _4481_/Q sky130_fd_sc_hd__dfrtp_1
X_3432_ _4127_/A _4129_/A vssd1 vssd1 vccd1 vccd1 _3432_/Y sky130_fd_sc_hd__xnor2_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ _3696_/A vssd1 vssd1 vccd1 vccd1 _3363_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_2202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_3960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3505__A _3519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2314_ _4575_/Q _2314_/B vssd1 vssd1 vccd1 vccd1 _4575_/D sky130_fd_sc_hd__xor2_1
XFILLER_6_1501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _4004_/A _3491_/B vssd1 vssd1 vccd1 vccd1 _3294_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_26_2174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3224__B _3444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2245_ _4529_/Q _4528_/Q _2248_/A vssd1 vssd1 vccd1 vccd1 _2245_/Y sky130_fd_sc_hd__nor3_1
X_5033_ _5033_/A vssd1 vssd1 vccd1 vccd1 _5033_/X sky130_fd_sc_hd__clkbuf_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2639__A1 _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2176_ _2176_/A vssd1 vssd1 vccd1 vccd1 _2176_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3240__A _3947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout169_A _3861_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4817_ _5007_/CLK _4817_/D _3452_/Y vssd1 vssd1 vccd1 vccd1 _4817_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_3133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_3756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4071__A _4071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4748_ _3416_/Y _4748_/D fanout233/X vssd1 vssd1 vccd1 vccd1 _4748_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4679_ _4719_/CLK _4679_/D fanout255/X vssd1 vssd1 vccd1 vccd1 _4679_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput37 _5034_/X vssd1 vssd1 vccd1 vccd1 cclk_I[2] sky130_fd_sc_hd__buf_2
XFILLER_11_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput48 _5045_/X vssd1 vssd1 vccd1 vccd1 cclk_Q[5] sky130_fd_sc_hd__buf_2
Xoutput59 _5056_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_Q[0] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3415__A _3903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_2826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4419__CLK _3899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_3389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_2583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4246__A _4249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4569__CLK _3855_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_3077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_2737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3325__A _4065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_2544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_2314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3044__B _4962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2030_ _4420_/Q _4419_/Q vssd1 vssd1 vccd1 vccd1 _2030_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_5_2290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_2121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_2165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_3133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3981_ _4446_/Q vssd1 vssd1 vccd1 vccd1 _4445_/D sky130_fd_sc_hd__inv_2
XFILLER_17_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_4121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2932_ _2932_/A vssd1 vssd1 vccd1 vccd1 _2932_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_3177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2863_ _2916_/A _2863_/B vssd1 vssd1 vccd1 vccd1 _2864_/B sky130_fd_sc_hd__nand2_1
XFILLER_15_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4602_ _3333_/Y _4602_/D _3700_/Y vssd1 vssd1 vccd1 vccd1 _4602_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2404__A _4619_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1814_ _4283_/Q _4282_/Q _1778_/D _1811_/B vssd1 vssd1 vccd1 vccd1 _1815_/B sky130_fd_sc_hd__a31o_1
XFILLER_12_2741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2794_ _4839_/D _4840_/Q vssd1 vssd1 vccd1 vccd1 _2795_/B sky130_fd_sc_hd__and2b_1
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4533_ _4533_/CLK _4533_/D fanout209/X vssd1 vssd1 vccd1 vccd1 _4533_/Q sky130_fd_sc_hd__dfrtp_4
X_1745_ _5006_/Q vssd1 vssd1 vccd1 vccd1 _5005_/D sky130_fd_sc_hd__inv_2
X_4464_ input26/X _4464_/D fanout198/X vssd1 vssd1 vccd1 vccd1 _4464_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1676_ _4888_/Q vssd1 vssd1 vccd1 vccd1 _4889_/D sky130_fd_sc_hd__inv_2
XFILLER_29_3983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1962__B _4397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3415_ _3903_/A _3420_/B vssd1 vssd1 vccd1 vccd1 _3415_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4395_ _4402_/CLK _4395_/D fanout185/X vssd1 vssd1 vccd1 vccd1 _4395_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_3869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3235__A _3738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3346_ _4065_/A _3543_/B vssd1 vssd1 vccd1 vccd1 _3346_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_3_3621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _3287_/A vssd1 vssd1 vccd1 vccd1 _3277_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5016_ _3570_/Y _5016_/D _3578_/Y vssd1 vssd1 vccd1 vccd1 _5016_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4711__CLK _4712_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2228_ _4521_/Q _2228_/B vssd1 vssd1 vccd1 vccd1 _4521_/D sky130_fd_sc_hd__xnor2_1
XFILLER_2_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2159_ _4488_/Q _2135_/D _2152_/B vssd1 vssd1 vccd1 vccd1 _2160_/B sky130_fd_sc_hd__a21bo_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_2229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4861__CLK _4865_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_3829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_2630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_2663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_2685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_2852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_4003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_4014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_2770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_2842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4833__RESET_B fanout237/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_2728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_3131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2984__A _4946_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4391__CLK _4429_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input14_A comp_high_Q[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3260__20_A _3264__22/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f__0625_ clkbuf_0__0625_/X vssd1 vssd1 vccd1 vccd1 _3654__84/A sky130_fd_sc_hd__clkbuf_16
XFILLER_2_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2208__B _4523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_4029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_2730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_2785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_4008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_3224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
+ _4891_/Q _2956_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3749_/A fanout187/X vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_29_2545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output82_A _5079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1782__B _4289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3055__A _5024_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4734__CLK _4943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4180_ _4737_/Q vssd1 vssd1 vccd1 vccd1 _4736_/D sky130_fd_sc_hd__inv_2
XFILLER_4_3941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_2205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_TE_B
+ _2545_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2894__A _4931_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3131_ _3131_/A vssd1 vssd1 vccd1 vccd1 _3133_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3062_ _4994_/Q _4993_/Q _4992_/Q _3098_/A vssd1 vssd1 vccd1 vccd1 _3085_/B sky130_fd_sc_hd__or4_2
XFILLER_20_3777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3502__B _3556_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4884__CLK _4920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2013_ _4462_/D _4404_/Q _4402_/Q vssd1 vssd1 vccd1 vccd1 _2013_/Y sky130_fd_sc_hd__nor3_1
XFILLER_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3182__69_A _3189__72/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3964_ _4411_/Q vssd1 vssd1 vccd1 vccd1 _4412_/D sky130_fd_sc_hd__inv_2
XFILLER_32_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_2983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2915_ _4896_/Q _2891_/D _2908_/B vssd1 vssd1 vccd1 vccd1 _2916_/B sky130_fd_sc_hd__a21bo_1
XFILLER_18_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3875__D _3875_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_2847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3895_ _3895_/A _3895_/B vssd1 vssd1 vccd1 vccd1 _4368_/D sky130_fd_sc_hd__xnor2_1
XFILLER_31_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2134__A _4491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_2137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2846_ _4859_/Q _2846_/B vssd1 vssd1 vccd1 vccd1 _4859_/D sky130_fd_sc_hd__xnor2_1
XFILLER_12_3283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2777_ _4814_/Q _4813_/Q vssd1 vssd1 vccd1 vccd1 _2777_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__1973__A _4392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout120/X fanout249/X vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_GATE_N _5048_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4516_ _2294_/B1 _4516_/D _3287_/Y vssd1 vssd1 vccd1 vccd1 _4516_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout201_A fanout202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1728_ _4971_/Q vssd1 vssd1 vccd1 vccd1 _4972_/D sky130_fd_sc_hd__inv_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_3633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4447_ _3932_/A _4447_/D _3243_/Y vssd1 vssd1 vccd1 vccd1 _4447_/Q sky130_fd_sc_hd__dfrtp_4
X_1659_ _4873_/Q vssd1 vssd1 vccd1 vccd1 _4872_/D sky130_fd_sc_hd__inv_2
XFILLER_28_2077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_2932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_3677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4378_ _4378_/CLK _4378_/D fanout219/X vssd1 vssd1 vccd1 vccd1 _4378_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_input6_A comp_high_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _3947_/A _3438_/B vssd1 vssd1 vccd1 vccd1 _3329_/Y sky130_fd_sc_hd__xnor2_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
+ _4949_/Q _3051_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_2460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4607__CLK _3861_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_2925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_2324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2044__A _2143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_2368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1883__A _1909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_2693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4757__CLK _2631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_3132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_2683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5090__A _5090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_3813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4287__CLK _4288_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_2413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2700_ _4834_/D _4776_/Q vssd1 vssd1 vccd1 vccd1 _2701_/B sky130_fd_sc_hd__xnor2_1
XFILLER_12_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2631_ _2631_/A _2631_/B _2631_/C vssd1 vssd1 vccd1 vccd1 _2631_/X sky130_fd_sc_hd__and3_1
X_3179__68 _3189__72/A vssd1 vssd1 vccd1 vccd1 _3179__68/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2562_ _4706_/Q _2562_/B vssd1 vssd1 vccd1 vccd1 _2562_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_3137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4301_ _3898_/B _4301_/D _3779__120/Y vssd1 vssd1 vccd1 vccd1 _4301_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2493_ _2493_/A _2493_/B vssd1 vssd1 vccd1 vccd1 _4669_/D sky130_fd_sc_hd__xnor2_1
XFILLER_29_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4232_ _4822_/Q vssd1 vssd1 vccd1 vccd1 _4821_/D sky130_fd_sc_hd__inv_2
XFILLER_26_3986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4163_ _4702_/Q vssd1 vssd1 vccd1 vccd1 _4703_/D sky130_fd_sc_hd__clkinv_2
XFILLER_25_1549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3513__A _3519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3114_ _3114_/A _4998_/Q vssd1 vssd1 vccd1 vccd1 _4998_/D sky130_fd_sc_hd__xor2_1
XFILLER_3_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4094_ _4606_/Q vssd1 vssd1 vccd1 vccd1 _4605_/D sky130_fd_sc_hd__inv_2
XANTENNA__3232__B _3889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3045_ _4964_/Q _4963_/Q vssd1 vssd1 vccd1 vccd1 _3045_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_20_2873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_3913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1968__A _4397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout151_A _4920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4996_ _5047_/A _4996_/D fanout242/X vssd1 vssd1 vccd1 vccd1 _4996_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_3957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4063__B _4063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3947_ _3947_/A _3947_/B vssd1 vssd1 vccd1 vccd1 _4380_/D sky130_fd_sc_hd__xnor2_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout128/X fanout246/X vssd1 vssd1 vccd1 vccd1 _5077_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_14_3389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_2081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3421__39 _3425__41/A vssd1 vssd1 vccd1 vccd1 _3421__39/Y sky130_fd_sc_hd__inv_2
X_3878_ _3870_/Y _4131_/A vssd1 vssd1 vccd1 vccd1 _3878_/X sky130_fd_sc_hd__and2b_1
XFILLER_14_2699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2829_ _4857_/Q _4856_/Q _2829_/C vssd1 vssd1 vccd1 vccd1 _2829_/X sky130_fd_sc_hd__and3_1
XANTENNA__2799__A _3877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3407__B _3440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4425__RESET_B fanout195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_3305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3732__95 _3732__95/A vssd1 vssd1 vccd1 vccd1 _3732__95/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_3349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_2626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_TE_B
+ _2538_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2039__A _4466_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_3456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_3890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1965__A1 _4392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2502__A _2566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3317__B _3889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3763__103 _3765__105/A vssd1 vssd1 vccd1 vccd1 _3763__103/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_2609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_2300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3198__6_A _3199__7/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3333__A _3925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_2125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output45_A _5042_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2891__B _4895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4850_ _4852_/CLK _4850_/D _3476__46/Y vssd1 vssd1 vccd1 vccd1 _4850_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_2032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_2043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4922__CLK _4981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3801_ _4299_/Q vssd1 vssd1 vccd1 vccd1 _4298_/D sky130_fd_sc_hd__inv_2
X_4781_ _5007_/CLK _4781_/D _3431_/Y vssd1 vssd1 vccd1 vccd1 _4781_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1993_ _4396_/Q _1993_/B vssd1 vssd1 vccd1 vccd1 _1993_/X sky130_fd_sc_hd__and2b_1
XFILLER_11_3529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3663_ _3669_/A vssd1 vssd1 vccd1 vccd1 _3663_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3508__A _4127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2412__A _2412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2614_ _4731_/Q _4730_/Q vssd1 vssd1 vccd1 vccd1 _2614_/Y sky130_fd_sc_hd__xnor2_4
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
+ _4710_/Q _2611_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_3594_ _3597_/A vssd1 vssd1 vccd1 vccd1 _3594_/Y sky130_fd_sc_hd__inv_2
X_2545_ _4699_/Q _4698_/Q vssd1 vssd1 vccd1 vccd1 _2545_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__4302__CLK _3899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_2014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_2266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2476_ _4667_/Q _4666_/Q vssd1 vssd1 vccd1 vccd1 _2476_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_5_2119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_2288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4215_ _4787_/Q vssd1 vssd1 vccd1 vccd1 _4788_/D sky130_fd_sc_hd__inv_2
XFILLER_29_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3243__A _3255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout199_A fanout221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4146_ _4687_/Q vssd1 vssd1 vccd1 vccd1 _4686_/D sky130_fd_sc_hd__inv_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_2979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ _4571_/Q vssd1 vssd1 vccd1 vccd1 _4572_/D sky130_fd_sc_hd__inv_2
XFILLER_0_2742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_2681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3028_ _3028_/A vssd1 vssd1 vccd1 vccd1 _3028_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4979_ _4131_/B _4979_/D _3548_/Y vssd1 vssd1 vccd1 vccd1 _4979_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_2846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout240 fanout241/X vssd1 vssd1 vccd1 vccd1 fanout240/X sky130_fd_sc_hd__buf_2
XANTENNA__4249__A _4249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3769__108_A _3770__109/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout251 fanout252/X vssd1 vssd1 vccd1 vccd1 fanout251/X sky130_fd_sc_hd__buf_2
XFILLER_1_3229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_2675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
+ _4768_/Q _2708_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_21_2445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_2539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4945__CLK _2807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_2341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_3253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3328__A _3340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4347__RESET_B fanout195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4325__CLK _5040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_2883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_3118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_2312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2330_ _4581_/Q _2305_/D _2322_/B vssd1 vssd1 vccd1 vccd1 _2331_/B sky130_fd_sc_hd__a21bo_1
X_2261_ _4559_/D _4518_/Q vssd1 vssd1 vccd1 vccd1 _2262_/D sky130_fd_sc_hd__xnor2_1
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
+ _4425_/Q _2102_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__3063__A _4991_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2115__A1 _3892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4000_ _4123_/B vssd1 vssd1 vccd1 vccd1 _4000_/Y sky130_fd_sc_hd__clkinv_4
X_2192_ _4496_/Q _2192_/B vssd1 vssd1 vccd1 vccd1 _4496_/D sky130_fd_sc_hd__xor2_1
XFILLER_1_3763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3510__B _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4902_ _4905_/CLK _4902_/D fanout231/X vssd1 vssd1 vccd1 vccd1 _4902_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4833_ input30/X _4833_/D fanout237/X vssd1 vssd1 vccd1 vccd1 _4834_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_11_4027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_3473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4764_ _4811_/CLK _4764_/D fanout250/X vssd1 vssd1 vccd1 vccd1 _4764_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1976_ _1973_/X _1974_/Y _1975_/X vssd1 vssd1 vccd1 vccd1 _1977_/B sky130_fd_sc_hd__o21a_1
XFILLER_11_3359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4770__RESET_B fanout253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_2051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3715_ _3721_/A vssd1 vssd1 vccd1 vccd1 _3715_/Y sky130_fd_sc_hd__inv_2
X_4695_ _3386_/Y _4695_/D _3674_/Y vssd1 vssd1 vccd1 vccd1 _4695_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3238__A _4004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3646_ _4195_/A vssd1 vssd1 vccd1 vccd1 _3646_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_3834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3577_ _3588_/A vssd1 vssd1 vccd1 vccd1 _3587_/A sky130_fd_sc_hd__buf_6
XFILLER_28_3889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2528_ _4741_/D _4683_/Q _4681_/Q vssd1 vssd1 vccd1 vccd1 _2528_/Y sky130_fd_sc_hd__nor3_1
XFILLER_9_2052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_2096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3163__63 _3169__65/A vssd1 vssd1 vccd1 vccd1 _3163__63/Y sky130_fd_sc_hd__inv_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2459_ _2464_/C _2459_/B vssd1 vssd1 vccd1 vccd1 _2459_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_2951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_2765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4129_ _4129_/A _4129_/B vssd1 vssd1 vccd1 vccd1 _4657_/D sky130_fd_sc_hd__xor2_1
XANTENNA__3701__A _4071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3420__B _3420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3082__A2 _3058_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4858__RESET_B fanout228/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
+ _4483_/Q _2201_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_16_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2036__B _4430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_3871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4440__RESET_B fanout198/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_2293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4498__CLK _4248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_2704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_2715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3611__A _3616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_4016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_4038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1830_ _1777_/C _1826_/Y _1823_/X vssd1 vssd1 vccd1 vccd1 _1831_/B sky130_fd_sc_hd__o21ai_1
XFILLER_15_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_2912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_3094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_2945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_4082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1761_ _4247_/Y _1761_/B _1761_/C vssd1 vssd1 vccd1 vccd1 _1763_/B sky130_fd_sc_hd__or3_2
XANTENNA__3058__A _4989_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3500_ _5062_/A vssd1 vssd1 vccd1 vccd1 _3519_/A sky130_fd_sc_hd__buf_6
XFILLER_10_3381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4480_ _3892_/A _4480_/D _3267__23/Y vssd1 vssd1 vccd1 vccd1 _4480_/Q sky130_fd_sc_hd__dfrtp_1
X_1692_ _4920_/Q vssd1 vssd1 vccd1 vccd1 _4921_/D sky130_fd_sc_hd__inv_2
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_GATE_N
+ _3576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3431_ _3445_/A vssd1 vssd1 vccd1 vccd1 _3431_/Y sky130_fd_sc_hd__inv_2
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2897__A _4895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3362_ _3895_/A _3372_/B vssd1 vssd1 vccd1 vccd1 _3362_/Y sky130_fd_sc_hd__xnor2_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ _2996_/A _2361_/B _2361_/C vssd1 vssd1 vccd1 vccd1 _2314_/B sky130_fd_sc_hd__and3_1
XFILLER_6_2236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3293_/Y sky130_fd_sc_hd__inv_2
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_3847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _5040_/A vssd1 vssd1 vccd1 vccd1 _5032_/X sky130_fd_sc_hd__buf_2
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _4526_/Q _2244_/B vssd1 vssd1 vccd1 vccd1 _4526_/D sky130_fd_sc_hd__xnor2_1
XFILLER_26_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2175_ _4491_/Q _2175_/B vssd1 vssd1 vccd1 vccd1 _4491_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__3521__A _5062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout144/X fanout215/X vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__3240__B _3438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4951__RESET_B fanout208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4269__RESET_B _4359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4816_ _3451_/Y _4816_/D _3640_/Y vssd1 vssd1 vccd1 vccd1 _4816_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout231_A fanout235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4747_ input21/X _4747_/D fanout222/X vssd1 vssd1 vccd1 vccd1 _4747_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1959_ _4388_/Q _4387_/Q vssd1 vssd1 vccd1 vccd1 _1959_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_11_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4678_ _4717_/CLK _4678_/D fanout255/X vssd1 vssd1 vccd1 vccd1 _4678_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_3642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput38 _5035_/X vssd1 vssd1 vccd1 vccd1 cclk_I[3] sky130_fd_sc_hd__buf_2
XFILLER_28_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput49 _5046_/X vssd1 vssd1 vccd1 vccd1 cclk_Q[6] sky130_fd_sc_hd__buf_2
XFILLER_28_2952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_3539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3415__B _3420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_2770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3431__A _3445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_2595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__0641_ clkbuf_0__0641_/X vssd1 vssd1 vccd1 vccd1 _3784__125/A sky130_fd_sc_hd__clkbuf_16
XFILLER_17_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4246__B _4250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4252__A1 _4126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_4082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_2333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_3089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_4118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_TE_B
+ _2613_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_3428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2213__C _4524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3606__A _5062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3771__110_A _3776__115/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2510__A _4674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3325__B _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_3049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_2326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_3937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_3891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3341__A _3895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_2177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4709__RESET_B fanout247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3980_ _4443_/Q vssd1 vssd1 vccd1 vccd1 _4444_/D sky130_fd_sc_hd__inv_2
XANTENNA__3313__25_A _3365__31/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_3145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2931_ _4899_/Q _2931_/B vssd1 vssd1 vccd1 vccd1 _4899_/D sky130_fd_sc_hd__xnor2_1
XFILLER_15_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_4133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_4144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4362__RESET_B fanout202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2862_ _2861_/Y _2817_/C _4865_/Q vssd1 vssd1 vccd1 vccd1 _2863_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_3443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_2319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4601_ _4981_/CLK _4601_/D _3332_/Y vssd1 vssd1 vccd1 vccd1 _4601_/Q sky130_fd_sc_hd__dfrtp_1
X_1813_ _4280_/Q _1813_/B vssd1 vssd1 vccd1 vccd1 _4280_/D sky130_fd_sc_hd__xnor2_1
XFILLER_15_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_TE_B
+ _3051_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2793_ _2793_/A vssd1 vssd1 vccd1 vccd1 _2795_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_2753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5019__CLK input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4532_ _4532_/CLK _4532_/D fanout211/X vssd1 vssd1 vccd1 vccd1 _4532_/Q sky130_fd_sc_hd__dfstp_1
X_1744_ _5003_/Q vssd1 vssd1 vccd1 vccd1 _5004_/D sky130_fd_sc_hd__inv_2
X_4463_ input26/X _4463_/D fanout198/X vssd1 vssd1 vccd1 vccd1 _4464_/D sky130_fd_sc_hd__dfrtp_1
X_1675_ _4889_/Q vssd1 vssd1 vccd1 vccd1 _4888_/D sky130_fd_sc_hd__inv_2
XANTENNA__3516__A _3934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3414_ _3414_/A vssd1 vssd1 vccd1 vccd1 _3414_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2420__A _2566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4394_ _4429_/CLK _4394_/D fanout188/X vssd1 vssd1 vccd1 vccd1 _4394_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_1608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3345_ _3361_/A vssd1 vssd1 vccd1 vccd1 _3345_/Y sky130_fd_sc_hd__inv_2
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout158/X fanout205/X vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__dlrtn_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3276_ _3935_/A _3440_/B vssd1 vssd1 vccd1 vccd1 _3276_/Y sky130_fd_sc_hd__xnor2_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5015_ _3930_/X _5015_/D _3569_/Y vssd1 vssd1 vccd1 vccd1 _5015_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_6_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2227_ _2218_/C _2226_/X _2173_/X vssd1 vssd1 vccd1 vccd1 _2228_/B sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout181_A _5057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3251__A _3255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2158_ _4486_/Q _2158_/B vssd1 vssd1 vccd1 vccd1 _4486_/D sky130_fd_sc_hd__xnor2_1
XFILLER_17_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_2208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2089_ _4438_/Q _2089_/B vssd1 vssd1 vccd1 vccd1 _4438_/D sky130_fd_sc_hd__xnor2_1
XFILLER_35_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_3554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5063_/A fanout251/X vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_17_1996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_2263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3426__A _3896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_4048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_3419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4536__CLK _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_2657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2984__B _4945_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_2370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_4100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_2497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_3129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4686__CLK _5007_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f__0624_ clkbuf_0__0624_/X vssd1 vssd1 vccd1 vccd1 _3656_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_31_4008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_2428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2208__C _4522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_2742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5088__A _5088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2505__A _2566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_2797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_2005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_2027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_2049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_3236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3336__A _3340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2240__A _2327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3130_ _5026_/Q _5025_/D vssd1 vssd1 vccd1 vccd1 _3131_/A sky130_fd_sc_hd__and2b_1
XFILLER_20_3723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2894__B _4905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3061_ _5024_/D _4998_/Q _4996_/Q _4995_/Q vssd1 vssd1 vccd1 vccd1 _3098_/A sky130_fd_sc_hd__or4_1
XFILLER_20_3767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2012_ _4462_/D _4404_/Q _4402_/Q vssd1 vssd1 vccd1 vccd1 _2012_/X sky130_fd_sc_hd__and3_1
XFILLER_23_1499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2227__B1 _2173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3963_ _4412_/Q vssd1 vssd1 vccd1 vccd1 _4411_/D sky130_fd_sc_hd__inv_2
X_2914_ _4894_/Q _2914_/B vssd1 vssd1 vccd1 vccd1 _4894_/D sky130_fd_sc_hd__xnor2_1
XFILLER_14_2826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3894_ _4368_/Q vssd1 vssd1 vccd1 vccd1 _3895_/A sky130_fd_sc_hd__buf_12
XFILLER_31_3863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4409__CLK _4063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_2296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2845_ _2916_/A _2845_/B vssd1 vssd1 vccd1 vccd1 _2846_/B sky130_fd_sc_hd__nand2_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_2149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2776_ _3114_/A _4812_/Q vssd1 vssd1 vccd1 vccd1 _4812_/D sky130_fd_sc_hd__xor2_1
X_4515_ _3286_/Y _4515_/D _3723_/Y vssd1 vssd1 vccd1 vccd1 _4515_/Q sky130_fd_sc_hd__dfrtp_1
X_1727_ _4972_/Q vssd1 vssd1 vccd1 vccd1 _4971_/D sky130_fd_sc_hd__inv_2
XFILLER_12_1860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3246__A _3917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2150__A _2178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4559__CLK input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4446_ _3242_/Y _4446_/D _3745_/Y vssd1 vssd1 vccd1 vccd1 _4446_/Q sky130_fd_sc_hd__dfrtp_4
X_1658_ _4870_/Q vssd1 vssd1 vccd1 vccd1 _4871_/D sky130_fd_sc_hd__inv_2
XFILLER_8_2117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_2911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4377_ _4658_/CLK _4377_/D fanout212/X vssd1 vssd1 vccd1 vccd1 _4377_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3328_ _3340_/A vssd1 vssd1 vccd1 vccd1 _3328_/Y sky130_fd_sc_hd__inv_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_3485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_2784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2466__B1 _2465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4284__RESET_B fanout194/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout119/X fanout248/X vssd1 vssd1 vccd1 vccd1 _5078_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_3649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_2472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_2661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_4042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_3216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_2559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3258__18 _3262__21/A vssd1 vssd1 vccd1 vccd1 _4471_/CLK sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_0__1637__A _3194_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_2203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2235__A _4526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_3137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2630_ _2464_/C _2456_/Y _4063_/B vssd1 vssd1 vccd1 vccd1 _2631_/C sky130_fd_sc_hd__a21o_1
XFILLER_31_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2561_ _4707_/Q _4706_/Q _2561_/C vssd1 vssd1 vccd1 vccd1 _2561_/X sky130_fd_sc_hd__and3_1
XFILLER_29_2310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3066__A _3066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4300_ _3914_/A _4300_/D _3158__58/Y vssd1 vssd1 vccd1 vccd1 _4300_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_3149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_2343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2492_ _2490_/X _2491_/Y _1975_/X vssd1 vssd1 vccd1 vccd1 _2493_/B sky130_fd_sc_hd__o21a_1
XFILLER_29_3099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4231_ _4819_/Q vssd1 vssd1 vccd1 vccd1 _4820_/D sky130_fd_sc_hd__inv_2
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4162_ _4703_/Q vssd1 vssd1 vccd1 vccd1 _4702_/D sky130_fd_sc_hd__inv_2
XANTENNA__3161__61_A _3169__65/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3113_ _4997_/Q _3113_/B vssd1 vssd1 vccd1 vccd1 _4997_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_3625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4093_ _4603_/Q vssd1 vssd1 vccd1 vccd1 _4604_/D sky130_fd_sc_hd__inv_2
XFILLER_3_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3044_ _3114_/A _4962_/Q vssd1 vssd1 vccd1 vccd1 _4962_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_3669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_4003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_4036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_4047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_4058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4995_ _5047_/A _4995_/D fanout242/X vssd1 vssd1 vccd1 vccd1 _4995_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_3493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_3969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2145__A _4485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3946_ _3946_/A vssd1 vssd1 vccd1 vccd1 _3947_/A sky130_fd_sc_hd__buf_12
XFILLER_14_3357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout144_A _5059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4063__C _4063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3877_ _3877_/A _4131_/A vssd1 vssd1 vccd1 vccd1 _3925_/B sky130_fd_sc_hd__nor2_4
XFILLER_34_2093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2828_ _4854_/Q _2828_/B vssd1 vssd1 vccd1 vccd1 _4854_/D sky130_fd_sc_hd__xor2_1
XANTENNA__4381__CLK _3845_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3575__55 _3656_/A vssd1 vssd1 vccd1 vccd1 _5031_/CLK sky130_fd_sc_hd__inv_2
X_2759_ _4806_/Q _2759_/B vssd1 vssd1 vccd1 vccd1 _4806_/D sky130_fd_sc_hd__xnor2_1
XFILLER_30_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_4143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4429_ _4429_/CLK _4429_/D fanout194/X vssd1 vssd1 vccd1 vccd1 _4429_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_8_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3704__A _4071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3201__9_A _3201__9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_GATE_N _4359_/CLK
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_2570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_2567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4724__CLK _1765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_2111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4874__CLK _4187_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3708__93 _3732__95/A vssd1 vssd1 vccd1 vccd1 _3708__93/Y sky130_fd_sc_hd__inv_2
XFILLER_26_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3157__57_A _3159__59/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3614__A _3616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_2251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3333__B _3442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_2367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_2137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2891__C _4894_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_2000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3800_ _4296_/Q vssd1 vssd1 vccd1 vccd1 _4297_/D sky130_fd_sc_hd__inv_2
X_4780_ _3430_/Y _4780_/D _3651_/Y vssd1 vssd1 vccd1 vccd1 _4780_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1992_ _4397_/Q _1992_/B vssd1 vssd1 vccd1 vccd1 _1993_/B sky130_fd_sc_hd__nor2_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3731_ _4010_/A vssd1 vssd1 vccd1 vccd1 _3731_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3662_ _3669_/A vssd1 vssd1 vccd1 vccd1 _3662_/Y sky130_fd_sc_hd__inv_2
X_2613_ _4729_/Q _4728_/Q vssd1 vssd1 vccd1 vccd1 _2613_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__3508__B _4129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3593_ _3597_/A vssd1 vssd1 vccd1 vccd1 _3593_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2544_ _4697_/Q _4696_/Q vssd1 vssd1 vccd1 vccd1 _2544_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_26_3740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4905__RESET_B fanout231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2475_ _4665_/Q _4664_/Q vssd1 vssd1 vccd1 vccd1 _2475_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_29_2195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4214_ _4788_/Q vssd1 vssd1 vccd1 vccd1 _4787_/D sky130_fd_sc_hd__clkinv_2
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5056_/A fanout193/X vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_22_3648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4145_ _4684_/Q vssd1 vssd1 vccd1 vccd1 _4685_/D sky130_fd_sc_hd__inv_2
XFILLER_20_4084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4076_ _4572_/Q vssd1 vssd1 vccd1 vccd1 _4571_/D sky130_fd_sc_hd__clkinv_2
X_3027_ _4956_/Q _3027_/B vssd1 vssd1 vccd1 vccd1 _4956_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_3499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4747__CLK input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_3733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4978_ _3547_/Y _4978_/D _3590_/Y vssd1 vssd1 vccd1 vccd1 _4978_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_3777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4897__CLK _4905_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_2442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3929_ _3929_/A vssd1 vssd1 vccd1 vccd1 _4124_/B sky130_fd_sc_hd__inv_2
XANTENNA__2603__A _2680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
+ _4868_/Q _2887_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__2041__C _4431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4646__RESET_B _3684_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_4078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3434__A _4065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout230 input33/X vssd1 vssd1 vccd1 vccd1 fanout230/X sky130_fd_sc_hd__clkbuf_4
Xfanout241 fanout257/X vssd1 vssd1 vccd1 vccd1 fanout241/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4277__CLK _4281_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4249__B _4250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_2560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout252 fanout253/X vssd1 vssd1 vccd1 vccd1 fanout252/X sky130_fd_sc_hd__buf_2
XFILLER_25_2571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf _4314_/Q _1919_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_21_2435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_3010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_2353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_3221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_2542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3609__A _3616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2513__A _4675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2060__A1 _4431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3344__A _4127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2260_ _4531_/Q _2260_/B vssd1 vssd1 vccd1 vccd1 _4531_/D sky130_fd_sc_hd__xnor2_1
XFILLER_26_2379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2115__A2 _3899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2191_ _3066_/A _2191_/B _2191_/C _2191_/D vssd1 vssd1 vccd1 vccd1 _2192_/B sky130_fd_sc_hd__and4_1
XFILLER_1_3753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_3775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4901_ _4901_/CLK _4901_/D fanout232/X vssd1 vssd1 vccd1 vccd1 _4901_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_3029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2919__A_N _4897_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4832_ _3467_/Y _4832_/D _3631_/Y vssd1 vssd1 vccd1 vccd1 _4832_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_3452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_4039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_3305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_1_0_0_clk_master_A clkbuf_0_clk_master/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4763_ _4803_/CLK _4763_/D fanout247/X vssd1 vssd1 vccd1 vccd1 _4763_/Q sky130_fd_sc_hd__dfrtp_4
X_1975_ _2858_/A vssd1 vssd1 vccd1 vccd1 _1975_/X sky130_fd_sc_hd__buf_12
XANTENNA__3519__A _3519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3714_ _3721_/A vssd1 vssd1 vccd1 vccd1 _3714_/Y sky130_fd_sc_hd__inv_2
X_4694_ _4920_/CLK _4694_/D _3385_/Y vssd1 vssd1 vccd1 vccd1 _4694_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_31_2063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3238__B _3491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3645_ _4195_/A vssd1 vssd1 vccd1 vccd1 _3645_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3576_ _3576_/A vssd1 vssd1 vccd1 vccd1 _3576_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3000__B1 _2143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout107_A _4905_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2527_ _4741_/D _4683_/Q _4681_/Q vssd1 vssd1 vccd1 vccd1 _2527_/X sky130_fd_sc_hd__and3_1
XFILLER_0_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_3401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3254__A _3891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_2064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2458_ _3908_/A _2807_/A vssd1 vssd1 vccd1 vccd1 _2459_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_3445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2389_ _2387_/X _2388_/Y _1975_/X vssd1 vssd1 vccd1 vccd1 _2390_/B sky130_fd_sc_hd__o21a_1
XFILLER_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4128_ _4657_/Q vssd1 vssd1 vccd1 vccd1 _4129_/A sky130_fd_sc_hd__buf_12
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout136/X fanout238/X vssd1 vssd1 vccd1 vccd1 _5084_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4059_ _4563_/Q _4564_/Q vssd1 vssd1 vccd1 vccd1 _4126_/A sky130_fd_sc_hd__xnor2_4
XFILLER_20_2490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3429__A _3445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4898__RESET_B fanout232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3148__B _3148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_4107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_4046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_4068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3164__A _3945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_2666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4912__CLK _5007_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_3091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_2495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_2014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_3062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_2069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3339__A _3903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_3669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2243__A _2327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1760_ _1760_/A vssd1 vssd1 vccd1 vccd1 _1760_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_2957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3058__B _4988_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1691_ _4921_/Q vssd1 vssd1 vccd1 vccd1 _4920_/D sky130_fd_sc_hd__inv_2
XANTENNA__1792__B1 _1791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3430_ _4189_/A _4190_/A vssd1 vssd1 vccd1 vccd1 _3430_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__2897__B _4894_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3361_ _3361_/A vssd1 vssd1 vccd1 vccd1 _3361_/Y sky130_fd_sc_hd__inv_2
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2312_ _4577_/Q _2316_/B _2318_/A vssd1 vssd1 vccd1 vccd1 _2361_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__4592__CLK _4188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3292_ _4065_/A _3543_/B vssd1 vssd1 vccd1 vccd1 _3292_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_3_3826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5031_/CLK _5031_/D fanout226/X vssd1 vssd1 vccd1 vccd1 _5031_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_26_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2243_ _2327_/A _2243_/B vssd1 vssd1 vccd1 vccd1 _2244_/B sky130_fd_sc_hd__nand2_2
XFILLER_22_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2174_ _2134_/D _2172_/Y _2173_/X vssd1 vssd1 vccd1 vccd1 _2175_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__2418__A _2418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
+ _4614_/Q _2440_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4815_ _4187_/Y _4815_/D _3450_/Y vssd1 vssd1 vccd1 vccd1 _4815_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_30_3725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3249__A _3255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4991__RESET_B fanout242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout224_A fanout230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4746_ input21/X _4746_/D fanout222/X vssd1 vssd1 vccd1 vccd1 _4747_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_33_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1958_ _4386_/Q _4385_/Q vssd1 vssd1 vccd1 vccd1 _1958_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_11_2445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4677_ _4717_/CLK _4677_/D fanout254/X vssd1 vssd1 vccd1 vccd1 _4677_/Q sky130_fd_sc_hd__dfrtp_1
X_1889_ _4319_/Q _4318_/Q _1857_/D _1886_/B vssd1 vssd1 vccd1 vccd1 _1890_/B sky130_fd_sc_hd__a31o_1
XFILLER_28_3610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1992__A _4397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4935__CLK _5030_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput39 _5036_/X vssd1 vssd1 vccd1 vccd1 cclk_I[4] sky130_fd_sc_hd__buf_2
X_3559_ _3571_/A vssd1 vssd1 vccd1 vccd1 _3559_/Y sky130_fd_sc_hd__inv_2
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3684_/A fanout217/X vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_0_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3371__34_A _3469__42/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_4059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_3275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3712__A _3721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_3369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__0640_ clkbuf_0__0640_/X vssd1 vssd1 vccd1 vccd1 _3776__115/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__4315__CLK _5040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_3625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_2913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4252__A2 _4248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_3046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_A
+ _4764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_4094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3206__13 _3262__21/A vssd1 vssd1 vccd1 vccd1 _4380_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_3934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_3371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4465__CLK input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_2209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_3967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_2091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
+ _4672_/Q _2542_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__2510__B _2510_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_2463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_3905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_3949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3622__A _4256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3341__B _3372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2238__A _4524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_2095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_3834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2930_ _2890_/D _2929_/Y _2858_/X vssd1 vssd1 vccd1 vccd1 _2931_/B sky130_fd_sc_hd__o21ai_1
XFILLER_18_3889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_3157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2861_ _2861_/A vssd1 vssd1 vccd1 vccd1 _2861_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_2478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_2489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4600_ _3331_/Y _4600_/D _3701_/Y vssd1 vssd1 vccd1 vccd1 _4600_/Q sky130_fd_sc_hd__dfrtp_1
X_1812_ _1779_/D _1811_/X _3109_/A vssd1 vssd1 vccd1 vccd1 _1813_/B sky130_fd_sc_hd__o21ai_1
X_2792_ _4840_/Q _4839_/D vssd1 vssd1 vccd1 vccd1 _2793_/A sky130_fd_sc_hd__and2b_1
XFILLER_34_1777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3602__76 _3654__84/A vssd1 vssd1 vccd1 vccd1 _3602__76/Y sky130_fd_sc_hd__inv_2
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1743_ _5004_/Q vssd1 vssd1 vccd1 vccd1 _5003_/D sky130_fd_sc_hd__inv_2
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_2765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4531_ _4532_/CLK _4531_/D fanout212/X vssd1 vssd1 vccd1 vccd1 _4531_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_29_3930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1674_ _4886_/Q vssd1 vssd1 vccd1 vccd1 _4887_/D sky130_fd_sc_hd__inv_2
X_4462_ input26/X _4462_/D fanout199/X vssd1 vssd1 vccd1 vccd1 _4463_/D sky130_fd_sc_hd__dfrtp_1
XANTENNA__3516__B _3933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3413_ _3912_/A _3446_/B vssd1 vssd1 vccd1 vccd1 _3413_/Y sky130_fd_sc_hd__xnor2_1
X_4393_ _4402_/CLK _4393_/D fanout190/X vssd1 vssd1 vccd1 vccd1 _4393_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_2249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3344_ _4127_/A _4129_/A vssd1 vssd1 vccd1 vccd1 _3344_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_7_3770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_2056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3275_ _3287_/A vssd1 vssd1 vccd1 vccd1 _3275_/Y sky130_fd_sc_hd__inv_2
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3532__A _3588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4338__CLK _3899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _3568_/Y _5014_/D _3579_/Y vssd1 vssd1 vccd1 vccd1 _5014_/Q sky130_fd_sc_hd__dfrtp_1
X_2226_ _4522_/Q _2226_/B vssd1 vssd1 vccd1 vccd1 _2226_/X sky130_fd_sc_hd__and2b_1
XFILLER_3_3689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_4081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_2966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2157_ _2178_/A _2157_/B vssd1 vssd1 vccd1 vccd1 _2158_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_4012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout174_A _4121_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_4056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2088_ _2178_/A _2088_/B vssd1 vssd1 vccd1 vccd1 _2089_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4488__CLK _5042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_4078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1987__A _2061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_2810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4729_ _3405_/Y _4729_/D _3664_/Y vssd1 vssd1 vccd1 vccd1 _4729_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_2876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_4141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[1\].w1.ro_block_I.ro_pol.tribuf.t_buf_TE_B _2130_/Y vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_4027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2787__A_N _4836_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3426__B _3904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3442__A _3924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2058__A _2061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_4112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__0623_ clkbuf_0__0623_/X vssd1 vssd1 vccd1 vccd1 _3470_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_2_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3683__90 _3683__90/A vssd1 vssd1 vccd1 vccd1 _3683__90/Y sky130_fd_sc_hd__inv_2
XFILLER_16_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_2607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5055_/A fanout244/X vssd1 vssd1 vccd1 vccd1 _5079_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3617__A _5062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_TE_B
+ _2714_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_3860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_3893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3352__A _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3060_ _4986_/Q _4985_/Q _3068_/C _3071_/A vssd1 vssd1 vccd1 vccd1 _3112_/B sky130_fd_sc_hd__a31o_1
XFILLER_27_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2011_ _4400_/Q _2011_/B vssd1 vssd1 vccd1 vccd1 _4400_/D sky130_fd_sc_hd__xnor2_1
XFILLER_18_3631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2227__A1 _2218_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_A
+ _4897_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3962_ _4409_/Q vssd1 vssd1 vccd1 vccd1 _4410_/D sky130_fd_sc_hd__inv_2
XFILLER_18_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4780__CLK _3430_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2913_ _2916_/A _2913_/B vssd1 vssd1 vccd1 vccd1 _2914_/B sky130_fd_sc_hd__nand2_1
XFILLER_14_2805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3893_ _4367_/Q _3895_/B vssd1 vssd1 vccd1 vccd1 _4367_/D sky130_fd_sc_hd__xnor2_1
XFILLER_17_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4333__D _4333_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2844_ _4860_/Q _2819_/D _2837_/B vssd1 vssd1 vccd1 vccd1 _2845_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__2134__C _4489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_2562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2775_ _4811_/Q _2775_/B vssd1 vssd1 vccd1 vccd1 _4811_/D sky130_fd_sc_hd__xor2_1
XANTENNA__3527__A _3916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2431__A _4652_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4514_ _3899_/A _4514_/D _3285_/Y vssd1 vssd1 vccd1 vccd1 _4514_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1973__C _1973_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1726_ _4969_/Q vssd1 vssd1 vccd1 vccd1 _4970_/D sky130_fd_sc_hd__inv_2
X_3153__117 _3784__125/A vssd1 vssd1 vccd1 vccd1 _3153__117/Y sky130_fd_sc_hd__inv_2
XANTENNA__3246__B _3444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4445_ _4063_/B _4445_/D _3241_/Y vssd1 vssd1 vccd1 vccd1 _4445_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_3782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4376_ _4376_/CLK _4376_/D fanout214/X vssd1 vssd1 vccd1 vccd1 _4376_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3327_ _4004_/A _3491_/B vssd1 vssd1 vccd1 vccd1 _3327_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_25_2967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2466__A1 _2470_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2209_ _4519_/Q vssd1 vssd1 vccd1 vccd1 _2221_/A sky130_fd_sc_hd__inv_2
XFILLER_19_3417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2466__B2 _4131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
+ _4433_/Q _2094_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2606__A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_4020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3437__A _3445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_2673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2341__A _2412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_2684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_4054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2060__B1_N _2053_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_4076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_3364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_2580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2154__B1 _2003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4653__CLK input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3172__A _3777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5009__CLK _1765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3900__A _3900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[0\].w1.ro_block_Q.ro_pol.tribuf.t_buf _2108_/X _1956_/Y vssd1
+ vssd1 vccd1 vccd1 _5090_/A sky130_fd_sc_hd__ebufn_8
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5099__A _5099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2516__A _4676_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0__1653__A _3470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_3149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3347__A _3361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_3023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2560_ _4704_/Q _2560_/B vssd1 vssd1 vccd1 vccd1 _4704_/D sky130_fd_sc_hd__xor2_1
XFILLER_5_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_3078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2491_ _4670_/Q _2491_/B vssd1 vssd1 vccd1 vccd1 _2491_/Y sky130_fd_sc_hd__nor2_1
X_4230_ _4820_/Q vssd1 vssd1 vccd1 vccd1 _4819_/D sky130_fd_sc_hd__inv_2
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_3819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4161_ _4700_/Q vssd1 vssd1 vccd1 vccd1 _4701_/D sky130_fd_sc_hd__inv_2
XFILLER_7_2151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_3773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3112_ _3112_/A _3112_/B _3112_/C _3112_/D vssd1 vssd1 vccd1 vccd1 _3113_/B sky130_fd_sc_hd__and4_1
X_4092_ _4604_/Q vssd1 vssd1 vccd1 vccd1 _4603_/D sky130_fd_sc_hd__inv_2
XFILLER_0_3637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3043_ _4961_/Q _3043_/B vssd1 vssd1 vccd1 vccd1 _4961_/D sky130_fd_sc_hd__xor2_1
XFILLER_3_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_2853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1968__C _4395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4994_ _5047_/A _4994_/D fanout239/X vssd1 vssd1 vccd1 vccd1 _4994_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_14_3325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3945_ _3945_/A _3947_/B vssd1 vssd1 vccd1 vccd1 _4379_/D sky130_fd_sc_hd__xnor2_1
XFILLER_18_2771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4526__CLK _5042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3876_ _3876_/A vssd1 vssd1 vccd1 vccd1 _4131_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout137_A _5060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2827_ _2996_/A _2875_/B _2875_/C vssd1 vssd1 vccd1 vccd1 _2828_/B sky130_fd_sc_hd__and3_1
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout180/X fanout188/X vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_14_1956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3257__A _5057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2161__A _4487_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0__0625_ _3601_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0625_/X sky130_fd_sc_hd__clkbuf_16
X_2758_ _2719_/D _2757_/Y _2687_/X vssd1 vssd1 vccd1 vccd1 _2759_/B sky130_fd_sc_hd__o21ai_1
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4676__CLK _4717_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1709_ _4937_/Q _1709_/B vssd1 vssd1 vccd1 vccd1 _4938_/D sky130_fd_sc_hd__xnor2_1
X_2689_ _4770_/Q _2689_/B vssd1 vssd1 vccd1 vccd1 _4770_/D sky130_fd_sc_hd__xnor2_1
XFILLER_21_4008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4428_ _4429_/CLK _4428_/D fanout194/X vssd1 vssd1 vccd1 vccd1 _4428_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_2742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_2983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4359_ _4359_/CLK _4359_/D fanout195/X vssd1 vssd1 vccd1 vccd1 _4359_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3884__A0 _3882_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3720__A _3721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4288__SET_B fanout199/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_3723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1965__A3 _1973_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3167__A _3933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_2517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_0__1648__A _3368_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_2274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_3957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_2149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_2081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__1638_ clkbuf_0__1638_/X vssd1 vssd1 vccd1 vccd1 _3262__21/A sky130_fd_sc_hd__clkbuf_16
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3770__109 _3770__109/A vssd1 vssd1 vccd1 vccd1 _3770__109/Y sky130_fd_sc_hd__inv_2
XFILLER_15_3645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[6\].w1.ro_block_Q.ro_pol.tribuf.t_buf _3129_/X _2981_/Y vssd1
+ vssd1 vccd1 vccd1 _5090_/A sky130_fd_sc_hd__ebufn_8
XFILLER_15_2911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1991_ _4394_/Q _1991_/B vssd1 vssd1 vccd1 vccd1 _4394_/D sky130_fd_sc_hd__xnor2_1
XFILLER_13_4070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3730_ _4010_/A vssd1 vssd1 vccd1 vccd1 _3730_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_2988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3661_ _3669_/A vssd1 vssd1 vccd1 vccd1 _3661_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2612_ _4727_/Q _4726_/Q vssd1 vssd1 vccd1 vccd1 _2612_/Y sky130_fd_sc_hd__xnor2_1
X_3592_ _3597_/A vssd1 vssd1 vccd1 vccd1 _3592_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2543_ _4695_/Q _4694_/Q vssd1 vssd1 vccd1 vccd1 _2543_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__2848__A_N _4861_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2474_ _4663_/Q _4662_/Q vssd1 vssd1 vccd1 vccd1 _2474_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_29_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2118__B1 _3888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4213_ _4785_/Q vssd1 vssd1 vccd1 vccd1 _4786_/D sky130_fd_sc_hd__inv_2
XFILLER_25_2049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_2915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4144_ _4685_/Q vssd1 vssd1 vccd1 vccd1 _4684_/D sky130_fd_sc_hd__inv_2
XFILLER_4_3581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_4096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_3362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4075_ _4569_/Q vssd1 vssd1 vccd1 vccd1 _4570_/D sky130_fd_sc_hd__inv_2
XANTENNA__3540__A _3550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3026_ _2987_/D _3025_/Y _1791_/X vssd1 vssd1 vccd1 vccd1 _3027_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_3489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout254_A fanout255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4977_ _5013_/CLK _4977_/D _3546_/Y vssd1 vssd1 vccd1 vccd1 _4977_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_3133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1995__A _4395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3928_ _3934_/A _3933_/A vssd1 vssd1 vccd1 vccd1 _3929_/A sky130_fd_sc_hd__xnor2_4
XFILLER_10_2307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3859_ _4369_/Q vssd1 vssd1 vccd1 vccd1 _3904_/A sky130_fd_sc_hd__buf_6
XFILLER_20_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3715__A _3721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_4068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3434__B _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout220 fanout221/X vssd1 vssd1 vccd1 vccd1 fanout220/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_3126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5048_/A fanout191/X vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__dlrtn_1
Xfanout231 fanout235/X vssd1 vssd1 vccd1 vccd1 fanout231/X sky130_fd_sc_hd__buf_4
Xfanout242 fanout257/X vssd1 vssd1 vccd1 vccd1 fanout242/X sky130_fd_sc_hd__buf_4
XFILLER_21_3137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout253 fanout256/X vssd1 vssd1 vccd1 vccd1 fanout253/X sky130_fd_sc_hd__clkbuf_4
XFILLER_19_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4615__RESET_B fanout232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_2519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3450__A _3466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2066__A _4431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout128/X fanout243/X vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__dlrtn_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_3277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2596__B1 _2518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2060__A2 _2036_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4991__CLK _5047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3625__A _4256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3344__B _4129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3063__C _4989_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2190_ _4555_/D _4482_/Q vssd1 vssd1 vccd1 vccd1 _2191_/D sky130_fd_sc_hd__xnor2_1
XFILLER_1_3721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4371__CLK _3598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3360__A _3903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4900_ _4901_/CLK _4900_/D fanout232/X vssd1 vssd1 vccd1 vccd1 _4900_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4831_ _4852_/CLK _4831_/D _3466_/Y vssd1 vssd1 vccd1 vccd1 _4831_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2704__A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4762_ _4803_/CLK _4762_/D fanout245/X vssd1 vssd1 vccd1 vccd1 _4762_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1974_ _4391_/Q _1974_/B vssd1 vssd1 vccd1 vccd1 _1974_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3713_ _3721_/A vssd1 vssd1 vccd1 vccd1 _3713_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_2616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_A
+ _4397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4693_ _3384_/Y _4693_/D _3675_/Y vssd1 vssd1 vccd1 vccd1 _4693_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_2638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3644_ _4195_/A vssd1 vssd1 vccd1 vccd1 _3644_/Y sky130_fd_sc_hd__inv_2
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
+ _4984_/Q _3122_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__3535__A _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_2021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2526_ _4679_/Q _2526_/B vssd1 vssd1 vccd1 vccd1 _4679_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__3254__B _3889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2457_ _2468_/A _4124_/B vssd1 vssd1 vccd1 vccd1 _2457_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4714__CLK _4717_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2388_ _4613_/Q _2388_/B vssd1 vssd1 vccd1 vccd1 _2388_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4127_ _4127_/A _4129_/B vssd1 vssd1 vccd1 vccd1 _4656_/D sky130_fd_sc_hd__xor2_1
XANTENNA__3270__A _3287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4058_ _4552_/Q vssd1 vssd1 vccd1 vccd1 _4553_/D sky130_fd_sc_hd__inv_2
XANTENNA__4864__CLK _4865_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3009_ _4953_/Q _4952_/Q _2988_/D _3006_/B vssd1 vssd1 vccd1 vccd1 _3010_/B sky130_fd_sc_hd__a31o_1
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_2516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2036__D _2036_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_GATE_N
+ _5063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_2148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_4119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3659_/A fanout240/X vssd1 vssd1 vccd1 vccd1 _5076_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_4_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2987__C _4954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3445__A _3445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4867__RESET_B fanout226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4394__CLK _4429_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2287__C_N _3900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3180__A _3904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_2059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3339__B _3420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_2925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_2936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1690_ _4918_/Q vssd1 vssd1 vccd1 vccd1 _4919_/D sky130_fd_sc_hd__inv_2
XANTENNA__3355__A _3361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3360_ _3903_/A _3420_/B vssd1 vssd1 vccd1 vccd1 _3360_/Y sky130_fd_sc_hd__xnor2_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2311_ _4580_/Q _4579_/Q _4578_/Q _2322_/B vssd1 vssd1 vccd1 vccd1 _2316_/B sky130_fd_sc_hd__or4_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _4564_/Q vssd1 vssd1 vccd1 vccd1 _3543_/B sky130_fd_sc_hd__buf_12
XFILLER_26_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5030_/CLK _5030_/D fanout224/X vssd1 vssd1 vccd1 vccd1 _5030_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2242_ _4527_/Q _2207_/D _2235_/B vssd1 vssd1 vccd1 vccd1 _2243_/B sky130_fd_sc_hd__a21bo_1
XFILLER_6_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4186__A _4189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2173_ _2858_/A vssd1 vssd1 vccd1 vccd1 _2173_/X sky130_fd_sc_hd__buf_6
XANTENNA__3090__A _3109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3776__115 _3776__115/A vssd1 vssd1 vccd1 vccd1 _3776__115/Y sky130_fd_sc_hd__inv_2
XFILLER_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_2825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4814_ _3449_/Y _4814_/D _3641_/Y vssd1 vssd1 vccd1 vccd1 _4814_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_3261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2434__A _2608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4267__CLK _3846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4745_ input21/X _4745_/D fanout222/X vssd1 vssd1 vccd1 vccd1 _4746_/D sky130_fd_sc_hd__dfrtp_1
X_1957_ _4384_/Q _4383_/Q vssd1 vssd1 vccd1 vccd1 _1957_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4676_ _4717_/CLK _4676_/D fanout253/X vssd1 vssd1 vccd1 vccd1 _4676_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout217_A fanout219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1888_ _4316_/Q _1888_/B vssd1 vssd1 vccd1 vccd1 _4316_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__3265__A _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4960__RESET_B fanout212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_4141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3558_ _4249_/A _4250_/A vssd1 vssd1 vccd1 vccd1 _3558_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_26_4091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_3699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2732__B1 _1975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4278__RESET_B fanout201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2509_ _2480_/D _2508_/X _2344_/X vssd1 vssd1 vccd1 vccd1 _2510_/B sky130_fd_sc_hd__o21ai_2
XFILLER_2_4027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3489_ _4065_/A _3543_/B vssd1 vssd1 vccd1 vccd1 _3489_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_22_3221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_2603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_2553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_2925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_2313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_TE_B
+ _2781_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_3361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2344__A _2858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_2671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_2693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3175__A _3917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_3215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2909__A_N _4894_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_2453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3903__A _3903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_2339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_3893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_3879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_2424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2254__A _4559_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_2446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2860_ _4863_/Q _2860_/B vssd1 vssd1 vccd1 vccd1 _4863_/D sky130_fd_sc_hd__xnor2_1
XFILLER_16_3581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_3445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1811_ _4281_/Q _1811_/B vssd1 vssd1 vccd1 vccd1 _1811_/X sky130_fd_sc_hd__and2b_1
X_2791_ _2791_/A vssd1 vssd1 vccd1 vccd1 _2791_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4530_ _4532_/CLK _4530_/D fanout211/X vssd1 vssd1 vccd1 vccd1 _4530_/Q sky130_fd_sc_hd__dfrtp_1
X_1742_ _5001_/Q vssd1 vssd1 vccd1 vccd1 _5002_/D sky130_fd_sc_hd__inv_2
XFILLER_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4461_ input26/X _4461_/D fanout199/X vssd1 vssd1 vccd1 vccd1 _4462_/D sky130_fd_sc_hd__dfrtp_4
X_3366__32 _3366__32/A vssd1 vssd1 vccd1 vccd1 _3366__32/Y sky130_fd_sc_hd__inv_2
X_1673_ _4887_/Q vssd1 vssd1 vccd1 vccd1 _4886_/D sky130_fd_sc_hd__inv_2
XANTENNA__3085__A _4991_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3412_ _3414_/A vssd1 vssd1 vccd1 vccd1 _3412_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_3828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4392_ _4402_/CLK _4392_/D fanout187/X vssd1 vssd1 vccd1 vccd1 _4392_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4371__RESET_B fanout214/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_2002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _3361_/A vssd1 vssd1 vccd1 vccd1 _3343_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _3947_/A _3438_/B vssd1 vssd1 vccd1 vccd1 _3274_/Y sky130_fd_sc_hd__xnor2_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5013_/CLK _5013_/D _3567_/Y vssd1 vssd1 vccd1 vccd1 _5013_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2225_ _4523_/Q _2225_/B vssd1 vssd1 vccd1 vccd1 _2226_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_2873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2429__A _2566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf _4276_/Q _1851_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_1_4093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2156_ _4488_/Q _4487_/Q _2135_/D _2153_/B vssd1 vssd1 vccd1 vccd1 _2157_/B sky130_fd_sc_hd__a31o_1
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2087_ _4466_/D _4440_/Q vssd1 vssd1 vccd1 vccd1 _2088_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout167_A _3865_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_2600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_2677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4902__CLK _4905_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2989_ _4948_/Q vssd1 vssd1 vccd1 vccd1 _3001_/A sky130_fd_sc_hd__inv_2
XFILLER_30_2822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_2221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4728_ _5013_/CLK _4728_/D _3404_/Y vssd1 vssd1 vccd1 vccd1 _4728_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_2276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
+ _4803_/Q _2779_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_4659_ _4659_/CLK _4659_/D fanout211/X vssd1 vssd1 vccd1 vccd1 _4659_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_3513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3723__A _4010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3442__B _3442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_3189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4432__CLK _5033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3530__53_A _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4582__CLK _4590_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_2154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_3249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_2515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_2537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_3023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_3067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3633__A _3642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_2125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_2294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_3725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3352__B _3440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
+ _4861_/Q _2879_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_23_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2010_ _1961_/C _2006_/Y _2003_/X vssd1 vssd1 vccd1 vccd1 _2011_/B sky130_fd_sc_hd__o21ai_1
XFILLER_18_3610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3961_ _4410_/Q vssd1 vssd1 vccd1 vccd1 _4409_/D sky130_fd_sc_hd__inv_2
XFILLER_17_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2912_ _4896_/Q _4895_/Q _2891_/D _2909_/B vssd1 vssd1 vccd1 vccd1 _2913_/B sky130_fd_sc_hd__a31o_1
XFILLER_16_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3892_ _3892_/A _3892_/B _3901_/B vssd1 vssd1 vccd1 vccd1 _3895_/B sky130_fd_sc_hd__or3_2
XFILLER_18_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1986__A1 _4395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2843_ _4858_/Q _2843_/B vssd1 vssd1 vccd1 vccd1 _4858_/D sky130_fd_sc_hd__xnor2_1
XFILLER_30_2107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_3275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__0641_ _3777_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0641_/X sky130_fd_sc_hd__clkbuf_16
X_2774_ _3112_/A _2774_/B _2774_/C _2774_/D vssd1 vssd1 vccd1 vccd1 _2775_/B sky130_fd_sc_hd__and4_1
XFILLER_34_1597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3527__B _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4513_ _3284_/Y _4513_/D _3724_/Y vssd1 vssd1 vccd1 vccd1 _4513_/Q sky130_fd_sc_hd__dfrtp_2
X_1725_ _4970_/Q vssd1 vssd1 vccd1 vccd1 _4969_/D sky130_fd_sc_hd__inv_2
XFILLER_12_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_3750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4305__CLK _3892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4444_ _3240_/Y _4444_/D _3746_/Y vssd1 vssd1 vccd1 vccd1 _4444_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_2014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_3888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4375_ _3598_/A _4375_/D fanout214/X vssd1 vssd1 vccd1 vccd1 _4375_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_2924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_4083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _3340_/A vssd1 vssd1 vccd1 vccd1 _3326_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4455__CLK _3899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_3371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
+ _4518_/Q _2273_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3257_ _5057_/A vssd1 vssd1 vccd1 vccd1 _3257_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_2731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_2742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2208_ _4524_/Q _4523_/Q _4522_/Q _2208_/D vssd1 vssd1 vccd1 vccd1 _2218_/C sky130_fd_sc_hd__and4_2
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3188_ _3885_/A _3886_/A vssd1 vssd1 vccd1 vccd1 _3188_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_6_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2139_ _4493_/Q _4492_/Q _4491_/Q _2176_/A vssd1 vssd1 vccd1 vccd1 _2162_/B sky130_fd_sc_hd__or4_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_4010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout157/X fanout203/X vssd1 vssd1 vccd1 vccd1 _5082_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_10_3905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_4076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3718__A _3721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2622__A _2622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_3260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3453__A _4127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_2592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_2517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2069__A _2178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4948__CLK _4962_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_2191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input12_A comp_high_Q[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1701__A _4248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_3816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
+ _4576_/Q _2371_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_31_3117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4328__CLK _4063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2532__A _2566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_2861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3187__71 _3189__72/A vssd1 vssd1 vccd1 vccd1 _3187__71/Y sky130_fd_sc_hd__inv_2
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2490_ _4671_/Q _4670_/Q _2490_/C vssd1 vssd1 vccd1 vccd1 _2490_/X sky130_fd_sc_hd__and3_1
XANTENNA_output80_A _5077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4478__CLK _1952_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3363__A _3696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4160_ _4701_/Q vssd1 vssd1 vccd1 vccd1 _4700_/D sky130_fd_sc_hd__inv_2
XFILLER_7_2163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_clk_master clkbuf_3_1_0_clk_master/A vssd1 vssd1 vccd1 vccd1 _4359_/CLK
+ sky130_fd_sc_hd__clkbuf_8
X_3111_ _5024_/D _4983_/Q vssd1 vssd1 vccd1 vccd1 _3112_/D sky130_fd_sc_hd__xnor2_1
XFILLER_7_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4091_ _4601_/Q vssd1 vssd1 vccd1 vccd1 _4602_/D sky130_fd_sc_hd__inv_2
X_3042_ _3112_/A _3042_/B _3042_/C _3042_/D vssd1 vssd1 vccd1 vccd1 _3043_/B sky130_fd_sc_hd__and4_1
XFILLER_3_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_4141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4993_ _5047_/A _4993_/D fanout242/X vssd1 vssd1 vccd1 vccd1 _4993_/Q sky130_fd_sc_hd__dfrtp_1
X_3944_ _4131_/B _3944_/B vssd1 vssd1 vccd1 vccd1 _3947_/B sky130_fd_sc_hd__nand2_2
XFILLER_14_2614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2081__B1 _2003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3875_ _3899_/A _3901_/A _3901_/B _3875_/D vssd1 vssd1 vccd1 vccd1 _3876_/A sky130_fd_sc_hd__or4_1
XANTENNA__3538__A _3550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2826_ _4856_/Q _2830_/B _2832_/A vssd1 vssd1 vccd1 vccd1 _2875_/C sky130_fd_sc_hd__o21ai_1
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__0624_ _3600_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0624_/X sky130_fd_sc_hd__clkbuf_16
X_2757_ _4808_/Q _4807_/Q _2760_/A vssd1 vssd1 vccd1 vccd1 _2757_/Y sky130_fd_sc_hd__nor3_1
XFILLER_25_4101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2384__A1 _4613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1708_ _4938_/Q _1709_/B vssd1 vssd1 vccd1 vccd1 _4937_/D sky130_fd_sc_hd__xnor2_1
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_3641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2688_ _2647_/D _2686_/Y _2687_/X vssd1 vssd1 vccd1 vccd1 _2689_/B sky130_fd_sc_hd__o21ai_1
XFILLER_25_3433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4427_ _4429_/CLK _4427_/D fanout194/X vssd1 vssd1 vccd1 vccd1 _4427_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_3527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3273__A _3287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4358_ _4359_/CLK _4358_/D fanout186/X vssd1 vssd1 vccd1 vccd1 _4358_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_5_2826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3884__A1 _3888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input4_A comp_high_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3309_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3309_/Y sky130_fd_sc_hd__inv_2
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _5040_/A _4289_/D fanout190/X vssd1 vssd1 vccd1 vccd1 _4289_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_3273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[4\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf _2790_/A _2642_/Y vssd1
+ vssd1 vccd1 vccd1 _5091_/A sky130_fd_sc_hd__ebufn_8
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3749_/A fanout187/X vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__dlrtn_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3653__83 _3655__85/A vssd1 vssd1 vccd1 vccd1 _3653__83/Y sky130_fd_sc_hd__inv_2
XFILLER_32_3437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_A
+ _4711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3448__A _3466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4620__CLK _4623_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_3219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4770__CLK _4812_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_2325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout120/X fanout249/X vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_20_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2527__A _4741_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__1637_ clkbuf_0__1637_/X vssd1 vssd1 vccd1 vccd1 _3201__9/A sky130_fd_sc_hd__clkbuf_16
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_2057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xnet199_2 _3600_/A vssd1 vssd1 vccd1 vccd1 _1935_/A sky130_fd_sc_hd__inv_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1990_ _2061_/A _1990_/B vssd1 vssd1 vccd1 vccd1 _1991_/B sky130_fd_sc_hd__nand2_1
XFILLER_14_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_2809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3358__A _3912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_GATE_N _5048_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2262__A _3066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3660_ _3669_/A vssd1 vssd1 vccd1 vccd1 _3660_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_2279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2611_ _4725_/Q _4724_/Q vssd1 vssd1 vccd1 vccd1 _2611_/Y sky130_fd_sc_hd__xnor2_2
X_3591_ _3597_/A vssd1 vssd1 vccd1 vccd1 _3591_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2542_ _4693_/Q _4692_/Q vssd1 vssd1 vccd1 vccd1 _2542_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_5_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4189__A _4189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2473_ _4661_/Q _4660_/Q vssd1 vssd1 vccd1 vccd1 _2473_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__3093__A _3109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2118__A1 _3892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4212_ _4786_/Q vssd1 vssd1 vccd1 vccd1 _4785_/D sky130_fd_sc_hd__inv_2
XFILLER_29_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_3869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4143_ _4666_/Q vssd1 vssd1 vccd1 vccd1 _4667_/D sky130_fd_sc_hd__inv_2
XANTENNA__1877__B1 _1823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4074_ _4570_/Q vssd1 vssd1 vccd1 vccd1 _4569_/D sky130_fd_sc_hd__inv_2
XFILLER_0_3457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3025_ _4958_/Q _4957_/Q _3028_/A vssd1 vssd1 vccd1 vccd1 _3025_/Y sky130_fd_sc_hd__nor3_1
XFILLER_3_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4985__RESET_B fanout234/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_2673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2841__A2 _4859_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout247_A fanout257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4976_ _3545_/Y _4976_/D _3591_/Y vssd1 vssd1 vccd1 vccd1 _4976_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4643__CLK _3861_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3927_ _4377_/Q vssd1 vssd1 vccd1 vccd1 _3933_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_14_3189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3268__A _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_2455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2172__A _4493_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3858_ _4370_/Q vssd1 vssd1 vccd1 vccd1 _3896_/A sky130_fd_sc_hd__buf_6
XFILLER_10_2319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2809_ _2809_/A1 _2802_/Y _3914_/B vssd1 vssd1 vccd1 vccd1 _2809_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_2780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3789_ _4271_/Q vssd1 vssd1 vccd1 vccd1 _4270_/D sky130_fd_sc_hd__inv_2
XANTENNA__4793__CLK _4943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_4014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout210 fanout213/X vssd1 vssd1 vccd1 vccd1 fanout210/X sky130_fd_sc_hd__buf_4
Xfanout221 input33/X vssd1 vssd1 vccd1 vccd1 fanout221/X sky130_fd_sc_hd__buf_4
XFILLER_5_2612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_3285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout232 fanout234/X vssd1 vssd1 vccd1 vccd1 fanout232/X sky130_fd_sc_hd__buf_4
Xfanout243 fanout245/X vssd1 vssd1 vccd1 vccd1 fanout243/X sky130_fd_sc_hd__buf_2
Xfanout254 fanout255/X vssd1 vssd1 vccd1 vccd1 fanout254/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_2645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3469__42 _3469__42/A vssd1 vssd1 vccd1 vccd1 _4843_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__3731__A _4010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_2509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_2448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_2391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_3201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3178__A _3912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3472__44_A _3528__52/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3906__A _3914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[6\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf_A _3128_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_2348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout128/X fanout246/X vssd1 vssd1 vccd1 vccd1 _5077_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_8_2280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3063__D _3085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4516__CLK _2294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3641__A _3642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3360__B _3420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4666__CLK _2470_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
+ _4395_/Q _2025_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_15_3421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4830_ _3465_/Y _4830_/D _3633_/Y vssd1 vssd1 vccd1 vccd1 _4830_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_4008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4761_ _4809_/CLK _4761_/D fanout254/X vssd1 vssd1 vccd1 vccd1 _4761_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1973_ _4392_/Q _4391_/Q _1973_/C vssd1 vssd1 vccd1 vccd1 _1973_/X sky130_fd_sc_hd__and3_1
XANTENNA__3088__A _4989_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3712_ _3721_/A vssd1 vssd1 vccd1 vccd1 _3712_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4692_ _5013_/CLK _4692_/D _3383_/Y vssd1 vssd1 vccd1 vccd1 _4692_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_18_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3643_ _3643_/A vssd1 vssd1 vccd1 vccd1 _4195_/A sky130_fd_sc_hd__buf_8
XFILLER_11_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_3837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3535__B _3556_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2525_ _2478_/C _2521_/Y _2518_/X vssd1 vssd1 vccd1 vccd1 _2526_/B sky130_fd_sc_hd__o21ai_1
XFILLER_6_3611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_4115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2456_ _2807_/A _3922_/A vssd1 vssd1 vccd1 vccd1 _2456_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_3414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1819__B1_N _1810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2387_ _4614_/Q _4613_/Q _2387_/C vssd1 vssd1 vccd1 vccd1 _2387_/X sky130_fd_sc_hd__and3_1
XFILLER_9_1387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3551__A _3924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout197_A fanout198/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4126_ _4126_/A _4248_/C vssd1 vssd1 vccd1 vccd1 _4129_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4057_ _4553_/Q vssd1 vssd1 vccd1 vccd1 _4552_/D sky130_fd_sc_hd__inv_2
XANTENNA__2167__A _2178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3008_ _4950_/Q _3008_/B vssd1 vssd1 vccd1 vccd1 _4950_/D sky130_fd_sc_hd__xnor2_1
XFILLER_24_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4959_ _4962_/CLK _4959_/D fanout212/X vssd1 vssd1 vccd1 vccd1 _4959_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_3852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_2285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3726__A _4010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_2602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_3071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_3007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3461__A _3934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_2370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4007__A1 _3935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_2617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_3086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_2374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3058__D _3058_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3636__A _3642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_2683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2310_ _4583_/Q _4582_/Q _4581_/Q _2333_/B vssd1 vssd1 vccd1 vccd1 _2322_/B sky130_fd_sc_hd__or4_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3290_/Y sky130_fd_sc_hd__inv_2
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ _4525_/Q _2241_/B vssd1 vssd1 vccd1 vccd1 _4525_/D sky130_fd_sc_hd__xnor2_1
XFILLER_22_2009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_3789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4577__RESET_B fanout226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2172_ _4493_/Q _4492_/Q _2176_/A vssd1 vssd1 vccd1 vccd1 _2172_/Y sky130_fd_sc_hd__nor3_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4186__B _4190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4813_ _4247_/Y _4813_/D _3448_/Y vssd1 vssd1 vccd1 vccd1 _4813_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_3885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_3273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1956_ _4382_/Q _4381_/Q vssd1 vssd1 vccd1 vccd1 _1956_/Y sky130_fd_sc_hd__xnor2_2
X_4744_ input21/X input5/X fanout229/X vssd1 vssd1 vccd1 vccd1 _4745_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_33_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_2583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4675_ _4717_/CLK _4675_/D fanout253/X vssd1 vssd1 vccd1 vccd1 _4675_/Q sky130_fd_sc_hd__dfrtp_4
X_1887_ _1858_/D _1886_/X _1823_/X vssd1 vssd1 vccd1 vccd1 _1888_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__3546__A _3550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3626_ _4256_/A vssd1 vssd1 vccd1 vccd1 _3626_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout112_A _3576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3265__B _3886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3557_ _3571_/A vssd1 vssd1 vccd1 vccd1 _3557_/Y sky130_fd_sc_hd__inv_2
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2508_ _4675_/Q _2508_/B vssd1 vssd1 vccd1 vccd1 _2508_/X sky130_fd_sc_hd__and2b_1
XFILLER_24_2808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3488_ _3498_/A vssd1 vssd1 vccd1 vccd1 _3488_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_4039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4831__CLK _4852_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2439_ _4636_/Q _4635_/Q vssd1 vssd1 vccd1 vccd1 _2439_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__3281__A _3287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_2795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4109_ _4635_/Q vssd1 vssd1 vccd1 vccd1 _4636_/D sky130_fd_sc_hd__inv_2
XFILLER_0_3051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5089_ _5089_/A vssd1 vssd1 vccd1 vccd1 _5089_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4981__CLK _4981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_2937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_2683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3456__A _3466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4361__CLK _4472_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2971__A1 _3929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2360__A _4648_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_2981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3175__B _3444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3903__B _3904_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1704__A _3556_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4670__RESET_B fanout242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_6_0_clk_master clkbuf_3_7_0_clk_master/A vssd1 vssd1 vccd1 vccd1 _4472_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_21_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2535__A _3066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_4114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_4136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3016__A_N _4954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2254__B _4533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_2458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_3593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1810_ _4282_/Q _1810_/B vssd1 vssd1 vccd1 vccd1 _1811_/B sky130_fd_sc_hd__nor2_1
XFILLER_15_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2790_ _2790_/A _2790_/B vssd1 vssd1 vccd1 vccd1 _2791_/A sky130_fd_sc_hd__or2_1
XFILLER_12_3457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4704__CLK _4718_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1741_ _5002_/Q vssd1 vssd1 vccd1 vccd1 _5001_/D sky130_fd_sc_hd__inv_2
XFILLER_15_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_3921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4460_ _3256_/Y _4460_/D _3737_/Y vssd1 vssd1 vccd1 vccd1 _4460_/Q sky130_fd_sc_hd__dfrtp_4
X_1672_ _4884_/Q vssd1 vssd1 vccd1 vccd1 _4885_/D sky130_fd_sc_hd__inv_2
XANTENNA__3085__B _3085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3411_ _3917_/A _3444_/B vssd1 vssd1 vccd1 vccd1 _3411_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_25_3807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4854__CLK _4865_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4391_ _4429_/CLK _4391_/D fanout194/X vssd1 vssd1 vccd1 vccd1 _4391_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_29_3998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3342_ _3696_/A vssd1 vssd1 vccd1 vccd1 _3361_/A sky130_fd_sc_hd__buf_6
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3273_ _3287_/A vssd1 vssd1 vccd1 vccd1 _3273_/Y sky130_fd_sc_hd__inv_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _3566_/Y _5012_/D _3580_/Y vssd1 vssd1 vccd1 vccd1 _5012_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _4520_/Q _2224_/B vssd1 vssd1 vccd1 vccd1 _4520_/D sky130_fd_sc_hd__xnor2_1
XFILLER_22_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4347__D _4347_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2155_ _4485_/Q _2155_/B vssd1 vssd1 vccd1 vccd1 _4485_/D sky130_fd_sc_hd__xnor2_1
XFILLER_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2086_ _4437_/Q _2086_/B vssd1 vssd1 vccd1 vccd1 _4437_/D sky130_fd_sc_hd__xnor2_1
XFILLER_1_2681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2650__B1 _2661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_3546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2988_ _4953_/Q _4952_/Q _4951_/Q _2988_/D vssd1 vssd1 vccd1 vccd1 _2998_/C sky130_fd_sc_hd__and4_1
XFILLER_17_1966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_2391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4727_ _3403_/Y _4727_/D _3665_/Y vssd1 vssd1 vccd1 vccd1 _4727_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1939_ _3892_/B _3899_/A _3901_/A _3845_/Y vssd1 vssd1 vccd1 vccd1 _1939_/X sky130_fd_sc_hd__o211a_1
XFILLER_30_2856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3276__A _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3708__93_A _3732__95/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4658_ _4658_/CLK _4658_/D fanout211/X vssd1 vssd1 vccd1 vccd1 _4658_/Q sky130_fd_sc_hd__dfrtp_1
X_3609_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3609_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_3525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4589_ _5043_/A _4589_/D fanout222/X vssd1 vssd1 vccd1 vccd1 _4589_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__3902__A0 _3898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3574__54_A _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4428__RESET_B fanout194/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_2456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_2745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3186__A _3891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2090__A _4466_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout144/X fanout215/X vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
+ _4961_/Q _3054_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3914__A _3914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_3737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3418__37 _3469__42/A vssd1 vssd1 vccd1 vccd1 _4752_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_3666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3960_ _4407_/Q vssd1 vssd1 vccd1 vccd1 _4408_/D sky130_fd_sc_hd__inv_2
XFILLER_1_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_2211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2911_ _4893_/Q _2911_/B vssd1 vssd1 vccd1 vccd1 _4893_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__2632__B1 _3898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3891_ _3891_/A _3891_/B vssd1 vssd1 vccd1 vccd1 _4366_/D sky130_fd_sc_hd__xnor2_1
XFILLER_31_3833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2842_ _2916_/A _2842_/B vssd1 vssd1 vccd1 vccd1 _2843_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_3877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__0640_ _3766_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0640_/X sky130_fd_sc_hd__clkbuf_16
X_2773_ _4838_/D _4797_/Q vssd1 vssd1 vccd1 vccd1 _2774_/D sky130_fd_sc_hd__xnor2_1
XFILLER_30_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1724_ _4967_/Q vssd1 vssd1 vccd1 vccd1 _4968_/D sky130_fd_sc_hd__inv_2
X_4512_ _3914_/A _4512_/D _3283_/Y vssd1 vssd1 vccd1 vccd1 _4512_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4443_ _4063_/C _4443_/D _3239_/Y vssd1 vssd1 vccd1 vccd1 _4443_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_3845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4374_ _4374_/CLK _4374_/D fanout208/X vssd1 vssd1 vccd1 vccd1 _4374_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_2059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3543__B _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ _4065_/A _3543_/B vssd1 vssd1 vccd1 vccd1 _3325_/Y sky130_fd_sc_hd__xnor2_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3885_/A _3886_/A vssd1 vssd1 vccd1 vccd1 _3256_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_23_3383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2207_ _4527_/Q _4526_/Q _4525_/Q _2207_/D vssd1 vssd1 vccd1 vccd1 _2208_/D sky130_fd_sc_hd__and4_1
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2138_ _4555_/D _4497_/Q _4495_/Q _4494_/Q vssd1 vssd1 vccd1 vccd1 _2176_/A sky130_fd_sc_hd__or4_2
XFILLER_3_2798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2175__A _4491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2069_ _2178_/A _2069_/B vssd1 vssd1 vccd1 vccd1 _2070_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_3154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_3619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_4044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_4055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_2339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2622__B _2622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_2030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_TE_B _1916_/Y vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_3272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3453__B _4129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_2220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__1653_ clkbuf_0__1653_/X vssd1 vssd1 vccd1 vccd1 _3528__52/A sky130_fd_sc_hd__clkbuf_16
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1701__B _4248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3423__40 _3425__41/A vssd1 vssd1 vccd1 vccd1 _3423__40/Y sky130_fd_sc_hd__inv_2
XFILLER_13_3541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout158/X fanout205/X vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_31_2406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3644__A _4195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_2357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_3979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output73_A _5070_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3110_ _4996_/Q _3110_/B vssd1 vssd1 vccd1 vccd1 _4996_/D sky130_fd_sc_hd__xnor2_1
XFILLER_24_3681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_2175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4090_ _4602_/Q vssd1 vssd1 vccd1 vccd1 _4601_/D sky130_fd_sc_hd__inv_2
XFILLER_7_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5063_/A fanout251/X vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__dlrtn_1
X_3041_ _5020_/D _4947_/Q vssd1 vssd1 vccd1 vccd1 _3042_/D sky130_fd_sc_hd__xnor2_1
XFILLER_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_2877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_3441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_4028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4992_ _4997_/CLK _4992_/D fanout237/X vssd1 vssd1 vccd1 vccd1 _4992_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_18_3485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3943_ _4131_/A _4131_/C vssd1 vssd1 vccd1 vccd1 _3944_/B sky130_fd_sc_hd__nor2_1
XFILLER_34_2030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3819__A _4333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2723__A _4838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3267__23_A _3365__31/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_3641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3874_ _3897_/A _3908_/A vssd1 vssd1 vccd1 vccd1 _3875_/D sky130_fd_sc_hd__nand2_4
XFILLER_12_3051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2825_ _4859_/Q _4858_/Q _4857_/Q _2837_/B vssd1 vssd1 vccd1 vccd1 _2830_/B sky130_fd_sc_hd__or4_1
XFILLER_31_2940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3179__68_A _3189__72/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0__0623_ _3598_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0623_/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__4773__RESET_B fanout253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2756_ _4805_/Q _2756_/B vssd1 vssd1 vccd1 vccd1 _4805_/D sky130_fd_sc_hd__xnor2_1
XFILLER_25_4113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1707_ _1705_/Y _4190_/B _2977_/A vssd1 vssd1 vccd1 vccd1 _1709_/B sky130_fd_sc_hd__mux2_1
X_2687_ _2858_/A vssd1 vssd1 vccd1 vccd1 _2687_/X sky130_fd_sc_hd__buf_8
XANTENNA__3554__A _3571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4426_ _5033_/A _4426_/D fanout197/X vssd1 vssd1 vccd1 vccd1 _4426_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_2700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3193__75 _3193__75/A vssd1 vssd1 vccd1 vccd1 _4357_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_3697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4357_ _4357_/CLK _4357_/D fanout186/X vssd1 vssd1 vccd1 vccd1 _4357_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3308_ _3895_/A _3372_/B vssd1 vssd1 vccd1 vccd1 _3308_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_25_2777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _4288_/CLK _4288_/D fanout199/X vssd1 vssd1 vccd1 vccd1 _4288_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_25_2788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3239_ _3255_/A vssd1 vssd1 vccd1 vccd1 _3239_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_2562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_3205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
+ _4707_/Q _2614_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3729__A _4010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_A
+ _4392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwrapper_cell_loop\[1\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf _2278_/A _2129_/Y vssd1
+ vssd1 vccd1 vccd1 _5091_/A sky130_fd_sc_hd__ebufn_8
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3464__A _3466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_3163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_3005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_3843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2808__A _3877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3629__81 _3655__85/A vssd1 vssd1 vccd1 vccd1 _3629__81/Y sky130_fd_sc_hd__inv_2
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3639__A _3642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_2069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_3961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3358__B _3446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4445__CLK _4063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2610_ _4723_/Q _4722_/Q vssd1 vssd1 vccd1 vccd1 _2610_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_13_2670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3590_ _3597_/A vssd1 vssd1 vccd1 vccd1 _3590_/Y sky130_fd_sc_hd__inv_2
X_2541_ _4691_/Q _4690_/Q vssd1 vssd1 vccd1 vccd1 _2541_/Y sky130_fd_sc_hd__xnor2_2
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
+ _4765_/Q _2711_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__4595__CLK _4916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_2143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2472_ _4003_/C _2472_/B vssd1 vssd1 vccd1 vccd1 _5067_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__4189__B _4190_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout119/X fanout248/X vssd1 vssd1 vccd1 vccd1 _5078_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_6_3837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2118__A2 _3875_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4211_ _4783_/Q vssd1 vssd1 vccd1 vccd1 _4784_/D sky130_fd_sc_hd__inv_2
XFILLER_25_2029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_4021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4142_ _4667_/Q vssd1 vssd1 vccd1 vccd1 _4666_/D sky130_fd_sc_hd__inv_2
XFILLER_4_3550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4073_ _4567_/Q vssd1 vssd1 vccd1 vccd1 _4568_/D sky130_fd_sc_hd__inv_2
XFILLER_0_2713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_3386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3024_ _4955_/Q _3024_/B vssd1 vssd1 vccd1 vccd1 _4955_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_2724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4975_ _2809_/A1 _4975_/D _3544_/Y vssd1 vssd1 vccd1 vccd1 _4975_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3549__A _3934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_2412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3926_ _4378_/Q vssd1 vssd1 vccd1 vccd1 _3934_/A sky130_fd_sc_hd__buf_8
XFILLER_20_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout142_A _2285_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3268__B _3886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2172__B _4492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3857_ _3909_/A vssd1 vssd1 vccd1 vccd1 _3857_/Y sky130_fd_sc_hd__clkinv_2
X_2808_ _3877_/A _4063_/B _4063_/C _4064_/A vssd1 vssd1 vccd1 vccd1 _2808_/X sky130_fd_sc_hd__or4_1
X_3788_ _4268_/Q vssd1 vssd1 vccd1 vccd1 _4269_/D sky130_fd_sc_hd__inv_2
XFILLER_31_2792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2739_ _2730_/C _2738_/X _2687_/X vssd1 vssd1 vccd1 vccd1 _2740_/B sky130_fd_sc_hd__o21ai_2
XFILLER_27_3529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3284__A _3903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_2806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_4026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_4037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3166__64 _3169__65/A vssd1 vssd1 vccd1 vccd1 _3166__64/Y sky130_fd_sc_hd__inv_2
XFILLER_27_2839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout200 fanout221/X vssd1 vssd1 vccd1 vccd1 fanout200/X sky130_fd_sc_hd__clkbuf_2
X_4409_ _4063_/B _4409_/D _3219_/Y vssd1 vssd1 vccd1 vccd1 _4409_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_3106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout211 fanout212/X vssd1 vssd1 vccd1 vccd1 fanout211/X sky130_fd_sc_hd__buf_4
Xfanout222 fanout223/X vssd1 vssd1 vccd1 vccd1 fanout222/X sky130_fd_sc_hd__clkbuf_4
Xfanout233 fanout234/X vssd1 vssd1 vccd1 vccd1 fanout233/X sky130_fd_sc_hd__buf_2
XFILLER_5_3358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_2624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout244 fanout245/X vssd1 vssd1 vccd1 vccd1 fanout244/X sky130_fd_sc_hd__buf_2
Xfanout255 fanout256/X vssd1 vssd1 vccd1 vccd1 fanout255/X sky130_fd_sc_hd__clkbuf_4
XFILLER_28_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4318__CLK _4324_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4468__CLK input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_3213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_3956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3459__A _3946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2363__A _2608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3178__B _3446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4624__RESET_B fanout236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_2821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3906__B _3908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3194__A _3470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_2305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_3695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_3709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_4112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_TE_B
+ _2025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4760_ _3426_/Y _4760_/D _3653__83/Y vssd1 vssd1 vccd1 vccd1 _4760_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1972_ _4389_/Q _1972_/B vssd1 vssd1 vccd1 vccd1 _4389_/D sky130_fd_sc_hd__xor2_1
XFILLER_15_2743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3088__B _3088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3711_ _5058_/A vssd1 vssd1 vccd1 vccd1 _3721_/A sky130_fd_sc_hd__buf_6
XFILLER_31_2033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4691_ _3382_/Y _4691_/D _3676_/Y vssd1 vssd1 vccd1 vccd1 _4691_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3642_ _3642_/A vssd1 vssd1 vccd1 vccd1 _3642_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3573_ _3576_/A vssd1 vssd1 vccd1 vccd1 _3573_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_3849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2524_ _4678_/Q _2524_/B vssd1 vssd1 vccd1 vccd1 _4678_/D sky130_fd_sc_hd__xnor2_1
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_GATE_N _5056_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2455_ _3658_/Y _3684_/Y vssd1 vssd1 vccd1 vccd1 _2455_/Y sky130_fd_sc_hd__nor2_2
XFILLER_6_2900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_3426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2386_ _4611_/Q _2386_/B vssd1 vssd1 vccd1 vccd1 _4611_/D sky130_fd_sc_hd__xor2_1
XANTENNA__3551__B _3923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2511__A2 _4676_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4125_ _4125_/A vssd1 vssd1 vccd1 vccd1 _4248_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4056_ _4550_/Q vssd1 vssd1 vccd1 vccd1 _4551_/D sky130_fd_sc_hd__inv_2
XFILLER_0_3277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_2460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3007_ _2998_/C _3006_/X _2858_/X vssd1 vssd1 vccd1 vccd1 _3008_/B sky130_fd_sc_hd__o21ai_1
XFILLER_20_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3279__A _3287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2183__A _4555_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4958_ _4958_/CLK _4958_/D fanout218/X vssd1 vssd1 vccd1 vccd1 _4958_/Q sky130_fd_sc_hd__dfrtp_2
X_3909_ _3909_/A vssd1 vssd1 vccd1 vccd1 _3910_/A sky130_fd_sc_hd__buf_2
X_4889_ _3499_/Y _4889_/D _3616_/Y vssd1 vssd1 vccd1 vccd1 _4889_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_4027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__1638_ _3205_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__1638_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_2614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3742__A _3748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwrapper_cell_loop\[3\].w1.ro_block_I.ro_pol.tribuf.t_buf _2628_/X _2475_/Y vssd1
+ vssd1 vccd1 vccd1 _5088_/A sky130_fd_sc_hd__ebufn_8
XFILLER_5_3188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3461__B _3933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2358__A _2412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_2476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_GATE_N
+ fanout128/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4290__CLK _4063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
+ _4526_/Q _2265_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4805__RESET_B fanout253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2805__B _2805_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_2629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_2175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2093__A _2608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _4359_/CLK fanout193/X vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__dlrtn_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_4075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3917__A _3917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3369__33_A _3469__42/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_2113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3652__A _4195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ _2327_/A _2240_/B vssd1 vssd1 vccd1 vccd1 _2241_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4633__CLK _5013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2171_ _4490_/Q _2171_/B vssd1 vssd1 vccd1 vccd1 _4490_/D sky130_fd_sc_hd__xnor2_1
XFILLER_1_3553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_3481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1900__A _1909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4783__CLK _1765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4812_ _4812_/CLK _4812_/D fanout252/X vssd1 vssd1 vccd1 vccd1 _4812_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_3241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_3717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_3285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4743_ input29/X _4743_/D fanout212/X vssd1 vssd1 vccd1 vccd1 _4743_/Q sky130_fd_sc_hd__dfrtp_1
X_1955_ _3931_/A _1955_/B vssd1 vssd1 vccd1 vccd1 _5064_/A sky130_fd_sc_hd__xnor2_4
XFILLER_11_3149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2731__A _4799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4674_ _4709_/CLK _4674_/D fanout247/X vssd1 vssd1 vccd1 vccd1 _4674_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1886_ _4317_/Q _1886_/B vssd1 vssd1 vccd1 vccd1 _1886_/X sky130_fd_sc_hd__and2b_1
XANTENNA__3185__70_A _3189__72/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3625_ _4256_/A vssd1 vssd1 vccd1 vccd1 _3625_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_3613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_3635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout105_A _3135_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3556_ _3556_/A _3556_/B vssd1 vssd1 vccd1 vccd1 _3556_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2507_ _4676_/Q _2507_/B vssd1 vssd1 vccd1 vccd1 _2508_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3320__29_A _3365__31/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3487_ _4127_/A _4129_/A vssd1 vssd1 vccd1 vccd1 _3487_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_2978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3562__A _4127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2438_ _4634_/Q _4633_/Q vssd1 vssd1 vccd1 vccd1 _2438_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_9_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_3245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2178__A _2178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_2544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2369_ _4602_/Q _4601_/Q vssd1 vssd1 vccd1 vccd1 _2369_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_5_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4108_ _4636_/Q vssd1 vssd1 vccd1 vccd1 _4635_/D sky130_fd_sc_hd__clkinv_2
XFILLER_2_1915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5088_ _5088_/A vssd1 vssd1 vccd1 vccd1 _5088_/X sky130_fd_sc_hd__buf_4
XFILLER_0_3063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2906__A _2916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4039_ _4535_/Q vssd1 vssd1 vccd1 vccd1 _4534_/D sky130_fd_sc_hd__inv_2
XFILLER_25_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4287__RESET_B fanout195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_2949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_3341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3737__A _5057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4506__CLK _3932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2971__A2 _4063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_3134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_2400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2184__B1 _2173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4656__CLK _3598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_1_0_w0.cclk_I clkbuf_0_w0.cclk_I/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_w0.cclk_I/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_27_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_2308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2487__A1 _4670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2088__A _2178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2239__A1 _4527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2816__A _4927_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_3837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_3469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3647__A _4195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_2893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2551__A _4710_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1740_ _4999_/Q vssd1 vssd1 vccd1 vccd1 _5000_/D sky130_fd_sc_hd__inv_2
XFILLER_11_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout136/X fanout238/X vssd1 vssd1 vccd1 vccd1 _5084_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__2411__A1 _4620_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1671_ _4885_/Q vssd1 vssd1 vccd1 vccd1 _4884_/D sky130_fd_sc_hd__inv_2
XANTENNA__3599__1_A _3470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3410_ _3414_/A vssd1 vssd1 vccd1 vccd1 _3410_/Y sky130_fd_sc_hd__inv_2
X_4390_ _4429_/CLK _4390_/D fanout194/X vssd1 vssd1 vccd1 vccd1 _4390_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_3977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3911__A1 _3914_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3341_ _3895_/A _3372_/B vssd1 vssd1 vccd1 vccd1 _3341_/Y sky130_fd_sc_hd__xnor2_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3382__A _4004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _4004_/A _3491_/B vssd1 vssd1 vccd1 vccd1 _3272_/Y sky130_fd_sc_hd__xnor2_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _2809_/A1 _5011_/D _3565_/Y vssd1 vssd1 vccd1 vccd1 _5011_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _2327_/A _2223_/B vssd1 vssd1 vccd1 vccd1 _2224_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4798__RESET_B fanout245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2154_ _2145_/C _2153_/X _2003_/X vssd1 vssd1 vccd1 vccd1 _2155_/B sky130_fd_sc_hd__o21ai_1
XFILLER_3_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2085_ _2083_/X _2084_/Y _2003_/X vssd1 vssd1 vccd1 vccd1 _2086_/B sky130_fd_sc_hd__o21ai_1
XFILLER_17_3303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4380__RESET_B fanout210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4529__CLK _4532_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2650__A1 _4764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_2657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_3525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2987_ _4956_/Q _4955_/Q _4954_/Q _2987_/D vssd1 vssd1 vccd1 vccd1 _2988_/D sky130_fd_sc_hd__and4_1
XFILLER_15_3093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3557__A _3571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout222_A fanout223/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2461__A _2631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_2835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4726_ _4916_/CLK _4726_/D _3402_/Y vssd1 vssd1 vccd1 vccd1 _4726_/Q sky130_fd_sc_hd__dfrtp_1
X_1938_ _1936_/X _1937_/Y _3845_/Y _1952_/A1 vssd1 vssd1 vccd1 vccd1 _1938_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_28_4100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3276__B _3440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4679__CLK _4719_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4657_ _4657_/CLK _4657_/D fanout222/X vssd1 vssd1 vccd1 vccd1 _4657_/Q sky130_fd_sc_hd__dfrtp_4
X_1869_ _4312_/Q _1869_/B vssd1 vssd1 vccd1 vccd1 _1869_/Y sky130_fd_sc_hd__nor2_1
X_3608_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3608_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_3443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4588_ _4590_/CLK _4588_/D fanout229/X vssd1 vssd1 vccd1 vccd1 _4588_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_8_3537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3539_ _4189_/A _4190_/A vssd1 vssd1 vccd1 vccd1 _3539_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_28_3498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1805__A _3114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3292__A _4065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_2560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2469__A1 _2631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2469__B2 _2468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_2374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_2713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_A
+ _4674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_2724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_2757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3467__A _3905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3186__B _3889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2090__B _4425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3914__B _3914_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_2241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_3946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_3705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_2368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4891__RESET_B fanout236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_4070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2910_ _2901_/C _2909_/X _2858_/X vssd1 vssd1 vccd1 vccd1 _2911_/B sky130_fd_sc_hd__o21ai_1
XFILLER_16_4081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3684_/A fanout216/X vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__2632__A1 _3914_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3890_ _4366_/Q vssd1 vssd1 vccd1 vccd1 _3891_/A sky130_fd_sc_hd__clkbuf_16
X_2841_ _4860_/Q _4859_/Q _2819_/D _2838_/B vssd1 vssd1 vccd1 vccd1 _2842_/B sky130_fd_sc_hd__a31o_1
XFILLER_31_3845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3197__5 _3199__7/A vssd1 vssd1 vccd1 vccd1 _4364_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4821__CLK _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3377__A _3393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_3889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2772_ _4810_/Q _2772_/B vssd1 vssd1 vccd1 vccd1 _4810_/D sky130_fd_sc_hd__xnor2_1
XFILLER_12_3277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2396__B1 _2344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4511_ _3282_/Y _4511_/D _3725_/Y vssd1 vssd1 vccd1 vccd1 _4511_/Q sky130_fd_sc_hd__dfrtp_2
X_1723_ _4968_/Q vssd1 vssd1 vccd1 vccd1 _4967_/D sky130_fd_sc_hd__inv_2
XFILLER_12_1831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4442_ _3238_/Y _4442_/D _3747_/Y vssd1 vssd1 vccd1 vccd1 _4442_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4971__CLK _4248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4373_ _4472_/CLK _4373_/D fanout204/X vssd1 vssd1 vccd1 vccd1 _4373_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4001__A _4001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3324_ _3340_/A vssd1 vssd1 vccd1 vccd1 _3324_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_2937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3255_/A vssd1 vssd1 vccd1 vccd1 _3255_/Y sky130_fd_sc_hd__inv_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ _4529_/Q _4528_/Q _2206_/C vssd1 vssd1 vccd1 vccd1 _2207_/D sky130_fd_sc_hd__and3_1
XFILLER_3_3489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3186_ _3891_/A _3889_/A vssd1 vssd1 vccd1 vccd1 _3186_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_23_1971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2137_ _4485_/Q _4484_/Q _2145_/C _2148_/A vssd1 vssd1 vccd1 vccd1 _2191_/B sky130_fd_sc_hd__a31o_1
XANTENNA__2456__A _2807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout172_A _3892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4351__CLK input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2068_ _4434_/Q _4433_/Q _2035_/D _2064_/B vssd1 vssd1 vccd1 vccd1 _2069_/B sky130_fd_sc_hd__a31o_1
XANTENNA__2175__B _2175_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_2421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_3311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3287__A _3287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2191__A _3066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4709_ _4709_/CLK _4709_/D fanout247/X vssd1 vssd1 vccd1 vccd1 _4709_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf_TE_B
+ _2546_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3735__97 _3759__99/A vssd1 vssd1 vccd1 vccd1 _3735__97/Y sky130_fd_sc_hd__inv_2
XANTENNA__4649__RESET_B fanout208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3006__A_N _4951_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_2458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3750__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1701__C _4248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4844__CLK _5030_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_2229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4994__CLK _5047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3925__A _3925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_2419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_3947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_3513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3660__A _3669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_3557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3040_ _4960_/Q _3040_/B vssd1 vssd1 vccd1 vccd1 _4960_/D sky130_fd_sc_hd__xnor2_1
XFILLER_7_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4991_ _5047_/A _4991_/D fanout242/X vssd1 vssd1 vccd1 vccd1 _4991_/Q sky130_fd_sc_hd__dfrtp_4
X_3942_ _4124_/C vssd1 vssd1 vccd1 vccd1 _4131_/C sky130_fd_sc_hd__buf_2
XFILLER_18_2741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3873_ _3883_/A _3883_/B _3882_/A vssd1 vssd1 vccd1 vccd1 _3901_/B sky130_fd_sc_hd__nand3_4
XFILLER_20_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2824_ _4862_/Q _4861_/Q _4860_/Q _2847_/B vssd1 vssd1 vccd1 vccd1 _2837_/B sky130_fd_sc_hd__or4_1
XFILLER_12_3063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_2362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2755_ _2771_/A _2755_/B vssd1 vssd1 vccd1 vccd1 _2756_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1706_ _4938_/Q _4937_/Q vssd1 vssd1 vccd1 vccd1 _2977_/A sky130_fd_sc_hd__xnor2_4
XFILLER_25_4125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2686_ _4772_/Q _4771_/Q _2690_/A vssd1 vssd1 vccd1 vccd1 _2686_/Y sky130_fd_sc_hd__nor3_1
X_4425_ _5033_/A _4425_/D fanout195/X vssd1 vssd1 vccd1 vccd1 _4425_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_3654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_3582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_2942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4717__CLK _4717_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4742__RESET_B fanout212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4356_ _4356_/CLK _4356_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _4356_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3307_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3307_/Y sky130_fd_sc_hd__inv_2
X_4287_ _4288_/CLK _4287_/D fanout195/X vssd1 vssd1 vccd1 vccd1 _4287_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3570__A _3934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _4004_/A _3491_/B vssd1 vssd1 vccd1 vccd1 _3238_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4867__CLK _4905_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_2574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2186__A _2922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_2505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2914__A _4894_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_2126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_3737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_2159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3745__A _3748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4397__CLK _4402_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_3092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4483__RESET_B fanout202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_2211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_2255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3480__A _5062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_3877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2808__B _4063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_2037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5022__CLK input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_2215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3012__A1 _4953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf _4311_/Q _1922_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
X_2540_ _4689_/Q _4688_/Q vssd1 vssd1 vccd1 vccd1 _2540_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_26_3722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2471_ _3900_/A _2459_/Y _2801_/C _2470_/X _3929_/A vssd1 vssd1 vccd1 vccd1 _2472_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_5_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_2238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4210_ _4784_/Q vssd1 vssd1 vccd1 vccd1 _4783_/D sky130_fd_sc_hd__inv_2
XFILLER_25_2008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4141_ _4664_/Q vssd1 vssd1 vccd1 vccd1 _4665_/D sky130_fd_sc_hd__inv_2
XANTENNA__3390__A _3917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_TE_B
+ _2539_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3079__A1 _4989_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4072_ _4568_/Q vssd1 vssd1 vccd1 vccd1 _4567_/D sky130_fd_sc_hd__inv_2
XFILLER_23_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3023_ _3030_/A _3023_/B vssd1 vssd1 vccd1 vccd1 _3024_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_2883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_2686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4974_ _3543_/Y _4974_/D _3592_/Y vssd1 vssd1 vccd1 vccd1 _4974_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3549__B _3933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3925_ _3925_/A _3925_/B vssd1 vssd1 vccd1 vccd1 _4376_/D sky130_fd_sc_hd__xor2_1
XFILLER_18_2593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[5\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf_A _2962_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3856_ _4368_/Q _4367_/Q vssd1 vssd1 vccd1 vccd1 _3909_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__2172__C _2176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout135_A _3375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2807_ _2807_/A _2807_/B vssd1 vssd1 vccd1 vccd1 _2807_/X sky130_fd_sc_hd__or2_1
XANTENNA__4994__RESET_B fanout239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3787_ _4269_/Q vssd1 vssd1 vccd1 vccd1 _4268_/D sky130_fd_sc_hd__clkinv_2
XANTENNA__3565__A _3571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_2192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2738_ _4801_/Q _2738_/B vssd1 vssd1 vccd1 vccd1 _2738_/X sky130_fd_sc_hd__and2b_1
Xclkbuf_2_0_0_clk_master clkbuf_2_1_0_clk_master/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_clk_master/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_29_4080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3284__B _3420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2669_ _4767_/Q _4766_/Q _2648_/D _2666_/B vssd1 vssd1 vccd1 vccd1 _2670_/B sky130_fd_sc_hd__a31o_1
XFILLER_5_4049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_3473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4408_ _3218_/Y _4408_/D _3757_/Y vssd1 vssd1 vccd1 vccd1 _4408_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_2750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout201 fanout202/X vssd1 vssd1 vccd1 vccd1 fanout201/X sky130_fd_sc_hd__buf_4
XANTENNA__2569__A_N _4708_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout212 fanout213/X vssd1 vssd1 vccd1 vccd1 fanout212/X sky130_fd_sc_hd__buf_4
Xfanout223 fanout230/X vssd1 vssd1 vccd1 vccd1 fanout223/X sky130_fd_sc_hd__buf_2
XFILLER_21_3118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4339_ _3184_/Y _4339_/D _3767__106/Y vssd1 vssd1 vccd1 vccd1 _4339_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout234 fanout235/X vssd1 vssd1 vccd1 vccd1 fanout234/X sky130_fd_sc_hd__buf_4
Xfanout245 fanout247/X vssd1 vssd1 vccd1 vccd1 fanout245/X sky130_fd_sc_hd__buf_2
XFILLER_25_2564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_2406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_2575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout256 fanout257/X vssd1 vssd1 vccd1 vccd1 fanout256/X sky130_fd_sc_hd__clkbuf_4
XFILLER_25_1863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_2371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5029__RESET_B fanout223/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3459__B _3945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_2502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3475__A _3905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
+ _4896_/Q _2951_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_30_2281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_2113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_3641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_3882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout180/X fanout184/X vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_1_3757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_4124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2554__A _4745_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1971_ _2143_/A _2020_/B _2020_/C vssd1 vssd1 vccd1 vccd1 _1972_/B sky130_fd_sc_hd__and3_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _5058_/A vssd1 vssd1 vccd1 vccd1 _3710_/Y sky130_fd_sc_hd__inv_4
XFILLER_35_2181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_3781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4690_ _4916_/CLK _4690_/D _3381_/Y vssd1 vssd1 vccd1 vccd1 _4690_/Q sky130_fd_sc_hd__dfrtp_2
X_3641_ _3642_/A vssd1 vssd1 vccd1 vccd1 _3641_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_3191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_2799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3385__A _3393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3572_ _3924_/A _3923_/A vssd1 vssd1 vccd1 vccd1 _3572_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_6_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2523_ _2566_/A _2523_/B vssd1 vssd1 vccd1 vccd1 _2524_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_4117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_3613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_2046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2454_ _2454_/A vssd1 vssd1 vccd1 vccd1 _2454_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_3405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_3596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2385_ _2996_/A _2432_/B _2432_/C vssd1 vssd1 vccd1 vccd1 _2386_/B sky130_fd_sc_hd__and3_1
XFILLER_22_2715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4124_ _4131_/A _4124_/B _4124_/C _4124_/D vssd1 vssd1 vccd1 vccd1 _4125_/A sky130_fd_sc_hd__or4_1
XFILLER_22_2737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
+ _4954_/Q _3046_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_20_3162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput1 comp_high_I[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4055_ _4551_/Q vssd1 vssd1 vccd1 vccd1 _4550_/D sky130_fd_sc_hd__inv_2
X_3006_ _4951_/Q _3006_/B vssd1 vssd1 vccd1 vccd1 _3006_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_3289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2464__A _3875_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout252_A fanout253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4905__CLK _4905_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_90 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2183__B _4497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4957_ _4958_/CLK _4957_/D fanout218/X vssd1 vssd1 vccd1 vccd1 _4957_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_2855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3908_ _3908_/A vssd1 vssd1 vccd1 vccd1 _3914_/B sky130_fd_sc_hd__buf_4
X_4888_ _4943_/CLK _4888_/D _3498_/Y vssd1 vssd1 vccd1 vccd1 _4888_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_32_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_3280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_3865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3839_ _3839_/A _3883_/B vssd1 vssd1 vccd1 vccd1 _4356_/D sky130_fd_sc_hd__xnor2_1
XFILLER_14_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3295__A _3309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1808__A _3114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0__1637_ _3194_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__1637_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_27_3305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_2626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0_w0.cclk_I clkbuf_0_w0.cclk_I/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_w0.cclk_I/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_5_3134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3199__7_A _3199__7/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
+ _4611_/Q _2443_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_25_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4435__CLK _5033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2374__A _4652_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4585__CLK _4623_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1718__A _4945_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3933__A _3933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2170_ _2178_/A _2170_/B vssd1 vssd1 vccd1 vccd1 _2171_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_3471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_2842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4928__CLK input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_A
+ _4988_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2284__A _2284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4811_ _4811_/CLK _4811_/D fanout250/X vssd1 vssd1 vccd1 vccd1 _4811_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
+ _4669_/Q _2545_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4742_ input29/X _4742_/D fanout212/X vssd1 vssd1 vccd1 vccd1 _4743_/D sky130_fd_sc_hd__dfrtp_1
X_1954_ _3865_/Y _1951_/X _1953_/X _2287_/A _1938_/Y vssd1 vssd1 vccd1 vccd1 _1955_/B
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4586__RESET_B fanout231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_2574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4673_ _4718_/CLK _4673_/D fanout239/X vssd1 vssd1 vccd1 vccd1 _4673_/Q sky130_fd_sc_hd__dfrtp_4
X_1885_ _4318_/Q _1885_/B vssd1 vssd1 vccd1 vccd1 _1886_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4308__CLK _3845_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3624_ _4256_/A vssd1 vssd1 vccd1 vccd1 _3624_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_3603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4004__A _4004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3555_ _3571_/A vssd1 vssd1 vccd1 vccd1 _3555_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_4050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3526__51 _3528__52/A vssd1 vssd1 vccd1 vccd1 _3526__51/Y sky130_fd_sc_hd__inv_2
X_2506_ _4673_/Q _2506_/B vssd1 vssd1 vccd1 vccd1 _4673_/D sky130_fd_sc_hd__xnor2_1
XFILLER_26_4083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3486_ _3498_/A vssd1 vssd1 vccd1 vccd1 _3486_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1940__A1 _3882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3562__B _4129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_3382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2459__A _2464_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2437_ _4632_/Q _4631_/Q vssd1 vssd1 vccd1 vccd1 _2437_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_22_2501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3142__B1 _2468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2368_ _4600_/Q _4599_/Q vssd1 vssd1 vccd1 vccd1 _2368_/Y sky130_fd_sc_hd__xnor2_2
X_4107_ _4633_/Q vssd1 vssd1 vccd1 vccd1 _4634_/D sky130_fd_sc_hd__inv_2
XFILLER_22_1833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5087_ _5087_/A vssd1 vssd1 vccd1 vccd1 _5087_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2299_ _4570_/Q _4569_/Q vssd1 vssd1 vccd1 vccd1 _2299_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_22_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4038_ _4516_/Q vssd1 vssd1 vccd1 vccd1 _4517_/D sky130_fd_sc_hd__inv_2
XFILLER_0_3097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1810__B _1810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_4065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_4098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_3353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_3938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_2630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_2641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2922__A _2922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[4\].w1.ro_block_I.ro_pol_eve.tribuf.t_buf _2795_/A _2644_/Y vssd1
+ vssd1 vccd1 vccd1 _5089_/A sky130_fd_sc_hd__ebufn_8
XANTENNA__3753__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_2423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_3909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_2011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2487__A2 _2491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_2033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input28_A phi1b_dig_Q[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2239__A2 _4526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_2405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3928__A _3934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_3415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_2714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_2151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2551__B _4709_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1670_ _4882_/Q vssd1 vssd1 vccd1 vccd1 _4883_/D sky130_fd_sc_hd__inv_2
XANTENNA_output96_A _5093_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3663__A _3669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3340_ _3340_/A vssd1 vssd1 vccd1 vccd1 _3340_/Y sky130_fd_sc_hd__inv_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3382__B _3491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3287_/A vssd1 vssd1 vccd1 vccd1 _3271_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3207__14_A _3264__22/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _3564_/Y _5010_/D _3581_/Y vssd1 vssd1 vccd1 vccd1 _5010_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_6_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _4521_/Q _2218_/C _2219_/B vssd1 vssd1 vccd1 vccd1 _2223_/B sky130_fd_sc_hd__a21bo_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3528__52_A _3528__52/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2153_ _4486_/Q _2153_/B vssd1 vssd1 vccd1 vccd1 _2153_/X sky130_fd_sc_hd__and2b_1
XFILLER_3_2959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_4096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1911__A _4351_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2084_ _4466_/D _4440_/Q _4438_/Q vssd1 vssd1 vccd1 vccd1 _2084_/Y sky130_fd_sc_hd__nor3_1
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3375_/A fanout240/X vssd1 vssd1 vccd1 vccd1 _5076_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1989__A1 _4395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2650__A2 _4763_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_TE_B
+ _2614_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_GATE_N
+ _5063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_2669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2986_ _4958_/Q _4957_/Q _2986_/C vssd1 vssd1 vccd1 vccd1 _2987_/D sky130_fd_sc_hd__and3_1
XFILLER_34_2983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4725_ _3401_/Y _4725_/D _3666_/Y vssd1 vssd1 vccd1 vccd1 _4725_/Q sky130_fd_sc_hd__dfrtp_1
X_1937_ _3892_/B _3910_/A vssd1 vssd1 vccd1 vccd1 _1937_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__2461__B _3877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4656_ _3598_/A _4656_/D fanout225/X vssd1 vssd1 vccd1 vccd1 _4656_/Q sky130_fd_sc_hd__dfrtp_4
X_1868_ _4313_/Q _4312_/Q _1868_/C vssd1 vssd1 vccd1 vccd1 _1868_/X sky130_fd_sc_hd__and3_1
XFILLER_28_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3607_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3607_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4280__CLK _4281_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4587_ _4590_/CLK _4587_/D fanout227/X vssd1 vssd1 vccd1 vccd1 _4587_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2166__A1 _4491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3573__A _3576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1799_ _4279_/Q _1799_/B vssd1 vssd1 vccd1 vccd1 _1800_/B sky130_fd_sc_hd__nor2_1
XFILLER_28_3455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3538_ _3550_/A vssd1 vssd1 vccd1 vccd1 _3538_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_2826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3292__B _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_3043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2469__A2 _3908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_2572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2917__A _4895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_2397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4437__RESET_B fanout198/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3748__A _3748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_2769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_3161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3467__B _3913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_2471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4623__CLK _4623_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3483__A _4249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4773__CLK _4812_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
+ _4430_/Q _2097_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__3106__B1 _1791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2827__A _2996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_3613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4860__RESET_B fanout226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3658__A _5060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2840_ _4857_/Q _2840_/B vssd1 vssd1 vccd1 vccd1 _4857_/D sky130_fd_sc_hd__xnor2_1
XFILLER_31_3857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_3245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2771_ _2771_/A _2771_/B vssd1 vssd1 vccd1 vccd1 _2772_/B sky130_fd_sc_hd__nand2_1
X_4510_ _2286_/B _4510_/D _3281_/Y vssd1 vssd1 vccd1 vccd1 _4510_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_34_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1722_ _4965_/Q vssd1 vssd1 vccd1 vccd1 _4966_/D sky130_fd_sc_hd__inv_2
XFILLER_12_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_2566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4441_ _2809_/A1 _4441_/D _3236_/Y vssd1 vssd1 vccd1 vccd1 _4441_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_29_3753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_2006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3393__A _3393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4372_ _4372_/CLK _4372_/D fanout214/X vssd1 vssd1 vccd1 vccd1 _4372_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_3639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_4114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ _3340_/A vssd1 vssd1 vccd1 vccd1 _3323_/Y sky130_fd_sc_hd__inv_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_4086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3254_ _3891_/A _3889_/A vssd1 vssd1 vccd1 vccd1 _3254_/Y sky130_fd_sc_hd__xnor2_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _4559_/D _4533_/Q _4531_/Q _4530_/Q vssd1 vssd1 vccd1 vccd1 _2206_/C sky130_fd_sc_hd__and4_1
XFILLER_23_2673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4948__RESET_B fanout208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_2767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2136_ _4483_/Q vssd1 vssd1 vccd1 vccd1 _2148_/A sky130_fd_sc_hd__inv_2
XFILLER_23_1994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2067_ _3112_/A vssd1 vssd1 vccd1 vccd1 _2178_/A sky130_fd_sc_hd__buf_4
XFILLER_1_2491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout165_A _3869_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
+ _4488_/Q _2196_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_30_4002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3568__A _3946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2472__A _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_4068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2969_ _3576_/Y _3605_/Y vssd1 vssd1 vccd1 vccd1 _2969_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_2021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_2190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_3389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4708_ _4712_/CLK _4708_/D fanout247/X vssd1 vssd1 vccd1 vccd1 _4708_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4796__CLK _3446_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_4003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_4036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4639_ _4943_/CLK _4639_/D _3355_/Y vssd1 vssd1 vccd1 vccd1 _4639_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_4058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_2601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_2573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1701__D _4187_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2075__B1 _2003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4271__RESET_B _5048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2382__A _4619_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3925__B _3925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1726__A _4969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3941__A _3941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4519__CLK _4532_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2557__A _4709_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_2824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4359__RESET_B fanout195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4669__CLK _4718_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4990_ _4997_/CLK _4990_/D fanout236/X vssd1 vssd1 vccd1 vccd1 _4990_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_3919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3941_ _3941_/A _3941_/B vssd1 vssd1 vccd1 vccd1 _4124_/C sky130_fd_sc_hd__nand2_1
XANTENNA__3388__A _3925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_2753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_A
+ _4488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2292__A _4068_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3872_ _3888_/A _3872_/B vssd1 vssd1 vccd1 vccd1 _3901_/A sky130_fd_sc_hd__nand2_2
XFILLER_31_3632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_2628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2823_ _4865_/Q _4864_/Q _4863_/Q _2861_/A vssd1 vssd1 vccd1 vccd1 _2847_/B sky130_fd_sc_hd__or4_1
XFILLER_31_3665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2754_ _4806_/Q _2719_/D _2747_/B vssd1 vssd1 vccd1 vccd1 _2755_/B sky130_fd_sc_hd__a21bo_1
XFILLER_31_2975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1705_ _4248_/A _4248_/C vssd1 vssd1 vccd1 vccd1 _1705_/Y sky130_fd_sc_hd__nor2_1
X_2685_ _4769_/Q _2685_/B vssd1 vssd1 vccd1 vccd1 _4769_/D sky130_fd_sc_hd__xnor2_1
XFILLER_25_4137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4424_ _3234_/Y _4424_/D _3748_/Y vssd1 vssd1 vccd1 vccd1 _4424_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_3414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4355_ _4359_/CLK _4355_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _4355_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3851__A _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3306_ _3903_/A _3420_/B vssd1 vssd1 vccd1 vccd1 _3306_/Y sky130_fd_sc_hd__xnor2_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _5040_/A _4286_/D fanout194/X vssd1 vssd1 vccd1 vccd1 _4286_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3570__B _3933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _4005_/A vssd1 vssd1 vccd1 vccd1 _3491_/B sky130_fd_sc_hd__buf_12
XFILLER_23_3193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_2481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3168_ _3935_/A _3440_/B vssd1 vssd1 vccd1 vccd1 _3168_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4711__RESET_B fanout245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2119_ _3910_/A _3941_/A _3900_/A _3900_/B _3908_/A vssd1 vssd1 vccd1 vccd1 _2119_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3099_ _3098_/Y _3056_/C _4994_/Q vssd1 vssd1 vccd1 vccd1 _3100_/B sky130_fd_sc_hd__mux2_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3298__A _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2498__A_N _4672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_2252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_2452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_2486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_2245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4811__CLK _4811_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_2339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4068__S _4068_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_3889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2808__C _4063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input10_A comp_high_Q[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4961__CLK _4962_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2048__B1 _1975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2824__B _4861_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4742__D _4742_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_4041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_3941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_3985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_2227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3012__A2 _2988_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2220__B1 _1975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2470_ _2470_/A1 _2469_/X _2465_/X vssd1 vssd1 vccd1 vccd1 _2470_/X sky130_fd_sc_hd__o21a_1
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_4001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_2189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3671__A _4135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_4034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4140_ _4665_/Q vssd1 vssd1 vccd1 vccd1 _4664_/D sky130_fd_sc_hd__inv_2
XFILLER_22_2908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout157/X fanout204/X vssd1 vssd1 vccd1 vccd1 _5082_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_0_4117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_4045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3390__B _3444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4491__CLK _5042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4071_ _4071_/A vssd1 vssd1 vccd1 vccd1 _4562_/D sky130_fd_sc_hd__inv_2
XFILLER_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3079__A2 _4988_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3022_ _4956_/Q _2987_/D _3015_/B vssd1 vssd1 vccd1 vccd1 _3023_/B sky130_fd_sc_hd__a21bo_1
XFILLER_23_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4973_ _4248_/A _4973_/D _3542_/Y vssd1 vssd1 vccd1 vccd1 _4973_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4652__D _4652_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3924_ _3924_/A vssd1 vssd1 vccd1 vccd1 _3925_/A sky130_fd_sc_hd__buf_12
XFILLER_18_2572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3855_ _3892_/B vssd1 vssd1 vccd1 vccd1 _3855_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_31_3473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3846__A _3846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2806_ _3941_/B _2809_/A1 _2462_/Y _2457_/Y _4003_/C vssd1 vssd1 vccd1 vccd1 _2807_/B
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_0__1653_ _3470_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__1653_/X sky130_fd_sc_hd__clkbuf_16
X_3786_ _4266_/Q vssd1 vssd1 vccd1 vccd1 _4267_/D sky130_fd_sc_hd__inv_2
XANTENNA_fanout128_A _3632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_2171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2737_ _4802_/Q _2737_/B vssd1 vssd1 vccd1 vccd1 _2738_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_3441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2668_ _4764_/Q _2668_/B vssd1 vssd1 vccd1 vccd1 _4764_/D sky130_fd_sc_hd__xnor2_1
XFILLER_29_3391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4834__CLK input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4407_ _4063_/C _4407_/D _3217_/Y vssd1 vssd1 vccd1 vccd1 _4407_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_RESET_B fanout193/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3581__A _3587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_2510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2599_ _4745_/D _4719_/Q _4717_/Q vssd1 vssd1 vccd1 vccd1 _2599_/Y sky130_fd_sc_hd__nor3_1
XFILLER_25_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout202 fanout220/X vssd1 vssd1 vccd1 vccd1 fanout202/X sky130_fd_sc_hd__buf_4
XFILLER_25_2532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout213 fanout220/X vssd1 vssd1 vccd1 vccd1 fanout213/X sky130_fd_sc_hd__clkbuf_2
Xfanout224 fanout230/X vssd1 vssd1 vccd1 vccd1 fanout224/X sky130_fd_sc_hd__clkbuf_4
Xfanout235 input33/X vssd1 vssd1 vccd1 vccd1 fanout235/X sky130_fd_sc_hd__clkbuf_4
X_4338_ _3899_/A _4338_/D _3182__69/Y vssd1 vssd1 vccd1 vccd1 _4338_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout246 fanout247/X vssd1 vssd1 vccd1 vccd1 fanout246/X sky130_fd_sc_hd__buf_2
XFILLER_25_1820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input2_A comp_high_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout257 input33/X vssd1 vssd1 vccd1 vccd1 fanout257/X sky130_fd_sc_hd__clkbuf_4
X_4269_ _3846_/A _4269_/D _4359_/CLK vssd1 vssd1 vccd1 vccd1 _4269_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_1853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4984__CLK _4997_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2925__A _4897_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3756__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3421__39_A _3425__41/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3475__B _3913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_GATE_N _5056_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_2318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_3918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3491__A _4001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2819__B _4859_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_2042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_2294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_3697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2835__A _2916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_4136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_3582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1970_ _4391_/Q _1974_/B _1977_/A vssd1 vssd1 vccd1 vccd1 _2020_/C sky130_fd_sc_hd__o21ai_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4707__CLK _4718_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3666__A _3669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_3793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3640_ _3642_/A vssd1 vssd1 vccd1 vccd1 _3640_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3571_ _3571_/A vssd1 vssd1 vccd1 vccd1 _3571_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4857__CLK _4865_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3749_/A fanout187/X vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__dlrtn_1
X_2522_ _2521_/Y _2478_/C _4679_/Q vssd1 vssd1 vccd1 vccd1 _2523_/B sky130_fd_sc_hd__mux2_1
XFILLER_6_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_2014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_4129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2453_ _2453_/A _2453_/B vssd1 vssd1 vccd1 vccd1 _2454_/A sky130_fd_sc_hd__or2_1
XFILLER_6_3625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1914__A _2608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2384_ _4613_/Q _2388_/B _2390_/A vssd1 vssd1 vccd1 vccd1 _2432_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__4374__RESET_B fanout208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_2874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4647__D _4647_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4123_ _4123_/A _4123_/B vssd1 vssd1 vccd1 vccd1 _4124_/D sky130_fd_sc_hd__nand2_1
XFILLER_20_3141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput2 comp_high_I[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_2
X_4054_ _4548_/Q vssd1 vssd1 vccd1 vccd1 _4549_/D sky130_fd_sc_hd__clkinv_2
XFILLER_0_3246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_3174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3005_ _4952_/Q _3005_/B vssd1 vssd1 vccd1 vccd1 _3006_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_2484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2464__B _3941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_80 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_91 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_2801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4387__CLK _3845_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4956_ _4958_/CLK _4956_/D fanout218/X vssd1 vssd1 vccd1 vccd1 _4956_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout245_A fanout247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3907_ _3907_/A vssd1 vssd1 vccd1 vccd1 _3907_/Y sky130_fd_sc_hd__inv_2
X_4887_ _3497_/Y _4887_/D _3618_/Y vssd1 vssd1 vccd1 vccd1 _4887_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3576__A _3576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_2255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2480__A _4674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3838_ _3838_/A _3883_/B vssd1 vssd1 vccd1 vccd1 _4355_/D sky130_fd_sc_hd__xnor2_1
XFILLER_31_3292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout120/X fanout249/X vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_10_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2499__B1 _2344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_2581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3209__15 _3264__22/A vssd1 vssd1 vccd1 vccd1 _3209__15/Y sky130_fd_sc_hd__inv_2
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_3001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_2322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3486__A _3498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_2366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3933__B _3935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4810_ _4812_/CLK _4810_/D fanout251/X vssd1 vssd1 vccd1 vccd1 _4810_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4741_ input29/X _4741_/D fanout210/X vssd1 vssd1 vccd1 vccd1 _4742_/D sky130_fd_sc_hd__dfrtp_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1953_ _1948_/Y _1952_/Y _3845_/Y vssd1 vssd1 vccd1 vccd1 _1953_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3396__A _3414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1909__A _1909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4930__D input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4672_ _4718_/CLK _4672_/D fanout239/X vssd1 vssd1 vccd1 vccd1 _4672_/Q sky130_fd_sc_hd__dfrtp_4
X_1884_ _4315_/Q _1884_/B vssd1 vssd1 vccd1 vccd1 _4315_/D sky130_fd_sc_hd__xnor2_1
X_3369__33 _3469__42/A vssd1 vssd1 vccd1 vccd1 _3369__33/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3623_ _4256_/A vssd1 vssd1 vccd1 vccd1 _3623_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3554_ _3571_/A vssd1 vssd1 vccd1 vccd1 _3554_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4555__RESET_B fanout202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2505_ _2566_/A _2505_/B vssd1 vssd1 vccd1 vccd1 _2506_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_3411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3485_ _4189_/A _4190_/A vssd1 vssd1 vccd1 vccd1 _3485_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__1940__A2 _1952_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2436_ _4630_/Q _4629_/Q vssd1 vssd1 vccd1 vccd1 _2436_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_29_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_2732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3142__A1 _4064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_2671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_2682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2367_ _4598_/Q _4597_/Q vssd1 vssd1 vccd1 vccd1 _2367_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_6_3499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_3269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout195_A fanout196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4106_ _4634_/Q vssd1 vssd1 vccd1 vccd1 _4633_/D sky130_fd_sc_hd__inv_2
X_5086_ _5086_/A vssd1 vssd1 vccd1 vccd1 _5086_/X sky130_fd_sc_hd__clkbuf_2
X_2298_ _4568_/Q _4567_/Q vssd1 vssd1 vccd1 vccd1 _2298_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_22_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4037_ _4517_/Q vssd1 vssd1 vccd1 vccd1 _4516_/D sky130_fd_sc_hd__inv_2
XFILLER_25_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_4055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_4077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3632_/A fanout246/X vssd1 vssd1 vccd1 vccd1 _5077_/A sky130_fd_sc_hd__dlrtn_1
X_4939_ _4943_/CLK _4939_/D _3524__50/Y vssd1 vssd1 vccd1 vccd1 _4939_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_2085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_2973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_2995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf _4288_/Q _1854_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4402__CLK _4402_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_2518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_2170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4552__CLK _2294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_2297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[1\].w1.ro_block_I.ro_pol_eve.tribuf.t_buf _2283_/A _2131_/Y vssd1
+ vssd1 vccd1 vccd1 _5089_/A sky130_fd_sc_hd__ebufn_8
XFILLER_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2385__A _2996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
+ _4800_/Q _2782_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_12_4117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_3552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3928__B _3933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_3427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2551__C _4708_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3944__A _4131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output89_A _5086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3782__123 _3784__125/A vssd1 vssd1 vccd1 vccd1 _3782__123/Y sky130_fd_sc_hd__inv_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ _3287_/A vssd1 vssd1 vccd1 vccd1 _3270_/Y sky130_fd_sc_hd__inv_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _2221_/A _2221_/B vssd1 vssd1 vccd1 vccd1 _4519_/D sky130_fd_sc_hd__xnor2_1
XFILLER_3_3639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_4031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_2855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2152_ _4487_/Q _2152_/B vssd1 vssd1 vccd1 vccd1 _2153_/B sky130_fd_sc_hd__nor2_1
XFILLER_26_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2083_ _4466_/D _4440_/Q _4438_/Q vssd1 vssd1 vccd1 vccd1 _2083_/X sky130_fd_sc_hd__and3_1
XFILLER_35_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_3663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2650__A3 _2658_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3838__B _3883_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2985_ _5020_/D _4962_/Q _4960_/Q _4959_/Q vssd1 vssd1 vccd1 vccd1 _2986_/C sky130_fd_sc_hd__and4_1
XFILLER_21_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4660__D _4660_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_2973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4724_ _1765_/A _4724_/D _3400_/Y vssd1 vssd1 vccd1 vccd1 _4724_/Q sky130_fd_sc_hd__dfrtp_1
X_1936_ _3872_/B _3910_/A vssd1 vssd1 vccd1 vccd1 _1936_/X sky130_fd_sc_hd__or2_1
XANTENNA__4425__CLK _5033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4655_ _3363_/Y _4655_/D fanout229/X vssd1 vssd1 vccd1 vccd1 _4655_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1867_ _4310_/Q _1867_/B vssd1 vssd1 vccd1 vccd1 _4310_/D sky130_fd_sc_hd__xor2_1
X_3606_ _5062_/A vssd1 vssd1 vccd1 vccd1 _3616_/A sky130_fd_sc_hd__buf_6
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
+ _4858_/Q _2882_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_1798_ _4276_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _4276_/D sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout208_A fanout220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4586_ _4623_/CLK _4586_/D fanout231/X vssd1 vssd1 vccd1 vccd1 _4586_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_28_3445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_2805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3537_ _4249_/A _4250_/A vssd1 vssd1 vccd1 vccd1 _3537_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_2733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3523__49_A _3523__49/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4575__CLK _4590_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3468_ _5061_/A vssd1 vssd1 vccd1 vccd1 _3468_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2419_ _2418_/Y _2375_/C _4622_/Q vssd1 vssd1 vccd1 vccd1 _2420_/B sky130_fd_sc_hd__mux2_1
X_3399_ _4127_/A _4129_/A vssd1 vssd1 vccd1 vccd1 _3399_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_24_1929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1821__B _1821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4835__D _4835_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_4117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5069_ _5069_/A vssd1 vssd1 vccd1 vccd1 _5069_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_3883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3776__115_A _3776__115/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3202__10 _3201__9/A vssd1 vssd1 vccd1 vccd1 _4374_/CLK sky130_fd_sc_hd__inv_2
XFILLER_33_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4918__CLK _5013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_2519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_2792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3483__B _4250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_2221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_2265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2865__B1 _2858_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4745__D _4745_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_2982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_2935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_4094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2770_ _4838_/D _4812_/Q vssd1 vssd1 vccd1 vccd1 _2771_/B sky130_fd_sc_hd__xnor2_1
XFILLER_12_2534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_2545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1721_ _4966_/Q vssd1 vssd1 vccd1 vccd1 _4965_/D sky130_fd_sc_hd__inv_2
XFILLER_11_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3674__A _4135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_2589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4440_ _5033_/A _4440_/D fanout198/X vssd1 vssd1 vccd1 vccd1 _4440_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_3743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4371_ _3598_/A _4371_/D fanout214/X vssd1 vssd1 vccd1 vccd1 _4371_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_4043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _3696_/A vssd1 vssd1 vccd1 vccd1 _3340_/A sky130_fd_sc_hd__buf_6
XFILLER_3_4126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3255_/A vssd1 vssd1 vccd1 vccd1 _3253_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2204_ _2858_/A vssd1 vssd1 vccd1 vccd1 _2996_/A sky130_fd_sc_hd__buf_12
X_3184_ _3895_/A _3372_/B vssd1 vssd1 vccd1 vccd1 _3184_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_26_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_2685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2135_ _4488_/Q _4487_/Q _4486_/Q _2135_/D vssd1 vssd1 vccd1 vccd1 _2145_/C sky130_fd_sc_hd__and4_1
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_3193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2066_ _4431_/Q _2066_/B vssd1 vssd1 vccd1 vccd1 _4431_/D sky130_fd_sc_hd__xnor2_1
XFILLER_1_2481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4988__RESET_B fanout235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout158_A _5058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3568__B _3945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3680__87 _3683__90/A vssd1 vssd1 vccd1 vccd1 _3680__87/Y sky130_fd_sc_hd__inv_2
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2968_ _2968_/A vssd1 vssd1 vccd1 vccd1 _2968_/X sky130_fd_sc_hd__clkbuf_1
X_4707_ _4718_/CLK _4707_/D fanout247/X vssd1 vssd1 vccd1 vccd1 _4707_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1919_ _4335_/Q _4334_/Q vssd1 vssd1 vccd1 vccd1 _1919_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__2277__A_N _4556_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2899_ _2996_/A _2946_/B _2946_/C vssd1 vssd1 vccd1 vccd1 _2900_/B sky130_fd_sc_hd__and3_1
XANTENNA__3584__A _3587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf_TE_B
+ _2715_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_4015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4638_ _3354_/Y _4638_/D _3689_/Y vssd1 vssd1 vccd1 vccd1 _4638_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4569_ _3855_/Y _4569_/D _3316__27/Y vssd1 vssd1 vccd1 vccd1 _4569_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_2646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1832__A _4347_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2663__A _2680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3772__111 _3776__115/A vssd1 vssd1 vccd1 vccd1 _3772__111/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2382__B _4618_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_2589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4740__CLK input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3494__A _3498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_3905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4890__CLK _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_3949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3941__B _3941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_2145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_2095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2557__B _4708_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3669__A _3669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
+ _4619_/Q _2435_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3940_ _3940_/A vssd1 vssd1 vccd1 vccd1 _3941_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__3388__B _3442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_2765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3871_ _3941_/A vssd1 vssd1 vccd1 vccd1 _3877_/A sky130_fd_sc_hd__buf_4
XFILLER_31_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2822_ _4927_/D _4869_/Q _4867_/Q _4866_/Q vssd1 vssd1 vccd1 vccd1 _2861_/A sky130_fd_sc_hd__or4_2
XFILLER_31_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_3043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_2320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2753_ _4804_/Q _2753_/B vssd1 vssd1 vccd1 vccd1 _4804_/D sky130_fd_sc_hd__xnor2_1
XFILLER_12_2375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1704_ _3556_/B _1704_/B vssd1 vssd1 vccd1 vccd1 _4936_/D sky130_fd_sc_hd__xor2_1
XFILLER_9_3601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2684_ _2771_/A _2684_/B vssd1 vssd1 vccd1 vccd1 _2685_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_3623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4423_ _1952_/A1 _4423_/D _3233_/Y vssd1 vssd1 vccd1 vccd1 _4423_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_3645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_3426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_4070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_4081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4354_ _4354_/CLK _4354_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _4354_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_2966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_2725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3851__B _3886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3305_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3305_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_3380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4285_ _4288_/CLK _4285_/D fanout194/X vssd1 vssd1 vccd1 vccd1 _4285_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_3222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_2769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _3255_/A vssd1 vssd1 vccd1 vccd1 _3236_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_2471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4613__CLK _4623_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3167_ _3933_/A vssd1 vssd1 vccd1 vccd1 _3440_/B sky130_fd_sc_hd__buf_12
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5059_/A fanout215/X vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__dlrtn_1
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2118_ _3892_/B _3875_/D _3888_/A vssd1 vssd1 vccd1 vccd1 _2118_/X sky130_fd_sc_hd__o21a_1
X_3098_ _3098_/A vssd1 vssd1 vccd1 vccd1 _3098_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3579__A _3587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2057__A1 _4431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2483__A _4741_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2049_ _2049_/A _2049_/B vssd1 vssd1 vccd1 vccd1 _4426_/D sky130_fd_sc_hd__xnor2_1
XFILLER_23_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4751__RESET_B fanout223/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4763__CLK _4803_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3298__B _3440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_2264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_2431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_2486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3318__28 _3365__31/A vssd1 vssd1 vccd1 vccd1 _3318__28/Y sky130_fd_sc_hd__inv_2
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2658__A _4764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4293__CLK _3929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2808__D _4064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2296__A1 _3877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[4\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf_A _2790_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3489__A _4065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2393__A _4613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_2239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_TE_B
+ _2708_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_4024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2568__A _4709_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[5\].w1.ro_block_Q.ro_pol.tribuf.t_buf_A _2963_/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4070_ _4565_/Q _4070_/B vssd1 vssd1 vccd1 vccd1 _4566_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_3417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2287__B _3931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3079__A3 _3058_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3021_ _4954_/Q _3021_/B vssd1 vssd1 vccd1 vccd1 _4954_/D sky130_fd_sc_hd__xnor2_1
XFILLER_4_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_A
+ _4951_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_2655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3399__A _4127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4972_ _3541_/Y _4972_/D _3593_/Y vssd1 vssd1 vccd1 vccd1 _4972_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_3105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3923_ _3923_/A _3925_/B vssd1 vssd1 vccd1 vccd1 _4375_/D sky130_fd_sc_hd__xor2_1
XFILLER_14_2404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_3441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3854_ _3872_/B vssd1 vssd1 vccd1 vccd1 _3892_/B sky130_fd_sc_hd__buf_4
XFILLER_31_3452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3846__B _3883_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2805_ _4251_/Y _2805_/B vssd1 vssd1 vccd1 vccd1 _5097_/A sky130_fd_sc_hd__xnor2_1
XFILLER_34_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3785_ _4267_/Q vssd1 vssd1 vccd1 vccd1 _4266_/D sky130_fd_sc_hd__clkinv_2
XFILLER_30_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2736_ _4799_/Q _2736_/B vssd1 vssd1 vccd1 vccd1 _4799_/D sky130_fd_sc_hd__xnor2_1
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2667_ _2658_/C _2666_/X _2518_/X vssd1 vssd1 vccd1 vccd1 _2668_/B sky130_fd_sc_hd__o21ai_1
XFILLER_9_3453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4406_ _4064_/A _4406_/D _3758_/Y vssd1 vssd1 vccd1 vccd1 _4406_/Q sky130_fd_sc_hd__dfrtp_4
X_2598_ _4745_/D _4719_/Q _4717_/Q vssd1 vssd1 vccd1 vccd1 _2598_/X sky130_fd_sc_hd__and3_1
XFILLER_5_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout203 fanout204/X vssd1 vssd1 vccd1 vccd1 fanout203/X sky130_fd_sc_hd__buf_2
XFILLER_9_2763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout214 fanout219/X vssd1 vssd1 vccd1 vccd1 fanout214/X sky130_fd_sc_hd__buf_4
X_4337_ _3181_/Y _4337_/D _3768__107/Y vssd1 vssd1 vccd1 vccd1 _4337_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_8_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout225 fanout230/X vssd1 vssd1 vccd1 vccd1 fanout225/X sky130_fd_sc_hd__buf_2
Xfanout236 fanout257/X vssd1 vssd1 vccd1 vccd1 fanout236/X sky130_fd_sc_hd__buf_4
Xfanout247 fanout257/X vssd1 vssd1 vccd1 vccd1 fanout247/X sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
+ _4392_/Q _2028_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_5_2638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4268_ _3149_/Y _4268_/D _4359_/CLK vssd1 vssd1 vccd1 vccd1 _4268_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_3052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_3085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3219_ _3233_/A vssd1 vssd1 vccd1 vccd1 _3219_/Y sky130_fd_sc_hd__inv_2
X_4199_ _4755_/Q vssd1 vssd1 vccd1 vccd1 _4756_/D sky130_fd_sc_hd__inv_2
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_3049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5063_/A fanout252/X vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_32_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3491__B _3491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2388__A _4613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_2021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4673__RESET_B fanout239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3947__A _3947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_2757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_2014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3570_ _3934_/A _3933_/A vssd1 vssd1 vccd1 vccd1 _3570_/Y sky130_fd_sc_hd__xnor2_1
X_2521_ _2521_/A vssd1 vssd1 vccd1 vccd1 _2521_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1952__B1 _3900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2452_ _4653_/D _4654_/Q vssd1 vssd1 vccd1 vccd1 _2453_/B sky130_fd_sc_hd__and2b_1
XFILLER_6_3637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_4051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2383_ _4616_/Q _4615_/Q _4614_/Q _2394_/B vssd1 vssd1 vccd1 vccd1 _2388_/B sky130_fd_sc_hd__or4_1
XFILLER_4_4073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4122_ _4656_/Q vssd1 vssd1 vccd1 vccd1 _4127_/A sky130_fd_sc_hd__buf_12
XFILLER_22_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4053_ _4549_/Q vssd1 vssd1 vccd1 vccd1 _4548_/D sky130_fd_sc_hd__inv_2
Xinput3 comp_high_I[2] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_3186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3004_ _4949_/Q _3004_/B vssd1 vssd1 vccd1 vccd1 _4949_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_2546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2464__C _2464_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_81 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_92 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4955_ _4958_/CLK _4955_/D fanout218/X vssd1 vssd1 vccd1 vccd1 _4955_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_2813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3906_ _3914_/A _3908_/A vssd1 vssd1 vccd1 vccd1 _3907_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout140_A _2285_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_2223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4886_ _4981_/CLK _4886_/D _3496_/Y vssd1 vssd1 vccd1 vccd1 _4886_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_2857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout238_A fanout239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3837_ _4357_/Q _4358_/Q vssd1 vssd1 vccd1 vccd1 _3883_/B sky130_fd_sc_hd__xor2_4
XFILLER_14_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_3889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_4008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_4019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2719_ _4806_/Q _4805_/Q _4804_/Q _2719_/D vssd1 vssd1 vccd1 vccd1 _2720_/D sky130_fd_sc_hd__and4_1
XFILLER_27_3329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3592__A _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3699_ _4071_/A vssd1 vssd1 vccd1 vccd1 _3699_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4951__CLK _4962_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4838__D _4838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2499__A1 _2490_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_3941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2001__A _4397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1840__A _4347_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_2170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4331__CLK _3171_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout119/X fanout248/X vssd1 vssd1 vccd1 vccd1 _5078_/A sky130_fd_sc_hd__dlrtn_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_3068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_2919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_3491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4481__CLK _3268_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3318__28_A _3365__31/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_2105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4854__RESET_B fanout228/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2846__A _4859_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_2980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2662__A1 _4764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4824__CLK _3459_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3677__A _4135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4740_ input29/X _4740_/D fanout224/X vssd1 vssd1 vccd1 vccd1 _4741_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_15_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1952_ _1952_/A1 _3892_/B _3900_/A vssd1 vssd1 vccd1 vccd1 _1952_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_15_2543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4671_ _4709_/CLK _4671_/D fanout241/X vssd1 vssd1 vccd1 vccd1 _4671_/Q sky130_fd_sc_hd__dfrtp_4
X_1883_ _1909_/A _1883_/B vssd1 vssd1 vccd1 vccd1 _1884_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3622_ _4256_/A vssd1 vssd1 vccd1 vccd1 _3622_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3553_ _3588_/A vssd1 vssd1 vccd1 vccd1 _3571_/A sky130_fd_sc_hd__buf_6
XFILLER_26_4030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_2904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_4113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2504_ _4674_/Q _2480_/D _2497_/B vssd1 vssd1 vccd1 vccd1 _2505_/B sky130_fd_sc_hd__a21bo_1
X_3484_ _3498_/A vssd1 vssd1 vccd1 vccd1 _3484_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_3445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2435_ _4628_/Q _4627_/Q vssd1 vssd1 vccd1 vccd1 _2435_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_9_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3142__A2 _4188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2366_ _4596_/Q _4595_/Q vssd1 vssd1 vccd1 vccd1 _2366_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__4524__RESET_B fanout202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4105_ _4631_/Q vssd1 vssd1 vccd1 vccd1 _4632_/D sky130_fd_sc_hd__inv_2
X_5085_ _5085_/A vssd1 vssd1 vccd1 vccd1 _5085_/X sky130_fd_sc_hd__clkbuf_4
X_2297_ _3929_/A _2297_/B vssd1 vssd1 vccd1 vccd1 _5066_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout188_A fanout196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4036_ _4514_/Q vssd1 vssd1 vccd1 vccd1 _4515_/D sky130_fd_sc_hd__inv_2
XFILLER_25_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3587__A _3587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2491__A _4670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_2621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4938_ _4938_/CLK _4938_/D fanout217/X vssd1 vssd1 vccd1 vccd1 _4938_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4869_ _4905_/CLK _4869_/D fanout226/X vssd1 vssd1 vccd1 vccd1 _4869_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_2075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_3091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_2182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5042__A _5042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2385__B _2432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_2418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3497__A _3924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4997__CLK _4997_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_3439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_3936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4121__A _4188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _2218_/X _2219_/Y _1975_/X vssd1 vssd1 vccd1 vccd1 _2221_/B sky130_fd_sc_hd__o21a_1
XFILLER_6_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_2867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2151_ _4484_/Q _2151_/B vssd1 vssd1 vccd1 vccd1 _4484_/D sky130_fd_sc_hd__xnor2_1
XFILLER_1_4087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_4018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2082_ _4436_/Q _2082_/B vssd1 vssd1 vccd1 vccd1 _4436_/D sky130_fd_sc_hd__xnor2_1
XFILLER_1_3397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_TE_B
+ _2782_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_2941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2984_ _4946_/Q _4945_/Q vssd1 vssd1 vccd1 vccd1 _2984_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_30_3517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_3528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4723_ _3399_/Y _4723_/D _3667_/Y vssd1 vssd1 vccd1 vccd1 _4723_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1935_ _1935_/A _3737_/Y vssd1 vssd1 vccd1 vccd1 _1935_/Y sky130_fd_sc_hd__nor2_2
XFILLER_11_2215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4654_ input20/X _4654_/D fanout217/X vssd1 vssd1 vccd1 vccd1 _4654_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_4114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1866_ _2143_/A _1912_/B _1912_/C vssd1 vssd1 vccd1 vccd1 _1867_/B sky130_fd_sc_hd__and3_1
X_3605_ _5062_/A vssd1 vssd1 vccd1 vccd1 _3605_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_11_1525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4585_ _4623_/CLK _4585_/D fanout231/X vssd1 vssd1 vccd1 vccd1 _4585_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4776__RESET_B fanout253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1797_ _3114_/A _1797_/B vssd1 vssd1 vccd1 vccd1 _1798_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3536_ _3550_/A vssd1 vssd1 vccd1 vccd1 _3536_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout103_A _3135_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4705__RESET_B fanout242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3467_ _3905_/A _3913_/A vssd1 vssd1 vccd1 vccd1 _3467_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_GATE_N
+ fanout128/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _4359_/CLK fanout193/X vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_2_3106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2418_ _2418_/A vssd1 vssd1 vccd1 vccd1 _2418_/Y sky130_fd_sc_hd__inv_2
X_3398_ _3414_/A vssd1 vssd1 vccd1 vccd1 _3398_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_3139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_2405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2349_ _2412_/A _2349_/B vssd1 vssd1 vccd1 vccd1 _2350_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_2449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5068_ _5068_/A vssd1 vssd1 vccd1 vccd1 _5068_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_4129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4019_ _4499_/Q vssd1 vssd1 vccd1 vccd1 _4498_/D sky130_fd_sc_hd__inv_2
XFILLER_35_3417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_2451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5037__A _5045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_3905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input33_A rstb vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_2084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5025__CLK input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3166__64_A _3169__65/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_2947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_2237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3020__A _3030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_2671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_3269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_2693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1720_ _4963_/Q vssd1 vssd1 vccd1 vccd1 _4964_/D sky130_fd_sc_hd__inv_2
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
+ _4989_/Q _3117_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_12_1856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4370_ _4370_/CLK _4370_/D fanout217/X vssd1 vssd1 vccd1 vccd1 _4370_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_3608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_4022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3321_ _3891_/A _3889_/A vssd1 vssd1 vccd1 vccd1 _3321_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_25_2907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3092__B1_N _3085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_4138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3690__A _3695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _3895_/A _3372_/B vssd1 vssd1 vccd1 vccd1 _3252_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_26_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ _4517_/Q _4516_/Q vssd1 vssd1 vccd1 vccd1 _2203_/Y sky130_fd_sc_hd__xnor2_2
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_3387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3183_ _4367_/Q vssd1 vssd1 vccd1 vccd1 _3372_/B sky130_fd_sc_hd__buf_12
XFILLER_3_2736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2134_ _4491_/Q _4490_/Q _4489_/Q _2134_/D vssd1 vssd1 vccd1 vccd1 _2135_/D sky130_fd_sc_hd__and4_1
X_2065_ _2036_/D _2064_/X _2003_/X vssd1 vssd1 vccd1 vccd1 _2066_/B sky130_fd_sc_hd__o21ai_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_4059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2967_ _2967_/A _2967_/B vssd1 vssd1 vccd1 vccd1 _2968_/A sky130_fd_sc_hd__or2_1
XFILLER_30_2602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3865__A _3908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout220_A fanout221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1918_ _4333_/Q _4332_/Q vssd1 vssd1 vccd1 vccd1 _1918_/Y sky130_fd_sc_hd__xnor2_2
X_4706_ _4709_/CLK _4706_/D fanout241/X vssd1 vssd1 vccd1 vccd1 _4706_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__4542__CLK _3932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_3781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2898_ _4892_/Q _2902_/B _2904_/A vssd1 vssd1 vccd1 vccd1 _2946_/C sky130_fd_sc_hd__o21ai_1
XFILLER_30_2657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4637_ _3922_/X _4637_/D _3353_/Y vssd1 vssd1 vccd1 vccd1 _4637_/Q sky130_fd_sc_hd__dfrtp_1
X_1849_ _4299_/Q _4298_/Q vssd1 vssd1 vccd1 vccd1 _1849_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_28_3221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_2089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_3243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4568_ _3315_/Y _4568_/D _3709__94/Y vssd1 vssd1 vccd1 vccd1 _4568_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4692__CLK _5013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3519_ _3519_/A vssd1 vssd1 vccd1 vccd1 _3519_/Y sky130_fd_sc_hd__inv_2
X_4499_ _4126_/A _4499_/D _3731_/Y vssd1 vssd1 vccd1 vccd1 _4499_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_1830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_2586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_2597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_3072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1832__B _4289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3105__A _5024_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout136/X fanout238/X vssd1 vssd1 vccd1 vccd1 _5084_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_17_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_3670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_2546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_3917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4280__RESET_B fanout199/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_3516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
+ _4704_/Q _2617_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_3779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2557__C _4707_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4415__CLK _2286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3870_ _4362_/Q _4361_/Q vssd1 vssd1 vccd1 vccd1 _3870_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_35_3781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2821_ _4857_/Q _4856_/Q _2829_/C _2832_/A vssd1 vssd1 vccd1 vccd1 _2875_/B sky130_fd_sc_hd__a31o_1
XFILLER_31_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3685__A _3696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2752_ _2771_/A _2752_/B vssd1 vssd1 vccd1 vccd1 _2753_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_2966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1703_ _3556_/A _1704_/B vssd1 vssd1 vccd1 vccd1 _4935_/D sky130_fd_sc_hd__xor2_1
X_2683_ _4770_/Q _2647_/D _2675_/B vssd1 vssd1 vccd1 vccd1 _2684_/B sky130_fd_sc_hd__a21bo_1
XFILLER_12_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_3613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4422_ _3232_/Y _4422_/D _3750_/Y vssd1 vssd1 vccd1 vccd1 _4422_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_3585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4353_ input17/X _4353_/D fanout189/X vssd1 vssd1 vccd1 vccd1 _4353_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3304_ _3912_/A _3446_/B vssd1 vssd1 vccd1 vccd1 _3304_/Y sky130_fd_sc_hd__xnor2_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4284_ _4288_/CLK _4284_/D fanout194/X vssd1 vssd1 vccd1 vccd1 _4284_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3235_ _3738_/A vssd1 vssd1 vccd1 vccd1 _3255_/A sky130_fd_sc_hd__buf_6
XFILLER_7_2680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2117_ _2286_/B _2115_/X _2116_/X _3892_/A vssd1 vssd1 vccd1 vccd1 _2121_/A sky130_fd_sc_hd__o211a_1
XANTENNA_fanout170_A _3861_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3097_ _4992_/Q _3097_/B vssd1 vssd1 vccd1 vccd1 _4992_/D sky130_fd_sc_hd__xnor2_1
XFILLER_3_1887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4908__CLK _4247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2048_ _2046_/X _2047_/Y _1975_/X vssd1 vssd1 vccd1 vccd1 _2049_/B sky130_fd_sc_hd__o21a_1
XANTENNA__2057__A2 _4430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_2221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
+ _4762_/Q _2714_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_22_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_2276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3999_ _4001_/A _4005_/A vssd1 vssd1 vccd1 vccd1 _4123_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__3595__A _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_3177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_2476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3169__65 _3169__65/A vssd1 vssd1 vccd1 vccd1 _3169__65/Y sky130_fd_sc_hd__inv_2
XFILLER_30_2498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_3062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3684_/A fanout216/X vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__2939__A _4931_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1843__A _2143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2658__B _4763_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4438__CLK _5041_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_2499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[5\].w1.ro_block_Q.ro_pol.tribuf.t_buf _2963_/X _2812_/Y vssd1
+ vssd1 vccd1 vccd1 _5090_/A sky130_fd_sc_hd__ebufn_8
XFILLER_8_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__1632_ clkbuf_0__1632_/X vssd1 vssd1 vccd1 vccd1 _3189__72/A sky130_fd_sc_hd__clkbuf_16
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4588__CLK _4590_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5050__A _5058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3489__B _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4461__RESET_B fanout199/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4961__SET_B fanout208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_2114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_2208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_3725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2568__B _2568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_3471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_3313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_4058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf _4281_/Q _1846_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_27_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3478__47 _3528__52/A vssd1 vssd1 vccd1 vccd1 _3478__47/Y sky130_fd_sc_hd__inv_2
X_3020_ _3030_/A _3020_/B vssd1 vssd1 vccd1 vccd1 _3021_/B sky130_fd_sc_hd__nand2_1
XFILLER_3_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_2645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2584__A _2680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3399__B _4129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4971_ _4248_/B _4971_/D _3540_/Y vssd1 vssd1 vccd1 vccd1 _4971_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_3275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3922_ _3922_/A vssd1 vssd1 vccd1 vccd1 _3922_/X sky130_fd_sc_hd__buf_6
XFILLER_31_4143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3853_ _4366_/Q _4365_/Q vssd1 vssd1 vccd1 vccd1 _3872_/B sky130_fd_sc_hd__xnor2_2
XFILLER_14_2449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2804_ _3914_/B _2799_/Y _2800_/X _2803_/Y vssd1 vssd1 vccd1 vccd1 _2805_/B sky130_fd_sc_hd__a31o_1
XFILLER_31_2741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2735_ _2771_/A _2735_/B vssd1 vssd1 vccd1 vccd1 _2736_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_4072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2666_ _4765_/Q _2666_/B vssd1 vssd1 vccd1 vccd1 _2666_/X sky130_fd_sc_hd__and2b_1
XFILLER_12_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4405_ _2809_/A1 _4405_/D _3216_/Y vssd1 vssd1 vccd1 vccd1 _4405_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_3465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2597_ _4715_/Q _2597_/B vssd1 vssd1 vccd1 vccd1 _4715_/D sky130_fd_sc_hd__xnor2_1
Xfanout204 fanout207/X vssd1 vssd1 vccd1 vccd1 fanout204/X sky130_fd_sc_hd__clkbuf_2
X_4336_ _3914_/A _4336_/D _3179__68/Y vssd1 vssd1 vccd1 vccd1 _4336_/Q sky130_fd_sc_hd__dfrtp_2
Xclkbuf_1_0_2_clk_master clkbuf_1_0_2_clk_master/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clk_master/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_25_3279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout215 fanout217/X vssd1 vssd1 vccd1 vccd1 fanout215/X sky130_fd_sc_hd__buf_2
Xfanout226 fanout230/X vssd1 vssd1 vccd1 vccd1 fanout226/X sky130_fd_sc_hd__buf_4
XFILLER_5_2606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout237 fanout257/X vssd1 vssd1 vccd1 vccd1 fanout237/X sky130_fd_sc_hd__buf_2
XFILLER_25_2556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout248 fanout250/X vssd1 vssd1 vccd1 vccd1 fanout248/X sky130_fd_sc_hd__buf_2
XFILLER_5_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4267_ _3846_/A _4267_/D _5056_/A vssd1 vssd1 vccd1 vccd1 _4267_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_2409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3218_ _3947_/A _3438_/B vssd1 vssd1 vccd1 vccd1 _3218_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4730__CLK _4920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4198_ _4756_/Q vssd1 vssd1 vccd1 vccd1 _4755_/D sky130_fd_sc_hd__inv_2
XFILLER_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_2385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3149_ _3838_/A _3839_/A vssd1 vssd1 vccd1 vccd1 _3149_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4880__CLK _4916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_2349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_3938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5020__D _5020_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4901__RESET_B fanout232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3157__57 _3159__59/A vssd1 vssd1 vccd1 vccd1 _3157__57/Y sky130_fd_sc_hd__inv_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5045__A _5045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_2000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2910__B1 _2858_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_2987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5055_/A fanout244/X vssd1 vssd1 vccd1 vccd1 _5079_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_34_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_2725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_3161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_2769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4124__A _4131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4603__CLK _4943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2520_ _4677_/Q _2520_/B vssd1 vssd1 vccd1 vccd1 _4677_/D sky130_fd_sc_hd__xnor2_1
XFILLER_5_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1952__A1 _1952_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_4109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2579__A _4712_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2451_ _2451_/A vssd1 vssd1 vccd1 vccd1 _2453_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_26_3555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_3649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4753__CLK _3861_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2382_ _4619_/Q _4618_/Q _4617_/Q _2404_/B vssd1 vssd1 vccd1 vccd1 _2394_/B sky130_fd_sc_hd__or4_1
XFILLER_26_3588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
+ _4523_/Q _2268_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_29_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4121_ _4188_/B vssd1 vssd1 vccd1 vccd1 _4121_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_22_2729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4052_ _4546_/Q vssd1 vssd1 vccd1 vccd1 _4547_/D sky130_fd_sc_hd__inv_2
XFILLER_4_3395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_2650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_2661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput4 comp_high_I[3] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
X_3003_ _3030_/A _3003_/B vssd1 vssd1 vccd1 vccd1 _3004_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_3198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_GATE_N _4363_/CLK
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_82 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4954_ _4958_/CLK _4954_/D fanout218/X vssd1 vssd1 vccd1 vccd1 _4954_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_93 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3905_ _3905_/A vssd1 vssd1 vccd1 vccd1 _3912_/A sky130_fd_sc_hd__buf_12
XFILLER_14_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4885_ _3495_/Y _4885_/D _3619_/Y vssd1 vssd1 vccd1 vccd1 _4885_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_2235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_2869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3836_ _3883_/A vssd1 vssd1 vccd1 vccd1 _3846_/A sky130_fd_sc_hd__clkinv_2
XANTENNA_fanout133_A _4623_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2480__C _4672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4283__CLK _4288_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3873__A _3883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2718_ _4808_/Q _4807_/Q _2718_/C vssd1 vssd1 vccd1 vccd1 _2719_/D sky130_fd_sc_hd__and3_1
X_3698_ _4071_/A vssd1 vssd1 vccd1 vccd1 _3698_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1943__A1 _3882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2649_ _4762_/Q vssd1 vssd1 vccd1 vccd1 _2661_/A sky130_fd_sc_hd__inv_2
XFILLER_25_3021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_3273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3145__B1 _3139_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_2331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4319_ _4324_/CLK _4319_/D fanout189/X vssd1 vssd1 vccd1 vccd1 _4319_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_2364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_3964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3192__74_A _3193__75/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2120__A1 _3931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_2193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_2102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
+ _4581_/Q _2366_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4626__CLK _4626_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_4046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4776__CLK _4812_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2399__A _2412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_4142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4894__RESET_B fanout236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_3568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3023__A _3030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2662__A2 _2658_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1870__B1 _1791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1951_ _3882_/A _1951_/B _1951_/C vssd1 vssd1 vccd1 vccd1 _1951_/X sky130_fd_sc_hd__or3_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__0625_ clkbuf_0__0625_/X vssd1 vssd1 vccd1 vccd1 _3655__85/A sky130_fd_sc_hd__clkbuf_16
X_4670_ _4718_/CLK _4670_/D fanout242/X vssd1 vssd1 vccd1 vccd1 _4670_/Q sky130_fd_sc_hd__dfrtp_4
X_1882_ _4316_/Q _1858_/D _1875_/B vssd1 vssd1 vccd1 vccd1 _1883_/B sky130_fd_sc_hd__a21bo_1
XFILLER_19_1990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3621_ _4256_/A vssd1 vssd1 vccd1 vccd1 _3621_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3693__A _3695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3552_ _5028_/Q _5029_/Q vssd1 vssd1 vccd1 vccd1 _3552_/X sky130_fd_sc_hd__xor2_1
XFILLER_31_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2503_ _4672_/Q _2503_/B vssd1 vssd1 vccd1 vccd1 _4672_/D sky130_fd_sc_hd__xnor2_1
XFILLER_28_2916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3483_ _4249_/A _4250_/A vssd1 vssd1 vccd1 vccd1 _3483_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_2938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_3363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2434_ _2608_/A _4626_/Q vssd1 vssd1 vccd1 vccd1 _4626_/D sky130_fd_sc_hd__xor2_1
XFILLER_6_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_3457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2365_ _4594_/Q _4593_/Q vssd1 vssd1 vccd1 vccd1 _2365_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1941__A _3898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4104_ _4632_/Q vssd1 vssd1 vccd1 vccd1 _4631_/D sky130_fd_sc_hd__inv_2
XFILLER_0_3001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5084_ _5084_/A vssd1 vssd1 vccd1 vccd1 _5084_/X sky130_fd_sc_hd__buf_4
XFILLER_0_3023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2296_ _3877_/A _3907_/A _3932_/A _1937_/Y _2295_/Y vssd1 vssd1 vccd1 vccd1 _2297_/B
+ sky130_fd_sc_hd__o41a_1
X_4035_ _4515_/Q vssd1 vssd1 vccd1 vccd1 _4514_/D sky130_fd_sc_hd__inv_2
XANTENNA__2638__C1 _3875_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4564__RESET_B fanout223/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4649__CLK input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3868__A _3916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout250_A fanout256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4937_ _3598_/A _4937_/D fanout214/X vssd1 vssd1 vccd1 vccd1 _4937_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__2491__B _2491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_2190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4799__CLK _4811_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4868_ _4905_/CLK _4868_/D fanout231/X vssd1 vssd1 vccd1 vccd1 _4868_/Q sky130_fd_sc_hd__dfstp_1
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout180/X fanout184/X vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3819_ _4333_/Q vssd1 vssd1 vccd1 vccd1 _4332_/D sky130_fd_sc_hd__inv_2
XANTENNA__2169__A1 _4491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4799_ _4811_/CLK _4799_/D fanout247/X vssd1 vssd1 vccd1 vccd1 _4799_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_2953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3108__A _5024_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2012__A _4462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_2069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2385__C _2432_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2682__A _2922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3497__B _3923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_2474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5022__RESET_B fanout208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3018__A _4953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_4011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_2813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_4033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1761__A _4247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2150_ _2178_/A _2150_/B vssd1 vssd1 vccd1 vccd1 _2151_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_3321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_2879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2081_ _2034_/C _2077_/Y _2003_/X vssd1 vssd1 vccd1 vccd1 _2082_/B sky130_fd_sc_hd__o21ai_1
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_2570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_3329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3688__A _3695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4941__CLK _4943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2983_ _4944_/Q _4943_/Q vssd1 vssd1 vccd1 vccd1 _2983_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_15_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4722_ _5007_/CLK _4722_/D _3398_/Y vssd1 vssd1 vccd1 vccd1 _4722_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_12_3941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1934_ _1934_/A vssd1 vssd1 vccd1 vccd1 _1934_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_2986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_3963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1865_ _4312_/Q _1869_/B _1871_/A vssd1 vssd1 vccd1 vccd1 _1912_/C sky130_fd_sc_hd__o21ai_1
X_4653_ input20/X _4653_/D fanout217/X vssd1 vssd1 vccd1 vccd1 _4654_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_12_3996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4584_ _4623_/CLK _4584_/D fanout231/X vssd1 vssd1 vccd1 vccd1 _4584_/Q sky130_fd_sc_hd__dfrtp_2
X_1796_ _4277_/Q _1789_/C _1790_/B vssd1 vssd1 vccd1 vccd1 _1797_/B sky130_fd_sc_hd__a21bo_1
X_3535_ _3556_/A _3556_/B vssd1 vssd1 vccd1 vccd1 _3535_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_2713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4321__CLK _4324_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3466_ _3466_/A vssd1 vssd1 vccd1 vccd1 _3466_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_3002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_2779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2417_ _2922_/A vssd1 vssd1 vccd1 vccd1 _2566_/A sky130_fd_sc_hd__buf_6
XFILLER_6_3265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2767__A _4838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_2301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3397_ _4189_/A _4190_/A vssd1 vssd1 vccd1 vccd1 _3397_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_22_2323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2348_ _2347_/Y _2303_/C _4586_/Q vssd1 vssd1 vccd1 vccd1 _2349_/B sky130_fd_sc_hd__mux2_1
XANTENNA__2486__B _4672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5067_ _5067_/A vssd1 vssd1 vccd1 vccd1 _5067_/X sky130_fd_sc_hd__clkbuf_1
X_2279_ _2279_/A vssd1 vssd1 vccd1 vccd1 _2279_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4018_ _4480_/Q vssd1 vssd1 vccd1 vccd1 _4481_/D sky130_fd_sc_hd__inv_2
XFILLER_0_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xw0.ro_block_I.ro_pol.tribuf.t_buf _1934_/X _1772_/Y vssd1 vssd1 vccd1 vccd1 _5088_/A
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__3598__A _3598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1834__B1 _1823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5048_/A fanout191/X vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_33_1762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_3834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4814__CLK _3449_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3643_/A fanout245/X vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__5053__A _5061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4486__RESET_B fanout201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A phi1b_dig_Q[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_2890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3301__A _3309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_2205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_2959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3478__47_A _3528__52/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4344__CLK _3845_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output94_A _5091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2553__A1 _4707_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3255_/A vssd1 vssd1 vccd1 vccd1 _3251_/Y sky130_fd_sc_hd__inv_2
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2587__A _2680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _4515_/Q _4514_/Q vssd1 vssd1 vccd1 vccd1 _2202_/Y sky130_fd_sc_hd__xnor2_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2133_ _4493_/Q _4492_/Q _2133_/C vssd1 vssd1 vccd1 vccd1 _2134_/D sky130_fd_sc_hd__and3_1
XFILLER_1_2450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2064_ _4432_/Q _2064_/B vssd1 vssd1 vccd1 vccd1 _2064_/X sky130_fd_sc_hd__and2b_1
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_GATE_N
+ _5059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_2403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_4016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_4038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2966_ _4932_/D _4933_/Q vssd1 vssd1 vccd1 vccd1 _2967_/B sky130_fd_sc_hd__and2b_1
XFILLER_33_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4705_ _4718_/CLK _4705_/D fanout242/X vssd1 vssd1 vccd1 vccd1 _4705_/Q sky130_fd_sc_hd__dfrtp_1
X_1917_ _4331_/Q _4330_/Q vssd1 vssd1 vccd1 vccd1 _1917_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_15_2182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_2024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2897_ _4895_/Q _4894_/Q _4893_/Q _2908_/B vssd1 vssd1 vccd1 vccd1 _2902_/B sky130_fd_sc_hd__or4_1
XFILLER_11_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4636_ _3352_/Y _4636_/D _3690_/Y vssd1 vssd1 vccd1 vccd1 _4636_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout213_A fanout220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1848_ _4297_/Q _4296_/Q vssd1 vssd1 vccd1 vccd1 _1848_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_11_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_3233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4837__CLK input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1779_ _4280_/Q _4279_/Q _4278_/Q _1779_/D vssd1 vssd1 vccd1 vccd1 _1789_/C sky130_fd_sc_hd__and4_1
X_4567_ _2294_/B1 _4567_/D _3314__26/Y vssd1 vssd1 vccd1 vccd1 _4567_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4926__RESET_B fanout228/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3518_ _3924_/A _3923_/A vssd1 vssd1 vccd1 vccd1 _3518_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_3299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4498_ _4248_/A _4498_/D _3270_/Y vssd1 vssd1 vccd1 vccd1 _4498_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_3062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3449_ _4249_/A _4250_/A vssd1 vssd1 vccd1 vccd1 _3449_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__4987__CLK _4997_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf_A
+ _4961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_2153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_3983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_2164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5023__D input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4367__CLK _4472_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_2801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5048__A _5048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3375_/A fanout240/X vssd1 vssd1 vccd1 vccd1 _5076_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_26_3929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_3861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2557__D _2568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4127__A _4127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_3771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_3793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2820_ _4855_/Q vssd1 vssd1 vccd1 vccd1 _2832_/A sky130_fd_sc_hd__inv_2
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_TE_B _1917_/Y vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_2057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2751_ _4806_/Q _4805_/Q _2719_/D _2748_/B vssd1 vssd1 vccd1 vccd1 _2752_/B sky130_fd_sc_hd__a31o_1
XFILLER_12_2333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1702_ _4247_/A _1761_/C vssd1 vssd1 vccd1 vccd1 _1704_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2682_ _2922_/A vssd1 vssd1 vccd1 vccd1 _2771_/A sky130_fd_sc_hd__clkbuf_4
X_4421_ _2294_/B1 _4421_/D _3231_/Y vssd1 vssd1 vccd1 vccd1 _4421_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_3417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_2852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4352_ input17/X _4352_/D fanout189/X vssd1 vssd1 vccd1 vccd1 _4353_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_9_2935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3303_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3303_/Y sky130_fd_sc_hd__inv_2
X_4283_ _4288_/CLK _4283_/D fanout195/X vssd1 vssd1 vccd1 vccd1 _4283_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _3885_/A _3886_/A vssd1 vssd1 vccd1 vccd1 _3234_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_3_3246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[3\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf_A _2622_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_2451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3165_ _3947_/A _3438_/B vssd1 vssd1 vccd1 vccd1 _3165_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_3_1811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2116_ _3910_/A _3908_/A _1936_/X _1937_/Y _3898_/B vssd1 vssd1 vccd1 vccd1 _2116_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_3_2589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3096_ _3057_/D _3095_/Y _1791_/X vssd1 vssd1 vccd1 vccd1 _3097_/B sky130_fd_sc_hd__o21ai_1
X_2047_ _4427_/Q _2047_/B vssd1 vssd1 vccd1 vccd1 _2047_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_1899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout163_A _3939_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2057__A3 _2036_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_2233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_3991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3998_ _4471_/Q vssd1 vssd1 vccd1 vccd1 _4005_/A sky130_fd_sc_hd__buf_6
XFILLER_17_2288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_3145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2949_ _4907_/Q _4906_/Q vssd1 vssd1 vccd1 vccd1 _2949_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_30_3189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4619_ _4626_/CLK _4619_/D fanout233/X vssd1 vssd1 vccd1 vccd1 _4619_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_3113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5015__CLK _3930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2939__B _4905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2658__C _2658_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_2478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2020__A _3066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2296__A3 _3932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_3744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_3788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_2126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_3325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4532__CLK _4532_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4970_ _3539_/Y _4970_/D _3594_/Y vssd1 vssd1 vccd1 vccd1 _4970_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
+ _4893_/Q _2954_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_3921_ _3940_/A vssd1 vssd1 vccd1 vccd1 _3922_/A sky130_fd_sc_hd__inv_2
XANTENNA__4682__CLK _4718_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3419__38_A _3425__41/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3696__A _3696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3852_ _3888_/A vssd1 vssd1 vccd1 vccd1 _3892_/A sky130_fd_sc_hd__clkinv_2
XFILLER_32_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_2597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2803_ _4064_/A _2802_/Y _3914_/B vssd1 vssd1 vccd1 vccd1 _2803_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_2141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2734_ _4800_/Q _2730_/C _2731_/B vssd1 vssd1 vccd1 vccd1 _2735_/B sky130_fd_sc_hd__a21bo_1
XFILLER_34_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4518__RESET_B fanout219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2665_ _4766_/Q _2665_/B vssd1 vssd1 vccd1 vccd1 _2666_/B sky130_fd_sc_hd__nor2_1
XFILLER_29_3350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1944__A _3898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4404_ _4429_/CLK _4404_/D fanout189/X vssd1 vssd1 vccd1 vccd1 _4404_/Q sky130_fd_sc_hd__dfrtp_2
X_2596_ _2549_/C _2592_/Y _2518_/X vssd1 vssd1 vccd1 vccd1 _2597_/B sky130_fd_sc_hd__o21ai_1
XFILLER_25_3247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_2743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4335_ _3178_/Y _4335_/D _3769__108/Y vssd1 vssd1 vccd1 vccd1 _4335_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout205 fanout206/X vssd1 vssd1 vccd1 vccd1 fanout205/X sky130_fd_sc_hd__buf_2
XFILLER_29_2693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout216 fanout217/X vssd1 vssd1 vccd1 vccd1 fanout216/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout227 fanout230/X vssd1 vssd1 vccd1 vccd1 fanout227/X sky130_fd_sc_hd__buf_2
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout238 fanout239/X vssd1 vssd1 vccd1 vccd1 fanout238/X sky130_fd_sc_hd__buf_2
XFILLER_7_3190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout249 fanout250/X vssd1 vssd1 vccd1 vccd1 fanout249/X sky130_fd_sc_hd__buf_2
XFILLER_9_2798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4266_ _3883_/A _4266_/D _5056_/A vssd1 vssd1 vccd1 vccd1 _4266_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_1856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3217_ _3233_/A vssd1 vssd1 vccd1 vccd1 _3217_/Y sky130_fd_sc_hd__inv_2
X_4197_ _4753_/Q vssd1 vssd1 vccd1 vccd1 _4754_/D sky130_fd_sc_hd__clkinv_2
XFILLER_3_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3148_ _4248_/D _3148_/B vssd1 vssd1 vccd1 vccd1 _5071_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_3975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3079_ _4989_/Q _4988_/Q _3058_/D _3076_/B vssd1 vssd1 vccd1 vccd1 _3080_/B sky130_fd_sc_hd__a31o_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_A
+ _4430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_2085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3259__19_A _3262__21/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_2263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4405__CLK _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
+ _4951_/Q _3049_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4555__CLK input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_3689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5061__A _5061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_2966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_2977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2426__B1 _2344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__0641_ clkbuf_0__0641_/X vssd1 vssd1 vccd1 vccd1 _3781__122/A sky130_fd_sc_hd__clkbuf_16
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_2185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4611__RESET_B fanout231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1952__A2 _3892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2450_ _4654_/Q _4653_/D vssd1 vssd1 vccd1 vccd1 _2451_/A sky130_fd_sc_hd__and2b_1
XFILLER_9_2006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2579__B _2579_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2381_ _4622_/Q _4621_/Q _4620_/Q _2418_/A vssd1 vssd1 vccd1 vccd1 _2404_/B sky130_fd_sc_hd__or4_1
XFILLER_6_2927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4120_ _4656_/Q _4657_/Q vssd1 vssd1 vccd1 vccd1 _4188_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_3205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4051_ _4547_/Q vssd1 vssd1 vccd1 vccd1 _4546_/D sky130_fd_sc_hd__inv_2
XFILLER_7_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput5 comp_high_I[4] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_2673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3002_ _4950_/Q _2998_/C _2999_/B vssd1 vssd1 vccd1 vccd1 _3003_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_3249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_72 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_83 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4953_ _4958_/CLK _4953_/D fanout214/X vssd1 vssd1 vccd1 vccd1 _4953_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3904_ _3904_/A _3904_/B vssd1 vssd1 vccd1 vccd1 _4370_/D sky130_fd_sc_hd__xnor2_1
X_4884_ _4920_/CLK _4884_/D _3494_/Y vssd1 vssd1 vccd1 vccd1 _4884_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_2837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3835_ _3838_/A _3839_/A vssd1 vssd1 vccd1 vccd1 _3883_/A sky130_fd_sc_hd__xnor2_4
XFILLER_14_2247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4428__CLK _4429_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2480__D _2480_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_2561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3766_ _3777_/A vssd1 vssd1 vccd1 vccd1 _3766_/X sky130_fd_sc_hd__buf_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout126_A _5044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3873__B _3883_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2717_ _4838_/D _4812_/Q _4810_/Q _4809_/Q vssd1 vssd1 vccd1 vccd1 _2718_/C sky130_fd_sc_hd__and4_1
X_3697_ _4071_/A vssd1 vssd1 vccd1 vccd1 _3697_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4578__CLK _5043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_2608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2648_ _4767_/Q _4766_/Q _4765_/Q _2648_/D vssd1 vssd1 vccd1 vccd1 _2658_/C sky130_fd_sc_hd__and4_2
XANTENNA__3145__A1 _4064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2579_ _4712_/Q _2579_/B vssd1 vssd1 vccd1 vccd1 _2580_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_3077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4318_ _4324_/CLK _4318_/D fanout189/X vssd1 vssd1 vccd1 vccd1 _4318_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_5_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4249_ _4249_/A _4250_/B vssd1 vssd1 vccd1 vccd1 _4842_/D sky130_fd_sc_hd__xnor2_1
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_TE_B
+ _2026_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_4003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout157/X fanout203/X vssd1 vssd1 vccd1 vccd1 _5082_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_19_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_4058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_4069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_3357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3706__91_A _3732__95/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_2093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5056__A _5056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_4110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3304__A _3912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_2813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_2868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_4094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4863__RESET_B fanout226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3471__43 _3523__49/A vssd1 vssd1 vccd1 vccd1 _4845_/CLK sky130_fd_sc_hd__inv_2
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4135__A _4135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1950_ _3888_/A _3914_/A _1936_/X vssd1 vssd1 vccd1 vccd1 _1951_/C sky130_fd_sc_hd__a21oi_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__0624_ clkbuf_0__0624_/X vssd1 vssd1 vccd1 vccd1 _3777_/A sky130_fd_sc_hd__clkbuf_16
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1881_ _4314_/Q _1881_/B vssd1 vssd1 vccd1 vccd1 _4314_/D sky130_fd_sc_hd__xnor2_1
XFILLER_15_2567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3620_ _4256_/A vssd1 vssd1 vccd1 vccd1 _3620_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4720__CLK _4187_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3551_ _3924_/A _3923_/A vssd1 vssd1 vccd1 vccd1 _3551_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_3629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2502_ _2566_/A _2502_/B vssd1 vssd1 vccd1 vccd1 _2503_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_4043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3482_ _3498_/A vssd1 vssd1 vccd1 vccd1 _3482_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_4065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_3331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2433_ _4625_/Q _2433_/B vssd1 vssd1 vccd1 vccd1 _4625_/D sky130_fd_sc_hd__xor2_1
XANTENNA__4870__CLK _1700_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_2713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_3386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_3469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2364_ _4592_/Q _4591_/Q vssd1 vssd1 vccd1 vccd1 _2364_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_26_2674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1941__B _3914_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4103_ _4629_/Q vssd1 vssd1 vccd1 vccd1 _4630_/D sky130_fd_sc_hd__inv_2
X_2295_ _2288_/Y _2294_/Y _3932_/A vssd1 vssd1 vccd1 vccd1 _2295_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_22_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5083_ _5083_/A vssd1 vssd1 vccd1 vccd1 _5083_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3214__A _3848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4034_ _4512_/Q vssd1 vssd1 vccd1 vccd1 _4513_/D sky130_fd_sc_hd__inv_2
XFILLER_0_3057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_4003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
+ _4712_/Q _2609_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3868__B _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_2601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4936_ _4936_/CLK _4936_/D fanout224/X vssd1 vssd1 vccd1 vccd1 _4936_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout243_A fanout245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4867_ _4905_/CLK _4867_/D fanout226/X vssd1 vssd1 vccd1 vccd1 _4867_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_3622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_GATE_N _5056_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3818_ _4330_/Q vssd1 vssd1 vccd1 vccd1 _4331_/D sky130_fd_sc_hd__inv_2
X_4798_ _4811_/CLK _4798_/D fanout245/X vssd1 vssd1 vccd1 vccd1 _4798_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_2965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3749_ _3749_/A vssd1 vssd1 vccd1 vccd1 _3948_/A sky130_fd_sc_hd__buf_8
XFILLER_11_2987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_2416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_2223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_2245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_2278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2963__A _2963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3749_/A fanout187/X vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_28_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4743__CLK input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4274__RESET_B fanout199/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_3916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4893__CLK _4901_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_4001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_3559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_4023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_2825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1761__B _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_4045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3034__A _5020_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2080_ _4435_/Q _2080_/B vssd1 vssd1 vccd1 vccd1 _4435_/D sky130_fd_sc_hd__xnor2_1
XFILLER_1_3377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4273__CLK _3846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout120/X fanout249/X vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_1_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_3611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2982_ _4942_/Q _4941_/Q vssd1 vssd1 vccd1 vccd1 _2982_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4721_ _3397_/Y _4721_/D _3668_/Y vssd1 vssd1 vccd1 vccd1 _4721_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1933_ _1933_/A _1933_/B vssd1 vssd1 vccd1 vccd1 _1934_/A sky130_fd_sc_hd__or2_1
XFILLER_15_2353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_2818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
+ _4427_/Q _2100_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_4652_ input20/X _4652_/D fanout222/X vssd1 vssd1 vccd1 vccd1 _4653_/D sky130_fd_sc_hd__dfrtp_1
X_1864_ _4315_/Q _4314_/Q _4313_/Q _1875_/B vssd1 vssd1 vccd1 vccd1 _1869_/B sky130_fd_sc_hd__or4_1
XFILLER_15_2397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_2239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput30 phi1b_dig_Q[5] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_2
X_4583_ _4590_/CLK _4583_/D fanout227/X vssd1 vssd1 vccd1 vccd1 _4583_/Q sky130_fd_sc_hd__dfrtp_2
X_1795_ _2922_/A vssd1 vssd1 vccd1 vccd1 _3114_/A sky130_fd_sc_hd__buf_12
XFILLER_28_3415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3534_ _3550_/A vssd1 vssd1 vccd1 vccd1 _3534_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_2736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3465_ _3916_/A _3915_/A vssd1 vssd1 vccd1 vccd1 _3465_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_6_3233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2416_ _4620_/Q _2416_/B vssd1 vssd1 vccd1 vccd1 _4620_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__2859__B1 _2858_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3396_ _3414_/A vssd1 vssd1 vccd1 vccd1 _3396_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_3277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4616__CLK _4626_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_2554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2347_ _2347_/A vssd1 vssd1 vccd1 vccd1 _2347_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_2335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout193_A fanout196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_2346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2486__C _4671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5066_ _5066_/A vssd1 vssd1 vccd1 vccd1 _5066_/X sky130_fd_sc_hd__clkbuf_1
X_2278_ _2278_/A _2278_/B vssd1 vssd1 vccd1 vccd1 _2279_/A sky130_fd_sc_hd__or2_1
XFILLER_2_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4017_ _4481_/Q vssd1 vssd1 vccd1 vccd1 _4480_/D sky130_fd_sc_hd__inv_2
XFILLER_0_2153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3036__B1 _1791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4919_ _3514_/Y _4919_/D _3609_/Y vssd1 vssd1 vccd1 vccd1 _4919_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_1416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_2318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4296__CLK _3931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
+ _4485_/Q _2199_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_27_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input19_A phi1b_dig_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_2905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_2504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output87_A _5084_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4639__CLK _4943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2868__A _4927_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3903_/A _3420_/B vssd1 vssd1 vccd1 vccd1 _3250_/Y sky130_fd_sc_hd__xnor2_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_3417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3632_/A fanout246/X vssd1 vssd1 vccd1 vccd1 _5077_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_7_3597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _4513_/Q _4512_/Q vssd1 vssd1 vccd1 vccd1 _2201_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_23_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3181_ _3903_/A _3420_/B vssd1 vssd1 vccd1 vccd1 _3181_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4789__CLK _4920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2132_ _4555_/D _4497_/Q _4495_/Q _4494_/Q vssd1 vssd1 vccd1 vccd1 _2133_/C sky130_fd_sc_hd__and4_1
XFILLER_1_3141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3699__A _4071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2063_ _4433_/Q _2063_/B vssd1 vssd1 vccd1 vccd1 _2064_/B sky130_fd_sc_hd__nor2_1
XFILLER_1_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_4028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2965_ _2965_/A vssd1 vssd1 vccd1 vccd1 _2967_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_2773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4704_ _4718_/CLK _4704_/D fanout237/X vssd1 vssd1 vccd1 vccd1 _4704_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1916_ _4329_/Q _4328_/Q vssd1 vssd1 vccd1 vccd1 _1916_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_12_3761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2896_ _4898_/Q _4897_/Q _4896_/Q _2918_/B vssd1 vssd1 vccd1 vccd1 _2908_/B sky130_fd_sc_hd__or4_1
XFILLER_11_2047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4635_ _4920_/CLK _4635_/D _3351_/Y vssd1 vssd1 vccd1 vccd1 _4635_/Q sky130_fd_sc_hd__dfrtp_1
X_1847_ _4295_/Q _4294_/Q vssd1 vssd1 vccd1 vccd1 _1847_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_8_4018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout206_A fanout207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4566_ _4566_/CLK _4566_/D fanout211/X vssd1 vssd1 vccd1 vccd1 _4566_/Q sky130_fd_sc_hd__dfrtp_2
X_1778_ _4283_/Q _4282_/Q _4281_/Q _1778_/D vssd1 vssd1 vccd1 vccd1 _1779_/D sky130_fd_sc_hd__and4_1
X_3517_ _3519_/A vssd1 vssd1 vccd1 vccd1 _3517_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_3339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4497_ _4533_/CLK _4497_/D fanout210/X vssd1 vssd1 vccd1 vccd1 _4497_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_2638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_2408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3448_ _3466_/A vssd1 vssd1 vccd1 vccd1 _3448_/Y sky130_fd_sc_hd__inv_2
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ _3393_/A vssd1 vssd1 vccd1 vccd1 _3379_/Y sky130_fd_sc_hd__inv_2
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_2226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_2198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5049_ _5057_/A vssd1 vssd1 vccd1 vccd1 _5049_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3402__A _3414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_A
+ _4712_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_3683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2232__A1 _4524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_2846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_3861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_2294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_TE_B
+ _2101_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5064__A _5064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4931__CLK input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_3737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_4104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2471__A1 _3900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2471__B2 _3929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4311__CLK _4324_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2750_ _4803_/Q _2750_/B vssd1 vssd1 vccd1 vccd1 _4803_/D sky130_fd_sc_hd__xnor2_1
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_2946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1701_ _4248_/A _4248_/B _4248_/C _4187_/Y vssd1 vssd1 vccd1 vccd1 _1761_/C sky130_fd_sc_hd__or4_1
XANTENNA__4461__CLK input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2681_ _4768_/Q _2681_/B vssd1 vssd1 vccd1 vccd1 _4768_/D sky130_fd_sc_hd__xnor2_1
XFILLER_12_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf_TE_B
+ _2547_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4420_ _3230_/Y _4420_/D _3751_/Y vssd1 vssd1 vccd1 vccd1 _4420_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_3543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2598__A _4745_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4351_ input17/X _4351_/D fanout189/X vssd1 vssd1 vccd1 vccd1 _4352_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_7_4062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3302_ _3917_/A _3444_/B vssd1 vssd1 vccd1 vccd1 _3302_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_7_3361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4282_ _4288_/CLK _4282_/D fanout199/X vssd1 vssd1 vccd1 vccd1 _4282_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _3233_/A vssd1 vssd1 vccd1 vccd1 _3233_/Y sky130_fd_sc_hd__inv_2
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4377__RESET_B fanout212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ _3945_/A vssd1 vssd1 vccd1 vccd1 _3438_/B sky130_fd_sc_hd__buf_12
XFILLER_7_1981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2115_ _3892_/B _3899_/A _3900_/B vssd1 vssd1 vccd1 vccd1 _2115_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3095_ _4994_/Q _4993_/Q _3098_/A vssd1 vssd1 vccd1 vccd1 _3095_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__3222__A _3925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2046_ _4428_/Q _4427_/Q _2046_/C vssd1 vssd1 vccd1 vccd1 _2046_/X sky130_fd_sc_hd__and3_1
XFILLER_22_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout156_A _3922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3997_ _4470_/Q vssd1 vssd1 vccd1 vccd1 _4001_/A sky130_fd_sc_hd__buf_6
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_3878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2948_ _3114_/A _4905_/Q vssd1 vssd1 vccd1 vccd1 _4905_/D sky130_fd_sc_hd__xor2_1
XFILLER_30_3157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2879_ _4873_/Q _4872_/Q vssd1 vssd1 vccd1 vccd1 _2879_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_11_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3892__A _3892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4618_ _4626_/CLK _4618_/D fanout233/X vssd1 vssd1 vccd1 vccd1 _4618_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4549_ _3306_/Y _4549_/D _3713_/Y vssd1 vssd1 vccd1 vccd1 _4549_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_2330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_2413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_2205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_2374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_2385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_2045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4334__CLK _2286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4484__CLK _4533_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5059__A _5059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_4141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3307__A _3309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2211__A _4559_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_4005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_2811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_2603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_2614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_2877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3042__A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4827__CLK _4981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3920_ _3924_/A _3923_/A vssd1 vssd1 vccd1 vccd1 _3940_/A sky130_fd_sc_hd__xnor2_2
XFILLER_18_3277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2163__A_N _4489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3851_ _3885_/A _3886_/A vssd1 vssd1 vccd1 vccd1 _3888_/A sky130_fd_sc_hd__xnor2_4
XFILLER_35_3591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2802_ _2802_/A _2802_/B vssd1 vssd1 vccd1 vccd1 _2802_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4977__CLK _5013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2733_ _2733_/A _2733_/B vssd1 vssd1 vccd1 vccd1 _4798_/D sky130_fd_sc_hd__xnor2_1
XFILLER_12_2153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_2175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2664_ _4763_/Q _2664_/B vssd1 vssd1 vccd1 vccd1 _4763_/D sky130_fd_sc_hd__xnor2_1
X_4403_ _4429_/CLK _4403_/D fanout192/X vssd1 vssd1 vccd1 vccd1 _4403_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__1944__B _2286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2595_ _4714_/Q _2595_/B vssd1 vssd1 vccd1 vccd1 _4714_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__3217__A _3233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3762__102 _3765__105/A vssd1 vssd1 vccd1 vccd1 _3762__102/Y sky130_fd_sc_hd__inv_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_TE_B
+ _2094_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4334_ _2286_/B _4334_/D _3176__67/Y vssd1 vssd1 vccd1 vccd1 _4334_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_29_2683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout206 fanout207/X vssd1 vssd1 vccd1 vccd1 fanout206/X sky130_fd_sc_hd__clkbuf_2
Xfanout217 fanout219/X vssd1 vssd1 vccd1 vccd1 fanout217/X sky130_fd_sc_hd__clkbuf_4
XFILLER_9_2777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout228 fanout230/X vssd1 vssd1 vccd1 vccd1 fanout228/X sky130_fd_sc_hd__buf_4
XFILLER_25_1802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4265_ _4871_/Q vssd1 vssd1 vccd1 vccd1 _4870_/D sky130_fd_sc_hd__inv_2
Xfanout239 fanout241/X vssd1 vssd1 vccd1 vccd1 fanout239/X sky130_fd_sc_hd__buf_2
XFILLER_29_1993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1960__A _4462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3216_ _3233_/A vssd1 vssd1 vccd1 vccd1 _3216_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_2321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4196_ _4754_/Q vssd1 vssd1 vccd1 vccd1 _4753_/D sky130_fd_sc_hd__inv_2
XFILLER_23_2260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_3871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3147_ _4188_/B _3138_/X _3145_/Y _3146_/X vssd1 vssd1 vccd1 vccd1 _3148_/B sky130_fd_sc_hd__o22a_4
XFILLER_3_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_3893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3078_ _4986_/Q _3078_/B vssd1 vssd1 vccd1 vccd1 _4986_/D sky130_fd_sc_hd__xnor2_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2029_ _4418_/Q _4417_/Q vssd1 vssd1 vccd1 vccd1 _2029_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_32_3219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_2097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_2827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3773__112_A _3776__115/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_2210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_3843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2177__S _4493_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_3520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_3575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__0640_ clkbuf_0__0640_/X vssd1 vssd1 vccd1 vccd1 _3770__109/A sky130_fd_sc_hd__clkbuf_16
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_2_0_clk_master clkbuf_3_3_0_clk_master/A vssd1 vssd1 vccd1 vccd1 _4363_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_2197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_2039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5059_/A fanout215/X vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_5_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_3535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_3607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_2812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_4021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2380_ _4652_/D _4626_/Q _4624_/Q _4623_/Q vssd1 vssd1 vccd1 vccd1 _2418_/A sky130_fd_sc_hd__or4_2
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_4098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4050_ _4544_/Q vssd1 vssd1 vccd1 vccd1 _4545_/D sky130_fd_sc_hd__inv_2
XFILLER_4_2641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_A
+ _4861_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3001_ _3001_/A _3001_/B vssd1 vssd1 vccd1 vccd1 _4948_/D sky130_fd_sc_hd__xnor2_1
Xinput6 comp_high_I[5] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4952_ _4962_/CLK _4952_/D fanout210/X vssd1 vssd1 vccd1 vccd1 _4952_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_73 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5005__CLK _4187_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3500__A _5062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_84 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3903_ _3903_/A _3904_/B vssd1 vssd1 vccd1 vccd1 _4369_/D sky130_fd_sc_hd__xnor2_1
XFILLER_32_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4883_ _3493_/Y _4883_/D _3620_/Y vssd1 vssd1 vccd1 vccd1 _4883_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_32_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_2849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3834_ _4356_/Q vssd1 vssd1 vccd1 vccd1 _3839_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_3859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__1632_ _3172_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__1632_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_9_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1955__A _3931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_2573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4739__RESET_B _3658_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[2\].w1.ro_block_I.ro_pol.tribuf.t_buf _2454_/X _2300_/Y vssd1
+ vssd1 vccd1 vccd1 _5088_/A sky130_fd_sc_hd__ebufn_8
XANTENNA__3873__C _3882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2716_ _4796_/Q _4795_/Q vssd1 vssd1 vccd1 vccd1 _2716_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_31_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3696_ _3696_/A vssd1 vssd1 vccd1 vccd1 _4071_/A sky130_fd_sc_hd__buf_6
XANTENNA_fanout119_A _5062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2647_ _4770_/Q _4769_/Q _4768_/Q _2647_/D vssd1 vssd1 vccd1 vccd1 _2648_/D sky130_fd_sc_hd__and4_1
XANTENNA__3145__A2 _4248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2578_ _4709_/Q _2578_/B vssd1 vssd1 vccd1 vccd1 _4709_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4317_ _4324_/CLK _4317_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _4317_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_2574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_2344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4248_ _4248_/A _4248_/B _4248_/C _4248_/D vssd1 vssd1 vccd1 vccd1 _4250_/B sky130_fd_sc_hd__or4_2
X_3162__62 _3169__65/A vssd1 vssd1 vccd1 vccd1 _3162__62/Y sky130_fd_sc_hd__inv_2
XFILLER_21_2219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_3977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4179_ _4734_/Q vssd1 vssd1 vccd1 vccd1 _4735_/D sky130_fd_sc_hd__inv_2
XFILLER_28_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_2115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2408__A1 _4620_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3410__A _3414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_3049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_4037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3769__108 _3770__109/A vssd1 vssd1 vccd1 vccd1 _3769__108/Y sky130_fd_sc_hd__inv_2
XFILLER_10_3369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_2061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4522__CLK _4533_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_3844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_3877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_4122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4672__CLK _4718_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2696__A _4834_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3304__B _3446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout158/X fanout206/X vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_1_2825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5028__CLK _5030_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_3361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1759__B _5029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__0623_ clkbuf_0__0623_/X vssd1 vssd1 vccd1 vccd1 _3600_/A sky130_fd_sc_hd__clkbuf_16
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1880_ _1909_/A _1880_/B vssd1 vssd1 vccd1 vccd1 _1881_/B sky130_fd_sc_hd__nand2_1
XFILLER_15_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1775__A _2858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3550_ _3550_/A vssd1 vssd1 vccd1 vccd1 _3550_/Y sky130_fd_sc_hd__inv_2
X_2501_ _4674_/Q _4673_/Q _2480_/D _2498_/B vssd1 vssd1 vccd1 vccd1 _2502_/B sky130_fd_sc_hd__a31o_1
X_3481_ _3498_/A vssd1 vssd1 vccd1 vccd1 _3481_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_4077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2432_ _3066_/A _2432_/B _2432_/C _2432_/D vssd1 vssd1 vccd1 vccd1 _2433_/B sky130_fd_sc_hd__and4_2
XFILLER_29_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2335__B1 _2173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2363_ _2608_/A _4590_/Q vssd1 vssd1 vccd1 vccd1 _4590_/D sky130_fd_sc_hd__xor2_1
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
+ _4797_/Q _2785_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_4102_ _4630_/Q vssd1 vssd1 vccd1 vccd1 _4629_/D sky130_fd_sc_hd__inv_2
X_5082_ _5082_/A vssd1 vssd1 vccd1 vccd1 _5082_/X sky130_fd_sc_hd__clkbuf_1
X_2294_ _2286_/X _2293_/X _2294_/B1 vssd1 vssd1 vccd1 vccd1 _2294_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_26_1963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5063_/A fanout251/X vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_0_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3214__B _3847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4033_ _4513_/Q vssd1 vssd1 vccd1 vccd1 _4512_/D sky130_fd_sc_hd__inv_2
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3230__A _3895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4935_ _5030_/CLK _4935_/D fanout224/X vssd1 vssd1 vccd1 vccd1 _4935_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_2613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_2624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3200__8 _3201__9/A vssd1 vssd1 vccd1 vccd1 _4370_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_2012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_2181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2810__A1 _3914_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4866_ _5046_/A _4866_/D fanout228/X vssd1 vssd1 vccd1 vccd1 _4866_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout236_A fanout257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_3792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3817_ _4331_/Q vssd1 vssd1 vccd1 vccd1 _4330_/D sky130_fd_sc_hd__inv_2
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4797_ _4811_/CLK _4797_/D fanout249/X vssd1 vssd1 vccd1 vccd1 _4797_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_2933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3748_ _3748_/A vssd1 vssd1 vccd1 vccd1 _3748_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3679_ _4135_/A vssd1 vssd1 vccd1 vccd1 _3679_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_2371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3405__A _3947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_3835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
+ _4855_/Q _2885_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_2833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf _4316_/Q _1917_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_7_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2317__B1 _1975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3315__A _3891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_2837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_4057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3034__B _4962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_3345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5031__RESET_B fanout226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4904__SET_B fanout236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_3191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2981_ _4940_/Q _4939_/Q vssd1 vssd1 vccd1 vccd1 _2981_/Y sky130_fd_sc_hd__xnor2_4
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4187_/Y _4720_/D _3396_/Y vssd1 vssd1 vccd1 vccd1 _4720_/Q sky130_fd_sc_hd__dfrtp_1
X_1932_ _4352_/D _4353_/Q vssd1 vssd1 vccd1 vccd1 _1933_/B sky130_fd_sc_hd__and2b_1
XFILLER_34_2955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4651_ input20/X input4/X fanout222/X vssd1 vssd1 vccd1 vccd1 _4652_/D sky130_fd_sc_hd__dfrtp_4
X_1863_ _4318_/Q _4317_/Q _4316_/Q _1885_/B vssd1 vssd1 vccd1 vccd1 _1875_/B sky130_fd_sc_hd__or4_1
XFILLER_28_4106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput20 phi1b_dig_I[3] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_4117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput31 phi1b_dig_Q[6] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__buf_6
XFILLER_15_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4582_ _4590_/CLK _4582_/D fanout229/X vssd1 vssd1 vccd1 vccd1 _4582_/Q sky130_fd_sc_hd__dfrtp_2
X_1794_ _1839_/A vssd1 vssd1 vccd1 vccd1 _2922_/A sky130_fd_sc_hd__buf_12
X_3533_ _3550_/A vssd1 vssd1 vccd1 vccd1 _3533_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_2704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_3449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3464_ _3466_/A vssd1 vssd1 vccd1 vccd1 _3464_/Y sky130_fd_sc_hd__inv_2
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout119/X fanout248/X vssd1 vssd1 vccd1 vccd1 _5078_/A sky130_fd_sc_hd__dlrtn_1
X_2415_ _2376_/D _2414_/Y _2344_/X vssd1 vssd1 vccd1 vccd1 _2416_/B sky130_fd_sc_hd__o21ai_1
X_3395_ _3659_/A vssd1 vssd1 vccd1 vccd1 _3414_/A sky130_fd_sc_hd__buf_8
XANTENNA__3225__A _3233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_2533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_3109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_2461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_2544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2346_ _4584_/Q _2346_/B vssd1 vssd1 vccd1 vccd1 _4584_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_1821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_2566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5065_ _5065_/A vssd1 vssd1 vccd1 vccd1 _5065_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_2358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2277_ _4556_/D _4557_/Q vssd1 vssd1 vccd1 vccd1 _2278_/B sky130_fd_sc_hd__and2b_1
XFILLER_26_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout186_A fanout196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4016_ _4478_/Q vssd1 vssd1 vccd1 vccd1 _4479_/D sky130_fd_sc_hd__inv_2
XFILLER_25_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3895__A _3895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4918_ _5013_/CLK _4918_/D _3513_/Y vssd1 vssd1 vccd1 vccd1 _4918_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_4143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4849_ _3475_/Y _4849_/D _3629__81/Y vssd1 vssd1 vccd1 vccd1 _4849_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3135__A _3576_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2974__A _3877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4710__CLK _4712_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_2881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_TE_B
+ _2615_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_2917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_2939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_3807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4860__CLK _4865_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2214__A _4523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_4014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_3521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2553__A3 _2561_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _4511_/Q _4510_/Q vssd1 vssd1 vccd1 vccd1 _2200_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_3_3429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3180_ _3904_/A vssd1 vssd1 vccd1 vccd1 _3420_/B sky130_fd_sc_hd__buf_12
XFILLER_3_2706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_2886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_2645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2131_ _4481_/Q _4480_/Q vssd1 vssd1 vccd1 vccd1 _2131_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_1_3153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4390__CLK _4429_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2062_ _4430_/Q _2062_/B vssd1 vssd1 vccd1 vccd1 _4430_/D sky130_fd_sc_hd__xnor2_1
XFILLER_21_2380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf_TE_B
+ _3053_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_2741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2964_ _4933_/Q _4932_/D vssd1 vssd1 vccd1 vccd1 _2965_/A sky130_fd_sc_hd__and2b_1
XFILLER_34_3497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1915_ _4327_/Q _4326_/Q vssd1 vssd1 vccd1 vccd1 _1915_/Y sky130_fd_sc_hd__xnor2_4
Xclkbuf_1_0__f__1638_ clkbuf_0__1638_/X vssd1 vssd1 vccd1 vccd1 _3264__22/A sky130_fd_sc_hd__clkbuf_16
X_4703_ _3394_/Y _4703_/D _3669_/Y vssd1 vssd1 vccd1 vccd1 _4703_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_30_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_2785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2895_ _4901_/Q _4900_/Q _4899_/Q _2932_/A vssd1 vssd1 vccd1 vccd1 _2918_/B sky130_fd_sc_hd__or4_1
XFILLER_11_2004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2124__A _2286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1846_ _4293_/Q _4292_/Q vssd1 vssd1 vccd1 vccd1 _1846_/Y sky130_fd_sc_hd__xnor2_2
X_4634_ _3350_/Y _4634_/D _3691_/Y vssd1 vssd1 vccd1 vccd1 _4634_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2529__B1 _2518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4565_ _4658_/CLK _4565_/D fanout212/X vssd1 vssd1 vccd1 vccd1 _4565_/Q sky130_fd_sc_hd__dfrtp_2
X_1777_ _4285_/Q _4284_/Q _1777_/C vssd1 vssd1 vccd1 vccd1 _1778_/D sky130_fd_sc_hd__and3_4
XANTENNA__1963__A _4395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3516_ _3934_/A _3933_/A vssd1 vssd1 vccd1 vccd1 _3516_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_1_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4496_ _4532_/CLK _4496_/D fanout211/X vssd1 vssd1 vccd1 vccd1 _4496_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_28_2534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3447_ _3632_/A vssd1 vssd1 vccd1 vccd1 _3466_/A sky130_fd_sc_hd__buf_8
XFILLER_6_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
+ _4616_/Q _2438_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_28_1855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3378_ _4127_/A _4129_/A vssd1 vssd1 vccd1 vccd1 _3378_/Y sky130_fd_sc_hd__xnor2_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2329_ _2922_/A vssd1 vssd1 vccd1 vccd1 _2412_/A sky130_fd_sc_hd__buf_4
XFILLER_3_3996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5048_ _5048_/A vssd1 vssd1 vccd1 vccd1 _5048_/X sky130_fd_sc_hd__buf_2
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_GATE_N
+ _5063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_2505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_A
+ _4393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3009__A1 _4953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2768__B1 _2687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_7_0_clk_master clkbuf_3_7_0_clk_master/A vssd1 vssd1 vccd1 vccd1 _4658_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_11_3261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2969__A _3576_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1873__A _1909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2940__B1 _2858_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_2066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_4141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input31_A phi1b_dig_Q[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_2807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_2818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_2761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4676__RESET_B fanout253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
+ _4674_/Q _2540_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf_A
+ _4425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _4359_/CLK fanout190/X vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1700_ _1761_/B vssd1 vssd1 vccd1 vccd1 _1700_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_31_2958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2680_ _2680_/A _2680_/B vssd1 vssd1 vccd1 vccd1 _2681_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_2379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_3555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_3566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4350_ input17/X input1/X fanout191/X vssd1 vssd1 vccd1 vccd1 _4351_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_9_2904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3301_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3301_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4281_ _4281_/CLK _4281_/D fanout201/X vssd1 vssd1 vccd1 vccd1 _4281_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_29_2887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _3891_/A _3889_/A vssd1 vssd1 vccd1 vccd1 _3232_/Y sky130_fd_sc_hd__xnor2_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3503__A _3519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2114_ _3710_/Y _3737_/Y vssd1 vssd1 vccd1 vccd1 _2114_/Y sky130_fd_sc_hd__nor2_4
X_3094_ _4991_/Q _3094_/B vssd1 vssd1 vccd1 vccd1 _4991_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__3222__B _3442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2045_ _4425_/Q _2045_/B vssd1 vssd1 vccd1 vccd1 _4425_/D sky130_fd_sc_hd__xor2_1
XANTENNA__4346__RESET_B fanout195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_3813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_2246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout149_A _2114_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3996_ _4459_/Q vssd1 vssd1 vccd1 vccd1 _4460_/D sky130_fd_sc_hd__inv_2
XANTENNA__4286__CLK _5040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2947_ _4904_/Q _2947_/B vssd1 vssd1 vccd1 vccd1 _4904_/D sky130_fd_sc_hd__xor2_1
XFILLER_17_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_2435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_2446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2878_ _4871_/Q _4870_/Q vssd1 vssd1 vccd1 vccd1 _2878_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_15_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3892__B _3892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4617_ _4626_/CLK _4617_/D fanout234/X vssd1 vssd1 vccd1 vccd1 _4617_/Q sky130_fd_sc_hd__dfrtp_4
X_1829_ _4284_/Q _1829_/B vssd1 vssd1 vccd1 vccd1 _4284_/D sky130_fd_sc_hd__xnor2_1
XFILLER_12_2891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3574__54 _3656_/A vssd1 vssd1 vccd1 vccd1 _5029_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4548_ _2631_/A _4548_/D _3305_/Y vssd1 vssd1 vccd1 vccd1 _4548_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_3137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_2425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4479_ _3265_/Y _4479_/D _3734__96/Y vssd1 vssd1 vccd1 vccd1 _4479_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_3806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_3975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_2239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3413__A _3912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4629__CLK _4060_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_3470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4779__CLK _4187_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
+ _4389_/Q _2031_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_10_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2211__B _4533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3707__92 _3732__95/A vssd1 vssd1 vccd1 vccd1 _3707__92/Y sky130_fd_sc_hd__inv_2
XFILLER_24_3430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_4017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4857__RESET_B fanout228/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_2834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3323__A _3340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_A
+ _4526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_2533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1778__A _4283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3850_ _4363_/Q vssd1 vssd1 vccd1 vccd1 _3886_/A sky130_fd_sc_hd__buf_8
XFILLER_18_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2801_ _4003_/C _4131_/C _2801_/C vssd1 vssd1 vccd1 vccd1 _2802_/B sky130_fd_sc_hd__nand3_1
XFILLER_32_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_2891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_2733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout136/X fanout238/X vssd1 vssd1 vccd1 vccd1 _5084_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_31_3489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2732_ _2730_/X _2731_/Y _1975_/X vssd1 vssd1 vccd1 vccd1 _2733_/B sky130_fd_sc_hd__o21a_1
XFILLER_31_2777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_4114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2663_ _2680_/A _2663_/B vssd1 vssd1 vccd1 vccd1 _2664_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_4064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_4086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4402_ _4402_/CLK _4402_/D fanout189/X vssd1 vssd1 vccd1 vccd1 _4402_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2402__A _2412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_3205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2594_ _2680_/A _2594_/B vssd1 vssd1 vccd1 vccd1 _2595_/B sky130_fd_sc_hd__nand2_1
XANTENNA__1707__A1 _4190_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4333_ _3175_/Y _4333_/D _3770__109/Y vssd1 vssd1 vccd1 vccd1 _4333_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_3249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout207 fanout220/X vssd1 vssd1 vccd1 vccd1 fanout207/X sky130_fd_sc_hd__clkbuf_4
Xfanout218 fanout219/X vssd1 vssd1 vccd1 vccd1 fanout218/X sky130_fd_sc_hd__clkbuf_4
XFILLER_29_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4264_ _4852_/Q vssd1 vssd1 vccd1 vccd1 _4853_/D sky130_fd_sc_hd__inv_2
Xfanout229 fanout230/X vssd1 vssd1 vccd1 vccd1 fanout229/X sky130_fd_sc_hd__clkbuf_2
X_3215_ _3738_/A vssd1 vssd1 vccd1 vccd1 _3233_/A sky130_fd_sc_hd__buf_6
XFILLER_3_3056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4195_ _4195_/A vssd1 vssd1 vccd1 vccd1 _4748_/D sky130_fd_sc_hd__inv_2
XFILLER_7_2491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_3078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_2333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3233__A _3233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3146_ _4064_/A _4248_/B _3141_/Y _2468_/A vssd1 vssd1 vccd1 vccd1 _3146_/X sky130_fd_sc_hd__a31o_1
XFILLER_20_3883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3077_ _3068_/C _3076_/X _1791_/X vssd1 vssd1 vccd1 vccd1 _3078_/B sky130_fd_sc_hd__o21ai_1
XFILLER_23_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2028_ _4416_/Q _4415_/Q vssd1 vssd1 vccd1 vccd1 _2028_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_23_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4064__A _4064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4921__CLK _3516_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3979_ _4444_/Q vssd1 vssd1 vccd1 vccd1 _4443_/D sky130_fd_sc_hd__inv_2
XFILLER_10_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_2210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1946__A1 _3914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3408__A _3414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_GATE_N
+ _3375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_2161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4301__CLK _3898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2966__B _4933_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_2288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4950__RESET_B fanout210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2123__A1 _2294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_2935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4268__RESET_B _4359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4451__CLK _2286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_2842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3657__86_A _3683__90/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_RESET_B fanout193/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_3569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_2868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output62_A _5059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3000_ _2998_/X _2999_/Y _2143_/A vssd1 vssd1 vccd1 vccd1 _3001_/B sky130_fd_sc_hd__o21a_1
XFILLER_24_2592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4620__RESET_B fanout234/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput7 comp_high_I[6] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4951_ _4962_/CLK _4951_/D fanout208/X vssd1 vssd1 vccd1 vccd1 _4951_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_74 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3684_/A fanout216/X vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__dlrtn_1
XTAP_85 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3902_ _3898_/B _3900_/Y _3910_/B vssd1 vssd1 vccd1 vccd1 _3904_/B sky130_fd_sc_hd__mux2_4
X_4882_ _5013_/CLK _4882_/D _3492_/Y vssd1 vssd1 vccd1 vccd1 _4882_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_3220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3833_ _4355_/Q vssd1 vssd1 vccd1 vccd1 _3838_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_3827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2715_ _4794_/Q _4793_/Q vssd1 vssd1 vccd1 vccd1 _2715_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3695_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3695_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3228__A _3903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4324__CLK _4324_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2132__A _4555_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2646_ _4772_/Q _4771_/Q _2646_/C vssd1 vssd1 vccd1 vccd1 _2647_/D sky130_fd_sc_hd__and3_1
XFILLER_29_3193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2577_ _2680_/A _2577_/B vssd1 vssd1 vccd1 vccd1 _2578_/B sky130_fd_sc_hd__nand2_1
XANTENNA__1971__A _2143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4708__RESET_B fanout247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4316_ _4324_/CLK _4316_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _4316_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_29_2492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4474__CLK _1952_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_3956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4247_ _4247_/A vssd1 vssd1 vccd1 vccd1 _4247_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_19_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4361__RESET_B fanout202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4178_ _4735_/Q vssd1 vssd1 vccd1 vccd1 _4734_/D sky130_fd_sc_hd__inv_2
XFILLER_3_2163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3129_ _3129_/A vssd1 vssd1 vccd1 vccd1 _3129_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2408__A2 _4619_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_4005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_2636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2042__A _4430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_3856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4817__CLK _5007_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_4134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2153__A_N _4486_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4967__CLK _4247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_4030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_2848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3601__A _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output100_A _5097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_1_clk_master clkbuf_1_0_1_clk_master/A vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_2_clk_master/A
+ sky130_fd_sc_hd__clkbuf_8
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_2883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2500_ _4671_/Q _2500_/B vssd1 vssd1 vccd1 vccd1 _4671_/D sky130_fd_sc_hd__xnor2_1
X_3480_ _5062_/A vssd1 vssd1 vccd1 vccd1 _3498_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_13_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_4117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_4056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4497__CLK _4533_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2431_ _4652_/D _4611_/Q vssd1 vssd1 vccd1 vccd1 _2432_/D sky130_fd_sc_hd__xnor2_1
XFILLER_26_3333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1791__A _2858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_3219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2362_ _4589_/Q _2362_/B vssd1 vssd1 vccd1 vccd1 _4589_/D sky130_fd_sc_hd__xor2_1
XFILLER_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_2665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4101_ _4627_/Q vssd1 vssd1 vccd1 vccd1 _4628_/D sky130_fd_sc_hd__inv_2
XFILLER_6_2759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5081_ _5081_/A vssd1 vssd1 vccd1 vccd1 _5081_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_2518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2293_ _3899_/A _3898_/B _3908_/A _3941_/A vssd1 vssd1 vccd1 vccd1 _2293_/X sky130_fd_sc_hd__or4_1
XFILLER_24_3090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4032_ _4510_/Q vssd1 vssd1 vccd1 vccd1 _4511_/D sky130_fd_sc_hd__inv_2
XFILLER_26_1986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_2264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3511__A _3519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3230__B _3372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4934_ _3521_/Y _4934_/D fanout224/X vssd1 vssd1 vccd1 vccd1 _4934_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2127__A _3941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_3359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4865_ _4865_/CLK _4865_/D fanout226/X vssd1 vssd1 vccd1 vccd1 _4865_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_2193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1966__A _4462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3816_ _4328_/Q vssd1 vssd1 vccd1 vccd1 _4329_/D sky130_fd_sc_hd__inv_2
XANTENNA_fanout131_A _5043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A fanout230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4796_ _3446_/Y _4796_/D _3642_/Y vssd1 vssd1 vccd1 vccd1 _4796_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_2923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3747_ _3748_/A vssd1 vssd1 vccd1 vccd1 _3747_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5055_/A fanout244/X vssd1 vssd1 vccd1 vccd1 _5079_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_31_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3678_ _4135_/A vssd1 vssd1 vccd1 vccd1 _3678_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2797__A _3605_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2629_ _3631_/Y _3658_/Y vssd1 vssd1 vccd1 vccd1 _5044_/A sky130_fd_sc_hd__nor2_4
XFILLER_9_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3405__B _3438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_A
+ _4675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_2845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2014__B1 _2003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2565__A1 _4707_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_3653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_TE_B
+ _3120_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4283__RESET_B fanout195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2500__A _4671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3523__49 _3523__49/A vssd1 vssd1 vccd1 vccd1 _4938_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__3315__B _3889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_3302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_3241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_2849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_4069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_GATE_N _5048_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_2540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_A
+ _4707_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3331__A _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_3613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2980_ _4188_/B _2980_/B vssd1 vssd1 vccd1 vccd1 _5070_/A sky130_fd_sc_hd__xnor2_2
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1931_ _1931_/A vssd1 vssd1 vccd1 vccd1 _1933_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4650_ input28/X _4650_/D fanout207/X vssd1 vssd1 vccd1 vccd1 _4650_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_3955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1862_ _4321_/Q _4320_/Q _4319_/Q _1898_/A vssd1 vssd1 vccd1 vccd1 _1885_/B sky130_fd_sc_hd__or4_1
Xinput10 comp_high_Q[1] vssd1 vssd1 vccd1 vccd1 _4461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_3988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3601_ _3656_/A vssd1 vssd1 vccd1 vccd1 _3601_/X sky130_fd_sc_hd__buf_1
Xinput21 phi1b_dig_I[4] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_2
XFILLER_28_4129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1793_ _1793_/A _1793_/B vssd1 vssd1 vccd1 vccd1 _4275_/D sky130_fd_sc_hd__xnor2_1
Xinput32 phi1b_dig_Q[7] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_16
X_4581_ _4590_/CLK _4581_/D fanout227/X vssd1 vssd1 vccd1 vccd1 _4581_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3532_ _3588_/A vssd1 vssd1 vccd1 vccd1 _3550_/A sky130_fd_sc_hd__buf_6
XFILLER_28_3439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3463_ _3924_/A _3923_/A vssd1 vssd1 vccd1 vccd1 _3463_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__3506__A _4189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2414_ _4622_/Q _4621_/Q _2418_/A vssd1 vssd1 vccd1 vccd1 _2414_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__2410__A _4618_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3394_ _3903_/A _3420_/B vssd1 vssd1 vccd1 vccd1 _3394_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_22_3049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_2315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2345_ _2304_/D _2343_/Y _2344_/X vssd1 vssd1 vccd1 vccd1 _2346_/B sky130_fd_sc_hd__o21ai_1
XFILLER_6_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5064_ _5064_/A vssd1 vssd1 vccd1 vccd1 _5064_/X sky130_fd_sc_hd__clkbuf_1
X_2276_ _2276_/A vssd1 vssd1 vccd1 vccd1 _2278_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4015_ _4479_/Q vssd1 vssd1 vccd1 vccd1 _4478_/D sky130_fd_sc_hd__inv_2
XFILLER_0_2122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3241__A _3255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout179_A _3738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4512__CLK _3914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_2083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2492__B1 _1975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
+ _4986_/Q _3120_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_3877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_4111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3895__B _3895_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4917_ _3512_/Y _4917_/D _3610_/Y vssd1 vssd1 vccd1 vccd1 _4917_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4662__CLK _2470_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_2444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4848_ _3865_/Y _4848_/D _3474__45/Y vssd1 vssd1 vccd1 vccd1 _4848_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4779_ _4187_/Y _4779_/D _3429_/Y vssd1 vssd1 vccd1 vccd1 _4779_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3416__A _5060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2320__A _2327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_3611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_3791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_2044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_2055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4247__A _4247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_2929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_3977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_0__1632__A _3172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2214__B _4522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4464__RESET_B fanout198/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_2296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_4037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3326__A _3340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2230__A _2327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_3303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_2793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4535__CLK _3292_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2130_ _4479_/Q _4478_/Q vssd1 vssd1 vccd1 vccd1 _2130_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_1_3121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout180/X fanout184/X vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_21_3060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_3165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2061_ _2061_/A _2061_/B vssd1 vssd1 vccd1 vccd1 _2062_/B sky130_fd_sc_hd__nand2_1
XFILLER_1_2431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3061__A _5024_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_2475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_4133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_4144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_2497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_3465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2963_ _2963_/A vssd1 vssd1 vccd1 vccd1 _2963_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_2753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4702_ _2631_/A _4702_/D _3393_/Y vssd1 vssd1 vccd1 vccd1 _4702_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_1_0__f__1637_ clkbuf_0__1637_/X vssd1 vssd1 vccd1 vccd1 _3199__7/A sky130_fd_sc_hd__clkbuf_16
X_1914_ _2608_/A _4325_/Q vssd1 vssd1 vccd1 vccd1 _4325_/D sky130_fd_sc_hd__xor2_1
XFILLER_31_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_2163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2894_ _4931_/D _4905_/Q _4903_/Q _4902_/Q vssd1 vssd1 vccd1 vccd1 _2932_/A sky130_fd_sc_hd__or4_2
XFILLER_34_2797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_2174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_2639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4633_ _5013_/CLK _4633_/D _3349_/Y vssd1 vssd1 vccd1 vccd1 _4633_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_3796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1845_ _4291_/Q _4290_/Q vssd1 vssd1 vccd1 vccd1 _1845_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__2124__B _3941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_4009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4564_ _4564_/CLK _4564_/D fanout223/X vssd1 vssd1 vccd1 vccd1 _4564_/Q sky130_fd_sc_hd__dfrtp_4
X_1776_ _4347_/D _4289_/Q _4287_/Q _4286_/Q vssd1 vssd1 vccd1 vccd1 _1777_/C sky130_fd_sc_hd__and4_1
XFILLER_28_3225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3515_ _3519_/A vssd1 vssd1 vccd1 vccd1 _3515_/Y sky130_fd_sc_hd__inv_2
X_4495_ _4533_/CLK _4495_/D fanout205/X vssd1 vssd1 vccd1 vccd1 _4495_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3236__A _3255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3446_ _3905_/A _3446_/B vssd1 vssd1 vccd1 vccd1 _3446_/Y sky130_fd_sc_hd__xnor2_2
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3377_ _3393_/A vssd1 vssd1 vccd1 vccd1 _3377_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2328_ _4579_/Q _2328_/B vssd1 vssd1 vccd1 vccd1 _4579_/D sky130_fd_sc_hd__xnor2_1
XFILLER_23_3892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5047_ _5047_/A vssd1 vssd1 vccd1 vccd1 _5047_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2259_ _2327_/A _2259_/B vssd1 vssd1 vccd1 vccd1 _2260_/B sky130_fd_sc_hd__nand2_1
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3009__A2 _4952_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_2241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2969__B _3605_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3152__116 _3784__125/A vssd1 vssd1 vccd1 vccd1 _3152__116/Y sky130_fd_sc_hd__inv_2
XANTENNA__4558__CLK input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_2911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_2139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2985__A _5020_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input24_A phi1b_dig_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_4117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_2773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_2715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf_TE_B
+ _2716_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2225__A _4523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_3059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_2937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_2336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_2369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output92_A _5089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3056__A _4994_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3300_ _3925_/A _3442_/B vssd1 vssd1 vccd1 vccd1 _3300_/Y sky130_fd_sc_hd__xnor2_1
X_4280_ _4281_/CLK _4280_/D fanout199/X vssd1 vssd1 vccd1 vccd1 _4280_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_2949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_2899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_3205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _3233_/A vssd1 vssd1 vccd1 vccd1 _3231_/Y sky130_fd_sc_hd__inv_2
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _4363_/CLK fanout192/X vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_23_2487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2113_ _2113_/A vssd1 vssd1 vccd1 vccd1 _2113_/X sky130_fd_sc_hd__clkbuf_1
X_3093_ _3109_/A _3093_/B vssd1 vssd1 vccd1 vccd1 _3094_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_2498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2044_ _2143_/A _2091_/B _2091_/C vssd1 vssd1 vccd1 vccd1 _2045_/B sky130_fd_sc_hd__and3_1
XFILLER_23_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_3825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3995_ _4460_/Q vssd1 vssd1 vccd1 vccd1 _4459_/D sky130_fd_sc_hd__inv_2
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3643_/A fanout243/X vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__2135__A _4488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2946_ _3112_/A _2946_/B _2946_/C _2946_/D vssd1 vssd1 vccd1 vccd1 _2947_/B sky130_fd_sc_hd__and4_1
X_2877_ _3114_/A _4869_/Q vssd1 vssd1 vccd1 vccd1 _4869_/D sky130_fd_sc_hd__xor2_1
XANTENNA__3892__C _3901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4616_ _4626_/CLK _4616_/D fanout232/X vssd1 vssd1 vccd1 vccd1 _4616_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout211_A fanout212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1828_ _1909_/A _1828_/B vssd1 vssd1 vccd1 vccd1 _1829_/B sky130_fd_sc_hd__nand2_1
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf _4278_/Q _1849_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_30_1746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2789__B _4836_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4700__CLK _4852_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_3105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4547_ _3304_/Y _4547_/D _3714_/Y vssd1 vssd1 vccd1 vccd1 _4547_/Q sky130_fd_sc_hd__dfrtp_1
X_1759_ _5028_/Q _5029_/Q vssd1 vssd1 vccd1 vccd1 _1760_/A sky130_fd_sc_hd__xor2_1
XFILLER_25_3921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4478_ _1952_/A1 _4478_/D _3264__22/Y vssd1 vssd1 vccd1 vccd1 _4478_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_8_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_2448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3429_ _3445_/A vssd1 vssd1 vccd1 vccd1 _3429_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4850__CLK _4852_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_3998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_2161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3413__B _3446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
+ _4805_/Q _2777_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_2325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3262__21 _3262__21/A vssd1 vssd1 vccd1 vccd1 _3262__21/Y sky130_fd_sc_hd__inv_2
XFILLER_32_3947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_2369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2045__A _4425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1949__C1 _3892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5091__A _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2677__B1 _2518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4897__RESET_B fanout231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_4125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2800_ _3877_/A _4063_/B _4124_/D vssd1 vssd1 vccd1 vccd1 _2800_/X sky130_fd_sc_hd__or3_1
XFILLER_18_2589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_2881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2731_ _4799_/Q _2731_/B vssd1 vssd1 vccd1 vccd1 _2731_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_2745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1794__A _1839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_TE_B
+ _2265_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_4126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2662_ _4764_/Q _2658_/C _2659_/B vssd1 vssd1 vccd1 vccd1 _2663_/B sky130_fd_sc_hd__a21bo_1
XFILLER_12_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4401_ _4402_/CLK _4401_/D fanout188/X vssd1 vssd1 vccd1 vccd1 _4401_/Q sky130_fd_sc_hd__dfrtp_1
X_2593_ _2592_/Y _2549_/C _4715_/Q vssd1 vssd1 vccd1 vccd1 _2594_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_2713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_3217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4332_ _3931_/A _4332_/D _3173__66/Y vssd1 vssd1 vccd1 vccd1 _4332_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_2674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_2757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout208 fanout220/X vssd1 vssd1 vccd1 vccd1 fanout208/X sky130_fd_sc_hd__buf_4
XFILLER_29_1951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout219 fanout220/X vssd1 vssd1 vccd1 vccd1 fanout219/X sky130_fd_sc_hd__buf_2
X_4263_ _4853_/Q vssd1 vssd1 vccd1 vccd1 _4852_/D sky130_fd_sc_hd__inv_2
XFILLER_29_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3514__A _3946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2117__C1 _3892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3214_ _3848_/A _3847_/A vssd1 vssd1 vccd1 vccd1 _3214_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_5_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4194_ _4751_/Q _4194_/B vssd1 vssd1 vccd1 vccd1 _4752_/D sky130_fd_sc_hd__xor2_1
X_3145_ _4064_/A _4248_/B _3139_/Y vssd1 vssd1 vccd1 vccd1 _3145_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_2284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3659_/A fanout240/X vssd1 vssd1 vccd1 vccd1 _5076_/A sky130_fd_sc_hd__dlrtn_1
X_3076_ _4987_/Q _3076_/B vssd1 vssd1 vccd1 vccd1 _3076_/X sky130_fd_sc_hd__and2b_1
XFILLER_3_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2027_ _4414_/Q _4413_/Q vssd1 vssd1 vccd1 vccd1 _2027_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout161_A _4000_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_2011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4064__B _4064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3423__40_A _3425__41/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3978_ _4441_/Q vssd1 vssd1 vccd1 vccd1 _4442_/D sky130_fd_sc_hd__inv_2
X_2929_ _4901_/Q _4900_/Q _2932_/A vssd1 vssd1 vccd1 vccd1 _2929_/Y sky130_fd_sc_hd__nor3_1
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
+ _4520_/Q _2271_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_10_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1946__A2 _2286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_TE_B
+ _2709_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_2288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_2140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3424__A _3896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_3709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2123__A2 _3914_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4990__RESET_B fanout236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4746__CLK input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2831__B1 _2143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4896__CLK _4901_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5086__A _5086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2503__A _4672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3334__A _3340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
+ _4578_/Q _2369_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_4_3355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_A
+ _4989_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4276__CLK _4281_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_2621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput8 comp_high_I[7] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XFILLER_4_1964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4950_ _4962_/CLK _4950_/D fanout210/X vssd1 vssd1 vccd1 vccd1 _4950_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_75 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3901_ _3901_/A _3901_/B vssd1 vssd1 vccd1 vccd1 _3910_/B sky130_fd_sc_hd__nor2_1
XTAP_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4881_ _3491_/Y _4881_/D _3621_/Y vssd1 vssd1 vccd1 vccd1 _4881_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_2375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3832_ _4344_/Q vssd1 vssd1 vccd1 vccd1 _4345_/D sky130_fd_sc_hd__inv_2
XFILLER_14_2217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3509__A _3519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2413__A _4619_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2714_ _4792_/Q _4791_/Q vssd1 vssd1 vccd1 vccd1 _2714_/Y sky130_fd_sc_hd__xnor2_4
X_3694_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3694_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3228__B _3420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2132__B _4497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2645_ _4834_/D _4776_/Q _4774_/Q _4773_/Q vssd1 vssd1 vccd1 vccd1 _2646_/C sky130_fd_sc_hd__and4_1
XFILLER_31_1885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_3161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_3003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2576_ _4710_/Q _2551_/D _2568_/B vssd1 vssd1 vccd1 vccd1 _2577_/B sky130_fd_sc_hd__a21bo_1
XFILLER_9_3277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_2460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_2543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4619__CLK _4626_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4315_ _5040_/A _4315_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _4315_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_2313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3244__A _3925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4246_ _4249_/A _4250_/A vssd1 vssd1 vccd1 vccd1 _4247_/A sky130_fd_sc_hd__xnor2_4
XFILLER_25_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4177_ _4732_/Q vssd1 vssd1 vccd1 vccd1 _4733_/D sky130_fd_sc_hd__inv_2
XFILLER_25_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4769__CLK _4812_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3898__B _3898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3128_ _3128_/A _3128_/B vssd1 vssd1 vccd1 vccd1 _3129_/A sky130_fd_sc_hd__or2_1
XANTENNA__1699__A _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_2980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3059_ _4984_/Q vssd1 vssd1 vccd1 vccd1 _3071_/A sky130_fd_sc_hd__inv_2
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_4017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_4028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_3813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2977__B _2977_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4299__CLK _3914_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4489__RESET_B fanout201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_4020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_2799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_3341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_4086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_3374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_3249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3329__A _3947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3759__99 _3759__99/A vssd1 vssd1 vccd1 vccd1 _3759__99/Y sky130_fd_sc_hd__inv_2
XANTENNA__2233__A _2327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_2294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3048__B _4969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2583__A2 _4712_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_4107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_4129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_4068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2430_ _4624_/Q _2430_/B vssd1 vssd1 vccd1 vccd1 _4624_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_3417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_3367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2361_ _3066_/A _2361_/B _2361_/C _2361_/D vssd1 vssd1 vccd1 vccd1 _2362_/B sky130_fd_sc_hd__and4_1
XFILLER_26_2644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_3389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3064__A _4988_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4100_ _4628_/Q vssd1 vssd1 vccd1 vccd1 _4627_/D sky130_fd_sc_hd__inv_2
XFILLER_4_3141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5080_ _5080_/A vssd1 vssd1 vccd1 vccd1 _5080_/X sky130_fd_sc_hd__clkbuf_1
X_2292_ _4068_/S _2292_/B vssd1 vssd1 vccd1 vccd1 _5094_/A sky130_fd_sc_hd__xnor2_1
XFILLER_26_2688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3999__A _4001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4031_ _4511_/Q vssd1 vssd1 vccd1 vccd1 _4510_/D sky130_fd_sc_hd__inv_2
XFILLER_4_3185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4841__RESET_B fanout228/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_2210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_3990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_clk_master clkbuf_2_1_0_clk_master/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_clk_master/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_2337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_4028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4933_ input23/X _4933_/D fanout218/X vssd1 vssd1 vccd1 vccd1 _4933_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4864_ _4865_/CLK _4864_/D fanout228/X vssd1 vssd1 vccd1 vccd1 _4864_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_2659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3815_ _4329_/Q vssd1 vssd1 vccd1 vccd1 _4328_/D sky130_fd_sc_hd__inv_2
XFILLER_21_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4795_ _4852_/CLK _4795_/D _3445_/Y vssd1 vssd1 vccd1 vccd1 _4795_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3239__A _3255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2143__A _2143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3746_ _3748_/A vssd1 vssd1 vccd1 vccd1 _3746_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout124_A _4712_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_2372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4441__CLK _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3677_ _4135_/A vssd1 vssd1 vccd1 vccd1 _3677_/Y sky130_fd_sc_hd__inv_2
X_2628_ _2628_/A vssd1 vssd1 vccd1 vccd1 _2628_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_3085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2559_ _2996_/A _2606_/B _2606_/C vssd1 vssd1 vccd1 vccd1 _2560_/B sky130_fd_sc_hd__and3_1
XANTENNA__4591__CLK _4248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_0__0624__A _3600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4229_ _4817_/Q vssd1 vssd1 vccd1 vccd1 _4818_/D sky130_fd_sc_hd__inv_2
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3702__A _4071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3775__114 _3776__115/A vssd1 vssd1 vccd1 vccd1 _3775__114/Y sky130_fd_sc_hd__inv_2
XFILLER_15_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2798__C1 _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2053__A _4430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2565__A2 _2561_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2988__A _4953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4934__CLK _3521_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_3529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3612__A _3616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_2657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3331__B _3440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4314__CLK _4324_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_3193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__1653_ clkbuf_0__1653_/X vssd1 vssd1 vccd1 vccd1 _3523__49/A sky130_fd_sc_hd__clkbuf_16
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1930_ _4353_/Q _4352_/D vssd1 vssd1 vccd1 vccd1 _1931_/A sky130_fd_sc_hd__and2b_1
XFILLER_32_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4464__CLK input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1861_ _4351_/D _4325_/Q _4323_/Q _4322_/Q vssd1 vssd1 vccd1 vccd1 _1898_/A sky130_fd_sc_hd__or4_1
XFILLER_30_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3600_ _3600_/A vssd1 vssd1 vccd1 vccd1 _3600_/X sky130_fd_sc_hd__buf_1
XANTENNA__3204__12_A _3201__9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput11 comp_high_Q[2] vssd1 vssd1 vccd1 vccd1 _4554_/D sky130_fd_sc_hd__clkbuf_1
Xinput22 phi1b_dig_I[5] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_4
X_4580_ _4590_/CLK _4580_/D fanout227/X vssd1 vssd1 vccd1 vccd1 _4580_/Q sky130_fd_sc_hd__dfrtp_2
X_1792_ _1789_/X _1790_/Y _1791_/X vssd1 vssd1 vccd1 vccd1 _1793_/B sky130_fd_sc_hd__o21a_1
X_3211__16 _3264__22/A vssd1 vssd1 vccd1 vccd1 _3211__16/Y sky130_fd_sc_hd__inv_2
XANTENNA__4718__SET_B fanout242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput33 rstb vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_12
X_3531_ _3916_/A _3915_/A vssd1 vssd1 vccd1 vccd1 _3531_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_10_3691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3365__31 _3365__31/A vssd1 vssd1 vccd1 vccd1 _4659_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3462_ _3466_/A vssd1 vssd1 vccd1 vccd1 _3462_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3506__B _4190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2413_ _4619_/Q _2413_/B vssd1 vssd1 vccd1 vccd1 _4619_/D sky130_fd_sc_hd__xnor2_1
X_3393_ _3393_/A vssd1 vssd1 vccd1 vccd1 _3393_/Y sky130_fd_sc_hd__inv_2
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
+ _4397_/Q _2023_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout157/X fanout203/X vssd1 vssd1 vccd1 vccd1 _5082_/A sky130_fd_sc_hd__dlrtn_1
X_2344_ _2858_/A vssd1 vssd1 vccd1 vccd1 _2344_/X sky130_fd_sc_hd__buf_6
XFILLER_26_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5063_ _5063_/A vssd1 vssd1 vccd1 vccd1 _5063_/X sky130_fd_sc_hd__clkbuf_1
X_2275_ _4557_/Q _4556_/D vssd1 vssd1 vccd1 vccd1 _2276_/A sky130_fd_sc_hd__and2b_1
XFILLER_6_1856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4014_ _4476_/Q vssd1 vssd1 vccd1 vccd1 _4477_/D sky130_fd_sc_hd__inv_2
XFILLER_22_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1819__A1 _4283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_2040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_2292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2138__A _4555_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_3135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout241_A fanout257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4916_ _4916_/CLK _4916_/D _3511_/Y vssd1 vssd1 vccd1 vccd1 _4916_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4847_ _3473_/Y _4847_/D _3630__82/Y vssd1 vssd1 vccd1 vccd1 _4847_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_2478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4778_ _4247_/A _4778_/D _3652_/Y vssd1 vssd1 vccd1 vccd1 _4778_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_2743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_3488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_2765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3729_ _4010_/A vssd1 vssd1 vccd1 vccd1 _3729_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_2776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4763__RESET_B fanout247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3365__31_A _3365__31/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3371__34 _3469__42/A vssd1 vssd1 vccd1 vccd1 _3371__34/Y sky130_fd_sc_hd__inv_2
XFILLER_27_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2180__B1 _2173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_TE_B
+ _2783_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_3667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3432__A _4127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_2988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_4023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4487__CLK _5042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_2665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1994__B1 _1823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3607__A _3616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_2811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_2614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3342__A _3696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2060_ _4431_/Q _2036_/D _2053_/B vssd1 vssd1 vccd1 vccd1 _2061_/B sky130_fd_sc_hd__a21bo_1
XFILLER_1_3177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_A
+ _4489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1797__A _3114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2962_ _2962_/A _2962_/B vssd1 vssd1 vccd1 vccd1 _2963_/A sky130_fd_sc_hd__or2_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1913_ _4324_/Q _1913_/B vssd1 vssd1 vccd1 vccd1 _4324_/D sky130_fd_sc_hd__xor2_1
X_4701_ _3392_/Y _4701_/D _3671_/Y vssd1 vssd1 vccd1 vccd1 _4701_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_2765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2893_ _4893_/Q _4892_/Q _2901_/C _2904_/A vssd1 vssd1 vccd1 vccd1 _2946_/B sky130_fd_sc_hd__a31o_1
XFILLER_11_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4632_ _3348_/Y _4632_/D _3692_/Y vssd1 vssd1 vccd1 vccd1 _4632_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1844_ _4289_/Q _2608_/A vssd1 vssd1 vccd1 vccd1 _4289_/D sky130_fd_sc_hd__xor2_1
XFILLER_30_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4563_ _5030_/CLK _4563_/D fanout223/X vssd1 vssd1 vccd1 vccd1 _4563_/Q sky130_fd_sc_hd__dfrtp_4
X_1775_ _2858_/A vssd1 vssd1 vccd1 vccd1 _2143_/A sky130_fd_sc_hd__buf_12
XFILLER_11_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3749_/A fanout187/X vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__3517__A _3519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3514_ _3946_/A _3945_/A vssd1 vssd1 vccd1 vccd1 _3514_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__1963__C _4393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4494_ _5034_/A _4494_/D fanout202/X vssd1 vssd1 vccd1 vccd1 _4494_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_28_1802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2140__B _4489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3445_ _3445_/A vssd1 vssd1 vccd1 vccd1 _3445_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_3033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _3393_/A vssd1 vssd1 vccd1 vccd1 _3376_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2327_ _2327_/A _2327_/B vssd1 vssd1 vccd1 vccd1 _2328_/B sky130_fd_sc_hd__nand2_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3252__A _3895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5046_ _5046_/A vssd1 vssd1 vccd1 vccd1 _5046_/X sky130_fd_sc_hd__clkbuf_1
X_2258_ _4559_/D _4533_/Q vssd1 vssd1 vccd1 vccd1 _2259_/B sky130_fd_sc_hd__xnor2_1
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2189_ _4495_/Q _2189_/B vssd1 vssd1 vccd1 vccd1 _4495_/D sky130_fd_sc_hd__xnor2_1
XFILLER_22_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3009__A3 _2988_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_3697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1976__B1 _1975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_GATE_N
+ fanout128/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout120/X fanout249/X vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__3427__A _3632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2331__A _2412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_3793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2985__B _4962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_4129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input17_A phi1b_dig_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5089__A _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3337__A _3912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_2061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1783__C _4283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_2812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4502__CLK _4063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4614__RESET_B fanout234/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_2845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_4087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_4098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _3895_/A _3372_/B vssd1 vssd1 vccd1 vccd1 _3230_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_7_2630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4652__CLK input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2112_ _2112_/A _2112_/B vssd1 vssd1 vccd1 vccd1 _2113_/A sky130_fd_sc_hd__or2_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3092_ _4992_/Q _3057_/D _3085_/B vssd1 vssd1 vccd1 vccd1 _3093_/B sky130_fd_sc_hd__a21bo_1
XFILLER_23_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2043_ _4427_/Q _2047_/B _2049_/A vssd1 vssd1 vccd1 vccd1 _2091_/C sky130_fd_sc_hd__o21ai_1
XFILLER_1_2295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2416__A _4620_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3994_ _4457_/Q vssd1 vssd1 vccd1 vccd1 _4458_/D sky130_fd_sc_hd__inv_2
XFILLER_14_3837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2945_ _4931_/D _4890_/Q vssd1 vssd1 vccd1 vccd1 _2946_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__2135__B _4487_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2876_ _4868_/Q _2876_/B vssd1 vssd1 vccd1 vccd1 _4868_/D sky130_fd_sc_hd__xor2_1
XFILLER_30_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1827_ _1826_/Y _1777_/C _4285_/Q vssd1 vssd1 vccd1 vccd1 _1828_/B sky130_fd_sc_hd__mux2_1
X_4615_ _4626_/CLK _4615_/D fanout232/X vssd1 vssd1 vccd1 vccd1 _4615_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_2871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3247__A _3255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4546_ _4852_/CLK _4546_/D _3303_/Y vssd1 vssd1 vccd1 vccd1 _4546_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout204_A fanout207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1758_ _5017_/Q vssd1 vssd1 vccd1 vccd1 _5018_/D sky130_fd_sc_hd__inv_2
XFILLER_28_2322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4477_ _3263_/Y _4477_/D _3735__97/Y vssd1 vssd1 vccd1 vccd1 _4477_/Q sky130_fd_sc_hd__dfrtp_1
X_1689_ _4919_/Q vssd1 vssd1 vccd1 vccd1 _4918_/D sky130_fd_sc_hd__inv_2
XANTENNA__1990__A _2061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3428_ _3445_/A vssd1 vssd1 vccd1 vccd1 _3428_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
+ _4890_/Q _2957_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_24_1507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input9_A comp_high_Q[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3359_ _3361_/A vssd1 vssd1 vccd1 vccd1 _3359_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_3751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_2173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5029_ _5029_/CLK _5029_/D fanout223/X vssd1 vssd1 vccd1 vccd1 _5029_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3710__A _5058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4525__CLK _4533_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2061__A _2061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4675__CLK _4717_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2996__A _2996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_3673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0__1638__A _3205_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_2639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3620__A _4256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_2502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
+ _4948_/Q _3052_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_18_2546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_4137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_3414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4866__RESET_B fanout228/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2730_ _4800_/Q _4799_/Q _2730_/C vssd1 vssd1 vccd1 vccd1 _2730_/X sky130_fd_sc_hd__and3_1
XFILLER_9_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_2757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2661_ _2661_/A _2661_/B vssd1 vssd1 vccd1 vccd1 _4762_/D sky130_fd_sc_hd__xnor2_1
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4400_ _4402_/CLK _4400_/D fanout186/X vssd1 vssd1 vccd1 vccd1 _4400_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_4138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_3415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2592_ _2592_/A vssd1 vssd1 vccd1 vccd1 _2592_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_2631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4331_ _3171_/Y _4331_/D _3771__110/Y vssd1 vssd1 vccd1 vccd1 _4331_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_3229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_2725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4262_ _4850_/Q vssd1 vssd1 vccd1 vccd1 _4851_/D sky130_fd_sc_hd__inv_2
Xfanout209 fanout220/X vssd1 vssd1 vccd1 vccd1 fanout209/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_2769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3514__B _3945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4193_ _4752_/Q _4194_/B vssd1 vssd1 vccd1 vccd1 _4751_/D sky130_fd_sc_hd__xor2_1
XFILLER_23_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_2252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_3841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3144_ _3144_/A _3144_/B vssd1 vssd1 vccd1 vccd1 _5099_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_3935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3075_ _4988_/Q _3075_/B vssd1 vssd1 vccd1 vccd1 _3076_/B sky130_fd_sc_hd__nor2_1
XANTENNA__1969__B _4393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2026_ _4412_/Q _4411_/Q vssd1 vssd1 vccd1 vccd1 _2026_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout154_A _4981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_2023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4548__CLK _2631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3977_ _4442_/Q vssd1 vssd1 vccd1 vccd1 _4441_/D sky130_fd_sc_hd__inv_2
XANTENNA__1985__A _4392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_4070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_2370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_3970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_2392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2928_ _4898_/Q _2928_/B vssd1 vssd1 vccd1 vccd1 _4898_/D sky130_fd_sc_hd__xnor2_1
XFILLER_31_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4698__CLK _2807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2859_ _2818_/D _2857_/Y _2858_/X vssd1 vssd1 vccd1 vccd1 _2860_/B sky130_fd_sc_hd__o21ai_1
XFILLER_30_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4529_ _4532_/CLK _4529_/D fanout213/X vssd1 vssd1 vccd1 vccd1 _4529_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_8_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3705__A _4071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3314__26 _3365__31/A vssd1 vssd1 vccd1 vccd1 _3314__26/Y sky130_fd_sc_hd__inv_2
XANTENNA__3424__B _3904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3440__A _3934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4277__RESET_B fanout201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_4002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3615__A _3616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_2826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_3389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_2644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_3159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3320__29 _3365__31/A vssd1 vssd1 vccd1 vccd1 _3320__29/Y sky130_fd_sc_hd__inv_2
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_A
+ _4670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_2677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 comp_high_Q[0] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3350__A _3947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_76 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_4081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3900_ _3900_/A _3900_/B vssd1 vssd1 vccd1 vccd1 _3900_/Y sky130_fd_sc_hd__nand2_1
XTAP_87 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4880_ _4916_/CLK _4880_/D _3490_/Y vssd1 vssd1 vccd1 vccd1 _4880_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_3200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3831_ _4345_/Q vssd1 vssd1 vccd1 vccd1 _4344_/D sky130_fd_sc_hd__inv_2
XFILLER_18_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_2387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4840__CLK input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_2229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_3255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2713_ _4790_/Q _4789_/Q vssd1 vssd1 vccd1 vccd1 _2713_/Y sky130_fd_sc_hd__xnor2_4
X_3693_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3693_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2644_ _4760_/Q _4759_/Q vssd1 vssd1 vccd1 vccd1 _2644_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__4990__CLK _4997_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_3173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2575_ _4708_/Q _2575_/B vssd1 vssd1 vccd1 vccd1 _4708_/D sky130_fd_sc_hd__xnor2_1
XFILLER_29_2450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3525__A _3916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_3109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4314_ _4324_/CLK _4314_/D fanout191/X vssd1 vssd1 vccd1 vccd1 _4314_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3244__B _3442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4245_ _4843_/Q vssd1 vssd1 vccd1 vccd1 _4250_/A sky130_fd_sc_hd__buf_6
XFILLER_22_3947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3768__107_A _3770__109/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4176_ _4733_/Q vssd1 vssd1 vccd1 vccd1 _4732_/D sky130_fd_sc_hd__inv_2
XFILLER_0_3721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3127_ _5021_/D _5022_/Q vssd1 vssd1 vccd1 vccd1 _3128_/B sky130_fd_sc_hd__and2b_1
XFILLER_20_3693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1699__B _3556_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3058_ _4989_/Q _4988_/Q _4987_/Q _3058_/D vssd1 vssd1 vccd1 vccd1 _3068_/C sky130_fd_sc_hd__and4_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_4121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2009_ _4399_/Q _2009_/B vssd1 vssd1 vccd1 vccd1 _4399_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__4717__RESET_B fanout255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_2741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_2042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_2785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3435__A _3445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
+ _4709_/Q _2612_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_25_3582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_3665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4713__CLK _4717_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2993__B _4954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_2734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_2745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3170__A _3923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_4043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4863__CLK _4865_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2804__A1 _3914_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_3217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5097__A _5097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3329__B _3438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_4003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_3313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3345__A _3361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2360_ _4648_/D _4575_/Q vssd1 vssd1 vccd1 vccd1 _2361_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_2656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2291_ _2294_/B1 _3932_/A _2286_/X _2290_/X vssd1 vssd1 vccd1 vccd1 _2292_/B sky130_fd_sc_hd__o31a_1
XFILLER_26_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_2678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4393__CLK _4402_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4030_ _4508_/Q vssd1 vssd1 vccd1 vccd1 _4509_/D sky130_fd_sc_hd__inv_2
XFILLER_4_2430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3999__B _4005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3080__A _3109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_2255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4932_ input23/X _4932_/D fanout218/X vssd1 vssd1 vccd1 vccd1 _4933_/D sky130_fd_sc_hd__dfrtp_1
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
+ _4767_/Q _2709_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_33_3317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4863_ _4865_/CLK _4863_/D fanout226/X vssd1 vssd1 vccd1 vccd1 _4863_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_2184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3814_ _4326_/Q vssd1 vssd1 vccd1 vccd1 _4327_/D sky130_fd_sc_hd__clkinv_2
XANTENNA__2424__A _4652_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4794_ _3444_/Y _4794_/D _3644_/Y vssd1 vssd1 vccd1 vccd1 _4794_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3745_ _3748_/A vssd1 vssd1 vccd1 vccd1 _3745_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_2947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout117_A _4803_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3676_ _4135_/A vssd1 vssd1 vccd1 vccd1 _3676_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2627_ _2627_/A _2627_/B vssd1 vssd1 vccd1 vccd1 _2628_/A sky130_fd_sc_hd__or2_1
XFILLER_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3255__A _3255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4736__CLK _4852_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2558_ _4706_/Q _2562_/B _2564_/A vssd1 vssd1 vccd1 vccd1 _2606_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_3097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_2396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2489_ _4668_/Q _2489_/B vssd1 vssd1 vccd1 vccd1 _4668_/D sky130_fd_sc_hd__xor2_1
XFILLER_22_3755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_3849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4228_ _4818_/Q vssd1 vssd1 vccd1 vccd1 _4817_/D sky130_fd_sc_hd__inv_2
XANTENNA__4886__CLK _4981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4159_ _4698_/Q vssd1 vssd1 vccd1 vccd1 _4699_/D sky130_fd_sc_hd__inv_2
XANTENNA__3262__21_A _3262__21/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
+ _4439_/Q _2103_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_15_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4266__CLK _3883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2053__B _2053_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_2593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2988__B _4952_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3165__A _3947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_3677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_2807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4609__CLK _2470_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1860_ _4313_/Q _4312_/Q _1868_/C _1871_/A vssd1 vssd1 vccd1 vccd1 _1912_/B sky130_fd_sc_hd__a31o_1
XANTENNA__2244__A _4526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1791_ _2858_/A vssd1 vssd1 vccd1 vccd1 _1791_/X sky130_fd_sc_hd__buf_12
Xinput12 comp_high_Q[3] vssd1 vssd1 vccd1 vccd1 _4647_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput23 phi1b_dig_I[6] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_6
XFILLER_13_2070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput34 ud_en vssd1 vssd1 vccd1 vccd1 _1839_/A sky130_fd_sc_hd__buf_12
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
+ _4482_/Q _2202_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__4759__CLK _2631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3461_ _3934_/A _3933_/A vssd1 vssd1 vccd1 vccd1 _3461_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_26_3121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_2729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3075__A _4988_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2412_ _2412_/A _2412_/B vssd1 vssd1 vccd1 vccd1 _2413_/B sky130_fd_sc_hd__nand2_1
X_3392_ _3912_/A _3446_/B vssd1 vssd1 vccd1 vccd1 _3392_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_26_3165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2343_ _4586_/Q _4585_/Q _2347_/A vssd1 vssd1 vccd1 vccd1 _2343_/Y sky130_fd_sc_hd__nor3_1
XFILLER_26_2486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5062_ _5062_/A vssd1 vssd1 vccd1 vccd1 _5062_/X sky130_fd_sc_hd__clkbuf_1
X_2274_ _4553_/Q _4552_/Q vssd1 vssd1 vccd1 vccd1 _2274_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_6_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4013_ _4477_/Q vssd1 vssd1 vccd1 vccd1 _4476_/D sky130_fd_sc_hd__inv_2
XANTENNA__1819__A2 _1778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2138__B _4497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_3813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4915_ _3510_/Y _4915_/D _3611_/Y vssd1 vssd1 vccd1 vccd1 _4915_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4289__CLK _5040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_2424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4846_ _4852_/CLK _4846_/D _3472__44/Y vssd1 vssd1 vccd1 vccd1 _4846_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout234_A fanout235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_3445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4777_ _4247_/Y _4777_/D _3428_/Y vssd1 vssd1 vccd1 vccd1 _4777_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_2891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout158/X fanout205/X vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__dlrtn_1
X_1989_ _4395_/Q _1963_/D _1982_/B vssd1 vssd1 vccd1 vccd1 _1990_/B sky130_fd_sc_hd__a21bo_1
X_3728_ _4010_/A vssd1 vssd1 vccd1 vccd1 _3728_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_2788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3659_ _3659_/A vssd1 vssd1 vccd1 vccd1 _3669_/A sky130_fd_sc_hd__buf_6
XFILLER_28_3975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_2182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2180__A1 _2133_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3713__A _3721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_2068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3432__B _4129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2329__A _2922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_2873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_4002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_4013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4901__CLK _4901_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5063_/A fanout251/X vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_22_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_2265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_4142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_4028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3623__A _4256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_2626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_2637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4431__CLK _5033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3417__36 _3425__41/A vssd1 vssd1 vccd1 vccd1 _4750_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2961_ _4928_/D _4929_/Q vssd1 vssd1 vccd1 vccd1 _2962_/B sky130_fd_sc_hd__and2b_1
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4700_ _4852_/CLK _4700_/D _3391_/Y vssd1 vssd1 vccd1 vccd1 _4700_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1912_ _3066_/A _1912_/B _1912_/C _1912_/D vssd1 vssd1 vccd1 vccd1 _1913_/B sky130_fd_sc_hd__and4_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4581__CLK _4590_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2892_ _4891_/Q vssd1 vssd1 vccd1 vccd1 _2904_/A sky130_fd_sc_hd__inv_2
XFILLER_30_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_2007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4631_ _4916_/CLK _4631_/D _3347_/Y vssd1 vssd1 vccd1 vccd1 _4631_/Q sky130_fd_sc_hd__dfrtp_1
X_1843_ _2143_/A vssd1 vssd1 vccd1 vccd1 _2608_/A sky130_fd_sc_hd__buf_12
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1774_ _1839_/A vssd1 vssd1 vccd1 vccd1 _2858_/A sky130_fd_sc_hd__buf_12
X_4562_ _3311_/Y _4562_/D fanout222/X vssd1 vssd1 vccd1 vccd1 _4562_/Q sky130_fd_sc_hd__dfrtp_1
X_3513_ _3519_/A vssd1 vssd1 vccd1 vccd1 _3513_/Y sky130_fd_sc_hd__inv_2
X_4493_ _4533_/CLK _4493_/D fanout208/X vssd1 vssd1 vccd1 vccd1 _4493_/Q sky130_fd_sc_hd__dfrtp_4
X_3444_ _3916_/A _3444_/B vssd1 vssd1 vccd1 vccd1 _3444_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__2140__C _4488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _3375_/A vssd1 vssd1 vccd1 vccd1 _3393_/A sky130_fd_sc_hd__buf_8
XFILLER_6_2322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3533__A _3550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ _4581_/Q _4580_/Q _2305_/D _2323_/B vssd1 vssd1 vccd1 vccd1 _2327_/B sky130_fd_sc_hd__a31o_1
XFILLER_3_3955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3252__B _3372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5045_ _5045_/A vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__clkbuf_1
X_2257_ _4530_/Q _2257_/B vssd1 vssd1 vccd1 vccd1 _4530_/D sky130_fd_sc_hd__xnor2_1
XFILLER_2_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2188_ _2327_/A _2188_/B vssd1 vssd1 vccd1 vccd1 _2189_/B sky130_fd_sc_hd__nand2_1
XANTENNA__1988__A _4393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_TE_B
+ _2442_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4924__CLK _4943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_3529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_2221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_2265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4829_ _4943_/CLK _4829_/D _3464_/Y vssd1 vssd1 vccd1 vccd1 _4829_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_2563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4304__CLK _2294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_2014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_3603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4984__RESET_B fanout232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_3669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3443__A _3445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3102__B1 _1791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3524__50_A _3528__52/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout119/X fanout248/X vssd1 vssd1 vccd1 vccd1 _5078_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5019__RESET_B fanout214/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3618__A _4256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3337__B _3446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_2879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output78_A _5075_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3353__A _3361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_A
+ _4952_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_2445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2111_ _4467_/D _4468_/Q vssd1 vssd1 vccd1 vccd1 _2112_/B sky130_fd_sc_hd__and2b_1
X_3091_ _4990_/Q _3091_/B vssd1 vssd1 vccd1 vccd1 _4990_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__4947__CLK _4962_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2042_ _4430_/Q _4429_/Q _4428_/Q _2053_/B vssd1 vssd1 vccd1 vccd1 _2047_/B sky130_fd_sc_hd__or4_1
XFILLER_3_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_2227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3993_ _4458_/Q vssd1 vssd1 vccd1 vccd1 _4457_/D sky130_fd_sc_hd__inv_2
XFILLER_34_3275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2944_ _4903_/Q _2944_/B vssd1 vssd1 vccd1 vccd1 _4903_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__2135__C _4486_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2875_ _3112_/A _2875_/B _2875_/C _2875_/D vssd1 vssd1 vccd1 vccd1 _2876_/B sky130_fd_sc_hd__and4_1
XANTENNA__2432__A _3066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4614_ _4623_/CLK _4614_/D fanout234/X vssd1 vssd1 vccd1 vccd1 _4614_/Q sky130_fd_sc_hd__dfrtp_4
X_1826_ _1826_/A vssd1 vssd1 vccd1 vccd1 _1826_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwrapper_cell_loop\[4\].w1.ro_block_Q.ro_pol.tribuf.t_buf _2791_/X _2641_/Y vssd1
+ vssd1 vccd1 vccd1 _5090_/A sky130_fd_sc_hd__ebufn_8
X_4545_ _3302_/Y _4545_/D _3715_/Y vssd1 vssd1 vccd1 vccd1 _4545_/Q sky130_fd_sc_hd__dfrtp_1
X_1757_ _5018_/Q vssd1 vssd1 vccd1 vccd1 _5017_/D sky130_fd_sc_hd__inv_2
XFILLER_11_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4476_ _1952_/A1 _4476_/D _3262__21/Y vssd1 vssd1 vccd1 vccd1 _4476_/Q sky130_fd_sc_hd__dfrtp_1
X_1688_ _4916_/Q vssd1 vssd1 vccd1 vccd1 _4917_/D sky130_fd_sc_hd__inv_2
X_3427_ _3632_/A vssd1 vssd1 vccd1 vccd1 _3445_/A sky130_fd_sc_hd__buf_8
XFILLER_28_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_3809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3263__A _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3192__74 _3193__75/A vssd1 vssd1 vccd1 vccd1 _4356_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_2141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3358_ _3912_/A _3446_/B vssd1 vssd1 vccd1 vccd1 _3358_/Y sky130_fd_sc_hd__xnor2_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _4586_/Q _4585_/Q _4584_/Q _2347_/A vssd1 vssd1 vccd1 vccd1 _2333_/B sky130_fd_sc_hd__or4_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_2196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3289_ _5058_/A vssd1 vssd1 vccd1 vccd1 _3309_/A sky130_fd_sc_hd__buf_6
XFILLER_2_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5028_ _5030_/CLK _5028_/D fanout214/X vssd1 vssd1 vccd1 vccd1 _5028_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_2349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_3949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1949__A1 _3888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_2625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_2658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3438__A _3946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_3685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2126__A1 _3877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_2890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_2826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_2583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[6\].w1.ro_block_Q.ro_pol.tribuf.t_buf_A _3129_/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3628__80 _3655__85/A vssd1 vssd1 vccd1 vccd1 _3628__80/Y sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__0637_ clkbuf_0__0637_/X vssd1 vssd1 vccd1 vccd1 _3759__99/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__1778__D _1778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3348__A _4004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_2769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2660_ _2658_/X _2659_/Y _1975_/X vssd1 vssd1 vccd1 vccd1 _2661_/B sky130_fd_sc_hd__o21a_1
XFILLER_29_4045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_4056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2591_ _4713_/Q _2591_/B vssd1 vssd1 vccd1 vccd1 _4713_/D sky130_fd_sc_hd__xnor2_1
XFILLER_29_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4330_ _3932_/A _4330_/D _3169__65/Y vssd1 vssd1 vccd1 vccd1 _4330_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_2737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_2518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4261_ _4851_/Q vssd1 vssd1 vccd1 vccd1 _4850_/D sky130_fd_sc_hd__inv_2
XFILLER_29_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3083__A _3109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2117__A1 _2286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3212_ _3848_/A _3847_/A vssd1 vssd1 vccd1 vccd1 _3212_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_GATE_N
+ _3576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4192_ _4064_/B _4066_/B _4192_/S vssd1 vssd1 vccd1 vccd1 _4194_/B sky130_fd_sc_hd__mux2_1
XANTENNA__3682__89_A _3683__90/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3143_ _4248_/B _3138_/X _3140_/Y _3142_/X vssd1 vssd1 vccd1 vccd1 _3144_/B sky130_fd_sc_hd__o22a_2
XFILLER_23_2264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3074_ _4985_/Q _3074_/B vssd1 vssd1 vccd1 vccd1 _4985_/D sky130_fd_sc_hd__xnor2_1
XFILLER_1_2060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2025_ _4410_/Q _4409_/Q vssd1 vssd1 vccd1 vccd1 _2025_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__1969__C _4392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_3050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_2057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout147_A _4429_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3976_ _4423_/Q vssd1 vssd1 vccd1 vccd1 _4424_/D sky130_fd_sc_hd__inv_2
XFILLER_17_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_2202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2927_ _3030_/A _2927_/B vssd1 vssd1 vccd1 vccd1 _2928_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_2809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2858_ _2858_/A vssd1 vssd1 vccd1 vccd1 _2858_/X sky130_fd_sc_hd__buf_6
XFILLER_15_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4576__RESET_B fanout226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1809_ _4279_/Q _1809_/B vssd1 vssd1 vccd1 vccd1 _4279_/D sky130_fd_sc_hd__xnor2_1
X_2789_ _4835_/D _4836_/Q vssd1 vssd1 vccd1 vccd1 _2790_/B sky130_fd_sc_hd__and2b_1
XFILLER_2_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4528_ _4533_/CLK _4528_/D fanout209/X vssd1 vssd1 vccd1 vccd1 _4528_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_2131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4459_ _1952_/A1 _4459_/D _3255_/Y vssd1 vssd1 vccd1 vccd1 _4459_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_3753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5056_/A fanout190/X vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_8_2258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_2905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3721__A _3721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3440__B _3440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_3779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3168__A _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2072__A _2178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_3517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2800__A _3877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_2838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_2849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_4069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_2601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3631__A _5061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3350__B _3438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2247__A _4527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3474__45 _3528__52/A vssd1 vssd1 vccd1 vccd1 _3474__45/Y sky130_fd_sc_hd__inv_2
XFILLER_33_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_77 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_88 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_3089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3830_ _4342_/Q vssd1 vssd1 vccd1 vccd1 _4343_/D sky130_fd_sc_hd__inv_2
XFILLER_33_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_3966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_3977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_3999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2712_ _4788_/Q _4787_/Q vssd1 vssd1 vccd1 vccd1 _2712_/Y sky130_fd_sc_hd__xnor2_4
Xwrapper_cell_loop\[6\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf _3128_/A _2982_/Y vssd1
+ vssd1 vccd1 vccd1 _5091_/A sky130_fd_sc_hd__ebufn_8
X_3692_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3692_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3195__3 _3199__7/A vssd1 vssd1 vccd1 vccd1 _4360_/CLK sky130_fd_sc_hd__inv_2
X_2643_ _4758_/Q _4757_/Q vssd1 vssd1 vccd1 vccd1 _2643_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_29_3130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2132__D _4494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2574_ _2680_/A _2574_/B vssd1 vssd1 vccd1 vccd1 _2575_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_3185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4313_ _5040_/A _4313_/D fanout185/X vssd1 vssd1 vccd1 vccd1 _4313_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__3525__B _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_2473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_2567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4244_ _4842_/Q vssd1 vssd1 vccd1 vccd1 _4249_/A sky130_fd_sc_hd__buf_6
XFILLER_29_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4175_ _4730_/Q vssd1 vssd1 vccd1 vccd1 _4731_/D sky130_fd_sc_hd__inv_2
XFILLER_3_2133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3541__A _4127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3126_ _3126_/A vssd1 vssd1 vccd1 vccd1 _3128_/A sky130_fd_sc_hd__buf_2
XFILLER_3_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_2199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2157__A _2178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3057_ _4992_/Q _4991_/Q _4990_/Q _3057_/D vssd1 vssd1 vccd1 vccd1 _3058_/D sky130_fd_sc_hd__and4_2
XFILLER_3_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2008_ _2061_/A _2008_/B vssd1 vssd1 vccd1 vccd1 _2009_/B sky130_fd_sc_hd__nand2_1
XFILLER_14_4133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4665__CLK _3372_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3959_ _4408_/Q vssd1 vssd1 vccd1 vccd1 _4407_/D sky130_fd_sc_hd__inv_2
XFILLER_10_3329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_2753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_2628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_2797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_3804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3716__A _3721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2042__D _2053_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2964__A_N _4933_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_3677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout136/X fanout238/X vssd1 vssd1 vccd1 vccd1 _5084_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_24_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2993__C _4953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3451__A _4189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2501__A1 _4674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2067__A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_2517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_3598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4427__RESET_B fanout194/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_2263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3626__A _4256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_4037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_3325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4538__CLK _4063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_2729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2290_ _3941_/B _2288_/Y _2289_/X _1937_/Y vssd1 vssd1 vccd1 vccd1 _2290_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_29_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_2420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3361__A _3361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_2464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4688__CLK _1765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf _4313_/Q _1920_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XANTENNA__2256__B1 _2173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4931_ input23/X _4931_/D fanout225/X vssd1 vssd1 vccd1 vccd1 _4932_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_20_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4862_ _4865_/CLK _4862_/D fanout224/X vssd1 vssd1 vccd1 vccd1 _4862_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_3741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_2005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3813_ _4327_/Q vssd1 vssd1 vccd1 vccd1 _4326_/D sky130_fd_sc_hd__inv_2
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4793_ _4943_/CLK _4793_/D _3443_/Y vssd1 vssd1 vccd1 vccd1 _4793_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_3638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_2049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3744_ _3748_/A vssd1 vssd1 vccd1 vccd1 _3744_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_2959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3675_ _4135_/A vssd1 vssd1 vccd1 vccd1 _3675_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3536__A _3550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput100 _5097_/X vssd1 vssd1 vccd1 vccd1 sin_out[5] sky130_fd_sc_hd__buf_2
XFILLER_9_3021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2626_ _4746_/D _4747_/Q vssd1 vssd1 vccd1 vccd1 _2627_/B sky130_fd_sc_hd__and2b_1
XFILLER_9_3032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2557_ _4709_/Q _4708_/Q _4707_/Q _2568_/B vssd1 vssd1 vccd1 vccd1 _2562_/B sky130_fd_sc_hd__or4_2
XFILLER_9_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_2123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2488_ _2996_/A _2535_/B _2535_/C vssd1 vssd1 vccd1 vccd1 _2489_/B sky130_fd_sc_hd__and3_1
X_4227_ _4815_/Q vssd1 vssd1 vccd1 vccd1 _4816_/D sky130_fd_sc_hd__inv_2
XFILLER_22_3767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_2178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3271__A _3287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4158_ _4699_/Q vssd1 vssd1 vccd1 vccd1 _4698_/D sky130_fd_sc_hd__inv_2
XFILLER_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3109_ _3109_/A _3109_/B vssd1 vssd1 vccd1 vccd1 _3110_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_3585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4089_ _4599_/Q vssd1 vssd1 vccd1 vccd1 _4600_/D sky130_fd_sc_hd__inv_2
XFILLER_16_3516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2798__A1 _3929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_2447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2988__C _4951_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3446__A _3905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3165__B _3438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3684_/A fanout216/X vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_3441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3181__A _3903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_2795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_3605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
+ _4898_/Q _2949_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_1_1958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4679__RESET_B fanout255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2244__B _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_3947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_2369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_2661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1790_ _4276_/Q _1790_/B vssd1 vssd1 vccd1 vccd1 _1790_/Y sky130_fd_sc_hd__nor2_1
Xinput13 comp_high_Q[4] vssd1 vssd1 vccd1 vccd1 _4740_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput24 phi1b_dig_I[7] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_6
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3356__A _3917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3460_ _3466_/A vssd1 vssd1 vccd1 vccd1 _3460_/Y sky130_fd_sc_hd__inv_2
X_2411_ _4620_/Q _2376_/D _2404_/B vssd1 vssd1 vccd1 vccd1 _2412_/B sky130_fd_sc_hd__a21bo_1
XFILLER_26_3133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3391_ _3393_/A vssd1 vssd1 vccd1 vccd1 _3391_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_2421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2342_ _4583_/Q _2342_/B vssd1 vssd1 vccd1 vccd1 _4583_/D sky130_fd_sc_hd__xnor2_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5061_ _5061_/A vssd1 vssd1 vccd1 vccd1 _5061_/X sky130_fd_sc_hd__clkbuf_1
X_2273_ _4551_/Q _4550_/Q vssd1 vssd1 vccd1 vccd1 _2273_/Y sky130_fd_sc_hd__xnor2_1
X_4012_ _4474_/Q vssd1 vssd1 vccd1 vccd1 _4475_/D sky130_fd_sc_hd__inv_2
XFILLER_4_2261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_3803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4914_ _1765_/A _4914_/D _3509_/Y vssd1 vssd1 vccd1 vccd1 _4914_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4349__RESET_B fanout195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_4125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_2436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4845_ _4845_/CLK _4845_/D fanout218/X vssd1 vssd1 vccd1 vccd1 _4845_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4776_ _4812_/CLK _4776_/D fanout253/X vssd1 vssd1 vccd1 vccd1 _4776_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_3457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout227_A fanout230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1988_ _4393_/Q _1988_/B vssd1 vssd1 vccd1 vccd1 _4393_/D sky130_fd_sc_hd__xnor2_1
XFILLER_14_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_2745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3727_ _4010_/A vssd1 vssd1 vccd1 vccd1 _3727_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3266__A _3600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2170__A _2178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3658_ _5060_/A vssd1 vssd1 vccd1 vccd1 _3658_/Y sky130_fd_sc_hd__inv_2
X_2609_ _4721_/Q _4720_/Q vssd1 vssd1 vccd1 vccd1 _2609_/Y sky130_fd_sc_hd__xnor2_2
X_3589_ _3597_/A vssd1 vssd1 vccd1 vccd1 _3589_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_clk_master clkbuf_0_clk_master/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_clk_master/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_6_3761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_3625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_3575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_2896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_4047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_GATE_N _4359_/CLK
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4772__RESET_B fanout253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_4058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_3357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4383__CLK _3845_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_2981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
+ _4613_/Q _2441_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_12_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_2233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_4110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_4007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3904__A _3904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_2649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout190 fanout193/X vssd1 vssd1 vccd1 vccd1 fanout190/X sky130_fd_sc_hd__buf_2
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_4103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5055_/A fanout244/X vssd1 vssd1 vccd1 vccd1 _5079_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_34_4136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2255__A _4559_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2960_ _2960_/A vssd1 vssd1 vccd1 vccd1 _2962_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4442__RESET_B _3747_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4726__CLK _4916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_2280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1911_ _4351_/D _4310_/Q vssd1 vssd1 vccd1 vccd1 _1912_/D sky130_fd_sc_hd__xnor2_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2891_ _4896_/Q _4895_/Q _4894_/Q _2891_/D vssd1 vssd1 vccd1 vccd1 _2901_/C sky130_fd_sc_hd__and4_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_3891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4630_ _3346_/Y _4630_/D _3693_/Y vssd1 vssd1 vccd1 vccd1 _4630_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1842_ _4288_/Q _1842_/B vssd1 vssd1 vccd1 vccd1 _4288_/D sky130_fd_sc_hd__xor2_1
X_4561_ input19/X _4561_/D fanout213/X vssd1 vssd1 vccd1 vccd1 _4561_/Q sky130_fd_sc_hd__dfrtp_1
X_1773_ _4273_/Q _4272_/Q vssd1 vssd1 vccd1 vccd1 _1773_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__4876__CLK _4248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3512_ _4001_/A _4005_/A vssd1 vssd1 vccd1 vccd1 _3512_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_7_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4492_ _5042_/A _4492_/D fanout200/X vssd1 vssd1 vccd1 vccd1 _4492_/Q sky130_fd_sc_hd__dfrtp_2
X_3443_ _3445_/A vssd1 vssd1 vccd1 vccd1 _3443_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3173__66_A _3193__75/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2698__B1 _2687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _4368_/Q _4367_/Q vssd1 vssd1 vccd1 vccd1 _3374_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_3_3901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_3079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
+ _4671_/Q _2543_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2325_ _4578_/Q _2325_/B vssd1 vssd1 vccd1 vccd1 _4578_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5044_/A vssd1 vssd1 vccd1 vccd1 _5044_/X sky130_fd_sc_hd__clkbuf_1
X_2256_ _2254_/X _2255_/Y _2173_/X vssd1 vssd1 vccd1 vccd1 _2257_/B sky130_fd_sc_hd__o21ai_1
XFILLER_26_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_2080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2187_ _4555_/D _4497_/Q vssd1 vssd1 vccd1 vccd1 _2188_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout177_A _3857_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2405__A_N _4618_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2165__A _4488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_2233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3417__36_A _3425__41/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4828_ _3463_/Y _4828_/D _3634_/Y vssd1 vssd1 vccd1 vccd1 _4828_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_2277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4759_ _2631_/A _4759_/D _3425__41/Y vssd1 vssd1 vccd1 vccd1 _4759_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_27_2004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_3773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3724__A _4010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3734__96 _3759__99/A vssd1 vssd1 vccd1 vccd1 _3734__96/Y sky130_fd_sc_hd__inv_2
XFILLER_24_2925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_3580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_4084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4953__RESET_B fanout214/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4749__CLK _5030_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_3165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4899__CLK _4901_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_2486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_3504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_4001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_2085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3634__A _3642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4279__CLK _4281_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2110_ _2110_/A vssd1 vssd1 vccd1 vccd1 _2112_/A sky130_fd_sc_hd__clkbuf_1
X_3090_ _3109_/A _3090_/B vssd1 vssd1 vccd1 vccd1 _3091_/B sky130_fd_sc_hd__nand2_1
X_2041_ _4433_/Q _4432_/Q _4431_/Q _2063_/B vssd1 vssd1 vccd1 vccd1 _2053_/B sky130_fd_sc_hd__or4_2
XANTENNA__4623__RESET_B fanout236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_2253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3992_ _4455_/Q vssd1 vssd1 vccd1 vccd1 _4456_/D sky130_fd_sc_hd__inv_2
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_2531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2943_ _3030_/A _2943_/B vssd1 vssd1 vccd1 vccd1 _2944_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_3107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2874_ _4927_/D _4854_/Q vssd1 vssd1 vccd1 vccd1 _2875_/D sky130_fd_sc_hd__xnor2_1
XANTENNA_wrapper_cell_loop\[5\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf_TE_B _2813_/Y
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4613_ _4623_/CLK _4613_/D fanout231/X vssd1 vssd1 vccd1 vccd1 _4613_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1825_ _4283_/Q _1825_/B vssd1 vssd1 vccd1 vccd1 _4283_/D sky130_fd_sc_hd__xnor2_1
XFILLER_12_2851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2432__B _2432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4350__D input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4544_ _2807_/A _4544_/D _3301_/Y vssd1 vssd1 vccd1 vccd1 _4544_/Q sky130_fd_sc_hd__dfrtp_1
X_1756_ _5015_/Q vssd1 vssd1 vccd1 vccd1 _5016_/D sky130_fd_sc_hd__inv_2
XFILLER_8_3119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4475_ _3261_/Y _4475_/D _3736__98/Y vssd1 vssd1 vccd1 vccd1 _4475_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_2407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1687_ _4917_/Q vssd1 vssd1 vccd1 vccd1 _4916_/D sky130_fd_sc_hd__inv_2
XANTENNA__3544__A _3550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3426_ _3896_/A _3904_/A vssd1 vssd1 vccd1 vccd1 _3426_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_2368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3263__B _3886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3357_ _3361_/A vssd1 vssd1 vccd1 vccd1 _3357_/Y sky130_fd_sc_hd__inv_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _4648_/D _4590_/Q _4588_/Q _4587_/Q vssd1 vssd1 vccd1 vccd1 _2347_/A sky130_fd_sc_hd__or4_2
XFILLER_6_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3288_ _3891_/A _3889_/A vssd1 vssd1 vccd1 vccd1 _3288_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_2_2039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5027_ _3573_/Y _5027_/D fanout237/X vssd1 vssd1 vccd1 vccd1 _5027_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_6_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2239_ _4527_/Q _4526_/Q _2207_/D _2236_/B vssd1 vssd1 vccd1 vccd1 _2240_/B sky130_fd_sc_hd__a31o_1
XANTENNA__3096__B1 _1791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4364__RESET_B fanout199/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_3917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3719__A _3721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1949__A2 _3898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout180/X fanout184/X vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_2085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3438__B _3438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_2962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_2973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_4113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4421__CLK _2294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3454__A _3466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_3664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_3445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4571__CLK _3855_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_2849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input22_A phi1b_dig_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3901__B _3901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_3296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3087__B1 _1791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1702__A _4247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
+ _4432_/Q _2095_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_13_3861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3348__B _3491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_4107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2590_ _2550_/D _2589_/Y _2518_/X vssd1 vssd1 vccd1 vccd1 _2591_/B sky130_fd_sc_hd__o21ai_1
XANTENNA_output90_A _5087_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4260_ _4848_/Q vssd1 vssd1 vccd1 vccd1 _4849_/D sky130_fd_sc_hd__inv_2
XANTENNA__4914__CLK _1765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2494__B1_N _2491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4191_ _4752_/Q _4751_/Q vssd1 vssd1 vccd1 vccd1 _4192_/S sky130_fd_sc_hd__xnor2_2
X_3142_ _4064_/A _4188_/B _3141_/Y _2468_/A vssd1 vssd1 vccd1 vccd1 _3142_/X sky130_fd_sc_hd__a31o_1
XFILLER_7_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4195__A _4195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3073_ _3109_/A _3073_/B vssd1 vssd1 vccd1 vccd1 _3074_/B sky130_fd_sc_hd__nand2_1
X_2024_ _4408_/Q _4407_/Q vssd1 vssd1 vccd1 vccd1 _2024_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_18_3761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3975_ _4424_/Q vssd1 vssd1 vccd1 vccd1 _4423_/D sky130_fd_sc_hd__inv_2
XFILLER_17_2069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3539__A _4189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_3669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2926_ _4899_/Q _2890_/D _2918_/B vssd1 vssd1 vccd1 vccd1 _2927_/B sky130_fd_sc_hd__a21bo_1
XFILLER_30_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2857_ _4865_/Q _4864_/Q _2861_/A vssd1 vssd1 vccd1 vccd1 _2857_/Y sky130_fd_sc_hd__nor3_1
XFILLER_30_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1808_ _3114_/A _1808_/B vssd1 vssd1 vccd1 vccd1 _1809_/B sky130_fd_sc_hd__nand2_1
X_2788_ _2788_/A vssd1 vssd1 vccd1 vccd1 _2790_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4527_ _5034_/A _4527_/D fanout203/X vssd1 vssd1 vccd1 vccd1 _4527_/Q sky130_fd_sc_hd__dfrtp_2
X_1739_ _5000_/Q vssd1 vssd1 vccd1 vccd1 _4999_/D sky130_fd_sc_hd__inv_2
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3274__A _3947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4458_ _3254_/Y _4458_/D _3739_/Y vssd1 vssd1 vccd1 vccd1 _4458_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
+ _4490_/Q _2194_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_3409_ _3925_/A _3442_/B vssd1 vssd1 vccd1 vccd1 _3409_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_2198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4389_ _4429_/CLK _4389_/D fanout192/X vssd1 vssd1 vccd1 vccd1 _4389_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3449__A _4249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2353__A _4648_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3168__B _3440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _4363_/CLK fanout191/X vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_30_3460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_TE_B
+ _2095_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4937__CLK _3598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2800__B _4063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3184__A _3895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_4059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3643_/A fanout243/X vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__4286__RESET_B fanout194/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_3106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3912__A _3912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2528__A _4741_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4317__CLK _4324_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_2392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_3035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_4061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_78 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_89 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4467__CLK input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_2209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3359__A _3361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2711_ _4786_/Q _4785_/Q vssd1 vssd1 vccd1 vccd1 _2711_/Y sky130_fd_sc_hd__xnor2_4
X_3691_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3691_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2642_ _4756_/Q _4755_/Q vssd1 vssd1 vccd1 vccd1 _2642_/Y sky130_fd_sc_hd__xnor2_2
X_2573_ _4710_/Q _4709_/Q _2551_/D _2569_/B vssd1 vssd1 vccd1 vccd1 _2574_/B sky130_fd_sc_hd__a31o_1
XANTENNA__3094__A _4991_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4312_ _5040_/A _4312_/D fanout185/X vssd1 vssd1 vccd1 vccd1 _4312_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__3373__35_A _3469__42/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_3905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4243_ _4831_/Q vssd1 vssd1 vccd1 vccd1 _4832_/D sky130_fd_sc_hd__inv_2
XFILLER_9_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[3\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf _2622_/A _2474_/Y vssd1
+ vssd1 vccd1 vccd1 _5091_/A sky130_fd_sc_hd__ebufn_8
XFILLER_22_3949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4174_ _4731_/Q vssd1 vssd1 vccd1 vccd1 _4730_/D sky130_fd_sc_hd__inv_2
XANTENNA__3541__B _4129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_2145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3125_ _5022_/Q _5021_/D vssd1 vssd1 vccd1 vccd1 _3126_/A sky130_fd_sc_hd__and2b_1
XFILLER_23_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_2950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3056_ _4994_/Q _4993_/Q _3056_/C vssd1 vssd1 vccd1 vccd1 _3057_/D sky130_fd_sc_hd__and3_1
XFILLER_3_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_2109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2007_ _2006_/Y _1961_/C _4400_/Q vssd1 vssd1 vccd1 vccd1 _2008_/B sky130_fd_sc_hd__mux2_1
XANTENNA_fanout257_A input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_3411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3269__A _4469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2173__A _2858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3958_ _4405_/Q vssd1 vssd1 vccd1 vccd1 _4406_/D sky130_fd_sc_hd__clkinv_2
XFILLER_32_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_2765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2909_ _4894_/Q _2909_/B vssd1 vssd1 vccd1 vccd1 _2909_/X sky130_fd_sc_hd__and2b_1
X_3889_ _3889_/A _3891_/B vssd1 vssd1 vccd1 vccd1 _4365_/D sky130_fd_sc_hd__xnor2_1
XFILLER_8_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_3562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_2850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_4081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_2872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3451__B _4190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_2643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_3511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_3555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2083__A _4466_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_2821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_2220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2811__A _4126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_3897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3659_/A fanout241/X vssd1 vssd1 vccd1 vccd1 _5076_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__2789__A_N _4835_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3642__A _3642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_2371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2258__A _4559_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4930_ input23/X input7/X fanout236/X vssd1 vssd1 vccd1 vccd1 _4931_/D sky130_fd_sc_hd__dfrtp_4
Xclkbuf_1_1_2_clk_master clkbuf_1_1_2_clk_master/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clk_master/A
+ sky130_fd_sc_hd__clkbuf_8
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4861_ _4865_/CLK _4861_/D fanout224/X vssd1 vssd1 vccd1 vccd1 _4861_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_18_2153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_3753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_2175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_3021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3812_ _4308_/Q vssd1 vssd1 vccd1 vccd1 _4309_/D sky130_fd_sc_hd__inv_2
XFILLER_18_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4792_ _3442_/Y _4792_/D _3645_/Y vssd1 vssd1 vccd1 vccd1 _4792_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3743_ _3748_/A vssd1 vssd1 vccd1 vccd1 _3743_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3674_ _4135_/A vssd1 vssd1 vccd1 vccd1 _3674_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4890__RESET_B fanout237/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2625_ _2625_/A vssd1 vssd1 vccd1 vccd1 _2627_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput101 _5098_/X vssd1 vssd1 vccd1 vccd1 sin_out[6] sky130_fd_sc_hd__buf_2
XFILLER_12_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_2321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2556_ _4712_/Q _4711_/Q _4710_/Q _2579_/B vssd1 vssd1 vccd1 vccd1 _2568_/B sky130_fd_sc_hd__or4_2
XFILLER_9_2365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2487_ _4670_/Q _2491_/B _2493_/A vssd1 vssd1 vccd1 vccd1 _2535_/C sky130_fd_sc_hd__o21ai_1
XFILLER_26_3893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4226_ _4816_/Q vssd1 vssd1 vccd1 vccd1 _4815_/D sky130_fd_sc_hd__inv_2
XFILLER_22_3779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4157_ _4696_/Q vssd1 vssd1 vccd1 vccd1 _4697_/D sky130_fd_sc_hd__inv_2
XFILLER_21_1309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2168__A _4489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3108_ _5024_/D _4998_/Q vssd1 vssd1 vccd1 vccd1 _3109_/B sky130_fd_sc_hd__xnor2_1
X_4088_ _4600_/Q vssd1 vssd1 vccd1 vccd1 _4599_/D sky130_fd_sc_hd__inv_2
X_3039_ _3109_/A _3039_/B vssd1 vssd1 vccd1 vccd1 _3040_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_3528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_2139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3727__A _4010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2631__A _2631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2988__D _2988_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3446__B _3446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4560__RESET_B fanout210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_4143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2722__A2 _4799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3462__A _3466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
+ _4983_/Q _3123_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_8_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3181__B _3420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1710__A _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_0_clk_master_A clk_master vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_2640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4648__RESET_B fanout208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_2673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput14 comp_high_Q[5] vssd1 vssd1 vccd1 vccd1 _4833_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3637__A _3642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput25 phi1b_dig_Q[0] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3356__B _3444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_2971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2410_ _4618_/Q _2410_/B vssd1 vssd1 vccd1 vccd1 _4618_/D sky130_fd_sc_hd__xnor2_1
X_3390_ _3917_/A _3444_/B vssd1 vssd1 vccd1 vccd1 _3390_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_26_3145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2174__B1 _2173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_2505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2341_ _2412_/A _2341_/B vssd1 vssd1 vccd1 vccd1 _2342_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_3189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_2527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5060_ _5060_/A vssd1 vssd1 vccd1 vccd1 _5060_/X sky130_fd_sc_hd__clkbuf_1
X_2272_ _4549_/Q _4548_/Q vssd1 vssd1 vccd1 vccd1 _2272_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4011_ _4475_/Q vssd1 vssd1 vccd1 vccd1 _4474_/D sky130_fd_sc_hd__inv_2
XFILLER_22_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2138__D _4494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2229__A1 _4524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4913_ _3508_/Y _4913_/D _3612_/Y vssd1 vssd1 vccd1 vccd1 _4913_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_3859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_3149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4844_ _5030_/CLK _4844_/D fanout218/X vssd1 vssd1 vccd1 vccd1 _4844_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_4137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_3583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_3594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4775_ _4811_/CLK _4775_/D fanout250/X vssd1 vssd1 vccd1 vccd1 _4775_/Q sky130_fd_sc_hd__dfstp_1
X_1987_ _2061_/A _1987_/B vssd1 vssd1 vccd1 vccd1 _1988_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_2713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3547__A _3946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3726_ _4010_/A vssd1 vssd1 vccd1 vccd1 _3726_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout122_A _4709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3314__26_A _3365__31/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2608_ _2608_/A _4719_/Q vssd1 vssd1 vccd1 vccd1 _4719_/D sky130_fd_sc_hd__xor2_1
X_3588_ _3588_/A vssd1 vssd1 vccd1 vccd1 _3597_/A sky130_fd_sc_hd__buf_6
XFILLER_9_2140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf_A
+ _4947_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2539_ _4687_/Q _4686_/Q vssd1 vssd1 vccd1 vccd1 _2539_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3282__A _3912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_2820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_3637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4209_ _4781_/Q vssd1 vssd1 vccd1 vccd1 _4782_/D sky130_fd_sc_hd__inv_2
XFILLER_21_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_2613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4528__CLK _4533_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_2657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_3694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4741__RESET_B fanout210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3457__A _4004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2361__A _3066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_2223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_3719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_4122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4678__CLK _4717_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3904__B _3904_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_2742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_3329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1705__A _4248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_2560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout180 _3738_/A vssd1 vssd1 vccd1 vccd1 fanout180/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_3147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3920__A _3924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout191 fanout192/X vssd1 vssd1 vccd1 vccd1 fanout191/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_4115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2255__B _4533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1910_ _4323_/Q _1910_/B vssd1 vssd1 vccd1 vccd1 _4323_/D sky130_fd_sc_hd__xnor2_1
XFILLER_17_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2890_ _4899_/Q _4898_/Q _4897_/Q _2890_/D vssd1 vssd1 vccd1 vccd1 _2891_/D sky130_fd_sc_hd__and4_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_3723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1841_ _3066_/A _1841_/B _1841_/C _1841_/D vssd1 vssd1 vccd1 vccd1 _1842_/B sky130_fd_sc_hd__and4_1
XFILLER_19_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_2178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4482__RESET_B fanout208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3367__A _3895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4560_ input19/X _4560_/D fanout210/X vssd1 vssd1 vccd1 vccd1 _4561_/D sky130_fd_sc_hd__dfrtp_1
X_1772_ _4271_/Q _4270_/Q vssd1 vssd1 vccd1 vccd1 _1772_/Y sky130_fd_sc_hd__xnor2_2
X_3511_ _3519_/A vssd1 vssd1 vccd1 vccd1 _3511_/Y sky130_fd_sc_hd__inv_2
X_4491_ _5042_/A _4491_/D fanout200/X vssd1 vssd1 vccd1 vccd1 _4491_/Q sky130_fd_sc_hd__dfrtp_2
X_3765__105 _3765__105/A vssd1 vssd1 vccd1 vccd1 _3765__105/Y sky130_fd_sc_hd__inv_2
XFILLER_6_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3442_ _3924_/A _3442_/B vssd1 vssd1 vccd1 vccd1 _3442_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__2147__B1 _1975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _2315_/C _2323_/X _2173_/X vssd1 vssd1 vccd1 vccd1 _2325_/B sky130_fd_sc_hd__o21ai_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5043_/A vssd1 vssd1 vccd1 vccd1 _5043_/X sky130_fd_sc_hd__clkbuf_1
X_2255_ _4559_/D _4533_/Q _4531_/Q vssd1 vssd1 vccd1 vccd1 _2255_/Y sky130_fd_sc_hd__nor3_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_TE_B
+ _2616_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2186_ _2922_/A vssd1 vssd1 vccd1 vccd1 _2327_/A sky130_fd_sc_hd__buf_6
XFILLER_1_2980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_2911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_2933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4827_ _4981_/CLK _4827_/D _3462_/Y vssd1 vssd1 vccd1 vccd1 _4827_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__3277__A _3287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_2289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2181__A _4493_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4758_ _3424_/Y _4758_/D _3654__84/Y vssd1 vssd1 vccd1 vccd1 _4758_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4689_ _3380_/Y _4689_/D _3677_/Y vssd1 vssd1 vccd1 vccd1 _4689_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4970__CLK _3539_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_3362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_3445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf_TE_B
+ _3054_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_2661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3740__A _3748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4350__CLK input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4993__RESET_B fanout242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf _4275_/Q _1852_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_16_3133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_3609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout157/X fanout203/X vssd1 vssd1 vccd1 vccd1 _5082_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_9_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_2443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2091__A _3066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3915__A _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_4057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
+ _4802_/Q _2780_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_7_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_3137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5028__RESET_B fanout214/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_2508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_3091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3650__A _4195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2040_ _4436_/Q _4435_/Q _4434_/Q _2077_/A vssd1 vssd1 vccd1 vccd1 _2063_/B sky130_fd_sc_hd__or4_1
XFILLER_5_2390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_2221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_2182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_2265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3991_ _4456_/Q vssd1 vssd1 vccd1 vccd1 _4455_/D sky130_fd_sc_hd__inv_2
XFILLER_34_2510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2942_ _4931_/D _4905_/Q vssd1 vssd1 vccd1 vccd1 _2943_/B sky130_fd_sc_hd__xnor2_1
XFILLER_34_3277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_2407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2873_ _4867_/Q _2873_/B vssd1 vssd1 vccd1 vccd1 _4867_/D sky130_fd_sc_hd__xnor2_1
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3097__A _4992_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_3553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4612_ _4626_/CLK _4612_/D fanout234/X vssd1 vssd1 vccd1 vccd1 _4612_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1824_ _1778_/D _1822_/Y _1823_/X vssd1 vssd1 vccd1 vccd1 _1825_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__2432__C _2432_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4993__CLK _5047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1755_ _5016_/Q vssd1 vssd1 vccd1 vccd1 _5015_/D sky130_fd_sc_hd__inv_2
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4543_ _3300_/Y _4543_/D _3716_/Y vssd1 vssd1 vccd1 vccd1 _4543_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_3048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1686_ _4914_/Q vssd1 vssd1 vccd1 vccd1 _4915_/D sky130_fd_sc_hd__inv_2
X_4474_ _1952_/A1 _4474_/D _3260__20/Y vssd1 vssd1 vccd1 vccd1 _4474_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_3914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_3925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _3917_/A _3444_/B vssd1 vssd1 vccd1 vccd1 _3356_/Y sky130_fd_sc_hd__xnor2_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_w0.cclk_I_A _1935_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2662__B1_N _2659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ _4578_/Q _4577_/Q _2315_/C _2318_/A vssd1 vssd1 vccd1 vccd1 _2361_/B sky130_fd_sc_hd__a31o_1
XFILLER_3_3765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_3693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3287_ _3287_/A vssd1 vssd1 vccd1 vccd1 _3287_/Y sky130_fd_sc_hd__inv_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3560__A _4189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4373__CLK _4472_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_2981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2238_ _4524_/Q _2238_/B vssd1 vssd1 vccd1 vccd1 _4524_/D sky130_fd_sc_hd__xnor2_1
X_5026_ input24/X _5026_/D fanout225/X vssd1 vssd1 vccd1 vccd1 _5026_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2176__A _2176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_A
+ _4431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2169_ _4491_/Q _2134_/D _2162_/B vssd1 vssd1 vccd1 vccd1 _2170_/B sky130_fd_sc_hd__a21bo_1
XFILLER_17_4143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
+ _4860_/Q _2880_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_3929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3162__62_A _3169__65/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_2097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_GATE_N
+ _5063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4716__CLK _4717_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3470__A _3470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_2530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3087__A1 _3058_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4866__CLK _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input15_A comp_high_Q[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3749_/A fanout187/X vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__dlrtn_1
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
+ _4532_/Q _2274_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_17_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_3553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_2841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_3840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_2896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_3407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3645__A _4195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4396__CLK _4402_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3210_ _3848_/A _3847_/A vssd1 vssd1 vccd1 vccd1 _3210_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_27_3092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4190_ _4190_/A _4190_/B vssd1 vssd1 vccd1 vccd1 _4750_/D sky130_fd_sc_hd__xnor2_1
XFILLER_25_1808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_2222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3141_ _3930_/X _4126_/A vssd1 vssd1 vccd1 vccd1 _3141_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_3833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3380__A _4065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3072_ _4986_/Q _3068_/C _3069_/B vssd1 vssd1 vccd1 vccd1 _3073_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_3949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout120/X fanout249/X vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__dlrtn_1
X_2023_ _4406_/Q _4405_/Q vssd1 vssd1 vccd1 vccd1 _2023_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_1_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3158__58_A _3159__59/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5021__CLK input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3974_ _4421_/Q vssd1 vssd1 vccd1 vccd1 _4422_/D sky130_fd_sc_hd__inv_2
XFILLER_12_4040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_3648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_GATE_N
+ _3632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3539__B _4190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2925_ _4897_/Q _2925_/B vssd1 vssd1 vccd1 vccd1 _4897_/D sky130_fd_sc_hd__xnor2_1
XFILLER_30_2237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2856_ _4862_/Q _2856_/B vssd1 vssd1 vccd1 vccd1 _4862_/D sky130_fd_sc_hd__xnor2_1
XFILLER_34_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
+ _4575_/Q _2372_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_1807_ _4280_/Q _1779_/D _1799_/B vssd1 vssd1 vccd1 vccd1 _1808_/B sky130_fd_sc_hd__a21bo_1
XFILLER_12_2671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2787_ _4836_/Q _4835_/D vssd1 vssd1 vccd1 vccd1 _2788_/A sky130_fd_sc_hd__and2b_1
XANTENNA__3555__A _3571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4526_ _5042_/A _4526_/D fanout202/X vssd1 vssd1 vccd1 vccd1 _4526_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout202_A fanout220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1738_ _4981_/Q vssd1 vssd1 vccd1 vccd1 _4982_/D sky130_fd_sc_hd__inv_2
XANTENNA__3274__B _3438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_2144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4457_ _2294_/B1 _4457_/D _3253_/Y vssd1 vssd1 vccd1 vccd1 _4457_/Q sky130_fd_sc_hd__dfrtp_1
X_1669_ _4883_/Q vssd1 vssd1 vccd1 vccd1 _4882_/D sky130_fd_sc_hd__inv_2
XFILLER_24_2008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3408_ _3414_/A vssd1 vssd1 vccd1 vccd1 _3408_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_3619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4388_ _3214_/Y _4388_/D _3759__99/Y vssd1 vssd1 vccd1 vccd1 _4388_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_input7_A comp_high_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _3903_/A _3420_/B vssd1 vssd1 vccd1 vccd1 _3339_/Y sky130_fd_sc_hd__xnor2_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3290__A _3309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4585__RESET_B fanout231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5009_ _1765_/A _5009_/D _3563_/Y vssd1 vssd1 vccd1 vccd1 _5009_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4269__CLK _3846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3449__B _4250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_2413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3465__A _3916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_4141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3184__B _3372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_2818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_3221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3912__B _3913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_2658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_2428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_2371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[1\].w1.ro_block_I.ro_pol.tribuf.t_buf _2284_/X _2130_/Y vssd1
+ vssd1 vccd1 vccd1 _5088_/A sky130_fd_sc_hd__ebufn_8
XFILLER_18_3047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_4073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_79 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_4095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_2368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_2379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2710_ _4784_/Q _4783_/Q vssd1 vssd1 vccd1 vccd1 _2710_/Y sky130_fd_sc_hd__xnor2_4
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout128/X fanout246/X vssd1 vssd1 vccd1 vccd1 _5077_/A sky130_fd_sc_hd__dlrtn_1
X_3690_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3690_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2641_ _4754_/Q _4753_/Q vssd1 vssd1 vccd1 vccd1 _2641_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__3375__A _3375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2572_ _2922_/A vssd1 vssd1 vccd1 vccd1 _2680_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_3007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4311_ _4324_/CLK _4311_/D fanout190/X vssd1 vssd1 vccd1 vccd1 _4311_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_2306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4242_ _4832_/Q vssd1 vssd1 vccd1 vccd1 _4831_/D sky130_fd_sc_hd__inv_2
XFILLER_25_2339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4173_ _4728_/Q vssd1 vssd1 vccd1 vccd1 _4729_/D sky130_fd_sc_hd__inv_2
XFILLER_3_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_2041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3124_ _5018_/Q _5017_/Q vssd1 vssd1 vccd1 vccd1 _3124_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_4_3893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_2085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3055_ _5024_/D _4998_/Q _4996_/Q _4995_/Q vssd1 vssd1 vccd1 vccd1 _3056_/C sky130_fd_sc_hd__and4_1
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_2995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2006_ _2006_/A vssd1 vssd1 vccd1 vccd1 _2006_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4411__CLK _3932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[0\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf _2107_/A _1957_/Y vssd1
+ vssd1 vccd1 vccd1 _5091_/A sky130_fd_sc_hd__ebufn_8
XFILLER_23_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout152_A _4920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_3445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_2711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3957_ _4406_/Q vssd1 vssd1 vccd1 vccd1 _4405_/D sky130_fd_sc_hd__inv_2
XFILLER_10_3309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_RESET_B fanout193/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2908_ _4895_/Q _2908_/B vssd1 vssd1 vccd1 vccd1 _2909_/B sky130_fd_sc_hd__nor2_1
XFILLER_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4561__CLK input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3888_ _3888_/A _3901_/B vssd1 vssd1 vccd1 vccd1 _3891_/B sky130_fd_sc_hd__or2_1
XFILLER_30_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2839_ _2829_/C _2838_/X _2687_/X vssd1 vssd1 vccd1 vccd1 _2840_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__3285__A _3287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_2490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__0637_ _3733_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0637_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4509_ _3280_/Y _4509_/D _3726_/Y vssd1 vssd1 vccd1 vccd1 _4509_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_3782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4766__RESET_B fanout255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_2840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_2079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2501__A3 _2480_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_3523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4904__CLK _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2973__B1 _3877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_2287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_2615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3923__A _3923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_3134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4436__RESET_B fanout198/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2258__B _4533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4434__CLK _5033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_2477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_2499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4860_ _4865_/CLK _4860_/D fanout226/X vssd1 vssd1 vccd1 vccd1 _4860_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4584__CLK _4623_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3811_ _4309_/Q vssd1 vssd1 vccd1 vccd1 _4308_/D sky130_fd_sc_hd__inv_2
X_4791_ _4981_/CLK _4791_/D _3441_/Y vssd1 vssd1 vccd1 vccd1 _4791_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3742_ _3748_/A vssd1 vssd1 vccd1 vccd1 _3742_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_3099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3673_ _4135_/A vssd1 vssd1 vccd1 vccd1 _3673_/Y sky130_fd_sc_hd__inv_2
X_2624_ _4747_/Q _4746_/D vssd1 vssd1 vccd1 vccd1 _2625_/A sky130_fd_sc_hd__and2b_1
Xoutput102 _5099_/X vssd1 vssd1 vccd1 vccd1 sin_out[7] sky130_fd_sc_hd__buf_2
XFILLER_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2555_ _4715_/Q _4714_/Q _4713_/Q _2592_/A vssd1 vssd1 vccd1 vccd1 _2579_/B sky130_fd_sc_hd__or4_2
XFILLER_25_2103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_3861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2486_ _4673_/Q _4672_/Q _4671_/Q _2497_/B vssd1 vssd1 vccd1 vccd1 _2491_/B sky130_fd_sc_hd__or4_2
XFILLER_5_2208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3552__B _5029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4225_ _4813_/Q vssd1 vssd1 vccd1 vccd1 _4814_/D sky130_fd_sc_hd__inv_2
XFILLER_25_2158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4156_ _4697_/Q vssd1 vssd1 vccd1 vccd1 _4696_/D sky130_fd_sc_hd__inv_2
XANTENNA__3211__16_A _3264__22/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3107_ _4995_/Q _3107_/B vssd1 vssd1 vccd1 vccd1 _4995_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_3554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4087_ _4597_/Q vssd1 vssd1 vccd1 vccd1 _4598_/D sky130_fd_sc_hd__inv_2
XFILLER_0_2842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4927__CLK input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3038_ _5020_/D _4962_/Q vssd1 vssd1 vccd1 vccd1 _3039_/B sky130_fd_sc_hd__xnor2_1
XFILLER_24_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_4090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_3865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4989_ _4997_/CLK _4989_/D fanout235/X vssd1 vssd1 vccd1 vccd1 _4989_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_3106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_3275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
+ _4394_/Q _2026_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__4307__CLK _3888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4947__RESET_B fanout208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_3636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_4111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3743__A _3748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4457__CLK _2294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_2742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_2617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_2939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2822__A _4927_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_3949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 comp_high_Q[6] vssd1 vssd1 vccd1 vccd1 _4926_/D sky130_fd_sc_hd__clkbuf_4
Xinput26 phi1b_dig_Q[1] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_2062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4617__RESET_B fanout234/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_3157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2340_ _4584_/Q _2304_/D _2333_/B vssd1 vssd1 vccd1 vccd1 _2341_/B sky130_fd_sc_hd__a21bo_1
XFILLER_26_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3372__B _3372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_2309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2271_ _4547_/Q _4546_/Q vssd1 vssd1 vccd1 vccd1 _2271_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_26_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4270__RESET_B _4359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4010_ _4010_/A vssd1 vssd1 vccd1 vccd1 _4469_/D sky130_fd_sc_hd__inv_2
XFILLER_4_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_2077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2229__A2 _4523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4912_ _5007_/CLK _4912_/D _3507_/Y vssd1 vssd1 vccd1 vccd1 _4912_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4843_ _4843_/CLK _4843_/D fanout226/X vssd1 vssd1 vccd1 vccd1 _4843_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4774_ _4812_/CLK _4774_/D fanout253/X vssd1 vssd1 vccd1 vccd1 _4774_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1986_ _4395_/Q _4394_/Q _1963_/D _1983_/B vssd1 vssd1 vccd1 vccd1 _1987_/B sky130_fd_sc_hd__a31o_1
XFILLER_11_2725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3547__B _3945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3725_ _4010_/A vssd1 vssd1 vccd1 vccd1 _3725_/Y sky130_fd_sc_hd__inv_2
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_TE_B
+ _3121_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3656_ _3656_/A vssd1 vssd1 vccd1 vccd1 _3656_/X sky130_fd_sc_hd__buf_1
XANTENNA_fanout115_A _4812_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2607_ _4718_/Q _2607_/B vssd1 vssd1 vccd1 vccd1 _4718_/D sky130_fd_sc_hd__xor2_1
XFILLER_27_2209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3587_ _3587_/A vssd1 vssd1 vccd1 vccd1 _3587_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3563__A _3571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3781__122 _3781__122/A vssd1 vssd1 vccd1 vccd1 _3781__122/Y sky130_fd_sc_hd__inv_2
XFILLER_27_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2538_ _4685_/Q _4684_/Q vssd1 vssd1 vccd1 vccd1 _2538_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__3282__B _3446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2179__A _4492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2469_ _2631_/A _3908_/A _2456_/Y _2461_/Y _2468_/A vssd1 vssd1 vccd1 vccd1 _2469_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_22_3555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4208_ _4782_/Q vssd1 vssd1 vccd1 vccd1 _4781_/D sky130_fd_sc_hd__inv_2
XFILLER_29_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4139_ _4662_/Q vssd1 vssd1 vccd1 vccd1 _4663_/D sky130_fd_sc_hd__inv_2
XFILLER_0_3373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_1_1_0_w0.cclk_I_A clkbuf_0_w0.cclk_I/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1979__A1 _4392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3738__A _3738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3457__B _3491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_4134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3473__A _3905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2156__A1 _4488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1705__B _4248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_3137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout170 _3861_/Y vssd1 vssd1 vccd1 vccd1 _3914_/A sky130_fd_sc_hd__buf_6
Xfanout181 _5057_/A vssd1 vssd1 vccd1 vccd1 _3738_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout192 fanout193/X vssd1 vssd1 vccd1 vccd1 fanout192/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3920__B _3923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_2353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3599__1 _3470_/A vssd1 vssd1 vccd1 vccd1 _3599__1/Y sky130_fd_sc_hd__inv_2
XFILLER_21_2386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout144/X fanout215/X vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_34_3437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__1632_ clkbuf_0__1632_/X vssd1 vssd1 vccd1 vccd1 _3193__75/A sky130_fd_sc_hd__clkbuf_16
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_2293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3648__A _4195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1840_ _4347_/D _4274_/Q vssd1 vssd1 vccd1 vccd1 _1841_/D sky130_fd_sc_hd__xnor2_1
XFILLER_19_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4869__RESET_B fanout226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3367__B _3372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_2482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1771_ _4269_/Q _4268_/Q vssd1 vssd1 vccd1 vccd1 _1771_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__4622__CLK _4626_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3510_ _4065_/A _3543_/B vssd1 vssd1 vccd1 vccd1 _3510_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_10_3481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_3219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4490_ _5034_/A _4490_/D fanout202/X vssd1 vssd1 vccd1 vccd1 _4490_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3441_ _3445_/A vssd1 vssd1 vccd1 vccd1 _3441_/Y sky130_fd_sc_hd__inv_2
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_GATE_N _4363_/CLK
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3383__A _3393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4772__CLK _4803_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _4368_/Q _3372_/B vssd1 vssd1 vccd1 vccd1 _3372_/Y sky130_fd_sc_hd__xnor2_4
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _4579_/Q _2323_/B vssd1 vssd1 vccd1 vccd1 _2323_/X sky130_fd_sc_hd__and2b_1
XFILLER_6_2336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5042_/A vssd1 vssd1 vccd1 vccd1 _5042_/X sky130_fd_sc_hd__clkbuf_1
X_2254_ _4559_/D _4533_/Q _4531_/Q vssd1 vssd1 vccd1 vccd1 _2254_/X sky130_fd_sc_hd__and3_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2185_ _4494_/Q _2185_/B vssd1 vssd1 vccd1 vccd1 _4494_/D sky130_fd_sc_hd__xnor2_1
Xwrapper_cell_loop\[6\].w1.ro_block_I.ro_pol_eve.tribuf.t_buf _3133_/A _2984_/Y vssd1
+ vssd1 vccd1 vccd1 _5089_/A sky130_fd_sc_hd__ebufn_8
XFILLER_4_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3558__A _4249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1830__B1 _1823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2462__A _3941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_2989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4826_ _3461_/Y _4826_/D _3635_/Y vssd1 vssd1 vccd1 vccd1 _4826_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout232_A fanout234/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_2680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4757_ _2631_/A _4757_/D _3423__40/Y vssd1 vssd1 vccd1 vccd1 _4757_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1969_ _4394_/Q _4393_/Q _4392_/Q _1982_/B vssd1 vssd1 vccd1 vccd1 _1974_/B sky130_fd_sc_hd__or4_2
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4688_ _1765_/A _4688_/D _3379_/Y vssd1 vssd1 vccd1 vccd1 _4688_/Q sky130_fd_sc_hd__dfrtp_1
X_3639_ _3642_/A vssd1 vssd1 vccd1 vccd1 _3639_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3293__A _3309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_3617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_4020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_4031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_3374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_3145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_2422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4645__CLK _2470_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3468__A _5061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_2455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4962__RESET_B fanout210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_2499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4795__CLK _4852_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_2656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3931__A _3931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout158/X fanout205/X vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_21_2161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_2194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_2208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3990_ _4453_/Q vssd1 vssd1 vccd1 vccd1 _4454_/D sky130_fd_sc_hd__inv_2
XFILLER_1_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_2500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3771__110 _3776__115/A vssd1 vssd1 vccd1 vccd1 _3771__110/Y sky130_fd_sc_hd__inv_2
XFILLER_14_3819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2941_ _4902_/Q _2941_/B vssd1 vssd1 vccd1 vccd1 _4902_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__2065__B1 _2003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3378__A _4127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1812__B1 _3109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2872_ _2916_/A _2872_/B vssd1 vssd1 vccd1 vccd1 _2873_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_2588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4611_ _4623_/CLK _4611_/D fanout231/X vssd1 vssd1 vccd1 vccd1 _4611_/Q sky130_fd_sc_hd__dfrtp_2
X_1823_ _2922_/A vssd1 vssd1 vccd1 vccd1 _1823_/X sky130_fd_sc_hd__buf_4
XFILLER_12_3598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4542_ _3932_/A _4542_/D _3299_/Y vssd1 vssd1 vccd1 vccd1 _4542_/Q sky130_fd_sc_hd__dfrtp_1
X_1754_ _5013_/Q vssd1 vssd1 vccd1 vccd1 _5014_/D sky130_fd_sc_hd__inv_2
X_4473_ _4473_/CLK _4473_/D fanout204/X vssd1 vssd1 vccd1 vccd1 _4473_/Q sky130_fd_sc_hd__dfrtp_1
X_1685_ _4915_/Q vssd1 vssd1 vccd1 vccd1 _4914_/D sky130_fd_sc_hd__inv_2
X_3424_ _3896_/A _3904_/A vssd1 vssd1 vccd1 vccd1 _3424_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_25_3937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_2359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ _3361_/A vssd1 vssd1 vccd1 vccd1 _3355_/Y sky130_fd_sc_hd__inv_2
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_2144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_3733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4518__CLK _4532_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2306_ _4576_/Q vssd1 vssd1 vccd1 vccd1 _2318_/A sky130_fd_sc_hd__inv_2
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5063_/A fanout251/X vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__dlrtn_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _3895_/A _3372_/B vssd1 vssd1 vccd1 vccd1 _3286_/Y sky130_fd_sc_hd__xnor2_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3560__B _4190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5025_ input24/X _5025_/D fanout225/X vssd1 vssd1 vccd1 vccd1 _5026_/D sky130_fd_sc_hd__dfrtp_1
XANTENNA__2457__A _2468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2237_ _2208_/D _2236_/X _2173_/X vssd1 vssd1 vccd1 vccd1 _2238_/B sky130_fd_sc_hd__o21ai_1
XFILLER_6_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2168_ _4489_/Q _2168_/B vssd1 vssd1 vccd1 vccd1 _4489_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__4668__CLK _4718_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2099_ _4452_/Q _4451_/Q vssd1 vssd1 vccd1 vccd1 _2099_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_35_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3288__A _3891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_3329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_2797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4809_ _4809_/CLK _4809_/D fanout255/X vssd1 vssd1 vccd1 vccd1 _4809_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3474__45_A _3528__52/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_3550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_2702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_2871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3751__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_3221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2295__B1 _3932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_4119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_2853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_4004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_2613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_2657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output76_A _5073_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3661__A _3669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3140_ _4064_/A _4188_/B _3139_/Y vssd1 vssd1 vccd1 vccd1 _3140_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_3917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_2256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3380__B _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4810__CLK _4812_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_2278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3071_ _3071_/A _3071_/B vssd1 vssd1 vccd1 vccd1 _4984_/D sky130_fd_sc_hd__xnor2_1
XFILLER_3_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2022_ _2608_/A _4404_/Q vssd1 vssd1 vccd1 vccd1 _4404_/D sky130_fd_sc_hd__xor2_1
XFILLER_23_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
+ _4991_/Q _3115_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_1_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4960__CLK _4962_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3973_ _4422_/Q vssd1 vssd1 vccd1 vccd1 _4421_/D sky130_fd_sc_hd__inv_2
XFILLER_34_3075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2924_ _3030_/A _2924_/B vssd1 vssd1 vccd1 vccd1 _2925_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_4085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_2959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2855_ _2916_/A _2855_/B vssd1 vssd1 vccd1 vccd1 _2856_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_3985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3836__A _3883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1806_ _4278_/Q _1806_/B vssd1 vssd1 vccd1 vccd1 _4278_/D sky130_fd_sc_hd__xnor2_1
XFILLER_12_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2786_ _4832_/Q _4831_/Q vssd1 vssd1 vccd1 vccd1 _2786_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_15_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4525_ _4533_/CLK _4525_/D fanout209/X vssd1 vssd1 vccd1 vccd1 _4525_/Q sky130_fd_sc_hd__dfrtp_2
X_1737_ _4982_/Q vssd1 vssd1 vccd1 vccd1 _4981_/D sky130_fd_sc_hd__inv_2
XFILLER_28_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_2112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_2123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4340__CLK _2294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout119/X fanout248/X vssd1 vssd1 vccd1 vccd1 _5078_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_29_3881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4456_ _3252_/Y _4456_/D _3740_/Y vssd1 vssd1 vccd1 vccd1 _4456_/Q sky130_fd_sc_hd__dfrtp_2
X_1668_ _4880_/Q vssd1 vssd1 vccd1 vccd1 _4881_/D sky130_fd_sc_hd__inv_2
XFILLER_5_3806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_2217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3407_ _3935_/A _3440_/B vssd1 vssd1 vccd1 vccd1 _3407_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_A
+ _4894_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4387_ _3845_/Y _4387_/D _3213__17/Y vssd1 vssd1 vccd1 vccd1 _4387_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_3609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3571__A _3571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3338_ _3340_/A vssd1 vssd1 vccd1 vccd1 _3338_/Y sky130_fd_sc_hd__inv_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2187__A _4555_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3269_ _4469_/Q vssd1 vssd1 vccd1 vccd1 _3287_/A sky130_fd_sc_hd__buf_6
XFILLER_3_2851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_2862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5008_ _3562_/Y _5008_/D _3582_/Y vssd1 vssd1 vccd1 vccd1 _5008_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4554__RESET_B fanout207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_3749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3746__A _3748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3465__B _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_4039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4833__CLK input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3481__A _3498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2504__A1 _4674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_3277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_3062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4983__CLK _4997_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_4041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2825__A _4859_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_3925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_2336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4462__D _4462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_2661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_TE_B
+ _2710_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_3259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_2536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
+ _4706_/Q _2615_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_13_3693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3656__A _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2640_ _4064_/A _2640_/B vssd1 vssd1 vccd1 vccd1 _5068_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__4363__CLK _4363_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2571_ _4707_/Q _2571_/B vssd1 vssd1 vccd1 vccd1 _4707_/D sky130_fd_sc_hd__xnor2_1
X_4310_ _4324_/CLK _4310_/D fanout194/X vssd1 vssd1 vccd1 vccd1 _4310_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_3249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4241_ _4829_/Q vssd1 vssd1 vccd1 vccd1 _4830_/D sky130_fd_sc_hd__inv_2
XFILLER_29_2498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1904__A _4351_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3391__A _3393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4172_ _4729_/Q vssd1 vssd1 vccd1 vccd1 _4728_/D sky130_fd_sc_hd__inv_2
XFILLER_7_2283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3123_ _5016_/Q _5015_/Q vssd1 vssd1 vccd1 vccd1 _3123_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_3_2125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_2097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3054_ _4982_/Q _4981_/Q vssd1 vssd1 vccd1 vccd1 _3054_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_3_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2005_ _4398_/Q _2005_/B vssd1 vssd1 vccd1 vccd1 _4398_/D sky130_fd_sc_hd__xnor2_1
XFILLER_35_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3956_ _4387_/Q vssd1 vssd1 vccd1 vccd1 _4388_/D sky130_fd_sc_hd__clkinv_2
XANTENNA__4706__CLK _4709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout145_A _3696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2907_ _4892_/Q _2907_/B vssd1 vssd1 vccd1 vccd1 _4892_/D sky130_fd_sc_hd__xnor2_1
XFILLER_34_2193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3887_ _4365_/Q vssd1 vssd1 vccd1 vccd1 _3889_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__3566__A _4001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2838_ _4858_/Q _2838_/B vssd1 vssd1 vccd1 vccd1 _2838_/X sky130_fd_sc_hd__and2b_1
XANTENNA__4856__CLK _4905_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2769_ _4809_/Q _2769_/B vssd1 vssd1 vccd1 vccd1 _4809_/D sky130_fd_sc_hd__xnor2_1
X_4508_ _3931_/A _4508_/D _3279_/Y vssd1 vssd1 vccd1 vccd1 _4508_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_3520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4439_ _5033_/A _4439_/D fanout195/X vssd1 vssd1 vccd1 vccd1 _4439_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_25_3575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
+ _4764_/Q _2712_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__2629__B _3658_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_3313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2645__A _4834_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2422__B1 _2344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_2391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2973__A1 _4064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2380__A _4652_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_2889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3923__B _3925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5011__CLK _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_2412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_2340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_3179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_2445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_2237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4729__CLK _3405_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_3711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5056_/A fanout190/X vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__dlrtn_1
X_3810_ _4306_/Q vssd1 vssd1 vccd1 vccd1 _4307_/D sky130_fd_sc_hd__inv_2
XFILLER_32_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4790_ _3440_/Y _4790_/D _3646_/Y vssd1 vssd1 vccd1 vccd1 _4790_/Q sky130_fd_sc_hd__dfrtp_4
X_3604__78 _3654__84/A vssd1 vssd1 vccd1 vccd1 _3604__78/Y sky130_fd_sc_hd__inv_2
X_3741_ _3748_/A vssd1 vssd1 vccd1 vccd1 _3741_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_2491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3386__A _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_2344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_2366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3672_ _4135_/A vssd1 vssd1 vccd1 vccd1 _3672_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2623_ _2623_/A vssd1 vssd1 vccd1 vccd1 _2623_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2554_ _4745_/D _4719_/Q _4717_/Q _4716_/Q vssd1 vssd1 vccd1 vccd1 _2592_/A sky130_fd_sc_hd__or4_1
XFILLER_6_3945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_3873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2485_ _4676_/Q _4675_/Q _4674_/Q _2507_/B vssd1 vssd1 vccd1 vccd1 _2497_/B sky130_fd_sc_hd__or4_1
XANTENNA_net199_2_A _3600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4010__A _4010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4224_ _4814_/Q vssd1 vssd1 vccd1 vccd1 _4813_/D sky130_fd_sc_hd__inv_2
XFILLER_2_3809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_3989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4155_ _4694_/Q vssd1 vssd1 vccd1 vccd1 _4695_/D sky130_fd_sc_hd__inv_2
XFILLER_25_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3106_ _3104_/X _3105_/Y _1791_/X vssd1 vssd1 vccd1 vccd1 _3107_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_2810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4086_ _4598_/Q vssd1 vssd1 vccd1 vccd1 _4597_/D sky130_fd_sc_hd__inv_2
XFILLER_23_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3037_ _4959_/Q _3037_/B vssd1 vssd1 vccd1 vccd1 _4959_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_4080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_3877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4988_ _4997_/CLK _4988_/D fanout235/X vssd1 vssd1 vccd1 vccd1 _4988_/Q sky130_fd_sc_hd__dfrtp_4
X_3939_ _4123_/A vssd1 vssd1 vccd1 vccd1 _3939_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__3296__A _3947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_4123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_3_0_clk_master clkbuf_3_3_0_clk_master/A vssd1 vssd1 vccd1 vccd1 _5048_/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_5_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_2958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4987__RESET_B fanout235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_3247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_2754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_2513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4740__D _4740_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput16 comp_high_Q[7] vssd1 vssd1 vccd1 vccd1 _5019_/D sky130_fd_sc_hd__buf_8
XFILLER_10_3641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput27 phi1b_dig_Q[2] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_2
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3934__A _3934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4401__CLK _4402_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2270_ _4545_/Q _4544_/Q vssd1 vssd1 vccd1 vccd1 _2270_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_6_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_2045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2285__A _3684_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4911_ _3506_/Y _4911_/D _3613_/Y vssd1 vssd1 vccd1 vccd1 _4911_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_2417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4842_ _5030_/CLK _4842_/D fanout224/X vssd1 vssd1 vccd1 vccd1 _4842_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_3585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4773_ _4812_/CLK _4773_/D fanout253/X vssd1 vssd1 vccd1 vccd1 _4773_/Q sky130_fd_sc_hd__dfrtp_1
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
+ _4525_/Q _2266_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1985_ _4392_/Q _1985_/B vssd1 vssd1 vccd1 vccd1 _4392_/D sky130_fd_sc_hd__xnor2_1
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout136/X fanout238/X vssd1 vssd1 vccd1 vccd1 _5084_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_15_2862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3724_ _4010_/A vssd1 vssd1 vccd1 vccd1 _3724_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4005__A _4005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3844__A _3848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2606_ _3112_/A _2606_/B _2606_/C _2606_/D vssd1 vssd1 vccd1 vccd1 _2607_/B sky130_fd_sc_hd__and4_1
X_3586_ _3587_/A vssd1 vssd1 vccd1 vccd1 _3586_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout108_A _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2537_ _2608_/A _4683_/Q vssd1 vssd1 vccd1 vccd1 _4683_/D sky130_fd_sc_hd__xor2_1
XFILLER_22_3501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_3681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2468_ _2468_/A _3929_/A vssd1 vssd1 vccd1 vccd1 _2801_/C sky130_fd_sc_hd__nand2_1
XFILLER_22_2800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4207_ _4779_/Q vssd1 vssd1 vccd1 vccd1 _4780_/D sky130_fd_sc_hd__inv_2
XFILLER_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2399_ _2412_/A _2399_/B vssd1 vssd1 vccd1 vccd1 _2400_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4138_ _4663_/Q vssd1 vssd1 vccd1 vccd1 _4662_/D sky130_fd_sc_hd__inv_2
XFILLER_28_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4069_ _4566_/Q _4070_/B vssd1 vssd1 vccd1 vccd1 _4565_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_2651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_3917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1979__A2 _1973_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_2951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4424__CLK _3234_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3754__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2156__A2 _4487_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3473__B _3913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
+ _4583_/Q _2364_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__4750__RESET_B fanout228/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_3191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_2799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout160 _4000_/Y vssd1 vssd1 vccd1 vccd1 _2809_/A1 sky130_fd_sc_hd__buf_12
XFILLER_1_3127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout171 _3855_/Y vssd1 vssd1 vccd1 vccd1 _2294_/B1 sky130_fd_sc_hd__buf_6
XFILLER_5_2573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout182 _4354_/Q vssd1 vssd1 vccd1 vccd1 _5057_/A sky130_fd_sc_hd__buf_4
Xfanout193 fanout196/X vssd1 vssd1 vccd1 vccd1 fanout193/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_2426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_2365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_4117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_2398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3929__A _3929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2833__A _2922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1770_ _4267_/Q _4266_/Q vssd1 vssd1 vccd1 vccd1 _1770_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3189__72 _3189__72/A vssd1 vssd1 vccd1 vccd1 _3189__72/Y sky130_fd_sc_hd__inv_2
XFILLER_10_3493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3664__A _3669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_2770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3440_ _3934_/A _3440_/B vssd1 vssd1 vccd1 vccd1 _3440_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_2508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4917__CLK _3512_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4838__RESET_B fanout231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_2210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2322_ _4580_/Q _2322_/B vssd1 vssd1 vccd1 vccd1 _2323_/B sky130_fd_sc_hd__nor2_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_TE_B
+ _2784_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_2243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5041_ _5041_/A vssd1 vssd1 vccd1 vccd1 _5041_/X sky130_fd_sc_hd__clkbuf_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2253_ _4529_/Q _2253_/B vssd1 vssd1 vccd1 vccd1 _4529_/D sky130_fd_sc_hd__xnor2_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1912__A _3066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_2050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2184_ _2182_/X _2183_/Y _2173_/X vssd1 vssd1 vccd1 vccd1 _2185_/B sky130_fd_sc_hd__o21ai_2
XFILLER_4_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3684_/A fanout216/X vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_20_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_3647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_2913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_3961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3558__B _4250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2462__B _3929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4825_ _4920_/CLK _4825_/D _3460_/Y vssd1 vssd1 vccd1 vccd1 _4825_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4447__CLK _3932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[3\].w1.ro_block_I.ro_pol_eve.tribuf.t_buf _2627_/A _2476_/Y vssd1
+ vssd1 vccd1 vccd1 _5089_/A sky130_fd_sc_hd__ebufn_8
XANTENNA__3032__B1 _1791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4756_ _3422_/Y _4756_/D _3655__85/Y vssd1 vssd1 vccd1 vccd1 _4756_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout225_A fanout230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1968_ _4397_/Q _4396_/Q _4395_/Q _1992_/B vssd1 vssd1 vccd1 vccd1 _1982_/B sky130_fd_sc_hd__or4_1
XFILLER_11_3279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4687_ _3378_/Y _4687_/D _3678_/Y vssd1 vssd1 vccd1 vccd1 _4687_/Q sky130_fd_sc_hd__dfrtp_2
X_1899_ _1898_/Y _1856_/C _4321_/Q vssd1 vssd1 vccd1 vccd1 _1900_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4597__CLK _3939_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3638_ _3642_/A vssd1 vssd1 vccd1 vccd1 _3638_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_3743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_4010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3569_ _3571_/A vssd1 vssd1 vccd1 vccd1 _3569_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_4115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_3414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_3386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_2713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_3469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2637__B _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_2685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4555__D _4555_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_2412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_2781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_3529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3484__A _3498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3931__B _4131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_2668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4465__D input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_2289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_3934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_3978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2940_ _2938_/X _2939_/Y _2858_/X vssd1 vssd1 vccd1 vccd1 _2941_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__2065__A1 _2036_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3198__6 _3199__7/A vssd1 vssd1 vccd1 vccd1 _4366_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__3378__B _4129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2871_ _4927_/D _4869_/Q vssd1 vssd1 vccd1 vccd1 _2872_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1822_ _4285_/Q _4284_/Q _1826_/A vssd1 vssd1 vccd1 vccd1 _1822_/Y sky130_fd_sc_hd__nor3_1
X_4610_ _3341_/Y _4610_/D _3695_/Y vssd1 vssd1 vccd1 vccd1 _4610_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_3577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4541_ _3298_/Y _4541_/D _3717_/Y vssd1 vssd1 vccd1 vccd1 _4541_/Q sky130_fd_sc_hd__dfrtp_2
X_1753_ _5014_/Q vssd1 vssd1 vccd1 vccd1 _5013_/D sky130_fd_sc_hd__inv_2
XFILLER_11_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3394__A _3903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4472_ _4472_/CLK _4472_/D fanout207/X vssd1 vssd1 vccd1 vccd1 _4472_/Q sky130_fd_sc_hd__dfrtp_1
X_1684_ _4912_/Q vssd1 vssd1 vccd1 vccd1 _4913_/D sky130_fd_sc_hd__inv_2
XANTENNA__4672__RESET_B fanout239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3354_ _3925_/A _3442_/B vssd1 vssd1 vccd1 vccd1 _3354_/Y sky130_fd_sc_hd__xnor2_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _4581_/Q _4580_/Q _4579_/Q _2305_/D vssd1 vssd1 vccd1 vccd1 _2315_/C sky130_fd_sc_hd__and4_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3285_ _3287_/A vssd1 vssd1 vccd1 vccd1 _3285_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_2167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5024_ input24/X _5024_/D fanout225/X vssd1 vssd1 vccd1 vccd1 _5025_/D sky130_fd_sc_hd__dfrtp_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ _4525_/Q _2236_/B vssd1 vssd1 vccd1 vccd1 _2236_/X sky130_fd_sc_hd__and2b_1
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_GATE_N _4359_/CLK
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_4101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2167_ _2178_/A _2167_/B vssd1 vssd1 vccd1 vccd1 _2168_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout175_A _1765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2098_ _4450_/Q _4449_/Q vssd1 vssd1 vccd1 vccd1 _2098_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_13_4009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3569__A _3571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3288__B _3889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_2033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4808_ _4809_/CLK _4808_/D fanout254/X vssd1 vssd1 vccd1 vccd1 _4808_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_1917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4739_ _3415_/Y _4739_/D _3658_/Y vssd1 vssd1 vccd1 vccd1 _4739_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5055_/A fanout244/X vssd1 vssd1 vccd1 vccd1 _5079_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__1817__A _1839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_2883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_2988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_2769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_3233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4612__CLK _4626_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_4109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3479__A _3905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_2810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_GATE_N
+ fanout128/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4762__CLK _4803_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_4016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_2669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3070_ _3068_/X _3069_/Y _2143_/A vssd1 vssd1 vccd1 vccd1 _3071_/B sky130_fd_sc_hd__o21a_1
XFILLER_7_1786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4292__CLK _4063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2021_ _4403_/Q _2021_/B vssd1 vssd1 vccd1 vccd1 _4403_/D sky130_fd_sc_hd__xor2_1
XFILLER_1_2042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3389__A _3393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2293__A _3899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_3775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3972_ _4419_/Q vssd1 vssd1 vccd1 vccd1 _4420_/D sky130_fd_sc_hd__clkinv_2
XFILLER_18_3797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2923_ _4899_/Q _4898_/Q _2890_/D _2919_/B vssd1 vssd1 vccd1 vccd1 _2924_/B sky130_fd_sc_hd__a31o_1
XFILLER_12_4053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_3931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_2386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2854_ _4863_/Q _2818_/D _2847_/B vssd1 vssd1 vccd1 vccd1 _2855_/B sky130_fd_sc_hd__a21bo_1
XFILLER_34_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1805_ _3114_/A _1805_/B vssd1 vssd1 vccd1 vccd1 _1806_/B sky130_fd_sc_hd__nand2_1
XFILLER_15_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2785_ _4830_/Q _4829_/Q vssd1 vssd1 vccd1 vccd1 _2785_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_30_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4524_ _5034_/A _4524_/D fanout202/X vssd1 vssd1 vccd1 vccd1 _4524_/Q sky130_fd_sc_hd__dfrtp_4
X_1736_ _4979_/Q vssd1 vssd1 vccd1 vccd1 _4980_/D sky130_fd_sc_hd__inv_2
XFILLER_9_3921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1667_ _4881_/Q vssd1 vssd1 vccd1 vccd1 _4880_/D sky130_fd_sc_hd__inv_2
X_4455_ _3899_/A _4455_/D _3251_/Y vssd1 vssd1 vccd1 vccd1 _4455_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3852__A _3888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3406_ _3414_/A vssd1 vssd1 vccd1 vccd1 _3406_/Y sky130_fd_sc_hd__inv_2
X_4386_ _3212_/Y _4386_/D _3760__100/Y vssd1 vssd1 vccd1 vccd1 _4386_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4635__CLK _4920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3337_ _3912_/A _3446_/B vssd1 vssd1 vccd1 vccd1 _3337_/Y sky130_fd_sc_hd__xnor2_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2468__A _2468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3268_ _3885_/A _3886_/A vssd1 vssd1 vccd1 vccd1 _3268_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__2187__B _4497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2219_ _4520_/Q _2219_/B vssd1 vssd1 vccd1 vccd1 _2219_/Y sky130_fd_sc_hd__nor2_1
X_5007_ _5007_/CLK _5007_/D _3561_/Y vssd1 vssd1 vccd1 vccd1 _5007_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_6_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4785__CLK _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4833__D _4833_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3299__A _3309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_2849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_2117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_2161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3156__56 _3159__59/A vssd1 vssd1 vccd1 vccd1 _3156__56/Y sky130_fd_sc_hd__inv_2
XFILLER_8_2741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_3245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2504__A2 _2480_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input20_A phi1b_dig_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_4031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_3904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_4086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_3915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_2651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_3249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_2673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4508__CLK _3931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3187__71_A _3189__72/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2570_ _2561_/C _2569_/X _2518_/X vssd1 vssd1 vccd1 vccd1 _2571_/B sky130_fd_sc_hd__o21ai_1
XFILLER_9_3217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3672__A _4135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4240_ _4830_/Q vssd1 vssd1 vccd1 vccd1 _4829_/D sky130_fd_sc_hd__inv_2
XFILLER_29_2477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4171_ _4726_/Q vssd1 vssd1 vccd1 vccd1 _4727_/D sky130_fd_sc_hd__clkinv_2
XFILLER_25_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_3610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3122_ _5014_/Q _5013_/Q vssd1 vssd1 vccd1 vccd1 _3122_/Y sky130_fd_sc_hd__xnor2_2
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout180/X fanout184/X vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_4_3873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_2065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3053_ _4980_/Q _4979_/Q vssd1 vssd1 vccd1 vccd1 _3053_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_23_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2004_ _1962_/D _2002_/Y _2003_/X vssd1 vssd1 vccd1 vccd1 _2005_/B sky130_fd_sc_hd__o21ai_1
XFILLER_23_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_2986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_4115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3955_ _4388_/Q vssd1 vssd1 vccd1 vccd1 _4387_/D sky130_fd_sc_hd__inv_2
XANTENNA__3847__A _3847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_2893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2906_ _2916_/A _2906_/B vssd1 vssd1 vccd1 vccd1 _2907_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3886_ _3886_/A _3886_/B vssd1 vssd1 vccd1 vccd1 _4364_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__3566__B _4005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_2036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2837_ _4859_/Q _2837_/B vssd1 vssd1 vccd1 vccd1 _2838_/B sky130_fd_sc_hd__nor2_1
XFILLER_34_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3202__10_A _3201__9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2768_ _2766_/X _2767_/Y _2687_/X vssd1 vssd1 vccd1 vccd1 _2769_/B sky130_fd_sc_hd__o21ai_1
XFILLER_12_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4507_ _3278_/Y _4507_/D _3727_/Y vssd1 vssd1 vccd1 vccd1 _4507_/Q sky130_fd_sc_hd__dfrtp_1
X_1719_ _4964_/Q vssd1 vssd1 vccd1 vccd1 _4963_/D sky130_fd_sc_hd__inv_2
X_2699_ _4773_/Q _2699_/B vssd1 vssd1 vccd1 vccd1 _4773_/D sky130_fd_sc_hd__xnor2_1
XFILLER_9_3751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3582__A _3587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4438_ _5041_/A _4438_/D fanout198/X vssd1 vssd1 vccd1 vccd1 _4438_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_28_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf _4310_/Q _1923_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_25_2831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_4051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_A
+ _4676_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4369_ _3598_/A _4369_/D fanout222/X vssd1 vssd1 vccd1 vccd1 _4369_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_2947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_4037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_3303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_3093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3757__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4704__RESET_B fanout237/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2661__A _2661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_2879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4800__CLK _4811_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3492__A _3498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4950__CLK _4962_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_3064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_A
+ _4708_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_2457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__1648_ clkbuf_0__1648_/X vssd1 vssd1 vccd1 vccd1 _3425__41/A sky130_fd_sc_hd__clkbuf_16
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4330__CLK _3932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_2145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3667__A _3669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2571__A _4707_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_2301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3740_ _3748_/A vssd1 vssd1 vccd1 vccd1 _3740_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3386__B _3440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_3079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4480__CLK _3892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3671_ _4135_/A vssd1 vssd1 vccd1 vccd1 _3671_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2622_ _2622_/A _2622_/B vssd1 vssd1 vccd1 vccd1 _2623_/A sky130_fd_sc_hd__or2_1
XFILLER_31_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2553_ _4707_/Q _4706_/Q _2561_/C _2564_/A vssd1 vssd1 vccd1 vccd1 _2606_/B sky130_fd_sc_hd__a31o_1
XFILLER_29_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2484_ _4679_/Q _4678_/Q _4677_/Q _2521_/A vssd1 vssd1 vccd1 vccd1 _2507_/B sky130_fd_sc_hd__or4_4
XFILLER_9_1612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
+ _4895_/Q _2952_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_25_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4648__D _4648_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4223_ _4795_/Q vssd1 vssd1 vccd1 vccd1 _4796_/D sky130_fd_sc_hd__inv_2
XFILLER_29_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_4141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4154_ _4695_/Q vssd1 vssd1 vccd1 vccd1 _4694_/D sky130_fd_sc_hd__inv_2
XFILLER_0_3501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _4363_/CLK fanout191/X vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__dlrtn_1
X_3105_ _5024_/D _4998_/Q _4996_/Q vssd1 vssd1 vccd1 vccd1 _3105_/Y sky130_fd_sc_hd__nor3_1
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4085_ _4595_/Q vssd1 vssd1 vccd1 vccd1 _4596_/D sky130_fd_sc_hd__clkinv_2
XFILLER_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_3495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3036_ _3034_/X _3035_/Y _1791_/X vssd1 vssd1 vccd1 vccd1 _3037_/B sky130_fd_sc_hd__o21ai_1
XFILLER_18_4070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout255_A fanout256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3643_/A fanout243/X vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_14_3233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4987_ _4997_/CLK _4987_/D fanout235/X vssd1 vssd1 vccd1 vccd1 _4987_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__3577__A _3588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4823__CLK _5013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3938_ _3946_/A _3945_/A vssd1 vssd1 vccd1 vccd1 _4123_/A sky130_fd_sc_hd__xnor2_4
XFILLER_14_2543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3296__B _3438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3869_ _3941_/A vssd1 vssd1 vccd1 vccd1 _3869_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_30_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4973__CLK _4248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1825__A _4283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_2926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_4135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_3384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2656__A _2996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_2799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5032__A _5040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4353__CLK input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
+ _4953_/Q _3047_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3487__A _4127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput17 phi1b_dig_I[0] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput28 phi1b_dig_Q[3] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_2
XFILLER_10_3653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_2698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_TE_B _1845_/Y vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1906__B1 _1823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_2414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2566__A _2566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2285__B _3710_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
+ _4625_/Q _2444_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_4_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_3807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4846__CLK _4852_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4626__RESET_B fanout236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4910_ _4187_/Y _4910_/D _3505_/Y vssd1 vssd1 vccd1 vccd1 _4910_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2634__A1 _4063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2634__B2 _3875_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4841_ _3468_/Y _4841_/D fanout228/X vssd1 vssd1 vccd1 vccd1 _4841_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_2407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3397__A _4189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4931__D _4931_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4772_ _4803_/CLK _4772_/D fanout253/X vssd1 vssd1 vccd1 vccd1 _4772_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4996__CLK _5047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1984_ _1973_/C _1983_/X _1823_/X vssd1 vssd1 vccd1 vccd1 _1985_/B sky130_fd_sc_hd__o21ai_1
XFILLER_33_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3723_ _4010_/A vssd1 vssd1 vccd1 vccd1 _3723_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_2197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3844__B _3847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2605_ _4745_/D _4704_/Q vssd1 vssd1 vccd1 vccd1 _2606_/D sky130_fd_sc_hd__xnor2_1
XFILLER_28_3947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3585_ _3587_/A vssd1 vssd1 vccd1 vccd1 _3585_/Y sky130_fd_sc_hd__inv_2
X_2536_ _4682_/Q _2536_/B vssd1 vssd1 vccd1 vccd1 _4682_/D sky130_fd_sc_hd__xor2_1
XFILLER_29_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2570__B1 _2518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_3693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2467_ _4131_/D _2467_/B vssd1 vssd1 vccd1 vccd1 _5095_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__3860__A _3896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4206_ _4780_/Q vssd1 vssd1 vccd1 vccd1 _4779_/D sky130_fd_sc_hd__inv_2
XFILLER_22_3557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2398_ _4617_/Q _4616_/Q _2377_/D _2395_/B vssd1 vssd1 vccd1 vccd1 _2399_/B sky130_fd_sc_hd__a31o_1
XFILLER_29_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4137_ _4660_/Q vssd1 vssd1 vccd1 vccd1 _4661_/D sky130_fd_sc_hd__inv_2
XFILLER_25_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3659_/A fanout240/X vssd1 vssd1 vccd1 vccd1 _5076_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_0_2630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4068_ _3944_/B _3947_/B _4068_/S vssd1 vssd1 vccd1 vccd1 _4070_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4367__RESET_B fanout207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3019_ _4956_/Q _4955_/Q _2987_/D _3016_/B vssd1 vssd1 vccd1 vccd1 _3020_/B sky130_fd_sc_hd__a31o_1
XFILLER_24_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_3653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5001__CLK _1700_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3100__A _3109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_3697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2389__B1 _1975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_2963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_2985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
+ _4668_/Q _2546_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_14_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1_1_clk_master clkbuf_1_1_1_clk_master/A vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_2_clk_master/A
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__4719__CLK _4719_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_3220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout150 _2114_/Y vssd1 vssd1 vccd1 vccd1 _5041_/A sky130_fd_sc_hd__clkbuf_2
Xfanout161 _4000_/Y vssd1 vssd1 vccd1 vccd1 _4916_/CLK sky130_fd_sc_hd__buf_6
Xfanout172 _3892_/A vssd1 vssd1 vccd1 vccd1 _1952_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__4869__CLK _4905_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout183 fanout186/X vssd1 vssd1 vccd1 vccd1 fanout183/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_2333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3709__94_A _3732__95/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout194 fanout196/X vssd1 vssd1 vccd1 vccd1 fanout194/X sky130_fd_sc_hd__buf_4
XFILLER_1_2416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_4129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3575__55_A _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3425__41 _3425__41/A vssd1 vssd1 vccd1 vccd1 _3425__41/Y sky130_fd_sc_hd__inv_2
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3010__A _3030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_3737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3945__A _3945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4399__CLK _4402_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3370_ _3895_/A _3372_/B vssd1 vssd1 vccd1 vccd1 _3370_/Y sky130_fd_sc_hd__xnor2_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2321_ _4577_/Q _2321_/B vssd1 vssd1 vccd1 vccd1 _4577_/D sky130_fd_sc_hd__xnor2_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_2255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2252_ _2206_/C _2248_/Y _2173_/X vssd1 vssd1 vccd1 vccd1 _2253_/B sky130_fd_sc_hd__o21ai_1
X_5040_ _5040_/A vssd1 vssd1 vccd1 vccd1 _5040_/X sky130_fd_sc_hd__buf_2
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4926__D _4926_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2183_ _4555_/D _4497_/Q _4495_/Q vssd1 vssd1 vccd1 vccd1 _2183_/Y sky130_fd_sc_hd__nor3_1
XFILLER_22_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_2062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_2950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4460__RESET_B _3737_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5024__CLK input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3839__B _3883_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_2925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_4084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_2958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4824_ _3459_/Y _4824_/D _3636_/Y vssd1 vssd1 vccd1 vccd1 _4824_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_3837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4755_ _2631_/A _4755_/D _3421__39/Y vssd1 vssd1 vccd1 vccd1 _4755_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1967_ _4400_/Q _4399_/Q _4398_/Q _2006_/A vssd1 vssd1 vccd1 vccd1 _1992_/B sky130_fd_sc_hd__or4_1
XANTENNA__3855__A _3892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout120_A _5062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout218_A fanout219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4686_ _5007_/CLK _4686_/D _3377_/Y vssd1 vssd1 vccd1 vccd1 _4686_/Q sky130_fd_sc_hd__dfrtp_2
X_1898_ _1898_/A vssd1 vssd1 vccd1 vccd1 _1898_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_3722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3637_ _3642_/A vssd1 vssd1 vccd1 vccd1 _3637_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_3827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3568_ _3946_/A _3945_/A vssd1 vssd1 vccd1 vccd1 _3568_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwrapper_cell_loop\[0\].w1.ro_block_I.ro_pol_eve.tribuf.t_buf _2112_/A _1959_/Y vssd1
+ vssd1 vccd1 vccd1 _5089_/A sky130_fd_sc_hd__ebufn_8
X_2519_ _2479_/D _2517_/Y _2518_/X vssd1 vssd1 vccd1 vccd1 _2520_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__3590__A _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3499_ _3916_/A _3915_/A vssd1 vssd1 vccd1 vccd1 _3499_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_2_3426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_2653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_2894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_2769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_2697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2934__A _3030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3655__85 _3655__85/A vssd1 vssd1 vccd1 vccd1 _3655__85/Y sky130_fd_sc_hd__inv_2
XFILLER_25_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_2192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_3792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_4049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_3359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_3129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_2406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4900__RESET_B fanout232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3005__A _4952_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf_TE_B
+ _2443_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_2235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_2513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_2070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_3501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4997__SET_B fanout232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2870_ _4866_/Q _2870_/B vssd1 vssd1 vccd1 vccd1 _4866_/D sky130_fd_sc_hd__xnor2_1
XFILLER_16_3692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_3545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1821_ _4282_/Q _1821_/B vssd1 vssd1 vccd1 vccd1 _4282_/D sky130_fd_sc_hd__xnor2_1
XFILLER_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3675__A _4135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4540_ _4063_/B _4540_/D _3297_/Y vssd1 vssd1 vccd1 vccd1 _4540_/Q sky130_fd_sc_hd__dfrtp_1
X_1752_ _5011_/Q vssd1 vssd1 vccd1 vccd1 _5012_/D sky130_fd_sc_hd__inv_2
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3394__B _3420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4471_ _4471_/CLK _4471_/D fanout212/X vssd1 vssd1 vccd1 vccd1 _4471_/Q sky130_fd_sc_hd__dfrtp_1
X_1683_ _4913_/Q vssd1 vssd1 vccd1 vccd1 _4912_/D sky130_fd_sc_hd__inv_2
X_3422_ _3896_/A _3904_/A vssd1 vssd1 vccd1 vccd1 _3422_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__2525__B1 _2518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3361_/A vssd1 vssd1 vccd1 vccd1 _3353_/Y sky130_fd_sc_hd__inv_2
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2304_ _4584_/Q _4583_/Q _4582_/Q _2304_/D vssd1 vssd1 vccd1 vccd1 _2305_/D sky130_fd_sc_hd__and4_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3903_/A _3420_/B vssd1 vssd1 vccd1 vccd1 _3284_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_26_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5023_ input24/X input8/X fanout240/X vssd1 vssd1 vccd1 vccd1 _5024_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_6_2179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2289__C1 _3941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2235_ _4526_/Q _2235_/B vssd1 vssd1 vccd1 vccd1 _2236_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
+ _4429_/Q _2098_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_2166_ _4491_/Q _4490_/Q _2134_/D _2163_/B vssd1 vssd1 vccd1 vccd1 _2167_/B sky130_fd_sc_hd__a31o_1
XFILLER_6_1489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2097_ _4448_/Q _4447_/Q vssd1 vssd1 vccd1 vccd1 _2097_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_17_3412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout168_A _3865_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_2700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2473__B _4660_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4807_ _4809_/CLK _4807_/D fanout254/X vssd1 vssd1 vccd1 vccd1 _4807_/Q sky130_fd_sc_hd__dfrtp_1
X_2999_ _4949_/Q _2999_/B vssd1 vssd1 vccd1 vccd1 _2999_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3585__A _3587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_2933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4738_ _2631_/A _4738_/D _3414_/Y vssd1 vssd1 vccd1 vccd1 _4738_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_2955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2764__B1 _2687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_2376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4669_ _4718_/CLK _4669_/D fanout242/X vssd1 vssd1 vccd1 vccd1 _4669_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_3613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_4117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1833__A _4347_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2664__A _4763_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5040__A _5040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4907__CLK _3502_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3479__B _3913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_2822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_2210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_2708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3495__A _3934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
+ _4487_/Q _2197_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_8_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_3305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_3972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4437__CLK _5041_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_3847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2020_ _3066_/A _2020_/B _2020_/C _2020_/D vssd1 vssd1 vccd1 vccd1 _2021_/B sky130_fd_sc_hd__and4_1
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_TE_B _1919_/Y vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2574__A _2680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4587__CLK _4590_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3971_ _4420_/Q vssd1 vssd1 vccd1 vccd1 _4419_/D sky130_fd_sc_hd__inv_2
XANTENNA__2293__B _3898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2922_ _2922_/A vssd1 vssd1 vccd1 vccd1 _3030_/A sky130_fd_sc_hd__buf_6
XFILLER_31_3921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_2939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2853_ _4861_/Q _2853_/B vssd1 vssd1 vccd1 vccd1 _4861_/D sky130_fd_sc_hd__xnor2_1
XFILLER_34_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1918__A _4333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1804_ _4280_/Q _4279_/Q _1779_/D _1800_/B vssd1 vssd1 vccd1 vccd1 _1805_/B sky130_fd_sc_hd__a31o_1
XFILLER_12_2641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2784_ _4828_/Q _4827_/Q vssd1 vssd1 vccd1 vccd1 _2784_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_34_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4523_ _4533_/CLK _4523_/D fanout209/X vssd1 vssd1 vccd1 vccd1 _4523_/Q sky130_fd_sc_hd__dfrtp_4
X_1735_ _4980_/Q vssd1 vssd1 vccd1 vccd1 _4979_/D sky130_fd_sc_hd__inv_2
XFILLER_29_3850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4893__RESET_B fanout232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4454_ _3250_/Y _4454_/D _3741_/Y vssd1 vssd1 vccd1 vccd1 _4454_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_3955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1666_ _4878_/Q vssd1 vssd1 vccd1 vccd1 _4879_/D sky130_fd_sc_hd__inv_2
XFILLER_9_3977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3405_ _3947_/A _3438_/B vssd1 vssd1 vccd1 vccd1 _3405_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_2169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4385_ _3845_/Y _4385_/D _3211__16/Y vssd1 vssd1 vccd1 vccd1 _4385_/Q sky130_fd_sc_hd__dfrtp_1
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout157/X fanout203/X vssd1 vssd1 vccd1 vccd1 _5082_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_28_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ _3340_/A vssd1 vssd1 vccd1 vccd1 _3336_/Y sky130_fd_sc_hd__inv_2
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2468__B _3929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5006_ _3560_/Y _5006_/D _3583_/Y vssd1 vssd1 vccd1 vccd1 _5006_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_2_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2218_ _4521_/Q _4520_/Q _2218_/C vssd1 vssd1 vccd1 vccd1 _2218_/X sky130_fd_sc_hd__and3_1
XFILLER_22_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2149_ _4485_/Q _2145_/C _2146_/B vssd1 vssd1 vccd1 vccd1 _2150_/B sky130_fd_sc_hd__a21bo_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_3718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_4121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_2405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_3442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_2438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1828__A _1909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_2752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_4100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_4094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4563__RESET_B fanout223/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2659__A _4763_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5035__A _5043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input13_A comp_high_Q[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_2630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_2685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_2516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output81_A _5078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4170_ _4727_/Q vssd1 vssd1 vccd1 vccd1 _4726_/D sky130_fd_sc_hd__inv_2
XFILLER_4_3841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3121_ _5012_/Q _5011_/Q vssd1 vssd1 vccd1 vccd1 _3121_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_7_2274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_2910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3052_ _4978_/Q _4977_/Q vssd1 vssd1 vccd1 vccd1 _3052_/Y sky130_fd_sc_hd__xnor2_2
X_2003_ _2922_/A vssd1 vssd1 vccd1 vccd1 _2003_/X sky130_fd_sc_hd__buf_6
XFILLER_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3954_ _4385_/Q vssd1 vssd1 vccd1 vccd1 _4386_/D sky130_fd_sc_hd__inv_2
XANTENNA__5021__RESET_B fanout207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_2883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2905_ _4893_/Q _2901_/C _2902_/B vssd1 vssd1 vccd1 vccd1 _2906_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__3847__B _3848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_3751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3885_ _3885_/A _3886_/B vssd1 vssd1 vccd1 vccd1 _4363_/D sky130_fd_sc_hd__xnor2_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2836_ _4856_/Q _2836_/B vssd1 vssd1 vccd1 vccd1 _4856_/D sky130_fd_sc_hd__xnor2_1
XFILLER_30_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_GATE_N
+ _5063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2767_ _4838_/D _4812_/Q _4810_/Q vssd1 vssd1 vccd1 vccd1 _2767_/Y sky130_fd_sc_hd__nor3_1
XFILLER_27_3809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3749_/A fanout187/X vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_12_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4506_ _3932_/A _4506_/D _3277_/Y vssd1 vssd1 vccd1 vccd1 _4506_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout200_A fanout221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1718_ _4945_/Q vssd1 vssd1 vccd1 vccd1 _4946_/D sky130_fd_sc_hd__inv_2
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2698_ _2696_/X _2697_/Y _2687_/X vssd1 vssd1 vccd1 vccd1 _2699_/B sky130_fd_sc_hd__o21ai_1
XFILLER_8_2016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4437_ _5041_/A _4437_/D fanout198/X vssd1 vssd1 vccd1 vccd1 _4437_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_3408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4368_ _4368_/CLK _4368_/D fanout204/X vssd1 vssd1 vccd1 vccd1 _4368_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input5_A comp_high_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _3891_/A _3889_/A vssd1 vssd1 vccd1 vccd1 _3319_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_3_3351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _3914_/B _4299_/D _3780__121/Y vssd1 vssd1 vccd1 vccd1 _4299_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3103__A _4994_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_3061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2942__A _4931_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4282__CLK _4288_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_4009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_2582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3209__15_A _3264__22/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xw0.ro_block_Q.ro_pol_eve.tribuf.t_buf _1928_/A _1771_/Y vssd1 vssd1 vccd1 vccd1 _5091_/A
+ sky130_fd_sc_hd__ebufn_8
XFILLER_2_2193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3013__A _3030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3948__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2852__A _2916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_3036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_2471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4625__CLK _5043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3670_ _5060_/A vssd1 vssd1 vccd1 vccd1 _4135_/A sky130_fd_sc_hd__buf_8
XFILLER_16_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2621_ _4742_/D _4743_/Q vssd1 vssd1 vccd1 vccd1 _2622_/B sky130_fd_sc_hd__and2b_1
XANTENNA__2177__A1 _2133_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4775__CLK _4811_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2552_ _4705_/Q vssd1 vssd1 vccd1 vccd1 _2564_/A sky130_fd_sc_hd__inv_2
XFILLER_6_3925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2483_ _4741_/D _4683_/Q _4681_/Q _4680_/Q vssd1 vssd1 vccd1 vccd1 _2521_/A sky130_fd_sc_hd__or4_1
XFILLER_9_2358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4222_ _4796_/Q vssd1 vssd1 vccd1 vccd1 _4795_/D sky130_fd_sc_hd__inv_2
XFILLER_29_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4153_ _4692_/Q vssd1 vssd1 vccd1 vccd1 _4693_/D sky130_fd_sc_hd__inv_2
XFILLER_29_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3104_ _5024_/D _4998_/Q _4996_/Q vssd1 vssd1 vccd1 vccd1 _3104_/X sky130_fd_sc_hd__and3_1
XFILLER_0_3524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4084_ _4596_/Q vssd1 vssd1 vccd1 vccd1 _4595_/D sky130_fd_sc_hd__inv_2
XFILLER_23_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3035_ _5020_/D _4962_/Q _4960_/Q vssd1 vssd1 vccd1 vccd1 _3035_/Y sky130_fd_sc_hd__nor3_1
XFILLER_20_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_2795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_3201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout150_A _2114_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4986_ _4997_/CLK _4986_/D fanout234/X vssd1 vssd1 vccd1 vccd1 _4986_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_3857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_3245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3937_ _4379_/Q vssd1 vssd1 vccd1 vccd1 _3945_/A sky130_fd_sc_hd__buf_12
XFILLER_10_3109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_3289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_3581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3868_ _3916_/A _3915_/A vssd1 vssd1 vccd1 vccd1 _3941_/A sky130_fd_sc_hd__xnor2_4
XFILLER_20_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2819_ _4860_/Q _4859_/Q _4858_/Q _2819_/D vssd1 vssd1 vccd1 vccd1 _2829_/C sky130_fd_sc_hd__and4_1
XANTENNA__3593__A _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3799_ _4297_/Q vssd1 vssd1 vccd1 vccd1 _4296_/D sky130_fd_sc_hd__inv_2
XFILLER_27_3606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4839__D _4839_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_4086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_TE_B
+ _2028_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_3249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1841__A _3066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout128/X fanout246/X vssd1 vssd1 vccd1 vccd1 _5077_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_25_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4648__CLK input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4996__RESET_B fanout242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4925__RESET_B _3605_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3487__B _4129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_2611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_3389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4798__CLK _4811_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput18 phi1b_dig_I[1] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput29 phi1b_dig_Q[4] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_2098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2159__A1 _4488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_2404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_3833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_2255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_2069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3678__A _4135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4840_ input22/X _4840_/D fanout227/X vssd1 vssd1 vccd1 vccd1 _4840_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2582__A _4710_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_4119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3397__B _4190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4771_ _4812_/CLK _4771_/D fanout253/X vssd1 vssd1 vccd1 vccd1 _4771_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1983_ _4393_/Q _1983_/B vssd1 vssd1 vccd1 vccd1 _1983_/X sky130_fd_sc_hd__and2b_1
X_3722_ _4469_/Q vssd1 vssd1 vccd1 vccd1 _4010_/A sky130_fd_sc_hd__buf_6
XFILLER_31_2165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_3915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2604_ _4717_/Q _2604_/B vssd1 vssd1 vccd1 vccd1 _4717_/D sky130_fd_sc_hd__xnor2_1
X_3584_ _3587_/A vssd1 vssd1 vccd1 vccd1 _3584_/Y sky130_fd_sc_hd__inv_2
X_2535_ _3066_/A _2535_/B _2535_/C _2535_/D vssd1 vssd1 vccd1 vccd1 _2536_/B sky130_fd_sc_hd__and4_1
XANTENNA__2570__A1 _2561_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2466_ _2470_/A1 _2463_/X _2465_/X _4131_/B vssd1 vssd1 vccd1 vccd1 _2467_/B sky130_fd_sc_hd__o22a_1
XFILLER_22_3525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4205_ _4777_/Q vssd1 vssd1 vccd1 vccd1 _4778_/D sky130_fd_sc_hd__inv_2
XANTENNA__3860__B _3904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_3569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2397_ _4614_/Q _2397_/B vssd1 vssd1 vccd1 vccd1 _4614_/D sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout198_A fanout221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_A
+ _4522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4136_ _4661_/Q vssd1 vssd1 vccd1 vccd1 _4660_/D sky130_fd_sc_hd__inv_2
XFILLER_0_3343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4067_ _4566_/Q _4565_/Q vssd1 vssd1 vccd1 vccd1 _4068_/S sky130_fd_sc_hd__xnor2_4
XFILLER_16_4019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3018_ _4953_/Q _3018_/B vssd1 vssd1 vccd1 vccd1 _4953_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_1930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3588__A _3588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4969_ _4187_/Y _4969_/D _3538_/Y vssd1 vssd1 vccd1 vccd1 _4969_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_14_3097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_3974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1836__A _4347_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_2702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2010__B1 _2003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4320__CLK _4324_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_3193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout140 _2285_/Y vssd1 vssd1 vccd1 vccd1 _5034_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_3035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout151 _4920_/CLK vssd1 vssd1 vccd1 vccd1 _4063_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_5_3287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout162 _5013_/CLK vssd1 vssd1 vccd1 vccd1 _4063_/C sky130_fd_sc_hd__buf_6
XFILLER_21_2312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5043__A _5043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout173 _4121_/Y vssd1 vssd1 vccd1 vccd1 _4248_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout184 fanout185/X vssd1 vssd1 vccd1 vccd1 fanout184/X sky130_fd_sc_hd__buf_2
Xfanout195 fanout196/X vssd1 vssd1 vccd1 vccd1 fanout195/X sky130_fd_sc_hd__clkbuf_4
XFILLER_25_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3498__A _3498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1824__B1 _1823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_clk_master clkbuf_2_3_0_clk_master/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clk_master/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_32_2474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2320_ _2327_/A _2320_/B vssd1 vssd1 vccd1 vccd1 _2321_/B sky130_fd_sc_hd__nand2_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4813__CLK _4247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2577__A _2680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2251_ _4528_/Q _2251_/B vssd1 vssd1 vccd1 vccd1 _4528_/D sky130_fd_sc_hd__xnor2_1
XFILLER_23_3889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2182_ _4555_/D _4497_/Q _4495_/Q vssd1 vssd1 vccd1 vccd1 _2182_/X sky130_fd_sc_hd__and3_1
XFILLER_1_3641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_4030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_3941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_4074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4823_ _5013_/CLK _4823_/D _3458_/Y vssd1 vssd1 vccd1 vccd1 _4823_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_3985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_3849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4754_ _3420_/Y _4754_/D _3657__86/Y vssd1 vssd1 vccd1 vccd1 _4754_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1966_ _4462_/D _4404_/Q _4402_/Q _4401_/Q vssd1 vssd1 vccd1 vccd1 _2006_/A sky130_fd_sc_hd__or4_1
XANTENNA__3775__114_A _3776__115/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
+ _4799_/Q _2783_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_2525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3705_ _4071_/A vssd1 vssd1 vccd1 vccd1 _3705_/Y sky130_fd_sc_hd__inv_2
X_4685_ _4248_/D _4685_/D _3679_/Y vssd1 vssd1 vccd1 vccd1 _4685_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_1982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1897_ _4319_/Q _1897_/B vssd1 vssd1 vccd1 vccd1 _4319_/D sky130_fd_sc_hd__xnor2_1
X_3636_ _3642_/A vssd1 vssd1 vccd1 vccd1 _3636_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout113_A _3588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3567_ _3571_/A vssd1 vssd1 vccd1 vccd1 _3567_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_3609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3871__A _3941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_4023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_4034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2518_ _2858_/A vssd1 vssd1 vccd1 vccd1 _2518_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3498_ _3498_/A vssd1 vssd1 vccd1 vccd1 _3498_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_2919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4493__CLK _4533_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2449_ _2449_/A vssd1 vssd1 vccd1 vccd1 _2449_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_2610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_2862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3680__87_A _3683__90/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4119_ _4645_/Q vssd1 vssd1 vccd1 vccd1 _4646_/D sky130_fd_sc_hd__inv_2
XFILLER_29_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5099_ _5099_/A vssd1 vssd1 vccd1 vccd1 _5099_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3111__A _5024_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_3462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_2469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_2182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5038__A _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_3305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4836__CLK input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_3338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
+ _4857_/Q _2883_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_2587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2397__A _4614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4986__CLK _4997_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_2120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3005__B _3005_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_2153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_3983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf _4318_/Q _1915_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_16_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[3\].w1.ro_block_Q.ro_pol.tribuf.t_buf _2623_/X _2473_/Y vssd1
+ vssd1 vccd1 vccd1 _5090_/A sky130_fd_sc_hd__ebufn_8
XANTENNA__3021__A _4954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_2525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2470__B1 _2465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1820_ _1909_/A _1820_/B vssd1 vssd1 vccd1 vccd1 _1821_/B sky130_fd_sc_hd__nand2_2
XFILLER_12_3557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1751_ _5012_/Q vssd1 vssd1 vccd1 vccd1 _5011_/D sky130_fd_sc_hd__inv_2
XFILLER_8_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4470_ _4658_/CLK _4470_/D fanout211/X vssd1 vssd1 vccd1 vccd1 _4470_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_3019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1682_ _4910_/Q vssd1 vssd1 vccd1 vccd1 _4911_/D sky130_fd_sc_hd__inv_2
XFILLER_32_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3691__A _3695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3352_ _3935_/A _3440_/B vssd1 vssd1 vccd1 vccd1 _3352_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_7_3861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _4586_/Q _4585_/Q _2303_/C vssd1 vssd1 vccd1 vccd1 _2304_/D sky130_fd_sc_hd__and3_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _3287_/A vssd1 vssd1 vccd1 vccd1 _3283_/Y sky130_fd_sc_hd__inv_2
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ input32/X _5022_/D fanout208/X vssd1 vssd1 vccd1 vccd1 _5022_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2234_ _4523_/Q _2234_/B vssd1 vssd1 vccd1 vccd1 _4523_/D sky130_fd_sc_hd__xnor2_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_2974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_3471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2165_ _4488_/Q _2165_/B vssd1 vssd1 vccd1 vccd1 _4488_/D sky130_fd_sc_hd__xnor2_1
X_2096_ _4446_/Q _4445_/Q vssd1 vssd1 vccd1 vccd1 _2096_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_17_2712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4709__CLK _4709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_3793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2770__A _4838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout230_A input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4806_ _4812_/CLK _4806_/D fanout256/X vssd1 vssd1 vccd1 vccd1 _4806_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_2789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2998_ _4950_/Q _4949_/Q _2998_/C vssd1 vssd1 vccd1 vccd1 _2998_/X sky130_fd_sc_hd__and3_1
XFILLER_30_2923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4859__CLK _4865_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1949_ _3888_/A _3898_/B _1948_/Y _3892_/B vssd1 vssd1 vccd1 vccd1 _1951_/B sky130_fd_sc_hd__o211a_1
X_4737_ _3413_/Y _4737_/D _3660_/Y vssd1 vssd1 vccd1 vccd1 _4737_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_3078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4668_ _4718_/CLK _4668_/D fanout242/X vssd1 vssd1 vccd1 vccd1 _4668_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_28_3531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3619_ _4256_/A vssd1 vssd1 vccd1 vccd1 _3619_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_3625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_4129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_3553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_3636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4599_ _4920_/CLK _4599_/D _3330_/Y vssd1 vssd1 vccd1 vccd1 _4599_/Q sky130_fd_sc_hd__dfrtp_1
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout144/X fanout215/X vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_6_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_TE_B
+ _2949_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1833__B _4289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_3213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_3163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_3257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2945__A _4931_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4389__CLK _4429_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2383__C _4614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf_TE_B
+ _2103_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_3270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2680__A _2680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3495__B _3933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_4029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_GATE_N _5048_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_2423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_A
+ _4671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_2445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_2309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_3859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2855__A _2916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3195__3_A _3199__7/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3970_ _4417_/Q vssd1 vssd1 vccd1 vccd1 _4418_/D sky130_fd_sc_hd__inv_2
XANTENNA__2293__C _3908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2921_ _4896_/Q _2921_/B vssd1 vssd1 vccd1 vccd1 _4896_/D sky130_fd_sc_hd__xnor2_1
XFILLER_34_2322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3686__A _3695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_3310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2852_ _2916_/A _2852_/B vssd1 vssd1 vccd1 vccd1 _2853_/B sky130_fd_sc_hd__nand2_1
XFILLER_12_4077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1803_ _4277_/Q _1803_/B vssd1 vssd1 vccd1 vccd1 _4277_/D sky130_fd_sc_hd__xnor2_1
X_2783_ _4826_/Q _4825_/Q vssd1 vssd1 vccd1 vccd1 _2783_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_12_2653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4522_ _4533_/CLK _4522_/D fanout209/X vssd1 vssd1 vccd1 vccd1 _4522_/Q sky130_fd_sc_hd__dfrtp_2
X_1734_ _4977_/Q vssd1 vssd1 vccd1 vccd1 _4978_/D sky130_fd_sc_hd__inv_2
XFILLER_12_1930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2210__A3 _2218_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4453_ _3914_/A _4453_/D _3249_/Y vssd1 vssd1 vccd1 vccd1 _4453_/Q sky130_fd_sc_hd__dfrtp_1
X_1665_ _4879_/Q vssd1 vssd1 vccd1 vccd1 _4878_/D sky130_fd_sc_hd__inv_2
XFILLER_9_3967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3404_ _3414_/A vssd1 vssd1 vccd1 vccd1 _3404_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_3809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4384_ _3210_/Y _4384_/D _3761__101/Y vssd1 vssd1 vccd1 vccd1 _4384_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3335_ _3917_/A _3444_/B vssd1 vssd1 vccd1 vccd1 _3335_/Y sky130_fd_sc_hd__xnor2_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _3600_/A vssd1 vssd1 vccd1 vccd1 _3266_/X sky130_fd_sc_hd__buf_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _4187_/Y _5005_/D _3559_/Y vssd1 vssd1 vccd1 vccd1 _5005_/Q sky130_fd_sc_hd__dfrtp_1
X_3778__119 _3781__122/A vssd1 vssd1 vccd1 vccd1 _3778__119/Y sky130_fd_sc_hd__inv_2
X_2217_ _4518_/Q _2217_/B vssd1 vssd1 vccd1 vccd1 _4518_/D sky130_fd_sc_hd__xor2_1
XFILLER_3_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout180_A _3738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4531__CLK _4532_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2148_ _2148_/A _2148_/B vssd1 vssd1 vccd1 vccd1 _4483_/D sky130_fd_sc_hd__xnor2_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2079_ _2178_/A _2079_/B vssd1 vssd1 vccd1 vccd1 _2080_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4681__CLK _4719_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3596__A _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_2417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
+ _4618_/Q _2436_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout158/X fanout206/X vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_17_1885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_2764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_2786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1844__A _4289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2659__B _2659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3761__101 _3765__105/A vssd1 vssd1 vccd1 vccd1 _3761__101/Y sky130_fd_sc_hd__inv_2
XFILLER_24_2502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5051__A _5059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_3321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2976__B2 _4126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_3641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5063_/A fanout251/X vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_13_3685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3169__65_A _3169__65/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4404__CLK _4429_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_2424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_2518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
+ _4676_/Q _2538_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_3120_ _5010_/Q _5009_/Q vssd1 vssd1 vccd1 vccd1 _3120_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__4554__CLK input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4273__RESET_B _5048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3051_ _4976_/Q _4975_/Q vssd1 vssd1 vccd1 vccd1 _3051_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_20_2922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2585__A _4711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2002_ _4400_/Q _4399_/Q _2006_/A vssd1 vssd1 vccd1 vccd1 _2002_/Y sky130_fd_sc_hd__nor3_1
XFILLER_14_4117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3953_ _4386_/Q vssd1 vssd1 vccd1 vccd1 _4385_/D sky130_fd_sc_hd__inv_2
XFILLER_14_2715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2904_ _2904_/A _2904_/B vssd1 vssd1 vccd1 vccd1 _4891_/D sky130_fd_sc_hd__xnor2_1
X_3884_ _3882_/Y _3888_/A _3884_/S vssd1 vssd1 vccd1 vccd1 _3886_/B sky130_fd_sc_hd__mux2_1
XFILLER_17_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_TE_B
+ _2096_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_3151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2835_ _2916_/A _2835_/B vssd1 vssd1 vccd1 vccd1 _2836_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2766_ _4838_/D _4812_/Q _4810_/Q vssd1 vssd1 vccd1 vccd1 _2766_/X sky130_fd_sc_hd__and3_1
X_1717_ _4946_/Q vssd1 vssd1 vccd1 vccd1 _4945_/D sky130_fd_sc_hd__inv_2
X_3528__52 _3528__52/A vssd1 vssd1 vccd1 vccd1 _3528__52/Y sky130_fd_sc_hd__inv_2
X_4505_ _3276_/Y _4505_/D _3728_/Y vssd1 vssd1 vccd1 vccd1 _4505_/Q sky130_fd_sc_hd__dfrtp_1
X_2697_ _4834_/D _4776_/Q _4774_/Q vssd1 vssd1 vccd1 vccd1 _2697_/Y sky130_fd_sc_hd__nor3_1
XFILLER_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4436_ _5041_/A _4436_/D fanout198/X vssd1 vssd1 vccd1 vccd1 _4436_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__2479__B _4676_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_4020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_2905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4367_ _4472_/CLK _4367_/D fanout207/X vssd1 vssd1 vccd1 vccd1 _4367_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_4075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _2286_/B _4298_/D _3157__57/Y vssd1 vssd1 vccd1 vccd1 _4298_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_2719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161__61 _3169__65/A vssd1 vssd1 vccd1 vccd1 _3161__61/Y sky130_fd_sc_hd__inv_2
XANTENNA__2495__A _2566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3249_ _3255_/A vssd1 vssd1 vccd1 vccd1 _3249_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_3305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_3316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2655__B1 _2661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_3505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2942__B _4905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1839__A _1839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_2361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_2203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_TE_B
+ _2542_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4427__CLK _4429_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5046__A _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4577__CLK _4590_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4713__RESET_B fanout255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_2540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
+ _4391_/Q _2029_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout119/X fanout248/X vssd1 vssd1 vccd1 vccd1 _5078_/A sky130_fd_sc_hd__dlrtn_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_2169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2620_ _2620_/A vssd1 vssd1 vccd1 vccd1 _2622_/A sky130_fd_sc_hd__clkbuf_2
X_3768__107 _3770__109/A vssd1 vssd1 vccd1 vccd1 _3768__107/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_2792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_3005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2551_ _4710_/Q _4709_/Q _4708_/Q _2551_/D vssd1 vssd1 vccd1 vccd1 _2561_/C sky130_fd_sc_hd__and4_2
XFILLER_9_2326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2482_ _4671_/Q _4670_/Q _2490_/C _2493_/A vssd1 vssd1 vccd1 vccd1 _2535_/B sky130_fd_sc_hd__a31o_1
XFILLER_29_2265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_3937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4221_ _4793_/Q vssd1 vssd1 vccd1 vccd1 _4794_/D sky130_fd_sc_hd__inv_2
XFILLER_25_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_3959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4152_ _4693_/Q vssd1 vssd1 vccd1 vccd1 _4692_/D sky130_fd_sc_hd__inv_2
XFILLER_7_2061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3103_ _4994_/Q _3103_/B vssd1 vssd1 vccd1 vccd1 _4994_/D sky130_fd_sc_hd__xnor2_1
X_4083_ _4593_/Q vssd1 vssd1 vccd1 vccd1 _4594_/D sky130_fd_sc_hd__inv_2
XFILLER_3_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_2993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3034_ _5020_/D _4962_/Q _4960_/Q vssd1 vssd1 vccd1 vccd1 _3034_/X sky130_fd_sc_hd__and3_1
XFILLER_23_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_3213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4985_ _4997_/CLK _4985_/D fanout234/X vssd1 vssd1 vccd1 vccd1 _4985_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3936_ _4380_/Q vssd1 vssd1 vccd1 vccd1 _3946_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_14_3257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3867_ _4373_/Q vssd1 vssd1 vccd1 vccd1 _3915_/A sky130_fd_sc_hd__buf_12
XANTENNA__3874__A _3897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2818_ _4863_/Q _4862_/Q _4861_/Q _2818_/D vssd1 vssd1 vccd1 vccd1 _2819_/D sky130_fd_sc_hd__and4_1
X_3798_ _4294_/Q vssd1 vssd1 vccd1 vccd1 _4295_/D sky130_fd_sc_hd__inv_2
XFILLER_14_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2749_ _2720_/D _2748_/X _2687_/X vssd1 vssd1 vccd1 vccd1 _2750_/B sky130_fd_sc_hd__o21ai_1
XFILLER_25_4043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_3561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_3414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4419_ _3899_/A _4419_/D _3229_/Y vssd1 vssd1 vccd1 vccd1 _4419_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_2713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_3217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3114__A _3114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_4003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_4025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_3313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput19 phi1b_dig_I[2] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_3845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_3889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2863__A _2916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4770_ _4812_/CLK _4770_/D fanout253/X vssd1 vssd1 vccd1 vccd1 _4770_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1982_ _4394_/Q _1982_/B vssd1 vssd1 vccd1 vccd1 _1983_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4742__CLK input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3721_ _3721_/A vssd1 vssd1 vccd1 vccd1 _3721_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_3891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3694__A _3695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3652_ _4195_/A vssd1 vssd1 vccd1 vccd1 _3652_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_3905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2603_ _2680_/A _2603_/B vssd1 vssd1 vccd1 vccd1 _2604_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4892__CLK _4901_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3583_ _3587_/A vssd1 vssd1 vccd1 vccd1 _3583_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_3949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2534_ _4741_/D _4668_/Q vssd1 vssd1 vccd1 vccd1 _2535_/D sky130_fd_sc_hd__xnor2_1
XFILLER_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_3723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_2134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2465_ _2289_/X _2464_/Y _3910_/A vssd1 vssd1 vccd1 vccd1 _2465_/X sky130_fd_sc_hd__a21o_2
XANTENNA__1942__A _3882_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_2167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4204_ _4778_/Q vssd1 vssd1 vccd1 vccd1 _4777_/D sky130_fd_sc_hd__clkinv_2
XFILLER_22_3537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2396_ _2387_/C _2395_/X _2344_/X vssd1 vssd1 vccd1 vccd1 _2397_/B sky130_fd_sc_hd__o21ai_1
XFILLER_26_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4135_ _4135_/A vssd1 vssd1 vccd1 vccd1 _4655_/D sky130_fd_sc_hd__inv_2
XFILLER_29_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4066_ _4564_/Q _4066_/B vssd1 vssd1 vccd1 vccd1 _4564_/D sky130_fd_sc_hd__xor2_1
XANTENNA__3869__A _3941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3017_ _2988_/D _3016_/X _2858_/X vssd1 vssd1 vccd1 vccd1 _3018_/B sky130_fd_sc_hd__o21ai_1
XFILLER_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2773__A _4838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_2593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4968_ _3537_/Y _4968_/D _3595_/Y vssd1 vssd1 vccd1 vccd1 _4968_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_3065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3919_ _4375_/Q vssd1 vssd1 vccd1 vccd1 _3923_/A sky130_fd_sc_hd__buf_8
X_4899_ _4901_/CLK _4899_/D fanout232/X vssd1 vssd1 vccd1 vccd1 _4899_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_2217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1836__B _4289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4376__RESET_B fanout214/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0__1648_ _3368_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__1648_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_27_3415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3109__A _3109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2013__A _4462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_2714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2948__A _3114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _4359_/CLK fanout190/X vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_25_3161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout130 _4748_/Q vssd1 vssd1 vccd1 vccd1 _5061_/A sky130_fd_sc_hd__buf_4
XFILLER_5_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2849__B1 _2687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_2460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout141 _2285_/Y vssd1 vssd1 vccd1 vccd1 _4533_/CLK sky130_fd_sc_hd__buf_2
Xfanout152 _4920_/CLK vssd1 vssd1 vccd1 vccd1 _4131_/B sky130_fd_sc_hd__buf_2
XFILLER_25_2471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4615__CLK _4626_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout163 _3939_/Y vssd1 vssd1 vccd1 vccd1 _5013_/CLK sky130_fd_sc_hd__buf_8
XFILLER_5_3299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout174 _4121_/Y vssd1 vssd1 vccd1 vccd1 _5007_/CLK sky130_fd_sc_hd__clkbuf_4
Xfanout185 fanout186/X vssd1 vssd1 vccd1 vccd1 fanout185/X sky130_fd_sc_hd__clkbuf_2
Xfanout196 fanout221/X vssd1 vssd1 vccd1 vccd1 fanout196/X sky130_fd_sc_hd__clkbuf_4
XFILLER_1_1717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4765__CLK _4811_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1824__A1 _1778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_3121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3026__B1 _1791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_A
+ _4953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4324__SET_B fanout194/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2858__A _2858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ _2327_/A _2250_/B vssd1 vssd1 vccd1 vccd1 _2251_/B sky130_fd_sc_hd__nand2_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4295__CLK _3941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2181_ _4493_/Q _2181_/B vssd1 vssd1 vccd1 vccd1 _4493_/D sky130_fd_sc_hd__xnor2_1
XFILLER_1_3653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3689__A _3695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_4042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3017__B1 _2858_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4822_ _3457_/Y _4822_/D _3637_/Y vssd1 vssd1 vccd1 vccd1 _4822_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_2239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_3205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_3997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4753_ _3861_/Y _4753_/D _3419__38/Y vssd1 vssd1 vccd1 vccd1 _4753_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_2662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1965_ _4392_/Q _4391_/Q _1973_/C _1977_/A vssd1 vssd1 vccd1 vccd1 _2020_/B sky130_fd_sc_hd__a31o_1
XFILLER_30_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1937__A _3892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3704_ _4071_/A vssd1 vssd1 vccd1 vccd1 _3704_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1896_ _1857_/D _1895_/Y _1823_/X vssd1 vssd1 vccd1 vccd1 _1897_/B sky130_fd_sc_hd__o21ai_1
X_4684_ _4187_/Y _4684_/D _3376_/Y vssd1 vssd1 vccd1 vccd1 _4684_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_1972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3635_ _3642_/A vssd1 vssd1 vccd1 vccd1 _3635_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_3746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout106_A _3135_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3566_ _4001_/A _4005_/A vssd1 vssd1 vccd1 vccd1 _3566_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_3779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2517_ _4679_/Q _4678_/Q _2521_/A vssd1 vssd1 vccd1 vccd1 _2517_/Y sky130_fd_sc_hd__nor3_1
XFILLER_2_4107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3497_ _3924_/A _3923_/A vssd1 vssd1 vccd1 vccd1 _3497_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_2_4129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2448_ _2448_/A _2448_/B vssd1 vssd1 vccd1 vccd1 _2449_/A sky130_fd_sc_hd__or2_1
XFILLER_22_3345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_2841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_2622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_3389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2379_ _4614_/Q _4613_/Q _2387_/C _2390_/A vssd1 vssd1 vccd1 vccd1 _2432_/B sky130_fd_sc_hd__a31o_1
XFILLER_6_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4788__CLK _3438_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4118_ _4646_/Q vssd1 vssd1 vccd1 vccd1 _4645_/D sky130_fd_sc_hd__inv_2
X_5098_ _5098_/A vssd1 vssd1 vccd1 vccd1 _5098_/X sky130_fd_sc_hd__clkbuf_1
X_4049_ _4545_/Q vssd1 vssd1 vccd1 vccd1 _4544_/D sky130_fd_sc_hd__inv_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_4142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_3441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2008__A _2061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4557__RESET_B fanout199/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_4029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_2500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_3317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5054__A _5062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_2638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf_TE_B
+ _2617_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout136/X fanout238/X vssd1 vssd1 vccd1 vccd1 _5084_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_5_3085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_3995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3302__A _3917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2470__A1 _2470_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_2261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1750_ _5009_/Q vssd1 vssd1 vccd1 vccd1 _5010_/D sky130_fd_sc_hd__inv_2
XFILLER_30_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_2879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1681_ _4911_/Q vssd1 vssd1 vccd1 vccd1 _4910_/D sky130_fd_sc_hd__inv_2
X_3420_ _3896_/A _3420_/B vssd1 vssd1 vccd1 vccd1 _3420_/Y sky130_fd_sc_hd__xnor2_1
X_3351_ _3361_/A vssd1 vssd1 vccd1 vccd1 _3351_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2588__A _4712_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2302_ _4648_/D _4590_/Q _4588_/Q _4587_/Q vssd1 vssd1 vccd1 vccd1 _2303_/C sky130_fd_sc_hd__and4_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _3912_/A _3446_/B vssd1 vssd1 vccd1 vccd1 _3282_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4930__CLK input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _2327_/A _2233_/B vssd1 vssd1 vccd1 vccd1 _2234_/B sky130_fd_sc_hd__nand2_1
X_5021_ input32/X _5021_/D fanout207/X vssd1 vssd1 vccd1 vccd1 _5022_/D sky130_fd_sc_hd__dfrtp_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2289__A1 _3898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2164_ _2135_/D _2163_/X _2003_/X vssd1 vssd1 vccd1 vccd1 _2165_/B sky130_fd_sc_hd__o21ai_1
XFILLER_17_4115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2095_ _4444_/Q _4443_/Q vssd1 vssd1 vccd1 vccd1 _2095_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__3212__A _3848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_2724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4310__CLK _4324_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_2014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_2757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4650__RESET_B fanout207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4805_ _4809_/CLK _4805_/D fanout253/X vssd1 vssd1 vccd1 vccd1 _4805_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_2047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2997_ _4947_/Q _2997_/B vssd1 vssd1 vccd1 vccd1 _4947_/D sky130_fd_sc_hd__xor2_1
XFILLER_9_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_2470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4736_ _4852_/CLK _4736_/D _3412_/Y vssd1 vssd1 vccd1 vccd1 _4736_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout223_A fanout230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1948_ _3888_/A _3900_/B vssd1 vssd1 vccd1 vccd1 _1948_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4667_ _3374_/Y _4667_/D _3680__87/Y vssd1 vssd1 vccd1 vccd1 _4667_/Q sky130_fd_sc_hd__dfrtp_1
X_1879_ _4316_/Q _4315_/Q _1858_/D _1876_/B vssd1 vssd1 vccd1 vccd1 _1880_/B sky130_fd_sc_hd__a31o_1
XANTENNA__3882__A _3882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3618_ _4256_/A vssd1 vssd1 vccd1 vccd1 _3618_/Y sky130_fd_sc_hd__inv_2
X_4598_ _3329_/Y _4598_/D _3702_/Y vssd1 vssd1 vccd1 vccd1 _4598_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_3648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_2925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3549_ _3934_/A _3933_/A vssd1 vssd1 vccd1 vccd1 _3549_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_8_2936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
+ _4988_/Q _3118_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_8_2947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_2897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5024__D _5024_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_2524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__0630_ clkbuf_0__0630_/X vssd1 vssd1 vccd1 vccd1 _3683__90/A sky130_fd_sc_hd__clkbuf_16
XFILLER_22_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_3801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_2857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4391__RESET_B fanout194/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_2109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4803__CLK _4803_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5049__A _5057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_2570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_4008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3706__91 _3732__95/A vssd1 vssd1 vccd1 vccd1 _3706__91/Y sky130_fd_sc_hd__inv_2
XFILLER_27_2363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_3827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_2249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_3781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_4001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2293__D _3941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2920_ _2891_/D _2919_/X _2858_/X vssd1 vssd1 vccd1 vccd1 _2921_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__2871__A _4927_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2851_ _4863_/Q _4862_/Q _2818_/D _2848_/B vssd1 vssd1 vccd1 vccd1 _2852_/B sky130_fd_sc_hd__a31o_1
XFILLER_12_3322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4483__CLK _5042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_2367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1802_ _1789_/C _1800_/X _3109_/A vssd1 vssd1 vccd1 vccd1 _1803_/B sky130_fd_sc_hd__o21ai_1
XFILLER_34_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2782_ _4824_/Q _4823_/Q vssd1 vssd1 vccd1 vccd1 _2782_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_2665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4521_ _4532_/CLK _4521_/D fanout211/X vssd1 vssd1 vccd1 vccd1 _4521_/Q sky130_fd_sc_hd__dfrtp_4
X_1733_ _4978_/Q vssd1 vssd1 vccd1 vccd1 _4977_/D sky130_fd_sc_hd__inv_2
XFILLER_15_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4452_ _3248_/Y _4452_/D _3742_/Y vssd1 vssd1 vccd1 vccd1 _4452_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_12_1986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1664_ _4876_/Q vssd1 vssd1 vccd1 vccd1 _4877_/D sky130_fd_sc_hd__inv_2
XFILLER_28_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3403_ _4004_/A _3491_/B vssd1 vssd1 vccd1 vccd1 _3403_/Y sky130_fd_sc_hd__xnor2_1
X_4383_ _3845_/Y _4383_/D _3209__15/Y vssd1 vssd1 vccd1 vccd1 _4383_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ _3340_/A vssd1 vssd1 vccd1 vccd1 _3334_/Y sky130_fd_sc_hd__inv_2
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _3885_/A _3886_/A vssd1 vssd1 vccd1 vccd1 _3265_/Y sky130_fd_sc_hd__xnor2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _3558_/Y _5004_/D _3584_/Y vssd1 vssd1 vccd1 vccd1 _5004_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_26_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2216_ _2996_/A _2262_/B _2262_/C vssd1 vssd1 vccd1 vccd1 _2217_/B sky130_fd_sc_hd__and3_1
X_2147_ _2145_/X _2146_/Y _1975_/X vssd1 vssd1 vccd1 vccd1 _2148_/B sky130_fd_sc_hd__o21a_1
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
+ _4718_/Q _2618_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA_fanout173_A _4121_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2078_ _2077_/Y _2034_/C _4436_/Q vssd1 vssd1 vccd1 vccd1 _2079_/B sky130_fd_sc_hd__mux2_1
XANTENNA__3877__A _3877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_4112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_2710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4719_ _4719_/CLK _4719_/D fanout255/X vssd1 vssd1 vccd1 vccd1 _4719_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5019__D _5019_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_4052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1844__B _2608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_2672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_2490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_2343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_4001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_4045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
+ _4761_/Q _2715_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_29_3137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_2160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_3602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_2013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_2182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_3613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_3646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3050_ _4974_/Q _4973_/Q vssd1 vssd1 vccd1 vccd1 _3050_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_20_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2585__B _2585_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2001_ _4397_/Q _2001_/B vssd1 vssd1 vccd1 vccd1 _4397_/D sky130_fd_sc_hd__xnor2_1
XFILLER_20_2956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5063_/A fanout244/X vssd1 vssd1 vccd1 vccd1 _5079_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_20_2989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3697__A _4071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3952_ _4383_/Q vssd1 vssd1 vccd1 vccd1 _4384_/D sky130_fd_sc_hd__inv_2
XFILLER_18_2841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2903_ _2901_/X _2902_/Y _2143_/A vssd1 vssd1 vccd1 vccd1 _2904_/B sky130_fd_sc_hd__o21a_1
XFILLER_17_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3883_ _3883_/A _3883_/B vssd1 vssd1 vccd1 vccd1 _3884_/S sky130_fd_sc_hd__nand2_1
XFILLER_31_3753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2834_ _4857_/Q _2829_/C _2830_/B vssd1 vssd1 vccd1 vccd1 _2835_/B sky130_fd_sc_hd__a21bo_1
XFILLER_31_3775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3630__82 _3654__84/A vssd1 vssd1 vccd1 vccd1 _3630__82/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2765_ _4808_/Q _2765_/B vssd1 vssd1 vccd1 vccd1 _4808_/D sky130_fd_sc_hd__xnor2_1
XFILLER_12_2473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4504_ _4063_/B _4504_/D _3275_/Y vssd1 vssd1 vccd1 vccd1 _4504_/Q sky130_fd_sc_hd__dfrtp_1
X_1716_ _4943_/Q vssd1 vssd1 vccd1 vccd1 _4944_/D sky130_fd_sc_hd__inv_2
X_2696_ _4834_/D _4776_/Q _4774_/Q vssd1 vssd1 vccd1 vccd1 _2696_/X sky130_fd_sc_hd__and3_1
XFILLER_9_3721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4435_ _5033_/A _4435_/D fanout197/X vssd1 vssd1 vccd1 vccd1 _4435_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_3765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2479__C _4675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4379__CLK _4472_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4366_ _4366_/CLK _4366_/D fanout200/X vssd1 vssd1 vccd1 vccd1 _4366_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_3568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_2834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_4054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_A
+ _4485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_4065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2776__A _3114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3317_ _3891_/A _3889_/A vssd1 vssd1 vccd1 vccd1 _3317_/Y sky130_fd_sc_hd__xnor2_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_4087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4297_ _3877_/A _4297_/D _3781__122/Y vssd1 vssd1 vccd1 vccd1 _4297_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _3912_/A _3446_/B vssd1 vssd1 vccd1 vccd1 _3248_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_27_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_GATE_N
+ fanout128/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2655__A1 _4763_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf _4280_/Q _1847_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5004__CLK _3558_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3400__A _3414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3683__90_A _3683__90/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_2827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_2849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_2226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2016__A _4462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1855__A _4351_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_2609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3312__24_A _3366__32/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_3128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5062__A _5062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_2449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_3862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3310__A _3891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_2359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1765__A _1765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4521__CLK _4532_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2550_ _4713_/Q _4712_/Q _4711_/Q _2550_/D vssd1 vssd1 vccd1 vccd1 _2551_/D sky130_fd_sc_hd__and4_1
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2481_ _4669_/Q vssd1 vssd1 vccd1 vccd1 _2493_/A sky130_fd_sc_hd__inv_2
XFILLER_29_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4220_ _4794_/Q vssd1 vssd1 vccd1 vccd1 _4793_/D sky130_fd_sc_hd__clkinv_2
XFILLER_29_2277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_3949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4671__CLK _4709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_2040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4151_ _4690_/Q vssd1 vssd1 vccd1 vccd1 _4691_/D sky130_fd_sc_hd__inv_2
XFILLER_29_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3102_ _3056_/C _3098_/Y _1791_/X vssd1 vssd1 vccd1 vccd1 _3103_/B sky130_fd_sc_hd__o21ai_1
XFILLER_20_3443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4494__RESET_B fanout202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4082_ _4594_/Q vssd1 vssd1 vccd1 vccd1 _4593_/D sky130_fd_sc_hd__inv_2
XFILLER_20_2731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3033_ _4958_/Q _3033_/B vssd1 vssd1 vccd1 vccd1 _4958_/D sky130_fd_sc_hd__xnor2_1
XFILLER_3_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4984_ _4997_/CLK _4984_/D fanout232/X vssd1 vssd1 vccd1 vccd1 _4984_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3220__A _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3935_ _3935_/A _3935_/B vssd1 vssd1 vccd1 vccd1 _4378_/D sky130_fd_sc_hd__xnor2_1
XFILLER_32_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout136_A _3375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3866_ _4374_/Q vssd1 vssd1 vccd1 vccd1 _3916_/A sky130_fd_sc_hd__buf_12
XANTENNA__3874__B _3908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2817_ _4865_/Q _4864_/Q _2817_/C vssd1 vssd1 vccd1 vccd1 _2818_/D sky130_fd_sc_hd__and3_1
XFILLER_14_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3797_ _4295_/Q vssd1 vssd1 vccd1 vccd1 _4294_/D sky130_fd_sc_hd__inv_2
XFILLER_14_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_2281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2748_ _4804_/Q _2748_/B vssd1 vssd1 vccd1 vccd1 _2748_/X sky130_fd_sc_hd__and2b_1
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_TE_B
+ _2199_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_4055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2679_ _4770_/Q _4769_/Q _2647_/D _2676_/B vssd1 vssd1 vccd1 vccd1 _2680_/B sky130_fd_sc_hd__a31o_1
X_4418_ _3228_/Y _4418_/D _3752_/Y vssd1 vssd1 vccd1 vccd1 _4418_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_3354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3770__109_A _3770__109/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4349_ input25/X _4349_/D fanout195/X vssd1 vssd1 vccd1 vccd1 _4349_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_2894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_2675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
+ _4522_/Q _2269_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_21_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_2602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_3369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_2012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4544__CLK _2807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5057__A _5057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_3107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4694__CLK _4920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_2428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_A
+ _4618_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3522__48 _3523__49/A vssd1 vssd1 vccd1 vccd1 _4936_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3305__A _3309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_2235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_2016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_2279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__1628_ clkbuf_0__1628_/X vssd1 vssd1 vccd1 vccd1 _3159__59/A sky130_fd_sc_hd__clkbuf_16
XFILLER_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1981_ _4391_/Q _1981_/B vssd1 vssd1 vccd1 vccd1 _4391_/D sky130_fd_sc_hd__xnor2_1
XFILLER_14_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3720_ _3721_/A vssd1 vssd1 vccd1 vccd1 _3720_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_2281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_3881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
+ _4580_/Q _2367_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_3651_ _4195_/A vssd1 vssd1 vccd1 vccd1 _3651_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_2189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2602_ _4745_/D _4719_/Q vssd1 vssd1 vccd1 vccd1 _2603_/B sky130_fd_sc_hd__xnor2_1
X_3582_ _3587_/A vssd1 vssd1 vccd1 vccd1 _3582_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2533_ _4681_/Q _2533_/B vssd1 vssd1 vccd1 vccd1 _4681_/D sky130_fd_sc_hd__xnor2_1
XFILLER_9_2102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_2124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4675__RESET_B fanout253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2464_ _3875_/D _3941_/B _2464_/C vssd1 vssd1 vccd1 vccd1 _2464_/Y sky130_fd_sc_hd__nand3_1
X_4203_ _4759_/Q vssd1 vssd1 vccd1 vccd1 _4760_/D sky130_fd_sc_hd__inv_2
XFILLER_6_3779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2395_ _4615_/Q _2395_/B vssd1 vssd1 vccd1 vccd1 _2395_/X sky130_fd_sc_hd__and2b_1
XANTENNA__3215__A _3738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4134_ _4658_/Q _4134_/B vssd1 vssd1 vccd1 vccd1 _4659_/D sky130_fd_sc_hd__xnor2_1
XFILLER_4_3481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4417__CLK _3914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4065_ _4065_/A _4066_/B vssd1 vssd1 vccd1 vccd1 _4563_/D sky130_fd_sc_hd__xor2_1
XFILLER_20_2561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3016_ _4954_/Q _3016_/B vssd1 vssd1 vccd1 vccd1 _3016_/X sky130_fd_sc_hd__and2b_1
XFILLER_3_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout253_A fanout256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4567__CLK _2294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4967_ _4247_/Y _4967_/D _3536_/Y vssd1 vssd1 vccd1 vccd1 _4967_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3885__A _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_2490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3918_ _4376_/Q vssd1 vssd1 vccd1 vccd1 _3924_/A sky130_fd_sc_hd__buf_8
XFILLER_31_4081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_3921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4898_ _4901_/CLK _4898_/D fanout232/X vssd1 vssd1 vccd1 vccd1 _4898_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3849_ _4364_/Q vssd1 vssd1 vccd1 vccd1 _3885_/A sky130_fd_sc_hd__buf_8
XFILLER_20_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_2726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2948__B _4905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout120 _5062_/A vssd1 vssd1 vccd1 vccd1 fanout120/X sky130_fd_sc_hd__clkbuf_2
Xfanout131 _5043_/A vssd1 vssd1 vccd1 vccd1 _4590_/CLK sky130_fd_sc_hd__buf_2
Xfanout142 _2285_/Y vssd1 vssd1 vccd1 vccd1 _4532_/CLK sky130_fd_sc_hd__buf_2
XFILLER_1_3109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout153 _3930_/X vssd1 vssd1 vccd1 vccd1 _4920_/CLK sky130_fd_sc_hd__buf_8
XFILLER_21_3048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout164 _2807_/A vssd1 vssd1 vccd1 vccd1 _4943_/CLK sky130_fd_sc_hd__buf_4
XFILLER_21_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout175 _1765_/A vssd1 vssd1 vccd1 vccd1 _4248_/A sky130_fd_sc_hd__buf_6
Xfanout186 fanout196/X vssd1 vssd1 vccd1 vccd1 fanout186/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout197 fanout198/X vssd1 vssd1 vccd1 vccd1 fanout197/X sky130_fd_sc_hd__clkbuf_4
XFILLER_25_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3160__60_A _3169__65/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _4363_/CLK fanout191/X vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_10_3442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_2741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2204__A _2858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3643_/A fanout243/X vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__dlrtn_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1762__B _1763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_3869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3035__A _5020_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2180_ _2133_/C _2176_/Y _2173_/X vssd1 vssd1 vccd1 vccd1 _2181_/B sky130_fd_sc_hd__o21ai_1
XFILLER_26_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2874__A _4927_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_2986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4821_ _2809_/A1 _4821_/D _3456_/Y vssd1 vssd1 vccd1 vccd1 _4821_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__3017__A1 _2988_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_2630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_3217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4752_ _4752_/CLK _4752_/D fanout223/X vssd1 vssd1 vccd1 vccd1 _4752_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1964_ _4390_/Q vssd1 vssd1 vccd1 vccd1 _1977_/A sky130_fd_sc_hd__inv_2
XFILLER_15_2674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3703_ _4071_/A vssd1 vssd1 vccd1 vccd1 _3703_/Y sky130_fd_sc_hd__inv_2
X_4683_ _4717_/CLK _4683_/D fanout255/X vssd1 vssd1 vccd1 vccd1 _4683_/Q sky130_fd_sc_hd__dfrtp_2
X_1895_ _4321_/Q _4320_/Q _1898_/A vssd1 vssd1 vccd1 vccd1 _1895_/Y sky130_fd_sc_hd__nor3_1
XFILLER_11_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4856__RESET_B fanout226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3634_ _3642_/A vssd1 vssd1 vccd1 vccd1 _3634_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2114__A _3710_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3565_ _3571_/A vssd1 vssd1 vccd1 vccd1 _3565_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_4003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2516_ _4676_/Q _2516_/B vssd1 vssd1 vccd1 vccd1 _4676_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3496_ _3498_/A vssd1 vssd1 vccd1 vccd1 _3496_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_3302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_4058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2447_ _4649_/D _4650_/Q vssd1 vssd1 vccd1 vccd1 _2448_/B sky130_fd_sc_hd__and2b_1
XFILLER_22_2601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_2770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2378_ _4612_/Q vssd1 vssd1 vccd1 vccd1 _2390_/A sky130_fd_sc_hd__inv_2
XFILLER_25_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4117_ _4643_/Q vssd1 vssd1 vccd1 vccd1 _4644_/D sky130_fd_sc_hd__inv_2
XFILLER_22_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5097_ _5097_/A vssd1 vssd1 vccd1 vccd1 _5097_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4048_ _4542_/Q vssd1 vssd1 vccd1 vccd1 _4543_/D sky130_fd_sc_hd__inv_2
XFILLER_33_4110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3156__56_A _3159__59/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_2741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_3751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2519__B1 _2518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4526__RESET_B fanout202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_3257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_2409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_3064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4732__CLK _4981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input29_A phi1b_dig_Q[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5070__A _5070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3302__B _3444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4882__CLK _5013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2758__B1 _2687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_2825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2222__A2 _2218_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1680_ _4908_/Q vssd1 vssd1 vccd1 vccd1 _4909_/D sky130_fd_sc_hd__inv_2
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3659_/A fanout240/X vssd1 vssd1 vccd1 vccd1 _5076_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_8_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4267__RESET_B _5056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.ro_block_I.ro_pol_eve.tribuf.t_buf _1933_/A _1773_/Y vssd1 vssd1 vccd1 vccd1 _5089_/A
+ sky130_fd_sc_hd__ebufn_8
X_3350_ _3947_/A _3438_/B vssd1 vssd1 vccd1 vccd1 _3350_/Y sky130_fd_sc_hd__xnor2_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2930__B1 _2858_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2301_ _4574_/Q _4573_/Q vssd1 vssd1 vccd1 vccd1 _2301_/Y sky130_fd_sc_hd__xnor2_2
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _3287_/A vssd1 vssd1 vccd1 vccd1 _3281_/Y sky130_fd_sc_hd__inv_2
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ input32/X _5020_/D fanout207/X vssd1 vssd1 vccd1 vccd1 _5021_/D sky130_fd_sc_hd__dfrtp_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2232_ _4524_/Q _2208_/D _2225_/B vssd1 vssd1 vccd1 vccd1 _2233_/B sky130_fd_sc_hd__a21bo_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2289__A2 _3941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2163_ _4489_/Q _2163_/B vssd1 vssd1 vccd1 vccd1 _2163_/X sky130_fd_sc_hd__and2b_1
XFILLER_1_3473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_4127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2094_ _4442_/Q _4441_/Q vssd1 vssd1 vccd1 vccd1 _2094_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__3212__B _3847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0_clk_master clkbuf_0_clk_master/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_clk_master/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_34_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_2736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_3773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1948__A _3888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4804_ _4809_/CLK _4804_/D fanout254/X vssd1 vssd1 vccd1 vccd1 _4804_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2996_ _2996_/A _3042_/B _3042_/C vssd1 vssd1 vccd1 vccd1 _2997_/B sky130_fd_sc_hd__and3_1
XFILLER_33_2059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2749__B1 _2687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_GATE_N _4363_/CLK
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4735_ _3411_/Y _4735_/D _3661_/Y vssd1 vssd1 vccd1 vccd1 _4735_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4605__CLK _4852_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1947_ _3870_/Y _1947_/B vssd1 vssd1 vccd1 vccd1 _5092_/A sky130_fd_sc_hd__xnor2_4
XFILLER_15_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4666_ _2470_/A1 _4666_/D _3373__35/Y vssd1 vssd1 vccd1 vccd1 _4666_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_TE_B
+ _3115_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1878_ _4313_/Q _1878_/B vssd1 vssd1 vccd1 vccd1 _4313_/D sky130_fd_sc_hd__xnor2_1
XFILLER_11_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3882__B _3888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3617_ _5062_/A vssd1 vssd1 vccd1 vccd1 _4256_/A sky130_fd_sc_hd__buf_6
X_4597_ _3939_/Y _4597_/D _3328_/Y vssd1 vssd1 vccd1 vccd1 _4597_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_2821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4755__CLK _2631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_4041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3548_ _3550_/A vssd1 vssd1 vccd1 vccd1 _3548_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_3599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_2865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_4096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3479_ _3905_/A _3913_/A vssd1 vssd1 vccd1 vccd1 _3479_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_22_3121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3403__A _4004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_2497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2019__A _4462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_2224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_2869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4285__CLK _4288_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4707__RESET_B fanout247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4360__RESET_B fanout198/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5065__A _5065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_A
+ _4799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_3098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_2228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_3793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_2302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_2335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2850_ _4860_/Q _2850_/B vssd1 vssd1 vccd1 vccd1 _4860_/D sky130_fd_sc_hd__xnor2_1
XFILLER_31_3946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1801_ _2858_/A vssd1 vssd1 vccd1 vccd1 _3109_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_12_3345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2781_ _4822_/Q _4821_/Q vssd1 vssd1 vccd1 vccd1 _2781_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_12_3389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_2081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4520_ _4532_/CLK _4520_/D fanout211/X vssd1 vssd1 vccd1 vccd1 _4520_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__4778__CLK _4247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1732_ _4975_/Q vssd1 vssd1 vccd1 vccd1 _4976_/D sky130_fd_sc_hd__inv_2
XFILLER_12_2677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1954__A1 _3865_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2599__A _4745_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4451_ _2286_/B _4451_/D _3247_/Y vssd1 vssd1 vccd1 vccd1 _4451_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_3914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1663_ _4877_/Q vssd1 vssd1 vccd1 vccd1 _4876_/D sky130_fd_sc_hd__inv_2
XFILLER_9_3925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3402_ _3414_/A vssd1 vssd1 vccd1 vccd1 _3402_/Y sky130_fd_sc_hd__inv_2
X_4382_ _3208_/Y _4382_/D _3762__102/Y vssd1 vssd1 vccd1 vccd1 _4382_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_4131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_4142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2903__B1 _2143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _3925_/A _3442_/B vssd1 vssd1 vccd1 vccd1 _3333_/Y sky130_fd_sc_hd__xnor2_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _4247_/Y _5003_/D _3557_/Y vssd1 vssd1 vccd1 vccd1 _5003_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_2762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2215_ _4520_/Q _2219_/B _2221_/A vssd1 vssd1 vccd1 vccd1 _2262_/C sky130_fd_sc_hd__o21ai_1
XFILLER_22_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3223__A _3233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2146_ _4484_/Q _2146_/B vssd1 vssd1 vccd1 vccd1 _2146_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_2889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2077_ _2077_/A vssd1 vssd1 vccd1 vccd1 _2077_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout166_A _3869_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3877__B _4131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2979_ _4248_/A _2975_/X _2978_/X vssd1 vssd1 vccd1 vccd1 _2980_/B sky130_fd_sc_hd__a21oi_4
XFILLER_11_2110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_3890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4718_ _4718_/CLK _4718_/D fanout242/X vssd1 vssd1 vccd1 vccd1 _4718_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_33_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_4114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_2165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4649_ input28/X _4649_/D fanout208/X vssd1 vssd1 vccd1 vccd1 _4650_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_2_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2302__A _4648_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[0\].w1.ro_block_I.ro_pol.tribuf.t_buf _2113_/X _1958_/Y vssd1
+ vssd1 vccd1 vccd1 _5088_/A sky130_fd_sc_hd__ebufn_8
XFILLER_8_2756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_2767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_2322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_4057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4959__RESET_B fanout212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_2319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_2010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_2508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4920__CLK _4920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_2098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_2964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_3149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3138__B1 _3941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3308__A _3895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_3822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4300__CLK _3914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_3658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_3669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3043__A _4961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2000_ _2061_/A _2000_/B vssd1 vssd1 vccd1 vccd1 _2001_/B sky130_fd_sc_hd__nand2_1
XFILLER_7_1598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_2968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3951_ _4384_/Q vssd1 vssd1 vccd1 vccd1 _4383_/D sky130_fd_sc_hd__inv_2
XFILLER_18_3565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2902_ _4892_/Q _2902_/B vssd1 vssd1 vccd1 vccd1 _2902_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3882_ _3882_/A _3888_/A vssd1 vssd1 vccd1 vccd1 _3882_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_14_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4282__RESET_B fanout199/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2833_ _2922_/A vssd1 vssd1 vccd1 vccd1 _2916_/A sky130_fd_sc_hd__buf_4
XFILLER_30_2018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_3787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2764_ _2718_/C _2760_/Y _2687_/X vssd1 vssd1 vccd1 vccd1 _2765_/B sky130_fd_sc_hd__o21ai_1
XFILLER_30_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4503_ _3274_/Y _4503_/D _3729_/Y vssd1 vssd1 vccd1 vccd1 _4503_/Q sky130_fd_sc_hd__dfrtp_1
X_1715_ _4944_/Q vssd1 vssd1 vccd1 vccd1 _4943_/D sky130_fd_sc_hd__inv_2
X_2695_ _4772_/Q _2695_/B vssd1 vssd1 vccd1 vccd1 _4772_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__3218__A _3947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3784__125 _3784__125/A vssd1 vssd1 vccd1 vccd1 _3784__125/Y sky130_fd_sc_hd__inv_2
XFILLER_9_3733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2122__A _4007_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4434_ _5033_/A _4434_/D fanout197/X vssd1 vssd1 vccd1 vccd1 _4434_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_29_3694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_3788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4365_ _4472_/CLK _4365_/D fanout200/X vssd1 vssd1 vccd1 vccd1 _4365_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_4033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _3931_/A _4296_/D _3156__56/Y vssd1 vssd1 vccd1 vccd1 _4296_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _3255_/A vssd1 vssd1 vccd1 vccd1 _3247_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_2631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_2581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3178_ _3912_/A _3446_/B vssd1 vssd1 vccd1 vccd1 _3178_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__2655__A2 _2659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3888__A _3888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2129_ _4477_/Q _4476_/Q vssd1 vssd1 vccd1 vccd1 _2129_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_TE_B
+ _2711_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4943__CLK _4943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3099__S _4994_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_2385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
+ _4892_/Q _2955_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_30_2596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3128__A _3128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4323__CLK _4324_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[6\].w1.ro_block_I.ro_pol.tribuf.t_buf _3134_/X _2983_/Y vssd1
+ vssd1 vccd1 vccd1 _5088_/A sky130_fd_sc_hd__ebufn_8
XANTENNA_input11_A comp_high_Q[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3310__B _3889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_4130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_3749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout157/X fanout203/X vssd1 vssd1 vccd1 vccd1 _5082_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2207__A _4527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_3473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1765__B _4248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_2201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3038__A _5020_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2480_ _4674_/Q _4673_/Q _4672_/Q _2480_/D vssd1 vssd1 vccd1 vccd1 _2490_/C sky130_fd_sc_hd__and4_1
XFILLER_29_2234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4816__CLK _3451_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_2109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2877__A _3114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
+ _4950_/Q _3050_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_4150_ _4691_/Q vssd1 vssd1 vccd1 vccd1 _4690_/D sky130_fd_sc_hd__inv_2
XFILLER_20_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput90 _5087_/X vssd1 vssd1 vccd1 vccd1 fb1_Q[7] sky130_fd_sc_hd__buf_2
X_3101_ _4993_/Q _3101_/B vssd1 vssd1 vccd1 vccd1 _4993_/D sky130_fd_sc_hd__xnor2_1
X_4081_ _4591_/Q vssd1 vssd1 vccd1 vccd1 _4592_/D sky130_fd_sc_hd__inv_2
XFILLER_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3032_ _2986_/C _3028_/Y _1791_/X vssd1 vssd1 vccd1 vccd1 _3033_/B sky130_fd_sc_hd__o21ai_1
XFILLER_20_2743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3501__A _3519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4463__RESET_B fanout198/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4983_ _4997_/CLK _4983_/D fanout234/X vssd1 vssd1 vccd1 vccd1 _4983_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3220__B _3440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3934_ _3934_/A vssd1 vssd1 vccd1 vccd1 _3935_/A sky130_fd_sc_hd__buf_12
XFILLER_18_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_GATE_N
+ _5059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_3540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3865_ _3908_/A vssd1 vssd1 vccd1 vccd1 _3865_/Y sky130_fd_sc_hd__inv_6
XFILLER_14_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2816_ _4927_/D _4869_/Q _4867_/Q _4866_/Q vssd1 vssd1 vccd1 vccd1 _2817_/C sky130_fd_sc_hd__and4_1
XFILLER_30_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3796_ _4292_/Q vssd1 vssd1 vccd1 vccd1 _4293_/D sky130_fd_sc_hd__inv_2
XFILLER_20_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_2861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout129_A _5061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_2883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2747_ _4805_/Q _2747_/B vssd1 vssd1 vccd1 vccd1 _2748_/B sky130_fd_sc_hd__nor2_1
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_A
+ _4948_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2573__A1 _4710_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2678_ _4767_/Q _2678_/B vssd1 vssd1 vccd1 vccd1 _4767_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__4496__CLK _4532_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4417_ _3914_/A _4417_/D _3227_/Y vssd1 vssd1 vccd1 vccd1 _4417_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_4078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_3585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_4089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4348_ input25/X _4348_/D fanout195/X vssd1 vssd1 vccd1 vccd1 _4349_/D sky130_fd_sc_hd__dfrtp_1
XANTENNA_input3_A comp_high_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4279_ _4281_/CLK _4279_/D fanout201/X vssd1 vssd1 vccd1 vccd1 _4279_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_2483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_2403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3411__A _3917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_GATE_N
+ fanout128/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3204__12 _3201__9/A vssd1 vssd1 vccd1 vccd1 _4378_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__1866__A _2143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_2046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_2923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4839__CLK input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_2967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2697__A _4834_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4989__CLK _4997_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_3753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_2175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_2028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4903__RESET_B fanout235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3749_/A fanout187/X vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3321__A _3891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3774__113 _3776__115/A vssd1 vssd1 vccd1 vccd1 _3774__113/Y sky130_fd_sc_hd__inv_2
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4369__CLK _3598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1980_ _2061_/A _1980_/B vssd1 vssd1 vccd1 vccd1 _1981_/B sky130_fd_sc_hd__nand2_1
XFILLER_19_2981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2252__B1 _2173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_2113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1776__A _4347_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_3893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3650_ _4195_/A vssd1 vssd1 vccd1 vccd1 _3650_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_2179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2601_ _4716_/Q _2601_/B vssd1 vssd1 vccd1 vccd1 _4716_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__2004__B1 _2003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3581_ _3587_/A vssd1 vssd1 vccd1 vccd1 _3581_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_3929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2532_ _2566_/A _2532_/B vssd1 vssd1 vccd1 vccd1 _2533_/B sky130_fd_sc_hd__nand2_1
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout120/X fanout250/X vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_6_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3364__30 _3366__32/A vssd1 vssd1 vccd1 vccd1 _4657_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_2053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_3725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2463_ _2631_/A _2631_/B _2461_/Y _2462_/Y vssd1 vssd1 vccd1 vccd1 _2463_/X sky130_fd_sc_hd__o22a_1
XFILLER_26_3664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_2930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4202_ _4760_/Q vssd1 vssd1 vccd1 vccd1 _4759_/D sky130_fd_sc_hd__inv_2
XFILLER_26_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2394_ _4616_/Q _2394_/B vssd1 vssd1 vccd1 vccd1 _2395_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_2985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4133_ _4659_/Q _4134_/B vssd1 vssd1 vccd1 vccd1 _4658_/D sky130_fd_sc_hd__xnor2_1
XFILLER_25_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_3493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4064_ _4064_/A _4064_/B vssd1 vssd1 vccd1 vccd1 _4066_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_2601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3015_ _4955_/Q _3015_/B vssd1 vssd1 vccd1 vccd1 _3016_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3231__A _3233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3682__89 _3683__90/A vssd1 vssd1 vccd1 vccd1 _3682__89/Y sky130_fd_sc_hd__inv_2
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4966_ _3535_/Y _4966_/D _3596_/Y vssd1 vssd1 vccd1 vccd1 _4966_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout246_A fanout247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_2322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3917_ _3917_/A _3917_/B vssd1 vssd1 vccd1 vccd1 _4374_/D sky130_fd_sc_hd__xnor2_1
XFILLER_33_2967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4897_ _4905_/CLK _4897_/D fanout231/X vssd1 vssd1 vccd1 vccd1 _4897_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3848_ _3848_/A _3848_/B vssd1 vssd1 vccd1 vccd1 _4360_/D sky130_fd_sc_hd__xnor2_1
XFILLER_20_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_3439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_4072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3406__A _3414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout110 _2969_/Y vssd1 vssd1 vccd1 vccd1 _5046_/A sky130_fd_sc_hd__buf_4
Xfanout121 _4841_/Q vssd1 vssd1 vccd1 vccd1 _5062_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_25_3185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout132 _2455_/Y vssd1 vssd1 vccd1 vccd1 _5043_/A sky130_fd_sc_hd__clkbuf_4
Xfanout143 fanout144/X vssd1 vssd1 vccd1 vccd1 _3684_/A sky130_fd_sc_hd__buf_2
Xfanout154 _4981_/CLK vssd1 vssd1 vccd1 vccd1 _3932_/A sky130_fd_sc_hd__buf_6
Xfanout165 _3869_/Y vssd1 vssd1 vccd1 vccd1 _2807_/A sky130_fd_sc_hd__buf_6
XFILLER_5_2556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout176 _4060_/Y vssd1 vssd1 vccd1 vccd1 _1765_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_5_2567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout187 fanout188/X vssd1 vssd1 vccd1 vccd1 fanout187/X sky130_fd_sc_hd__buf_2
XFILLER_1_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout198 fanout221/X vssd1 vssd1 vccd1 vccd1 fanout198/X sky130_fd_sc_hd__buf_4
XFILLER_21_2348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2964__B _4932_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_2280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3141__A _3930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_2200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_2709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_3101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2980__A _4188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_3719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
+ _4711_/Q _2610_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_32_2433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_3189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_2753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5017__CLK _3922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_2190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_2797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_2204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3035__B _4962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_3583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_3677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_2954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_3490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4820_ _3455_/Y _4820_/D _3638_/Y vssd1 vssd1 vccd1 vccd1 _4820_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _5030_/CLK _4751_/D fanout223/X vssd1 vssd1 vccd1 vccd1 _4751_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1963_ _4395_/Q _4394_/Q _4393_/Q _1963_/D vssd1 vssd1 vccd1 vccd1 _1973_/C sky130_fd_sc_hd__and4_1
XFILLER_14_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_3229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__0637_ clkbuf_0__0637_/X vssd1 vssd1 vccd1 vccd1 _3765__105/A sky130_fd_sc_hd__clkbuf_16
X_3702_ _4071_/A vssd1 vssd1 vccd1 vccd1 _3702_/Y sky130_fd_sc_hd__inv_2
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout128/X fanout246/X vssd1 vssd1 vccd1 vccd1 _5077_/A sky130_fd_sc_hd__dlrtn_1
X_4682_ _4718_/CLK _4682_/D fanout236/X vssd1 vssd1 vccd1 vccd1 _4682_/Q sky130_fd_sc_hd__dfstp_1
X_1894_ _4318_/Q _1894_/B vssd1 vssd1 vccd1 vccd1 _4318_/D sky130_fd_sc_hd__xnor2_1
XFILLER_11_2539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3633_ _3642_/A vssd1 vssd1 vccd1 vccd1 _3633_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2114__B _3737_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_3737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3564_ _4563_/Q _4564_/Q vssd1 vssd1 vccd1 vccd1 _3564_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_31_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2515_ _2566_/A _2515_/B vssd1 vssd1 vccd1 vccd1 _2516_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4896__RESET_B fanout232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3495_ _3934_/A _3933_/A vssd1 vssd1 vccd1 vccd1 _3495_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__3226__A _3912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
+ _4769_/Q _2707_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_2446_ _2446_/A vssd1 vssd1 vccd1 vccd1 _2448_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_3314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_3555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2377_ _4617_/Q _4616_/Q _4615_/Q _2377_/D vssd1 vssd1 vccd1 vccd1 _2387_/C sky130_fd_sc_hd__and4_1
XANTENNA_fanout196_A fanout221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4534__CLK _4248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4116_ _4644_/Q vssd1 vssd1 vccd1 vccd1 _4643_/D sky130_fd_sc_hd__inv_2
XFILLER_25_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5096_ _5096_/A vssd1 vssd1 vccd1 vccd1 _5096_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4047_ _4543_/Q vssd1 vssd1 vccd1 vccd1 _4542_/D sky130_fd_sc_hd__inv_2
XFILLER_0_2431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_4122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4684__CLK _4187_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3896__A _3896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_2406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4949_ _4962_/CLK _4949_/D fanout210/X vssd1 vssd1 vccd1 vccd1 _4949_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_2027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_2049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf_TE_B
+ _2785_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
+ _4426_/Q _2101_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_27_3269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_2618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_2281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_2239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_2041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_2962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4407__CLK _4063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_2594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_2012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4557__CLK input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2300_ _4572_/Q _4571_/Q vssd1 vssd1 vccd1 vccd1 _2300_/Y sky130_fd_sc_hd__xnor2_2
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3280_ _3917_/A _3444_/B vssd1 vssd1 vccd1 vccd1 _3280_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_27_3792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_2067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2231_ _4522_/Q _2231_/B vssd1 vssd1 vccd1 vccd1 _4522_/D sky130_fd_sc_hd__xnor2_1
XFILLER_1_4120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_2966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2162_ _4490_/Q _2162_/B vssd1 vssd1 vccd1 vccd1 _2163_/B sky130_fd_sc_hd__nor2_1
XFILLER_1_3441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2694__B1 _2687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_2988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_3485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2093_ _2608_/A _4440_/Q vssd1 vssd1 vccd1 vccd1 _4440_/D sky130_fd_sc_hd__xor2_1
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
+ _4484_/Q _2200_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_4_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_4139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_2773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4803_ _4803_/CLK _4803_/D fanout254/X vssd1 vssd1 vccd1 vccd1 _4803_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2995_ _4949_/Q _2999_/B _3001_/A vssd1 vssd1 vccd1 vccd1 _3042_/C sky130_fd_sc_hd__o21ai_1
X_4734_ _4943_/CLK _4734_/D _3410_/Y vssd1 vssd1 vccd1 vccd1 _4734_/Q sky130_fd_sc_hd__dfrtp_4
X_1946_ _3914_/A _2286_/B _1938_/Y _1941_/X _1945_/X vssd1 vssd1 vccd1 vccd1 _1947_/B
+ sky130_fd_sc_hd__a311oi_4
XFILLER_30_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_2336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1877_ _1868_/C _1876_/X _1823_/X vssd1 vssd1 vccd1 vccd1 _1878_/B sky130_fd_sc_hd__o21ai_1
X_4665_ _3372_/Y _4665_/D _3681__88/Y vssd1 vssd1 vccd1 vccd1 _4665_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_3501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3616_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3616_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout111_A _5063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4596_ _3327_/Y _4596_/D _3703_/Y vssd1 vssd1 vccd1 vccd1 _4596_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout209_A fanout220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3547_ _3946_/A _3945_/A vssd1 vssd1 vccd1 vccd1 _3547_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_6_4053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_3330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_2877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_3133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2429_ _2566_/A _2429_/B vssd1 vssd1 vccd1 vccd1 _2430_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_3385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_2421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_3177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3403__B _3491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5079_ _5079_/A vssd1 vssd1 vccd1 vccd1 _5079_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_3527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4250__A _4250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_2881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2912__A1 _4896_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_2025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2979__A1 _4248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_2314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_2347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1800_ _4278_/Q _1800_/B vssd1 vssd1 vccd1 vccd1 _1800_/X sky130_fd_sc_hd__and2b_1
XFILLER_12_3357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2780_ _4820_/Q _4819_/Q vssd1 vssd1 vccd1 vccd1 _2780_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_34_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1939__C1 _3845_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_2634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1731_ _4976_/Q vssd1 vssd1 vccd1 vccd1 _4975_/D sky130_fd_sc_hd__inv_2
XANTENNA__2600__B1 _2518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_2093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_3821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4488__RESET_B fanout201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4450_ _3246_/Y _4450_/D _3743_/Y vssd1 vssd1 vccd1 vccd1 _4450_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_3092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1662_ _4874_/Q vssd1 vssd1 vccd1 vccd1 _4875_/D sky130_fd_sc_hd__inv_2
XFILLER_32_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_3865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3401_ _4065_/A _3543_/B vssd1 vssd1 vccd1 vccd1 _3401_/Y sky130_fd_sc_hd__xnor2_1
X_4381_ _3845_/Y _4381_/D _3207__14/Y vssd1 vssd1 vccd1 vccd1 _4381_/Q sky130_fd_sc_hd__dfrtp_1
X_3332_ _3340_/A vssd1 vssd1 vccd1 vccd1 _3332_/Y sky130_fd_sc_hd__inv_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_TE_B
+ _2778_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _3885_/A _3886_/A vssd1 vssd1 vccd1 vccd1 _3263_/Y sky130_fd_sc_hd__xnor2_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2116__C1 _3898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3504__A _4249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5002_ _3556_/Y _5002_/D _3585_/Y vssd1 vssd1 vccd1 vccd1 _5002_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _4523_/Q _4522_/Q _4521_/Q _2225_/B vssd1 vssd1 vccd1 vccd1 _2219_/B sky130_fd_sc_hd__or4_2
X_3194_ _3470_/A vssd1 vssd1 vccd1 vccd1 _3194_/X sky130_fd_sc_hd__buf_1
XANTENNA__2667__B1 _2518_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_2774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2145_ _4485_/Q _4484_/Q _2145_/C vssd1 vssd1 vccd1 vccd1 _2145_/X sky130_fd_sc_hd__and3_1
XFILLER_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2076_ _4434_/Q _2076_/B vssd1 vssd1 vccd1 vccd1 _4434_/D sky130_fd_sc_hd__xnor2_1
XFILLER_1_2581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout159_A _4469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_3413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2978_ _4131_/C _2978_/B _2978_/C _2978_/D vssd1 vssd1 vccd1 vccd1 _2978_/X sky130_fd_sc_hd__and4b_1
XANTENNA__4722__CLK _5007_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3893__B _3895_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_2122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4717_ _4717_/CLK _4717_/D fanout255/X vssd1 vssd1 vccd1 vccd1 _4717_/Q sky130_fd_sc_hd__dfrtp_1
X_1929_ _1929_/A vssd1 vssd1 vccd1 vccd1 _1929_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4648_ input28/X _4648_/D fanout208/X vssd1 vssd1 vccd1 vccd1 _4649_/D sky130_fd_sc_hd__dfrtp_1
XANTENNA__3147__A1 _4188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4872__CLK _4247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_GATE_N _5056_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4579_ _4590_/CLK _4579_/D fanout227/X vssd1 vssd1 vccd1 vccd1 _4579_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_8_3469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3414__A _3414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3313__25 _3365__31/A vssd1 vssd1 vccd1 vccd1 _4566_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_1826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_2262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_2066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4928__RESET_B fanout214/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_3106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3308__B _3372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_3834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_3773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3324__A _3340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_2059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_4109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout144/X fanout215/X vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_3555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3950_ _4381_/Q vssd1 vssd1 vccd1 vccd1 _4382_/D sky130_fd_sc_hd__inv_2
XFILLER_18_2821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4745__CLK input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2901_ _4893_/Q _4892_/Q _2901_/C vssd1 vssd1 vccd1 vccd1 _2901_/X sky130_fd_sc_hd__and3_1
X_3881_ _4361_/Q _3881_/B vssd1 vssd1 vccd1 vccd1 _4362_/D sky130_fd_sc_hd__xnor2_1
XFILLER_17_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2832_ _2832_/A _2832_/B vssd1 vssd1 vccd1 vccd1 _4855_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__4669__RESET_B fanout242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_3165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__0630_ _3656_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0630_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_34_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_2442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4895__CLK _4901_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2763_ _4807_/Q _2763_/B vssd1 vssd1 vccd1 vccd1 _4807_/D sky130_fd_sc_hd__xnor2_1
X_4502_ _4063_/C _4502_/D _3273_/Y vssd1 vssd1 vccd1 vccd1 _4502_/Q sky130_fd_sc_hd__dfrtp_1
X_1714_ _4941_/Q vssd1 vssd1 vccd1 vccd1 _4942_/D sky130_fd_sc_hd__inv_2
X_2694_ _2646_/C _2690_/Y _2687_/X vssd1 vssd1 vccd1 vccd1 _2695_/B sky130_fd_sc_hd__o21ai_1
XFILLER_12_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3218__B _3438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3772__111_A _3776__115/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4433_ _5041_/A _4433_/D fanout197/X vssd1 vssd1 vccd1 vccd1 _4433_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_3745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_2950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4364_ _4364_/CLK _4364_/D fanout199/X vssd1 vssd1 vccd1 vccd1 _4364_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_2825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_A
+ _4613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_4045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3315_ _3891_/A _3889_/A vssd1 vssd1 vccd1 vccd1 _3315_/Y sky130_fd_sc_hd__xnor2_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4295_ _3941_/B _4295_/D _3782__123/Y vssd1 vssd1 vccd1 vccd1 _4295_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3234__A _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3246_ _3917_/A _3444_/B vssd1 vssd1 vccd1 vccd1 _3246_/Y sky130_fd_sc_hd__xnor2_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4275__CLK _4281_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3177_ _3913_/A vssd1 vssd1 vccd1 vccd1 _3446_/B sky130_fd_sc_hd__buf_12
XFILLER_26_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2128_ _4475_/Q _4474_/Q vssd1 vssd1 vccd1 vccd1 _2128_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__3888__B _3901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2792__B _4839_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4065__A _4065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2059_ _4429_/Q _2059_/B vssd1 vssd1 vccd1 vccd1 _4429_/D sky130_fd_sc_hd__xnor2_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_4091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_2829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_2397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_2542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3409__A _3925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2313__A _2996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3128__B _3128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_2460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4618__CLK _4626_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_2471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_2554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_2357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4768__CLK _4811_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_3121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_4142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2803__B1 _3914_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2207__B _4526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_3441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4762__RESET_B fanout245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3319__A _3891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2223__A _2327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3193__75_A _3193__75/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1765__C _4248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3038__B _4962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4298__CLK _2286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output72_A _5069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput80 _5077_/X vssd1 vssd1 vccd1 vccd1 fb1_I[5] sky130_fd_sc_hd__buf_2
Xoutput91 _5088_/X vssd1 vssd1 vccd1 vccd1 read_out_I[0] sky130_fd_sc_hd__buf_2
XFILLER_20_3401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3100_ _3109_/A _3100_/B vssd1 vssd1 vccd1 vccd1 _3101_/B sky130_fd_sc_hd__nand2_1
X_4080_ _4592_/Q vssd1 vssd1 vccd1 vccd1 _4591_/D sky130_fd_sc_hd__inv_2
XFILLER_23_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_3445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout158/X fanout205/X vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__dlrtn_1
X_3031_ _4957_/Q _3031_/B vssd1 vssd1 vccd1 vccd1 _4957_/D sky130_fd_sc_hd__xnor2_1
XFILLER_24_2891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_2755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_3341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4982_ _3551_/Y _4982_/D _3587_/Y vssd1 vssd1 vccd1 vccd1 _4982_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_RESET_B
+ fanout239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_2640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3933_ _3933_/A _3935_/B vssd1 vssd1 vccd1 vccd1 _4377_/D sky130_fd_sc_hd__xnor2_1
XFILLER_14_2515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3864_ _3905_/A _3913_/A vssd1 vssd1 vccd1 vccd1 _3908_/A sky130_fd_sc_hd__xnor2_4
XFILLER_18_1972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2815_ _4853_/Q _4852_/Q vssd1 vssd1 vccd1 vccd1 _2815_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_31_3585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3795_ _4293_/Q vssd1 vssd1 vccd1 vccd1 _4292_/D sky130_fd_sc_hd__inv_2
XANTENNA__3229__A _3233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2133__A _4493_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2746_ _4802_/Q _2746_/B vssd1 vssd1 vccd1 vccd1 _4802_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__2573__A2 _4709_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2677_ _2648_/D _2676_/X _2518_/X vssd1 vssd1 vccd1 vccd1 _2678_/B sky130_fd_sc_hd__o21ai_1
XFILLER_29_3470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4416_ _3226_/Y _4416_/D _3753_/Y vssd1 vssd1 vccd1 vccd1 _4416_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_3417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2787__B _4835_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_2852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_2863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4347_ input25/X _4347_/D fanout195/X vssd1 vssd1 vccd1 vccd1 _4348_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_8_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3576_/A fanout251/X vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__dlrtn_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4910__CLK _4187_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4278_ _4281_/CLK _4278_/D fanout201/X vssd1 vssd1 vccd1 vccd1 _4278_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3899__A _3899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3229_ _3233_/A vssd1 vssd1 vccd1 vccd1 _3229_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_2473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3411__B _3444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2308__A _4648_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_2459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_2361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4440__CLK _5033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4590__CLK _4590_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_3765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3321__B _3889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_2294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1776__B _4289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_2868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_2879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_3293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2600_ _2598_/X _2599_/Y _2518_/X vssd1 vssd1 vccd1 vccd1 _2601_/B sky130_fd_sc_hd__o21ai_1
XFILLER_31_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_2581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3580_ _3587_/A vssd1 vssd1 vccd1 vccd1 _3580_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2888__A _4931_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2531_ _4741_/D _4683_/Q vssd1 vssd1 vccd1 vccd1 _2532_/B sky130_fd_sc_hd__xnor2_1
XFILLER_13_1891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4933__CLK input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2462_ _3941_/B _3929_/A vssd1 vssd1 vccd1 vccd1 _2462_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_2065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_3737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4201_ _4757_/Q vssd1 vssd1 vccd1 vccd1 _4758_/D sky130_fd_sc_hd__clkinv_2
XFILLER_29_2087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2393_ _4613_/Q _2393_/B vssd1 vssd1 vccd1 vccd1 _4613_/D sky130_fd_sc_hd__xnor2_1
XFILLER_22_2806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4132_ _4005_/B _4131_/D _4131_/X vssd1 vssd1 vccd1 vccd1 _4134_/B sky130_fd_sc_hd__a21bo_1
XFILLER_26_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4063_ _4131_/A _4063_/B _4063_/C _4131_/C vssd1 vssd1 vccd1 vccd1 _4064_/B sky130_fd_sc_hd__or4_4
XFILLER_3_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_3275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3512__A _4001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3014_ _4952_/Q _3014_/B vssd1 vssd1 vccd1 vccd1 _4952_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4313__CLK _5040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3201__9 _3201__9/A vssd1 vssd1 vccd1 vccd1 _4372_/CLK sky130_fd_sc_hd__inv_2
X_4965_ _1700_/Y _4965_/D _3534_/Y vssd1 vssd1 vccd1 vccd1 _4965_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4613__RESET_B fanout231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_2913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_3901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3916_ _3916_/A vssd1 vssd1 vccd1 vccd1 _3917_/A sky130_fd_sc_hd__buf_12
XANTENNA_fanout141_A _2285_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4896_ _4901_/CLK _4896_/D fanout232/X vssd1 vssd1 vccd1 vccd1 _4896_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_3912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_2957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4463__CLK input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_2356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3847_ _3847_/A _3848_/B vssd1 vssd1 vccd1 vccd1 _4359_/D sky130_fd_sc_hd__xnor2_1
XFILLER_18_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_2209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_2670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2729_ _4797_/Q _2729_/B vssd1 vssd1 vccd1 vccd1 _4797_/D sky130_fd_sc_hd__xor2_1
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout119/X fanout248/X vssd1 vssd1 vccd1 vccd1 _5078_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_9_3361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout111 _5063_/A vssd1 vssd1 vccd1 vccd1 _5055_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_2671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout122 _4709_/CLK vssd1 vssd1 vccd1 vccd1 _4718_/CLK sky130_fd_sc_hd__buf_4
Xfanout133 _4623_/CLK vssd1 vssd1 vccd1 vccd1 _4626_/CLK sky130_fd_sc_hd__clkbuf_4
Xfanout144 _5059_/A vssd1 vssd1 vccd1 vccd1 fanout144/X sky130_fd_sc_hd__clkbuf_2
Xfanout155 _4981_/CLK vssd1 vssd1 vccd1 vccd1 _2468_/A sky130_fd_sc_hd__buf_2
Xfanout166 _3869_/Y vssd1 vssd1 vccd1 vccd1 _3931_/A sky130_fd_sc_hd__buf_8
XFILLER_25_2485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout177 _3857_/Y vssd1 vssd1 vccd1 vccd1 _3899_/A sky130_fd_sc_hd__buf_4
XFILLER_9_1992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout188 fanout196/X vssd1 vssd1 vccd1 vccd1 fanout188/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout199 fanout221/X vssd1 vssd1 vccd1 vccd1 fanout199/X sky130_fd_sc_hd__buf_4
XANTENNA__3422__A _3896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
+ _4811_/Q _2786_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__3141__B _4126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2482__A1 _4671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2980__B _2980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4806__CLK _4812_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4336__CLK _3914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3332__A _3340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_2966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_4012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4486__CLK _5042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1787__A _2143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_3809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4750_ _4750_/CLK _4750_/D fanout228/X vssd1 vssd1 vccd1 vccd1 _4750_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1962_ _4398_/Q _4397_/Q _4396_/Q _1962_/D vssd1 vssd1 vccd1 vccd1 _1963_/D sky130_fd_sc_hd__and4_1
XFILLER_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3701_ _4071_/A vssd1 vssd1 vccd1 vccd1 _3701_/Y sky130_fd_sc_hd__inv_2
X_4681_ _4719_/CLK _4681_/D fanout252/X vssd1 vssd1 vccd1 vccd1 _4681_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_30_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_2518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1893_ _1909_/A _1893_/B vssd1 vssd1 vccd1 vccd1 _1894_/B sky130_fd_sc_hd__nand2_1
XANTENNA__1984__B1 _1823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
+ _4854_/Q _2886_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA_wrapper_cell_loop\[6\].w1.ro_block_Q.ro_pol.tribuf.t_buf_TE_B _2981_/Y vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3632_ _3632_/A vssd1 vssd1 vccd1 vccd1 _3642_/A sky130_fd_sc_hd__buf_8
XFILLER_31_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3563_ _3571_/A vssd1 vssd1 vccd1 vccd1 _3563_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_4141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3507__A _3519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2514_ _4677_/Q _2479_/D _2507_/B vssd1 vssd1 vccd1 vccd1 _2515_/B sky130_fd_sc_hd__a21bo_1
XFILLER_6_3501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3494_ _3498_/A vssd1 vssd1 vccd1 vccd1 _3494_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_4016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf _4315_/Q _1918_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XANTENNA__3226__B _3446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2445_ _4650_/Q _4649_/D vssd1 vssd1 vccd1 vccd1 _2446_/A sky130_fd_sc_hd__and2b_1
XFILLER_29_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_3326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2376_ _4620_/Q _4619_/Q _4618_/Q _2376_/D vssd1 vssd1 vccd1 vccd1 _2377_/D sky130_fd_sc_hd__and4_1
XFILLER_25_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4115_ _4641_/Q vssd1 vssd1 vccd1 vccd1 _4642_/D sky130_fd_sc_hd__inv_2
XFILLER_20_3050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5095_ _5095_/A vssd1 vssd1 vccd1 vccd1 _5095_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4865__RESET_B fanout226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3242__A _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout189_A fanout196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4046_ _4540_/Q vssd1 vssd1 vccd1 vccd1 _4541_/D sky130_fd_sc_hd__inv_2
XFILLER_0_3177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4829__CLK _4943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_2393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_4134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4948_ _4962_/CLK _4948_/D fanout208/X vssd1 vssd1 vccd1 vccd1 _4948_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4979__CLK _4131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4879_ _3489_/Y _4879_/D _3622_/Y vssd1 vssd1 vccd1 vccd1 _4879_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_3753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__1628_ _3155_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__1628_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4359__CLK _4359_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4248__A _4248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2508__A_N _4675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2991__A _5020_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_2053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5079__A _5079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_2952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3327__A _4004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2231__A _4522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3185__70 _3189__72/A vssd1 vssd1 vccd1 vccd1 _3185__70/Y sky130_fd_sc_hd__inv_2
XFILLER_7_3843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_3624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2230_ _2327_/A _2230_/B vssd1 vssd1 vccd1 vccd1 _2231_/B sky130_fd_sc_hd__nand2_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2161_ _4487_/Q _2161_/B vssd1 vssd1 vccd1 vccd1 _4487_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__3062__A _4994_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4276__RESET_B fanout201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2092_ _4439_/Q _2092_/B vssd1 vssd1 vccd1 vccd1 _4439_/D sky130_fd_sc_hd__xor2_1
XFILLER_19_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_2680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _4359_/CLK fanout190/X vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__dlrtn_1
X_4802_ _4809_/CLK _4802_/D fanout254/X vssd1 vssd1 vccd1 vccd1 _4802_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2994_ _4952_/Q _4951_/Q _4950_/Q _3005_/B vssd1 vssd1 vccd1 vccd1 _2999_/B sky130_fd_sc_hd__or4_1
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4733_ _3409_/Y _4733_/D _3662_/Y vssd1 vssd1 vccd1 vccd1 _4733_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1945_ _1943_/X _2287_/A vssd1 vssd1 vccd1 vccd1 _1945_/X sky130_fd_sc_hd__and2b_1
XANTENNA__2125__B _2464_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_2315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_2495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4664_ _2470_/A1 _4664_/D _3371__34/Y vssd1 vssd1 vccd1 vccd1 _4664_/Q sky130_fd_sc_hd__dfrtp_1
X_1876_ _4314_/Q _1876_/B vssd1 vssd1 vccd1 vccd1 _1876_/X sky130_fd_sc_hd__and2b_1
XFILLER_11_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3615_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3615_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4595_ _4916_/CLK _4595_/D _3326_/Y vssd1 vssd1 vccd1 vccd1 _4595_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3237__A _4005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_A
+ _4895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2141__A _4487_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout104_A _3135_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3546_ _3550_/A vssd1 vssd1 vccd1 vccd1 _3546_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3477_ _3905_/A _3913_/A vssd1 vssd1 vccd1 vccd1 _3477_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_24_2709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1980__A _2061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2428_ _4652_/D _4626_/Q vssd1 vssd1 vccd1 vccd1 _2429_/B sky130_fd_sc_hd__xnor2_1
X_3191__73 _3193__75/A vssd1 vssd1 vccd1 vccd1 _4354_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_3145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_2580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4651__CLK input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_2444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2359_ _4588_/Q _2359_/B vssd1 vssd1 vccd1 vccd1 _4588_/D sky130_fd_sc_hd__xnor2_1
XFILLER_22_3189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_2538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_2488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5078_ _5078_/A vssd1 vssd1 vccd1 vccd1 _5078_/X sky130_fd_sc_hd__buf_2
XFILLER_2_1826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3471__43_A _3523__49/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4029_ _4509_/Q vssd1 vssd1 vccd1 vccd1 _4508_/D sky130_fd_sc_hd__inv_2
XANTENNA__5007__CLK _5007_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3700__A _4071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_2805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_3241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4007__S _4007_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4250__B _4250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3159__59 _3159__59/A vssd1 vssd1 vccd1 vccd1 _3159__59/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2051__A _2061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2912__A2 _4895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_2344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1890__A _1909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_3819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input34_A ud_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_3773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
+ _4615_/Q _2439_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_1_2048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3610__A _3616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_4048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_4059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_2359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_2771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1730_ _4973_/Q vssd1 vssd1 vccd1 vccd1 _4974_/D sky130_fd_sc_hd__inv_2
XFILLER_12_1901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_3800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1661_ _4875_/Q vssd1 vssd1 vccd1 vccd1 _4874_/D sky130_fd_sc_hd__inv_2
XFILLER_29_3833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3057__A _4992_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3400_ _3414_/A vssd1 vssd1 vccd1 vccd1 _3400_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4380_ _4380_/CLK _4380_/D fanout210/X vssd1 vssd1 vccd1 vccd1 _4380_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3331_ _3935_/A _3440_/B vssd1 vssd1 vccd1 vccd1 _3331_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4674__CLK _4709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5001_ _1700_/Y _5001_/D _3555_/Y vssd1 vssd1 vccd1 vccd1 _5001_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3504__B _4250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ _4526_/Q _4525_/Q _4524_/Q _2235_/B vssd1 vssd1 vccd1 vccd1 _2225_/B sky130_fd_sc_hd__or4_2
XANTENNA__2667__A1 _2658_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_2836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_2847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2144_ _4482_/Q _2144_/B vssd1 vssd1 vccd1 vccd1 _4482_/D sky130_fd_sc_hd__xor2_1
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2075_ _2035_/D _2074_/Y _2003_/X vssd1 vssd1 vccd1 vccd1 _2076_/B sky130_fd_sc_hd__o21ai_1
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3520__A _3916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_2593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3092__A1 _4992_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout136/X fanout238/X vssd1 vssd1 vccd1 vccd1 _5084_/A sky130_fd_sc_hd__dlrtn_1
X_2977_ _2977_/A _2977_/B vssd1 vssd1 vccd1 vccd1 _5098_/A sky130_fd_sc_hd__xor2_4
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
+ _4673_/Q _2541_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__1975__A _2858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_2281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4716_ _4717_/CLK _4716_/D fanout254/X vssd1 vssd1 vccd1 vccd1 _4716_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout221_A input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1928_ _1928_/A _1928_/B vssd1 vssd1 vccd1 vccd1 _1929_/A sky130_fd_sc_hd__or2_1
XFILLER_33_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4647_ input28/X _4647_/D fanout210/X vssd1 vssd1 vccd1 vccd1 _4648_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1859_ _4311_/Q vssd1 vssd1 vccd1 vccd1 _1871_/A sky130_fd_sc_hd__inv_2
XFILLER_28_4066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3147__A2 _3138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_4088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4578_ _5043_/A _4578_/D fanout228/X vssd1 vssd1 vccd1 vccd1 _4578_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__2355__B1 _2344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_2631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_3387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3529_ _3916_/A _3915_/A vssd1 vssd1 vccd1 vccd1 _3529_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_6_3150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_2697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_TE_B _1920_/Y vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_2302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_2379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3430__A _4189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_2900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xw0.ro_block_Q.ro_pol.tribuf.t_buf _1929_/X _1770_/Y vssd1 vssd1 vccd1 vccd1 _5090_/A
+ sky130_fd_sc_hd__ebufn_8
XFILLER_11_4081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_2406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2212__C _4527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5092__A _5092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3605__A _5062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3340__A _3340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2900_ _4890_/Q _2900_/B vssd1 vssd1 vccd1 vccd1 _4890_/D sky130_fd_sc_hd__xor2_1
XANTENNA__2226__A_N _4522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3880_ _4362_/Q _3881_/B vssd1 vssd1 vccd1 vccd1 _4361_/D sky130_fd_sc_hd__xnor2_1
X_2831_ _2829_/X _2830_/Y _2143_/A vssd1 vssd1 vccd1 vccd1 _2832_/B sky130_fd_sc_hd__o21a_1
XFILLER_31_3745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1795__A _2922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_2410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2762_ _2771_/A _2762_/B vssd1 vssd1 vccd1 vccd1 _2763_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4501_ _3272_/Y _4501_/D _3730_/Y vssd1 vssd1 vccd1 vccd1 _4501_/Q sky130_fd_sc_hd__dfrtp_1
X_1713_ _4942_/Q vssd1 vssd1 vccd1 vccd1 _4941_/D sky130_fd_sc_hd__inv_2
X_2693_ _4771_/Q _2693_/B vssd1 vssd1 vccd1 vccd1 _4771_/D sky130_fd_sc_hd__xnor2_1
XFILLER_12_2498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_3641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4432_ _5033_/A _4432_/D fanout197/X vssd1 vssd1 vccd1 vccd1 _4432_/Q sky130_fd_sc_hd__dfrtp_2
X_4363_ _4363_/CLK _4363_/D fanout200/X vssd1 vssd1 vccd1 vccd1 _4363_/Q sky130_fd_sc_hd__dfrtp_1
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
+ _4403_/Q _2032_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA__3515__A _3519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3684_/A fanout217/X vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__dlrtn_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4294_ _3932_/A _4294_/D _3154__118/Y vssd1 vssd1 vccd1 vccd1 _4294_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3234__B _3886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _3255_/A vssd1 vssd1 vccd1 vccd1 _3245_/Y sky130_fd_sc_hd__inv_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_2633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2127_ _3941_/B _2127_/B vssd1 vssd1 vccd1 vccd1 _5065_/A sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout171_A _3855_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3250__A _3903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2058_ _2061_/A _2058_/B vssd1 vssd1 vccd1 vccd1 _2059_/B sky130_fd_sc_hd__nand2_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3409__B _3442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4379__RESET_B fanout210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_2303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3144__B _3144_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__1642_ clkbuf_0__1642_/X vssd1 vssd1 vccd1 vccd1 _3366__32/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__4256__A _4256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2803__A1 _4064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3319__B _3889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3335__A _3917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput70 _5067_/X vssd1 vssd1 vccd1 vccd1 cos_out[3] sky130_fd_sc_hd__buf_2
Xoutput81 _5078_/X vssd1 vssd1 vccd1 vccd1 fb1_I[6] sky130_fd_sc_hd__buf_2
Xoutput92 _5089_/X vssd1 vssd1 vccd1 vccd1 read_out_I[1] sky130_fd_sc_hd__buf_2
XFILLER_20_3413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4712__CLK _4712_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3030_ _3030_/A _3030_/B vssd1 vssd1 vccd1 vccd1 _3031_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_3529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_2881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_2723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_4021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3707__92_A _3732__95/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4981_ _4981_/CLK _4981_/D _3550_/Y vssd1 vssd1 vccd1 vccd1 _4981_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_3807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_4098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4862__CLK _4865_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3932_ _3932_/A _3932_/B vssd1 vssd1 vccd1 vccd1 _3935_/B sky130_fd_sc_hd__nand2_4
XFILLER_17_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_2652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3863_ _4371_/Q vssd1 vssd1 vccd1 vccd1 _3913_/A sky130_fd_sc_hd__buf_6
XFILLER_20_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2814_ _4851_/Q _4850_/Q vssd1 vssd1 vccd1 vccd1 _2814_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_18_1984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3794_ _4290_/Q vssd1 vssd1 vccd1 vccd1 _4291_/D sky130_fd_sc_hd__inv_2
XFILLER_14_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2133__B _4492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2745_ _2771_/A _2745_/B vssd1 vssd1 vccd1 vccd1 _2746_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2676_ _4768_/Q _2676_/B vssd1 vssd1 vccd1 vccd1 _2676_/X sky130_fd_sc_hd__and2b_1
XANTENNA__4472__RESET_B fanout207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4415_ _2286_/B _4415_/D _3225_/Y vssd1 vssd1 vccd1 vccd1 _4415_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_3565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_3335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3245__A _3255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_2612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4346_ input25/X input9/X fanout195/X vssd1 vssd1 vccd1 vccd1 _4347_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_25_2623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_GATE_N
+ _3738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_A
+ _4395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4277_ _4281_/CLK _4277_/D fanout201/X vssd1 vssd1 vccd1 vccd1 _4277_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4392__CLK _4402_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3899__B _3914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3228_ _3903_/A _3420_/B vssd1 vssd1 vccd1 vccd1 _3228_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_GATE_N
+ _5063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_3339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_3604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5055_/A fanout244/X vssd1 vssd1 vccd1 vccd1 _5079_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_30_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3155__A _3777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_2133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2994__A _4952_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_3996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_2188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_3695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4983__RESET_B fanout234/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2234__A _4523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2530_ _4680_/Q _2530_/B vssd1 vssd1 vccd1 vccd1 _4680_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__2888__B _4905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_TE_B
+ _2029_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_2116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2461_ _2631_/A _3877_/A vssd1 vssd1 vccd1 vccd1 _2461_/Y sky130_fd_sc_hd__nand2_1
X_4200_ _4758_/Q vssd1 vssd1 vccd1 vccd1 _4757_/D sky130_fd_sc_hd__inv_2
XFILLER_6_3749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_4141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2392_ _2412_/A _2392_/B vssd1 vssd1 vccd1 vccd1 _2393_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4131_ _4131_/A _4131_/B _4131_/C _4131_/D vssd1 vssd1 vccd1 vccd1 _4131_/X sky130_fd_sc_hd__or4_1
XFILLER_20_3210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_3221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4062_ _4123_/B vssd1 vssd1 vccd1 vccd1 _4064_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3013_ _3030_/A _3013_/B vssd1 vssd1 vccd1 vccd1 _3014_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3512__B _4005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5018__RESET_B _3576_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2409__A _2412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4964_ _1760_/Y _4964_/D _3533_/Y vssd1 vssd1 vccd1 vccd1 _4964_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_3003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_3659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3915_ _3915_/A _3917_/B vssd1 vssd1 vccd1 vccd1 _4373_/D sky130_fd_sc_hd__xnor2_1
XFILLER_32_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4895_ _4901_/CLK _4895_/D fanout234/X vssd1 vssd1 vccd1 vccd1 _4895_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_14_3058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_4073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_3069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3846_ _3846_/A _3883_/B vssd1 vssd1 vccd1 vccd1 _3848_/B sky130_fd_sc_hd__nand2_2
XFILLER_31_3361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout134_A _2455_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_2368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3777_ _3777_/A vssd1 vssd1 vccd1 vccd1 _3777_/X sky130_fd_sc_hd__buf_1
XFILLER_10_1509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_2693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_2092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2728_ _2996_/A _2774_/B _2774_/C vssd1 vssd1 vccd1 vccd1 _2729_/B sky130_fd_sc_hd__and3_1
XFILLER_9_3351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2659_ _4763_/Q _2659_/B vssd1 vssd1 vccd1 vccd1 _2659_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_3384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_3226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout112 _3576_/A vssd1 vssd1 vccd1 vccd1 _5063_/A sky130_fd_sc_hd__buf_2
Xfanout123 _4719_/CLK vssd1 vssd1 vccd1 vccd1 _4717_/CLK sky130_fd_sc_hd__buf_2
X_4329_ _3168_/Y _4329_/D _3772__111/Y vssd1 vssd1 vccd1 vccd1 _4329_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout134 _2455_/Y vssd1 vssd1 vccd1 vccd1 _4623_/CLK sky130_fd_sc_hd__clkbuf_4
Xfanout145 _3696_/A vssd1 vssd1 vccd1 vccd1 _5059_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_2536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout156 _3922_/X vssd1 vssd1 vccd1 vccd1 _4981_/CLK sky130_fd_sc_hd__buf_8
Xfanout167 _3865_/Y vssd1 vssd1 vccd1 vccd1 _2286_/B sky130_fd_sc_hd__buf_6
XANTENNA__3703__A _4071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout178 _3857_/Y vssd1 vssd1 vccd1 vccd1 _2470_/A1 sky130_fd_sc_hd__buf_4
Xfanout189 fanout196/X vssd1 vssd1 vccd1 vccd1 fanout189/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3422__B _3904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2482__A2 _4670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4288__CLK _4288_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_4113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_3592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_3434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2989__A _4948_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1893__A _1909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
+ wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_2024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3613__A _3616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_2923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2890__C _4897_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1961_ _4400_/Q _4399_/Q _1961_/C vssd1 vssd1 vccd1 vccd1 _1962_/D sky130_fd_sc_hd__and3_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3700_ _4071_/A vssd1 vssd1 vccd1 vccd1 _3700_/Y sky130_fd_sc_hd__inv_2
X_4680_ _4719_/CLK _4680_/D fanout252/X vssd1 vssd1 vccd1 vccd1 _4680_/Q sky130_fd_sc_hd__dfrtp_1
X_1892_ _4319_/Q _1857_/D _1885_/B vssd1 vssd1 vccd1 vccd1 _1893_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__4900__CLK _4901_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1984__A1 _1973_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3631_ _5061_/A vssd1 vssd1 vccd1 vccd1 _3631_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__2899__A _2996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout180/X fanout185/X vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__dlrtn_1
X_3562_ _4127_/A _4129_/A vssd1 vssd1 vccd1 vccd1 _3562_/Y sky130_fd_sc_hd__xnor2_1
X_2513_ _4675_/Q _2513_/B vssd1 vssd1 vccd1 vccd1 _4675_/D sky130_fd_sc_hd__xnor2_1
X_3493_ _3946_/A _3945_/A vssd1 vssd1 vccd1 vccd1 _3493_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_6_3513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2444_ _4646_/Q _4645_/Q vssd1 vssd1 vccd1 vccd1 _2444_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_9_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_3557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_2773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2375_ _4622_/Q _4621_/Q _2375_/C vssd1 vssd1 vccd1 vccd1 _2376_/D sky130_fd_sc_hd__and3_1
XFILLER_6_2856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4114_ _4642_/Q vssd1 vssd1 vccd1 vccd1 _4641_/D sky130_fd_sc_hd__inv_2
XFILLER_9_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5094_ _5094_/A vssd1 vssd1 vccd1 vccd1 _5094_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3242__B _3440_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4045_ _4541_/Q vssd1 vssd1 vccd1 vccd1 _4540_/D sky130_fd_sc_hd__inv_2
XANTENNA__2139__A _4493_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_2361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_2372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_3109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_4_0_clk_master clkbuf_3_5_0_clk_master/A vssd1 vssd1 vccd1 vccd1 _5030_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__4430__CLK _5033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1978__A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4834__RESET_B fanout237/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4947_ _4962_/CLK _4947_/D fanout208/X vssd1 vssd1 vccd1 vccd1 _4947_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_3721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4580__CLK _4590_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_2154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4878_ _1765_/A _4878_/D _3488_/Y vssd1 vssd1 vccd1 vccd1 _4878_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_2799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_3765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3829_ _4343_/Q vssd1 vssd1 vccd1 vccd1 _4342_/D sky130_fd_sc_hd__inv_2
XFILLER_14_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2602__A _4745_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_3205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_3249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_2515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_3023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_2480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3433__A _3445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_2103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_2294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4248__B _4248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2991__B _4962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_2519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_2065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_2817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
+ _4985_/Q _3121_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_16_2997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3608__A _3616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2512__A _2566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3327__B _3491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2391__A1 _4614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3343__A _3361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_3669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_2957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2160_ _2178_/A _2160_/B vssd1 vssd1 vccd1 vccd1 _2161_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4453__CLK _3914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2091_ _3066_/A _2091_/B _2091_/C _2091_/D vssd1 vssd1 vccd1 vccd1 _2092_/B sky130_fd_sc_hd__and4_1
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_3429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4801_ _4809_/CLK _4801_/D fanout252/X vssd1 vssd1 vccd1 vccd1 _4801_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2993_ _4955_/Q _4954_/Q _4953_/Q _3015_/B vssd1 vssd1 vccd1 vccd1 _3005_/B sky130_fd_sc_hd__or4_2
XFILLER_30_3629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1944_ _3898_/B _2286_/B vssd1 vssd1 vccd1 vccd1 _2287_/A sky130_fd_sc_hd__nor2_1
X_4732_ _4981_/CLK _4732_/D _3408_/Y vssd1 vssd1 vccd1 vccd1 _4732_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_2474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_2939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4663_ _3370_/Y _4663_/D _3682__89/Y vssd1 vssd1 vccd1 vccd1 _4663_/Q sky130_fd_sc_hd__dfrtp_2
X_1875_ _4315_/Q _1875_/B vssd1 vssd1 vccd1 vccd1 _1876_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3518__A _3924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3614_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3614_/Y sky130_fd_sc_hd__inv_2
X_4594_ _3325_/Y _4594_/D _3704_/Y vssd1 vssd1 vccd1 vccd1 _4594_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_3525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_4000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3545_ _4001_/A _4005_/A vssd1 vssd1 vccd1 vccd1 _3545_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__2141__B _4486_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2427_ _4623_/Q _2427_/B vssd1 vssd1 vccd1 vccd1 _4623_/D sky130_fd_sc_hd__xnor2_1
XFILLER_9_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3253__A _3255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5048_/A fanout192/X vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_26_2592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2358_ _2412_/A _2358_/B vssd1 vssd1 vccd1 vccd1 _2359_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5077_ _5077_/A vssd1 vssd1 vccd1 vccd1 _5077_/X sky130_fd_sc_hd__buf_4
X_2289_ _3898_/B _3941_/B _3907_/A _3941_/A vssd1 vssd1 vccd1 vccd1 _2289_/X sky130_fd_sc_hd__a211o_1
XFILLER_6_1996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4028_ _4506_/Q vssd1 vssd1 vccd1 vccd1 _4507_/D sky130_fd_sc_hd__inv_2
XFILLER_0_2241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3643_/A fanout243/X vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_17_3974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3428__A _3445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4326__CLK _4063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_2861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_2301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4476__CLK _1952_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_2367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_2389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input27_A phi1b_dig_Q[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_4141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2507__A _4676_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_3451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_3484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1939__A1 _3892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_2647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3338__A _3340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1660_ _4872_/Q vssd1 vssd1 vccd1 vccd1 _4873_/D sky130_fd_sc_hd__inv_2
XANTENNA__3057__B _4991_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4819__CLK _1765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3330_ _3340_/A vssd1 vssd1 vccd1 vccd1 _3330_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_4134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2896__B _4897_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3261_ _3885_/A _3886_/A vssd1 vssd1 vccd1 vccd1 _3261_/Y sky130_fd_sc_hd__xnor2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3073__A _3109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5000_ _1760_/Y _5000_/D _3554_/Y vssd1 vssd1 vccd1 vccd1 _5000_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _4529_/Q _4528_/Q _4527_/Q _2248_/A vssd1 vssd1 vccd1 vccd1 _2235_/B sky130_fd_sc_hd__or4_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4969__CLK _4187_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_2743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2143_ _2143_/A _2191_/B _2191_/C vssd1 vssd1 vccd1 vccd1 _2144_/B sky130_fd_sc_hd__and3_1
XFILLER_23_2798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4497__RESET_B fanout210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2074_ _4436_/Q _4435_/Q _2077_/A vssd1 vssd1 vccd1 vccd1 _2074_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__3520__B _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2417__A _2922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_4127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2976_ _4131_/C _2972_/X _2975_/X _4126_/A vssd1 vssd1 vccd1 vccd1 _2977_/B sky130_fd_sc_hd__a2bb2o_2
XFILLER_30_3437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4715_ _4717_/CLK _4715_/D fanout254/X vssd1 vssd1 vccd1 vccd1 _4715_/Q sky130_fd_sc_hd__dfrtp_1
X_1927_ _4348_/D _4349_/Q vssd1 vssd1 vccd1 vccd1 _1928_/B sky130_fd_sc_hd__and2b_1
XFILLER_28_4001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3248__A _3912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_3893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_2758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2152__A _4487_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_4106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1858_ _4316_/Q _4315_/Q _4314_/Q _1858_/D vssd1 vssd1 vccd1 vccd1 _1868_/C sky130_fd_sc_hd__and4_1
XANTENNA_fanout214_A fanout219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4646_ _3362_/Y _4646_/D _3684_/Y vssd1 vssd1 vccd1 vccd1 _4646_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_4117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_3311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4499__CLK _4126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_4078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4577_ _4590_/CLK _4577_/D fanout226/X vssd1 vssd1 vccd1 vccd1 _4577_/Q sky130_fd_sc_hd__dfrtp_2
X_1789_ _4277_/Q _4276_/Q _1789_/C vssd1 vssd1 vccd1 vccd1 _1789_/X sky130_fd_sc_hd__and3_1
XFILLER_8_2715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_2643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_2529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3459_ _3946_/A _3945_/A vssd1 vssd1 vccd1 vccd1 _3459_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_28_1964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_2314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3711__A _5058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_4005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3659_/A fanout240/X vssd1 vssd1 vccd1 vccd1 _5076_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_22_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3430__B _4190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2327__A _2327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_2035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2062__A _4430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2997__A _4947_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_A
+ _4709_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf _4277_/Q _1850_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XFILLER_27_2153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_2247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4937__RESET_B fanout214/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_2938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3621__A _4256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_3513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2806__C1 _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_GATE_N _4363_/CLK
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_3568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_2845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2830_ _4856_/Q _2830_/B vssd1 vssd1 vccd1 vccd1 _2830_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
+ _4804_/Q _2778_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_31_3757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2761_ _2760_/Y _2718_/C _4808_/Q vssd1 vssd1 vccd1 vccd1 _2762_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4641__CLK _4852_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_3189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1712_ _4939_/Q vssd1 vssd1 vccd1 vccd1 _4940_/D sky130_fd_sc_hd__inv_2
X_4500_ _2809_/A1 _4500_/D _3271_/Y vssd1 vssd1 vccd1 vccd1 _4500_/Q sky130_fd_sc_hd__dfrtp_1
X_2692_ _2771_/A _2692_/B vssd1 vssd1 vccd1 vccd1 _2693_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_3631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4431_ _5033_/A _4431_/D fanout197/X vssd1 vssd1 vccd1 vccd1 _4431_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_12_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2700__A _4834_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4791__CLK _4981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4362_ _4362_/CLK _4362_/D fanout202/X vssd1 vssd1 vccd1 vccd1 _4362_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_29_3697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_4014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ _3929_/A _4293_/D _3783__124/Y vssd1 vssd1 vccd1 vccd1 _4293_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_3471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4678__RESET_B fanout255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _3925_/A _3442_/B vssd1 vssd1 vccd1 vccd1 _3244_/Y sky130_fd_sc_hd__xnor2_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3175_ _3917_/A _3444_/B vssd1 vssd1 vccd1 vccd1 _3175_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__3531__A _3916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2126_ _3877_/A _2121_/A _2123_/X _2125_/X vssd1 vssd1 vccd1 vccd1 _2127_/B sky130_fd_sc_hd__o31a_1
XFILLER_3_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3250__B _3420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_2380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_3012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2057_ _4431_/Q _4430_/Q _2036_/D _2054_/B vssd1 vssd1 vccd1 vccd1 _2058_/B sky130_fd_sc_hd__a31o_1
XANTENNA_fanout164_A _2807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_3922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_3381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2959_ _4929_/Q _4928_/D vssd1 vssd1 vccd1 vccd1 _2960_/A sky130_fd_sc_hd__and2b_1
XFILLER_13_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2576__A1 _4710_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_2555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4629_ _4060_/Y _4629_/D _3345_/Y vssd1 vssd1 vccd1 vccd1 _4629_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_30_1898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_3257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
+ _4862_/Q _2878_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_21_3904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_2337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4348__RESET_B fanout195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3196__4_A _3199__7/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3441__A _3445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4514__CLK _3899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4253__A1 _4248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_TE_B
+ _2097_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4664__CLK _2470_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_2499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_3815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3616__A _3616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_2309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
+ _4519_/Q _2272_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_29_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3335__B _3444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput60 _5057_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_Q[1] sky130_fd_sc_hd__buf_2
XFILLER_29_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput71 _5068_/X vssd1 vssd1 vccd1 vccd1 cos_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__4771__RESET_B fanout253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput82 _5079_/X vssd1 vssd1 vccd1 vccd1 fb1_I[7] sky130_fd_sc_hd__buf_2
Xoutput93 _5090_/X vssd1 vssd1 vccd1 vccd1 read_out_Q[0] sky130_fd_sc_hd__buf_2
XFILLER_7_2055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_3469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3351__A _3361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_RESET_B
+ fanout245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4980_ _3549_/Y _4980_/D _3589_/Y vssd1 vssd1 vccd1 vccd1 _4980_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_2620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_TE_B
+ _2543_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3931_ _3931_/A _4131_/A vssd1 vssd1 vccd1 vccd1 _3932_/B sky130_fd_sc_hd__nor2_1
XFILLER_18_3387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3862_ _4372_/Q vssd1 vssd1 vccd1 vccd1 _3905_/A sky130_fd_sc_hd__buf_8
XFILLER_20_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2813_ _4849_/Q _4848_/Q vssd1 vssd1 vccd1 vccd1 _2813_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3793_ _4291_/Q vssd1 vssd1 vccd1 vccd1 _4290_/D sky130_fd_sc_hd__inv_2
XFILLER_14_1827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_2230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2744_ _4803_/Q _2720_/D _2737_/B vssd1 vssd1 vccd1 vccd1 _2745_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__2133__C _2133_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2675_ _4769_/Q _2675_/B vssd1 vssd1 vccd1 vccd1 _2676_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_4037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4414_ _3224_/Y _4414_/D _3754_/Y vssd1 vssd1 vccd1 vccd1 _4414_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_3408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_2832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4345_ _3190_/Y _4345_/D _3763__103/Y vssd1 vssd1 vccd1 vccd1 _4345_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4276_ _4281_/CLK _4276_/D fanout201/X vssd1 vssd1 vccd1 vccd1 _4276_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4441__RESET_B _3236_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3227_ _3233_/A vssd1 vssd1 vccd1 vccd1 _3227_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_2431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3261__A _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
+ _4577_/Q _2370_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2109_ _4468_/Q _4467_/D vssd1 vssd1 vccd1 vccd1 _2110_/A sky130_fd_sc_hd__and2b_1
XFILLER_3_1774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3089_ _4992_/Q _4991_/Q _3057_/D _3086_/B vssd1 vssd1 vccd1 vccd1 _3090_/B sky130_fd_sc_hd__a31o_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk_master clk_master vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk_master/X sky130_fd_sc_hd__clkbuf_16
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2246__B1 _2173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2605__A _4745_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_2027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_2049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_2330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_2341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3436__A _4004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_3_0_w0.cclk_I clkbuf_2_3_0_w0.cclk_I/A vssd1 vssd1 vccd1 vccd1 _4288_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_24_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_2281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2994__B _4951_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_2145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_3745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3171__A _3925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2218__C _2218_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2237__B1 _2173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5098__A _5098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2515__A _2566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4952__RESET_B fanout210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3346__A _4065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2250__A _2327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2460_ _2456_/Y _2457_/Y _2459_/Y vssd1 vssd1 vccd1 vccd1 _2631_/B sky130_fd_sc_hd__a21o_1
XFILLER_6_3717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_4070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2391_ _4614_/Q _2387_/C _2388_/B vssd1 vssd1 vccd1 vccd1 _2392_/B sky130_fd_sc_hd__a21bo_1
X_4130_ _4659_/Q _4658_/Q vssd1 vssd1 vccd1 vccd1 _4131_/D sky130_fd_sc_hd__xnor2_1
XFILLER_9_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_3233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4061_ _4563_/Q vssd1 vssd1 vccd1 vccd1 _4065_/A sky130_fd_sc_hd__buf_12
XFILLER_0_3316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_2690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3012_ _4953_/Q _2988_/D _3005_/B vssd1 vssd1 vccd1 vccd1 _3013_/B sky130_fd_sc_hd__a21bo_1
XFILLER_20_3277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_2784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_2554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_2587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4963_ _1760_/A _4963_/D _3597_/Y vssd1 vssd1 vccd1 vccd1 _4963_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_3162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_3638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_3026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3914_ _3914_/A _3914_/B _3914_/C vssd1 vssd1 vccd1 vccd1 _3917_/B sky130_fd_sc_hd__or3_2
XANTENNA__2425__A _4652_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4894_ _4901_/CLK _4894_/D fanout236/X vssd1 vssd1 vccd1 vccd1 _4894_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_2937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3845_ _3882_/A vssd1 vssd1 vccd1 vccd1 _3845_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_14_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout127_A fanout128/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_4020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2727_ _4799_/Q _2731_/B _2733_/A vssd1 vssd1 vccd1 vccd1 _2774_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__3256__A _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2160__A _2178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_4086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2658_ _4764_/Q _4763_/Q _2658_/C vssd1 vssd1 vccd1 vccd1 _2658_/X sky130_fd_sc_hd__and3_1
X_2589_ _4715_/Q _4714_/Q _2592_/A vssd1 vssd1 vccd1 vccd1 _2589_/Y sky130_fd_sc_hd__nor3_1
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout157/X fanout203/X vssd1 vssd1 vccd1 vccd1 _5082_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_25_2421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout113 _3588_/A vssd1 vssd1 vccd1 vccd1 _3576_/A sky130_fd_sc_hd__buf_4
XFILLER_5_3249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout124 _4712_/CLK vssd1 vssd1 vccd1 vccd1 _4719_/CLK sky130_fd_sc_hd__clkbuf_2
X_4328_ _4063_/B _4328_/D _3166__64/Y vssd1 vssd1 vccd1 vccd1 _4328_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout135 _3375_/A vssd1 vssd1 vccd1 vccd1 _3659_/A sky130_fd_sc_hd__buf_2
XFILLER_9_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout146 _4562_/Q vssd1 vssd1 vccd1 vccd1 _3696_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_input1_A comp_high_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout157 _5058_/A vssd1 vssd1 vccd1 vccd1 fanout157/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout168 _3865_/Y vssd1 vssd1 vccd1 vccd1 _4852_/CLK sky130_fd_sc_hd__buf_6
Xfanout179 _3738_/A vssd1 vssd1 vccd1 vccd1 _3749_/A sky130_fd_sc_hd__clkbuf_2
X_4259_ _4849_/Q vssd1 vssd1 vccd1 vccd1 _4848_/D sky130_fd_sc_hd__inv_2
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_2283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2482__A3 _2490_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_2414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4702__CLK _2631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_3943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4852__CLK _4852_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_2161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_2036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_3553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_3597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_3471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1960_ _4462_/D _4404_/Q _4402_/Q _4401_/Q vssd1 vssd1 vccd1 vccd1 _1961_/C sky130_fd_sc_hd__and4_1
XFILLER_14_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1891_ _4317_/Q _1891_/B vssd1 vssd1 vccd1 vccd1 _4317_/D sky130_fd_sc_hd__xnor2_1
XFILLER_15_2656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2630__B1 _4063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_2391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3561_ _3571_/A vssd1 vssd1 vccd1 vccd1 _3561_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2512_ _2566_/A _2512_/B vssd1 vssd1 vccd1 vccd1 _2513_/B sky130_fd_sc_hd__nand2_1
X_3492_ _3498_/A vssd1 vssd1 vccd1 vccd1 _3492_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_3442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2443_ _4644_/Q _4643_/Q vssd1 vssd1 vccd1 vccd1 _2443_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_6_3525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_3464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_2824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2374_ _4652_/D _4626_/Q _4624_/Q _4623_/Q vssd1 vssd1 vccd1 vccd1 _2375_/C sky130_fd_sc_hd__and4_1
XFILLER_22_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_2785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_2868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4113_ _4639_/Q vssd1 vssd1 vccd1 vccd1 _4640_/D sky130_fd_sc_hd__inv_2
X_5093_ _5093_/A vssd1 vssd1 vccd1 vccd1 _5093_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4044_ _4538_/Q vssd1 vssd1 vccd1 vccd1 _4539_/D sky130_fd_sc_hd__inv_2
XANTENNA__2139__B _4492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_3413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
+ wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2155__A _4485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout244_A fanout245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4946_ _3531_/Y _4946_/D _3599__1/Y vssd1 vssd1 vccd1 vccd1 _4946_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4877_ _3487_/Y _4877_/D _3623_/Y vssd1 vssd1 vccd1 vccd1 _4877_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_3733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3828_ _4340_/Q vssd1 vssd1 vccd1 vccd1 _4341_/D sky130_fd_sc_hd__inv_2
XFILLER_14_2188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_3777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3738_/A fanout187/X vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_27_3217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3764__104 _3765__105/A vssd1 vssd1 vccd1 vccd1 _3764__104/Y sky130_fd_sc_hd__inv_2
XFILLER_27_2527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_3193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3714__A _3721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2688__B1 _2687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[2\].w1.ro_block_Q.ro_pol.tribuf.t_buf _2449_/X _2298_/Y vssd1
+ vssd1 vccd1 vccd1 _5090_/A sky130_fd_sc_hd__ebufn_8
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_2209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4248__C _4248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
+ _4396_/Q _2024_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_28_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn wrapper_cell_loop\[5\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout120/X fanout249/X vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_3611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_2211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_2976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_A
+ _4991_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2915__A1 _4896_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3624__A _4256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5030__CLK _5030_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_2903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_4134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3062__C _4992_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2090_ _4466_/D _4425_/Q vssd1 vssd1 vccd1 vccd1 _2091_/D sky130_fd_sc_hd__xnor2_1
XFILLER_5_2890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_4109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4800_ _4811_/CLK _4800_/D fanout250/X vssd1 vssd1 vccd1 vccd1 _4800_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3425__41_A _3425__41/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2992_ _4958_/Q _4957_/Q _4956_/Q _3028_/A vssd1 vssd1 vccd1 vccd1 _3015_/B sky130_fd_sc_hd__or4_1
X_4731_ _3407_/Y _4731_/D _3663_/Y vssd1 vssd1 vccd1 vccd1 _4731_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_2431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1943_ _3882_/A _3910_/A _3901_/A _1942_/Y _1936_/X vssd1 vssd1 vccd1 vccd1 _1943_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4898__CLK _4901_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4190__A _4190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2703__A _4834_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4662_ _2470_/A1 _4662_/D _3369__33/Y vssd1 vssd1 vccd1 vccd1 _4662_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4285__RESET_B fanout194/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1874_ _4312_/Q _1874_/B vssd1 vssd1 vccd1 vccd1 _4312_/D sky130_fd_sc_hd__xnor2_1
XFILLER_11_1605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3613_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3613_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3518__B _3923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4593_ _1765_/A _4593_/D _3324_/Y vssd1 vssd1 vccd1 vccd1 _4593_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3544_ _3550_/A vssd1 vssd1 vccd1 vccd1 _3544_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2141__C _4485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_4023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf_TE_B
+ _2618_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3475_ _3905_/A _3913_/A vssd1 vssd1 vccd1 vccd1 _3475_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_6_3333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3534__A _3550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2119__C1 _3908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2426_ _2424_/X _2425_/Y _2344_/X vssd1 vssd1 vccd1 vccd1 _2427_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__4278__CLK _4281_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_2665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2357_ _4648_/D _4590_/Q vssd1 vssd1 vccd1 vccd1 _2358_/B sky130_fd_sc_hd__xnor2_1
XFILLER_6_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout194_A fanout196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _5076_/A vssd1 vssd1 vccd1 vccd1 _5076_/X sky130_fd_sc_hd__buf_4
X_2288_ _2119_/X _2287_/X _3892_/B vssd1 vssd1 vccd1 vccd1 _2288_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_1986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4027_ _4507_/Q vssd1 vssd1 vccd1 vccd1 _4506_/D sky130_fd_sc_hd__inv_2
XFILLER_20_2181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_2531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4929_ input31/X _4929_/D fanout218/X vssd1 vssd1 vccd1 vccd1 _4929_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_3541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_2840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_3585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3444__A _3916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout128/X fanout246/X vssd1 vssd1 vccd1 vccd1 _5077_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_22_3681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_2028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_2197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_3007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2507__B _2507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_4028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_2030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3619__A _4256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1939__A2 _3899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2523__A _2566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1784__D _1810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output88_A _5085_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2896__C _4896_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3354__A _3925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2116__A2 _3908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2211_ _4559_/D _4533_/Q _4531_/Q _4530_/Q vssd1 vssd1 vccd1 vccd1 _2248_/A sky130_fd_sc_hd__or4_2
XFILLER_23_3478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2142_ _4484_/Q _2146_/B _2148_/A vssd1 vssd1 vccd1 vccd1 _2191_/C sky130_fd_sc_hd__o21ai_1
XFILLER_1_3241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_3191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2073_ _4433_/Q _2073_/B vssd1 vssd1 vccd1 vccd1 _4433_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__3077__B1 _1791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_3205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_3249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_4117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_4139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4466__RESET_B fanout198/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2975_ _2799_/B _2973_/X _2974_/Y _4131_/C vssd1 vssd1 vccd1 vccd1 _2975_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3529__A _3916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4714_ _4717_/CLK _4714_/D fanout254/X vssd1 vssd1 vccd1 vccd1 _4714_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1926_ _1926_/A vssd1 vssd1 vccd1 vccd1 _1928_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_11_2103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3248__B _3446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_2294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4645_ _2470_/A1 _4645_/D _3361_/Y vssd1 vssd1 vccd1 vccd1 _4645_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1857_ _4319_/Q _4318_/Q _4317_/Q _1857_/D vssd1 vssd1 vccd1 vccd1 _1858_/D sky130_fd_sc_hd__and4_1
XFILLER_28_4046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_4129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_3323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout207_A fanout220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4576_ _5043_/A _4576_/D fanout226/X vssd1 vssd1 vccd1 vccd1 _4576_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1788_ _4274_/Q _1788_/B vssd1 vssd1 vccd1 vccd1 _4274_/D sky130_fd_sc_hd__xor2_1
X_3527_ _3916_/A _3915_/A vssd1 vssd1 vccd1 vccd1 _3527_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_3389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_2655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3458_ _3466_/A vssd1 vssd1 vccd1 vccd1 _3458_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_3163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2409_ _2412_/A _2409_/B vssd1 vssd1 vccd1 vccd1 _2410_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_1976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_3196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_2210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3389_ _3393_/A vssd1 vssd1 vccd1 vccd1 _3389_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_2232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2608__A _2608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5059_ _5059_/A vssd1 vssd1 vccd1 vccd1 _5059_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_3305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2291__A1 _2294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_3051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3439__A _3445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_2946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4443__CLK _4063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3174__A _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4593__CLK _1765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2518__A _2858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_2860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
+ _4904_/Q _2958_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_2871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3349__A _3361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_3769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2760_ _2760_/A vssd1 vssd1 vccd1 vccd1 _2760_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1711_ _4940_/Q vssd1 vssd1 vccd1 vccd1 _4939_/D sky130_fd_sc_hd__inv_2
X_2691_ _2690_/Y _2646_/C _4772_/Q vssd1 vssd1 vccd1 vccd1 _2692_/B sky130_fd_sc_hd__mux2_1
XFILLER_12_2467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4430_ _5033_/A _4430_/D fanout197/X vssd1 vssd1 vccd1 vccd1 _4430_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_3654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4361_ _4472_/CLK _4361_/D fanout202/X vssd1 vssd1 vccd1 vccd1 _4361_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_3529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3084__A _4988_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_4026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4292_ _4063_/B _4292_/D _3153__117/Y vssd1 vssd1 vccd1 vccd1 _4292_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _3255_/A vssd1 vssd1 vccd1 vccd1 _3243_/Y sky130_fd_sc_hd__inv_2
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_3358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _3915_/A vssd1 vssd1 vccd1 vccd1 _3444_/B sky130_fd_sc_hd__buf_12
XFILLER_23_2574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_2585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_2657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3531__B _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2125_ _3901_/A _2464_/C _3900_/Y vssd1 vssd1 vccd1 vccd1 _2125_/X sky130_fd_sc_hd__or3b_1
XANTENNA__2428__A _4652_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4316__CLK _4324_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4647__RESET_B fanout210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2056_ _4428_/Q _2056_/B vssd1 vssd1 vccd1 vccd1 _4428_/D sky130_fd_sc_hd__xnor2_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_4061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout157_A _5058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4466__CLK input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_3809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2958_ _4925_/Q _4924_/Q vssd1 vssd1 vccd1 vccd1 _2958_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_30_3257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
+ _4947_/Q _3053_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_1909_ _1909_/A _1909_/B vssd1 vssd1 vccd1 vccd1 _1910_/B sky130_fd_sc_hd__nand2_1
X_2889_ _4901_/Q _4900_/Q _2889_/C vssd1 vssd1 vccd1 vccd1 _2890_/D sky130_fd_sc_hd__and3_1
XFILLER_11_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4628_ _3344_/Y _4628_/D _3694_/Y vssd1 vssd1 vccd1 vccd1 _4628_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_30_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_2_0_w0.cclk_I clkbuf_2_3_0_w0.cclk_I/A vssd1 vssd1 vccd1 vccd1 _4281_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_11_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4559_ input19/X _4559_/D fanout213/X vssd1 vssd1 vccd1 vccd1 _4560_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_2546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_3916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3722__A _4469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2338__A _2412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2290__A1_N _3941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_2309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3206__13_A _3262__21/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4959__CLK _4962_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_2743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2801__A _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_3827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_2238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_3849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput50 _5047_/X vssd1 vssd1 vccd1 vccd1 cclk_Q[7] sky130_fd_sc_hd__buf_2
Xoutput61 _5058_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_Q[2] sky130_fd_sc_hd__buf_2
XFILLER_8_3781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput72 _5069_/X vssd1 vssd1 vccd1 vccd1 cos_out[5] sky130_fd_sc_hd__buf_2
XFILLER_24_3551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput83 _5080_/X vssd1 vssd1 vccd1 vccd1 fb1_Q[0] sky130_fd_sc_hd__buf_2
Xoutput94 _5091_/X vssd1 vssd1 vccd1 vccd1 read_out_Q[1] sky130_fd_sc_hd__buf_2
XFILLER_7_2067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4339__CLK _3184_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3632__A _3632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_3437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_2714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3767__106_A _3770__109/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4489__CLK _5042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_3809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3930_ _4124_/B vssd1 vssd1 vccd1 vccd1 _3930_/X sky130_fd_sc_hd__buf_4
XFILLER_14_3219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2576__B1_N _2568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3861_ _3897_/A vssd1 vssd1 vccd1 vccd1 _3861_/Y sky130_fd_sc_hd__inv_6
XFILLER_32_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2812_ _4847_/Q _4846_/Q vssd1 vssd1 vccd1 vccd1 _2812_/Y sky130_fd_sc_hd__xnor2_2
X_3792_ _4272_/Q vssd1 vssd1 vccd1 vccd1 _4273_/D sky130_fd_sc_hd__inv_2
XANTENNA__2414__C _2418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2743_ _4801_/Q _2743_/B vssd1 vssd1 vccd1 vccd1 _4801_/D sky130_fd_sc_hd__xnor2_1
XFILLER_30_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_GATE_N _5056_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_4130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2674_ _4766_/Q _2674_/B vssd1 vssd1 vccd1 vccd1 _4766_/D sky130_fd_sc_hd__xnor2_1
XFILLER_29_3440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4413_ _3931_/A _4413_/D _3223_/Y vssd1 vssd1 vccd1 vccd1 _4413_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_3473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2514__B1_N _2507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4344_ _3845_/Y _4344_/D _3189__72/Y vssd1 vssd1 vccd1 vccd1 _4344_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_A
+ _4523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4899__RESET_B fanout232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_2866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3524__50 _3528__52/A vssd1 vssd1 vccd1 vccd1 _3524__50/Y sky130_fd_sc_hd__inv_2
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4275_ _4281_/CLK _4275_/D fanout199/X vssd1 vssd1 vccd1 vccd1 _4275_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3542__A _3550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3226_ _3912_/A _3446_/B vssd1 vssd1 vccd1 vccd1 _3226_/Y sky130_fd_sc_hd__xnor2_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3261__B _3886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_2382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2158__A _4486_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2494__A1 _4671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2108_ _2108_/A vssd1 vssd1 vccd1 vccd1 _2108_/X sky130_fd_sc_hd__clkbuf_1
X_3088_ _4989_/Q _3088_/B vssd1 vssd1 vccd1 vccd1 _4989_/D sky130_fd_sc_hd__xnor2_1
XFILLER_19_2407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1997__A _2061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2039_ _4466_/D _4440_/Q _4438_/Q _4437_/Q vssd1 vssd1 vccd1 vccd1 _2077_/A sky130_fd_sc_hd__or4_2
XFILLER_23_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3717__A _3721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3436__B _3491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout144/X fanout215/X vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_11_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_GATE_N
+ fanout128/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_2354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_3807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3452__A _3466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3530__53 _3656_/A vssd1 vssd1 vccd1 vccd1 _3530__53/Y sky130_fd_sc_hd__inv_2
XFILLER_24_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3171__B _3442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4631__CLK _4916_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1700__A _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4781__CLK _5007_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[5\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf _2962_/A _2813_/Y vssd1
+ vssd1 vccd1 vccd1 _5091_/A sky130_fd_sc_hd__ebufn_8
XFILLER_15_2805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_3241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_2297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_TE_B
+ _2200_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_2551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2531__A _4741_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3346__B _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_3613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_4110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_2912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2390_ _2390_/A _2390_/B vssd1 vssd1 vccd1 vccd1 _4612_/D sky130_fd_sc_hd__xnor2_1
XFILLER_29_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4992__RESET_B fanout237/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_GATE_N
+ _5063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_4082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3362__A _3895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4060_ _4126_/A vssd1 vssd1 vccd1 vccd1 _4060_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_20_3245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3011_ _4951_/Q _3011_/B vssd1 vssd1 vccd1 vccd1 _4951_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
+ _4708_/Q _2613_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_3_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_2599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2706__A _3114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4962_ _4962_/CLK _4962_/D fanout210/X vssd1 vssd1 vccd1 vccd1 _4962_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_3628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3913_ _3913_/A _3913_/B vssd1 vssd1 vccd1 vccd1 _4372_/D sky130_fd_sc_hd__xnor2_1
XFILLER_33_2905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4893_ _4901_/CLK _4893_/D fanout232/X vssd1 vssd1 vccd1 vccd1 _4893_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_14_3038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_3049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_3341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3844_ _3848_/A _3847_/A vssd1 vssd1 vccd1 vccd1 _3882_/A sky130_fd_sc_hd__xnor2_4
XFILLER_31_4086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__1642_ _3266_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__1642_/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__5027__RESET_B fanout237/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3537__A _4249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_2673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2726_ _4802_/Q _4801_/Q _4800_/Q _2737_/B vssd1 vssd1 vccd1 vccd1 _2731_/B sky130_fd_sc_hd__or4_2
XANTENNA__4504__CLK _4063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3256__B _3886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2657_ _4761_/Q _2657_/B vssd1 vssd1 vccd1 vccd1 _4761_/D sky130_fd_sc_hd__xor2_1
XFILLER_9_4098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2588_ _4712_/Q _2588_/B vssd1 vssd1 vccd1 vccd1 _4712_/D sky130_fd_sc_hd__xnor2_1
Xfanout103 _3135_/Y vssd1 vssd1 vccd1 vccd1 _4962_/CLK sky130_fd_sc_hd__buf_2
XANTENNA__2164__B1 _2003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4654__CLK input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout114 _4934_/Q vssd1 vssd1 vccd1 vccd1 _3588_/A sky130_fd_sc_hd__clkbuf_8
X_4327_ _3165_/Y _4327_/D _3773__112/Y vssd1 vssd1 vccd1 vccd1 _4327_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_2433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout125 _4709_/CLK vssd1 vssd1 vccd1 vccd1 _4712_/CLK sky130_fd_sc_hd__buf_2
XANTENNA__3272__A _4004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_2685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout136 _3375_/A vssd1 vssd1 vccd1 vccd1 fanout136/X sky130_fd_sc_hd__clkbuf_2
Xfanout147 _4429_/CLK vssd1 vssd1 vccd1 vccd1 _4402_/CLK sky130_fd_sc_hd__clkbuf_4
Xfanout158 _5058_/A vssd1 vssd1 vccd1 vccd1 fanout158/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4258_ _4846_/Q vssd1 vssd1 vccd1 vccd1 _4847_/D sky130_fd_sc_hd__inv_2
XFILLER_21_2319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout169 _3861_/Y vssd1 vssd1 vccd1 vccd1 _2631_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_25_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4189_ _4189_/A _4190_/B vssd1 vssd1 vccd1 vccd1 _4749_/D sky130_fd_sc_hd__xnor2_1
XFILLER_23_2190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_2295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_2237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
+ _4766_/Q _2710_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
Xwrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn wrapper_cell_loop\[1\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout158/X fanout205/X vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3447__A _3632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_2172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_3955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_2219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3780__121 _3781__122/A vssd1 vssd1 vccd1 vccd1 _3780__121/Y sky130_fd_sc_hd__inv_2
XFILLER_5_3751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1902__B1 _1823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_3565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3259__19 _3262__21/A vssd1 vssd1 vccd1 vccd1 _4473_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_3303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3576_/A fanout251/X vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_15_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2630__A1 _2464_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1890_ _1909_/A _1890_/B vssd1 vssd1 vccd1 vccd1 _1891_/B sky130_fd_sc_hd__nand2_1
XFILLER_15_2668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3357__A _3361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2261__A _4559_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3560_ _4189_/A _4190_/A vssd1 vssd1 vccd1 vccd1 _3560_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_31_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4677__CLK _4717_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2511_ _4677_/Q _4676_/Q _2479_/D _2508_/B vssd1 vssd1 vccd1 vccd1 _2512_/B sky130_fd_sc_hd__a31o_1
X_3491_ _4001_/A _3491_/B vssd1 vssd1 vccd1 vccd1 _3491_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2442_ _4642_/Q _4641_/Q vssd1 vssd1 vccd1 vccd1 _2442_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_6_3537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4188__A _4248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2373_ _4610_/Q _4609_/Q vssd1 vssd1 vccd1 vccd1 _2373_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_26_2764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4112_ _4640_/Q vssd1 vssd1 vccd1 vccd1 _4639_/D sky130_fd_sc_hd__inv_2
XFILLER_22_2628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5092_ _5092_/A vssd1 vssd1 vccd1 vccd1 _5092_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_3053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4043_ _4539_/Q vssd1 vssd1 vccd1 vccd1 _4538_/D sky130_fd_sc_hd__inv_2
XFILLER_20_3075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2139__C _4491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_4104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4945_ _2807_/A _4945_/D _3530__53/Y vssd1 vssd1 vccd1 vccd1 _4945_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_14_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_2281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_2123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4876_ _4248_/B _4876_/D _3486_/Y vssd1 vssd1 vccd1 vccd1 _4876_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_2757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout237_A fanout257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3827_ _4341_/Q vssd1 vssd1 vccd1 vccd1 _4340_/D sky130_fd_sc_hd__inv_2
XFILLER_21_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_2481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3758_ _3948_/A vssd1 vssd1 vccd1 vccd1 _3758_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2709_ _4782_/Q _4781_/Q vssd1 vssd1 vccd1 vccd1 _2709_/Y sky130_fd_sc_hd__xnor2_4
X_3689_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3689_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4843__RESET_B fanout226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
+ _4496_/Q _2203_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_5_3025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_3841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_2285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_3946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3730__A _4010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3264__22 _3264__22/A vssd1 vssd1 vccd1 vccd1 _3264__22/Y sky130_fd_sc_hd__inv_2
XFILLER_31_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3177__A _3913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
+ wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_A
+ _4672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_2587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4584__RESET_B fanout231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3709__94 _3732__95/A vssd1 vssd1 vccd1 vccd1 _3709__94/Y sky130_fd_sc_hd__inv_2
XANTENNA__3905__A _3905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_4030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_3638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_4052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_4063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3469__42_A _3469__42/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_4085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3640__A _3642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2991_ _5020_/D _4962_/Q _4960_/Q _4959_/Q vssd1 vssd1 vccd1 vccd1 _3028_/A sky130_fd_sc_hd__or4_2
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4730_ _4920_/CLK _4730_/D _3406_/Y vssd1 vssd1 vccd1 vccd1 _4730_/Q sky130_fd_sc_hd__dfrtp_4
X_1942_ _3882_/Y vssd1 vssd1 vccd1 vccd1 _1942_/Y sky130_fd_sc_hd__inv_2
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_2919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4661_ _3367_/Y _4661_/D _3683__90/Y vssd1 vssd1 vccd1 vccd1 _4661_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__4190__B _4190_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1873_ _1909_/A _1873_/B vssd1 vssd1 vccd1 vccd1 _1874_/B sky130_fd_sc_hd__nand2_1
X_3612_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3612_/Y sky130_fd_sc_hd__inv_2
X_4592_ _4188_/B _4592_/D _3705_/Y vssd1 vssd1 vccd1 vccd1 _4592_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3543_ _4563_/Q _3543_/B vssd1 vssd1 vccd1 vccd1 _3543_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_2804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2119__B1 _3900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
+ wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2425_ _4652_/D _4626_/Q _4624_/Q vssd1 vssd1 vccd1 vccd1 _2425_/Y sky130_fd_sc_hd__nor3_1
XFILLER_26_3273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_3389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2356_ _4587_/Q _2356_/B vssd1 vssd1 vccd1 vccd1 _4587_/D sky130_fd_sc_hd__xnor2_1
XFILLER_6_2655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_2677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5075_ _5075_/A vssd1 vssd1 vccd1 vccd1 _5075_/X sky130_fd_sc_hd__clkbuf_2
X_2287_ _2287_/A _3931_/A _3900_/A vssd1 vssd1 vccd1 vccd1 _2287_/X sky130_fd_sc_hd__or3b_1
XFILLER_22_2469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3550__A _3550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4026_ _4504_/Q vssd1 vssd1 vccd1 vccd1 _4505_/D sky130_fd_sc_hd__inv_2
XFILLER_0_2265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_2193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_3965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_2218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4842__CLK _5030_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4928_ input31/X _4928_/D fanout214/X vssd1 vssd1 vccd1 vccd1 _4929_/D sky130_fd_sc_hd__dfrtp_1
X_4859_ _4865_/CLK _4859_/D fanout224/X vssd1 vssd1 vccd1 vccd1 _4859_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_3553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4992__CLK _4997_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_2874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3725__A _4010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3444__B _3444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_2419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_clk_master clkbuf_2_3_0_clk_master/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clk_master/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_6_3890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_2143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_3660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3460__A _3466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_2741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_TE_B
+ _3116_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_2785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_2627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4765__RESET_B fanout256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_2362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_3869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3635__A _3642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_4103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_3413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3354__B _3442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4715__CLK _4717_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2210_ _4521_/Q _4520_/Q _2218_/C _2221_/A vssd1 vssd1 vccd1 vccd1 _2262_/B sky130_fd_sc_hd__a31o_1
XFILLER_3_3529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_2723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3190_ _3848_/A _3847_/A vssd1 vssd1 vccd1 vccd1 _3190_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_6_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_2817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2141_ _4487_/Q _4486_/Q _4485_/Q _2152_/B vssd1 vssd1 vccd1 vccd1 _2146_/B sky130_fd_sc_hd__or4_1
XFILLER_26_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3370__A _3895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2072_ _2178_/A _2072_/B vssd1 vssd1 vccd1 vccd1 _2073_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4865__CLK _4865_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_2574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2974_ _3877_/A _4124_/D vssd1 vssd1 vccd1 vccd1 _2974_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_1826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3529__B _3915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_2705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4713_ _4717_/CLK _4713_/D fanout255/X vssd1 vssd1 vccd1 vccd1 _4713_/Q sky130_fd_sc_hd__dfrtp_2
X_1925_ _4349_/Q _4348_/D vssd1 vssd1 vccd1 vccd1 _1926_/A sky130_fd_sc_hd__and2b_1
Xclkbuf_1_0__f__1648_ clkbuf_0__1648_/X vssd1 vssd1 vccd1 vccd1 _3469__42/A sky130_fd_sc_hd__clkbuf_16
XFILLER_34_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2433__B _2433_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_2727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4351__D _4351_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4644_ _3360_/Y _4644_/D _3686_/Y vssd1 vssd1 vccd1 vccd1 _4644_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_30_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1856_ _4321_/Q _4320_/Q _1856_/C vssd1 vssd1 vccd1 vccd1 _1857_/D sky130_fd_sc_hd__and3_1
XFILLER_11_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_1_0_w0.cclk_I clkbuf_2_1_0_w0.cclk_I/A vssd1 vssd1 vccd1 vccd1 _4324_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_28_4058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4575_ _4590_/CLK _4575_/D fanout225/X vssd1 vssd1 vccd1 vccd1 _4575_/Q sky130_fd_sc_hd__dfrtp_2
X_1787_ _2143_/A _1841_/B _1841_/C vssd1 vssd1 vccd1 vccd1 _1788_/B sky130_fd_sc_hd__and3_1
XANTENNA__3545__A _4001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3457_ _4004_/A _3491_/B vssd1 vssd1 vccd1 vccd1 _3457_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4395__CLK _4402_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2408_ _4620_/Q _4619_/Q _2376_/D _2405_/B vssd1 vssd1 vccd1 vccd1 _2409_/B sky130_fd_sc_hd__a31o_1
XFILLER_6_2441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3388_ _3925_/A _3442_/B vssd1 vssd1 vccd1 vccd1 _3388_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_2_3028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_2244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2339_ _4582_/Q _2339_/B vssd1 vssd1 vccd1 vccd1 _4582_/D sky130_fd_sc_hd__xnor2_1
XFILLER_22_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3280__A _3917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5058_ _5058_/A vssd1 vssd1 vccd1 vccd1 _5058_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4009_ _4472_/Q _4009_/B vssd1 vssd1 vccd1 vccd1 _4473_/D sky130_fd_sc_hd__xnor2_1
XFILLER_35_3317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2291__A2 _3932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5020__CLK input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_3085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_4073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_2958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_2969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_2671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3455__A _4065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4738__CLK _2631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xw0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5056_/A fanout190/X vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_3722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_2133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_2199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input32_A phi1b_dig_Q[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4888__CLK _4943_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3190__A _3848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1703__A _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2806__A1 _3941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2534__A _4741_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1710_ _3597_/A vssd1 vssd1 vccd1 vccd1 _4934_/D sky130_fd_sc_hd__inv_2
XFILLER_12_2446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2690_ _2690_/A vssd1 vssd1 vccd1 vccd1 _2690_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4360_ _4360_/CLK _4360_/D fanout198/X vssd1 vssd1 vccd1 vccd1 _4360_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_3508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_4080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3311_ _4469_/Q vssd1 vssd1 vccd1 vccd1 _3311_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4291_ _4003_/C _4291_/D _3784__125/Y vssd1 vssd1 vccd1 vccd1 _4291_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _3935_/A _3440_/B vssd1 vssd1 vccd1 vccd1 _3242_/Y sky130_fd_sc_hd__xnor2_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3264__22_A _3264__22/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2124_ _2286_/B _3941_/A vssd1 vssd1 vccd1 vccd1 _2464_/C sky130_fd_sc_hd__nand2_4
XFILLER_3_2669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2055_ _2046_/C _2054_/X _2003_/X vssd1 vssd1 vccd1 vccd1 _2056_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__3176__67_A _3189__72/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_4051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_4073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_3946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4616__RESET_B fanout232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2957_ _4923_/Q _4922_/Q vssd1 vssd1 vccd1 vccd1 _2957_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_17_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1908_ _4351_/D _4325_/Q vssd1 vssd1 vccd1 vccd1 _1909_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_2546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2888_ _4931_/D _4905_/Q _4903_/Q _4902_/Q vssd1 vssd1 vccd1 vccd1 _2889_/C sky130_fd_sc_hd__and4_1
XFILLER_11_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3732__95_A _3732__95/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4627_ _4248_/B _4627_/D _3343_/Y vssd1 vssd1 vccd1 vccd1 _4627_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1839_ _1839_/A vssd1 vssd1 vccd1 vccd1 _3066_/A sky130_fd_sc_hd__buf_12
XFILLER_28_3121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3275__A _3287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4558_ input19/X input3/X fanout206/X vssd1 vssd1 vccd1 vccd1 _4559_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_28_3165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3509_ _3519_/A vssd1 vssd1 vccd1 vccd1 _3509_/Y sky130_fd_sc_hd__inv_2
X_4489_ _5042_/A _4489_/D fanout201/X vssd1 vssd1 vccd1 vccd1 _4489_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_2475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_2486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_2558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_2497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_2074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3207__14 _3264__22/A vssd1 vssd1 vccd1 vccd1 _3207__14/Y sky130_fd_sc_hd__inv_2
XANTENNA__2354__A _4648_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_2457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3884__S _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4560__CLK input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_3191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput40 _5037_/X vssd1 vssd1 vccd1 vccd1 cclk_I[5] sky130_fd_sc_hd__buf_2
Xoutput51 _5048_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_I[0] sky130_fd_sc_hd__clkbuf_1
XFILLER_4_3613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput62 _5059_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_Q[3] sky130_fd_sc_hd__buf_2
XANTENNA__3913__A _3913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_4117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput73 _5070_/X vssd1 vssd1 vccd1 vccd1 cos_out[6] sky130_fd_sc_hd__buf_2
XFILLER_7_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput84 _5081_/X vssd1 vssd1 vccd1 vccd1 fb1_Q[1] sky130_fd_sc_hd__buf_2
Xoutput95 _5092_/X vssd1 vssd1 vccd1 vccd1 sin_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_2079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_2851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_4002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf_TE_B
+ _2712_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3522__48_A _3523__49/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3860_ _3896_/A _3904_/A vssd1 vssd1 vccd1 vccd1 _3897_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__2264__A _2608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4903__CLK _4905_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2811_ _4126_/A _2811_/B vssd1 vssd1 vccd1 vccd1 _5069_/A sky130_fd_sc_hd__xnor2_2
XFILLER_18_2699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3791_ _4273_/Q vssd1 vssd1 vccd1 vccd1 _4272_/D sky130_fd_sc_hd__inv_2
X_3213__17 _3264__22/A vssd1 vssd1 vccd1 vccd1 _3213__17/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3603__77 _3654__84/A vssd1 vssd1 vccd1 vccd1 _3603__77/Y sky130_fd_sc_hd__inv_2
XFILLER_12_2221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2742_ _2771_/A _2742_/B vssd1 vssd1 vccd1 vccd1 _2743_/B sky130_fd_sc_hd__nand2_1
X_3196__4 _3199__7/A vssd1 vssd1 vccd1 vccd1 _4362_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1766__A1 _4250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_4142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_2265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_2287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2673_ _2680_/A _2673_/B vssd1 vssd1 vccd1 vccd1 _2674_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_3502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3095__A _4994_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_2298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4412_ _3222_/Y _4412_/D _3755_/Y vssd1 vssd1 vccd1 vccd1 _4412_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_29_3452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_3305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_2751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4343_ _3188_/Y _4343_/D _3764__104/Y vssd1 vssd1 vccd1 vccd1 _4343_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4274_ _4281_/CLK _4274_/D fanout199/X vssd1 vssd1 vccd1 vccd1 _4274_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_3112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3225_ _3233_/A vssd1 vssd1 vccd1 vccd1 _3225_/Y sky130_fd_sc_hd__inv_2
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3140__B1 _3139_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_3961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_2394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2494__A2 _2490_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4433__CLK _5041_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2107_ _2107_/A _2107_/B vssd1 vssd1 vccd1 vccd1 _2108_/A sky130_fd_sc_hd__or2_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3087_ _3058_/D _3086_/X _1791_/X vssd1 vssd1 vccd1 vccd1 _3088_/B sky130_fd_sc_hd__o21ai_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2038_ _4428_/Q _4427_/Q _2046_/C _2049_/A vssd1 vssd1 vccd1 vccd1 _2091_/B sky130_fd_sc_hd__a31o_1
XFILLER_17_2121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_3732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4583__CLK _4590_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_2165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3989_ _4454_/Q vssd1 vssd1 vccd1 vccd1 _4453_/D sky130_fd_sc_hd__inv_2
XFILLER_10_3629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3373__35 _3469__42/A vssd1 vssd1 vccd1 vccd1 _3373__35/Y sky130_fd_sc_hd__inv_2
XFILLER_2_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3733__A _3777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_3872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2994__D _3005_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_3988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_2169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2349__A _2412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4926__CLK input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2084__A _4466_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3684_/A fanout217/X vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__dlrtn_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_3854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_3887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3908__A _3908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_A
+ _4954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_2574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3154__118 _3784__125/A vssd1 vssd1 vccd1 vccd1 _3154__118/Y sky130_fd_sc_hd__inv_2
XFILLER_6_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4306__CLK _1952_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_2014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapper_cell_loop\[2\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf _2448_/A _2299_/Y vssd1
+ vssd1 vccd1 vccd1 _5091_/A sky130_fd_sc_hd__ebufn_8
XFILLER_29_2025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_2108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_2047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_4061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_3669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_2935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_2946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_2957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4456__CLK _3252_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_2979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3362__B _3372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2259__A _2327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3010_ _3030_/A _3010_/B vssd1 vssd1 vccd1 vccd1 _3011_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_3257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_3498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_2545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4279__RESET_B fanout201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4961_ _4962_/CLK _4961_/D fanout208/X vssd1 vssd1 vccd1 vccd1 _4961_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_20_1899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_1_1_0_clk_master_A clkbuf_0_clk_master/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3912_ _3912_/A _3913_/B vssd1 vssd1 vccd1 vccd1 _4371_/D sky130_fd_sc_hd__xnor2_1
XFILLER_18_2441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2633__C1 _3929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4892_ _4901_/CLK _4892_/D fanout236/X vssd1 vssd1 vccd1 vccd1 _4892_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_14_2316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3843_ _4359_/Q vssd1 vssd1 vccd1 vccd1 _3847_/A sky130_fd_sc_hd__buf_4
XFILLER_18_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_4098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_2641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3537__B _4250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2936__B1 _2858_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2725_ _4805_/Q _4804_/Q _4803_/Q _2747_/B vssd1 vssd1 vccd1 vccd1 _2737_/B sky130_fd_sc_hd__or4_1
XFILLER_31_2685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_4033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2656_ _2996_/A _2704_/B _2704_/C vssd1 vssd1 vccd1 vccd1 _2657_/B sky130_fd_sc_hd__and3_1
XFILLER_9_3365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2587_ _2680_/A _2587_/B vssd1 vssd1 vccd1 vccd1 _2588_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3553__A _3588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout104 _3135_/Y vssd1 vssd1 vccd1 vccd1 _4958_/CLK sky130_fd_sc_hd__clkbuf_2
X_4326_ _4063_/C _4326_/D _3163__63/Y vssd1 vssd1 vccd1 vccd1 _4326_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout115 _4812_/CLK vssd1 vssd1 vccd1 vccd1 _4809_/CLK sky130_fd_sc_hd__buf_2
Xfanout126 _5044_/A vssd1 vssd1 vccd1 vccd1 _4709_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_25_2445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3272__B _3491_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout137 _5060_/A vssd1 vssd1 vccd1 vccd1 _3375_/A sky130_fd_sc_hd__buf_2
Xfanout148 _2114_/Y vssd1 vssd1 vccd1 vccd1 _4429_/CLK sky130_fd_sc_hd__clkbuf_4
X_4257_ _4847_/Q vssd1 vssd1 vccd1 vccd1 _4846_/D sky130_fd_sc_hd__inv_2
Xfanout159 _4469_/Q vssd1 vssd1 vccd1 vccd1 _5058_/A sky130_fd_sc_hd__buf_4
XFILLER_5_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4949__CLK _4962_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3208_ _3848_/A _3847_/A vssd1 vssd1 vccd1 vccd1 _3208_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_5_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4188_ _4248_/A _4188_/B _4248_/C vssd1 vssd1 vccd1 vccd1 _4190_/B sky130_fd_sc_hd__or3_4
XFILLER_28_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_2274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3526__51_A _3528__52/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3139_ _4124_/D _3136_/X _2978_/C vssd1 vssd1 vccd1 vccd1 _3139_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_16_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1801__A _2858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf _4312_/Q _1921_/Y vssd1
+ vssd1 vccd1 vccd1 w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D sky130_fd_sc_hd__ebufn_8
XANTENNA__3728__A _4010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3463__A _3924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4868__SET_B fanout231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2079__A _2178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_3785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4719__RESET_B fanout255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_4130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2807__A _2807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4372__RESET_B fanout214/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3366__32_A _3366__32/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output101_A _5098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_3662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_3673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3638__A _3642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_2972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_2994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_3709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2510_ _4674_/Q _2510_/B vssd1 vssd1 vccd1 vccd1 _4674_/D sky130_fd_sc_hd__xnor2_1
XFILLER_13_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3490_ _3498_/A vssd1 vssd1 vccd1 vccd1 _3490_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_4145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_3411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2441_ _4640_/Q _4639_/Q vssd1 vssd1 vccd1 vccd1 _2441_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_3455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_2732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2372_ _4608_/Q _4607_/Q vssd1 vssd1 vccd1 vccd1 _2372_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__4188__B _4188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4111_ _4637_/Q vssd1 vssd1 vccd1 vccd1 _4638_/D sky130_fd_sc_hd__inv_2
X_5091_ _5091_/A vssd1 vssd1 vccd1 vccd1 _5091_/X sky130_fd_sc_hd__buf_6
X_4042_ _4536_/Q vssd1 vssd1 vccd1 vccd1 _4537_/D sky130_fd_sc_hd__inv_2
XFILLER_22_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_3065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2139__D _2176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _5055_/A fanout244/X vssd1 vssd1 vccd1 vccd1 _5079_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_4_2583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2717__A _4838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_GATE_N
+ _3576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4944_ _3529_/Y _4944_/D _3602__76/Y vssd1 vssd1 vccd1 vccd1 _4944_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_2113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
+ _4897_/Q _2950_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[5\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_4875_ _3485_/Y _4875_/D _3624_/Y vssd1 vssd1 vccd1 vccd1 _4875_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3548__A _3550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_2769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3826_ _4338_/Q vssd1 vssd1 vccd1 vccd1 _4339_/D sky130_fd_sc_hd__inv_2
XFILLER_18_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout132_A _2455_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3757_ _3948_/A vssd1 vssd1 vccd1 vccd1 _3757_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4621__CLK _4626_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2708_ _4780_/Q _4779_/Q vssd1 vssd1 vccd1 vccd1 _2708_/Y sky130_fd_sc_hd__xnor2_4
X_3688_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3688_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2639_ _4003_/C _2631_/X _2636_/X _2638_/X vssd1 vssd1 vccd1 vccd1 _2640_/B sky130_fd_sc_hd__o31a_2
XANTENNA__2137__A1 _4485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3283__A _3287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4771__CLK _4812_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_2461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_3831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_2494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4309_ _3882_/A _4309_/D _3774__113/Y vssd1 vssd1 vccd1 vccd1 _4309_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_3925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1896__B1 _1823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_2347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_2013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_3657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3458__A _3466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_2522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wrapper_cell_loop\[6\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf_TE_B _2982_/Y
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_3825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
+ _4955_/Q _3045_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[6\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_4042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_2927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1887__B1 _1823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3921__A _3940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4553__RESET_B _3710_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2537__A _2608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2990_ _4950_/Q _4949_/Q _2998_/C _3001_/A vssd1 vssd1 vccd1 vccd1 _3042_/B sky130_fd_sc_hd__a31o_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1941_ _3898_/B _3914_/B _1941_/C vssd1 vssd1 vccd1 vccd1 _1941_/X sky130_fd_sc_hd__and3_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3368__A _3470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_2455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1872_ _4313_/Q _1868_/C _1869_/B vssd1 vssd1 vccd1 vccd1 _1873_/B sky130_fd_sc_hd__a21bo_1
X_4660_ _2470_/A1 _4660_/D _3366__32/Y vssd1 vssd1 vccd1 vccd1 _4660_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf_TE_B
+ _2786_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3611_ _3616_/A vssd1 vssd1 vccd1 vccd1 _3611_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_2_0_0_w0.cclk_I clkbuf_2_1_0_w0.cclk_I/A vssd1 vssd1 vccd1 vccd1 _5040_/A
+ sky130_fd_sc_hd__clkbuf_8
X_4591_ _4248_/B _4591_/D _3323_/Y vssd1 vssd1 vccd1 vccd1 _4591_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_7_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3542_ _3550_/A vssd1 vssd1 vccd1 vccd1 _3542_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_2827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
+ _4612_/Q _2442_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
X_3473_ _3905_/A _3913_/A vssd1 vssd1 vccd1 vccd1 _3473_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_2838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_4058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_4069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2424_ _4652_/D _4626_/Q _4624_/Q vssd1 vssd1 vccd1 vccd1 _2424_/X sky130_fd_sc_hd__and3_1
X_2355_ _2353_/X _2354_/Y _2344_/X vssd1 vssd1 vccd1 vccd1 _2356_/B sky130_fd_sc_hd__o21ai_1
XFILLER_6_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
+ wrapper_cell_loop\[2\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5074_ _5074_/A vssd1 vssd1 vccd1 vccd1 _5074_/X sky130_fd_sc_hd__clkbuf_1
X_2286_ _3910_/A _2286_/B _3931_/A vssd1 vssd1 vccd1 vccd1 _2286_/X sky130_fd_sc_hd__or3_1
XFILLER_4_3092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4025_ _4505_/Q vssd1 vssd1 vccd1 vccd1 _4504_/D sky130_fd_sc_hd__inv_2
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_3977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2055__B1 _2003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4927_ input31/X _4927_/D fanout214/X vssd1 vssd1 vccd1 vccd1 _4928_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_33_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3278__A _3925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2182__A _4555_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1802__B1 _3109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4858_ _4865_/CLK _4858_/D fanout228/X vssd1 vssd1 vccd1 vccd1 _4858_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3809_ _4307_/Q vssd1 vssd1 vccd1 vccd1 _4306_/D sky130_fd_sc_hd__inv_2
XFILLER_14_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4789_ _4920_/CLK _4789_/D _3439_/Y vssd1 vssd1 vccd1 vccd1 _4789_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_2853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_2337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3316__27 _3366__32/A vssd1 vssd1 vccd1 vccd1 _3316__27/Y sky130_fd_sc_hd__inv_2
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_2133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3741__A _3748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_2155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2357__A _4648_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ fanout180/X fanout184/X vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_28_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
+ _4670_/Q _2544_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[3\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2294__B1 _2294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4667__CLK _3374_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_3919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_2753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3188__A _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_2797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_2098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3916__A _3916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_2396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2966__A_N _4932_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_4115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173__66 _3193__75/A vssd1 vssd1 vccd1 vccd1 _3173__66/Y sky130_fd_sc_hd__inv_2
XANTENNA__3651__A _4195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_2735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2140_ _4490_/Q _4489_/Q _4488_/Q _2162_/B vssd1 vssd1 vccd1 vccd1 _2152_/B sky130_fd_sc_hd__or4_1
XFILLER_1_3254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3370__B _3372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2071_ _4434_/Q _2035_/D _2063_/B vssd1 vssd1 vccd1 vccd1 _2072_/B sky130_fd_sc_hd__a21bo_1
XFILLER_1_2531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2973_ _4064_/A _2462_/Y _2978_/B _3877_/A vssd1 vssd1 vccd1 vccd1 _2973_/X sky130_fd_sc_hd__a31o_1
XFILLER_34_2853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4712_ _4712_/CLK _4712_/D fanout256/X vssd1 vssd1 vccd1 vccd1 _4712_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1924_ _4345_/Q _4344_/Q vssd1 vssd1 vccd1 vccd1 _1924_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_30_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4643_ _3861_/Y _4643_/D _3359_/Y vssd1 vssd1 vccd1 vccd1 _4643_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_2138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1855_ _4351_/D _4325_/Q _4323_/Q _4322_/Q vssd1 vssd1 vccd1 vccd1 _1856_/C sky130_fd_sc_hd__and4_1
XFILLER_15_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1786_ _4276_/Q _1790_/B _1793_/A vssd1 vssd1 vccd1 vccd1 _1841_/C sky130_fd_sc_hd__o21ai_1
XFILLER_11_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4574_ _3321_/Y _4574_/D _3706__91/Y vssd1 vssd1 vccd1 vccd1 _4574_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3545__B _4005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3525_ _3916_/A _3915_/A vssd1 vssd1 vccd1 vccd1 _3525_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf_A
+ _4486_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_2729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3456_ _3466_/A vssd1 vssd1 vccd1 vccd1 _3456_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_3165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2407_ _4617_/Q _2407_/B vssd1 vssd1 vccd1 vccd1 _4617_/D sky130_fd_sc_hd__xnor2_1
XFILLER_2_3007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3387_ _3393_/A vssd1 vssd1 vccd1 vccd1 _3387_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3561__A _3571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_3992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2338_ _2412_/A _2338_/B vssd1 vssd1 vccd1 vccd1 _2339_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_2497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_2256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3280__B _3444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5057_ _5057_/A vssd1 vssd1 vccd1 vccd1 _5057_/X sky130_fd_sc_hd__clkbuf_1
X_2269_ _4543_/Q _4542_/Q vssd1 vssd1 vccd1 vccd1 _2269_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_35_4019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4008_ _4473_/Q _4009_/B vssd1 vssd1 vccd1 vccd1 _4472_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_1351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_2617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0_w0.cclk_I _1935_/Y vssd1 vssd1 vccd1 vccd1 clkbuf_0_w0.cclk_I/X sky130_fd_sc_hd__clkbuf_16
XFILLER_35_2639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_3638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_3075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_2937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2640__A _4064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[4\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf_TE_B
+ _2779_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3455__B _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_2145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_2156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3190__B _3847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input25_A phi1b_dig_Q[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2087__A _4466_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2806__A2 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_2815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_2149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xw0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _4363_/CLK fanout191/X vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__dlrtn_1
XANTENNA__4986__RESET_B fanout234/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3646__A _4195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4192__A0 _4064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output93_A _5090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_2911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_4131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3310_ _3891_/A _3889_/A vssd1 vssd1 vccd1 vccd1 _3310_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_29_2966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4290_ _4063_/C _4290_/D _3152__116/Y vssd1 vssd1 vccd1 vccd1 _4290_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_2808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn wrapper_cell_loop\[4\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3643_/A fanout243/X vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__dlrtn_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _3255_/A vssd1 vssd1 vccd1 vccd1 _3241_/Y sky130_fd_sc_hd__inv_2
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4832__CLK _3467_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3381__A _3393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_2762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3172_ _3777_/A vssd1 vssd1 vccd1 vccd1 _3172_/X sky130_fd_sc_hd__buf_1
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2123_ _2294_/B1 _3914_/B _3900_/B _2118_/X vssd1 vssd1 vccd1 vccd1 _2123_/X sky130_fd_sc_hd__o31a_1
XFILLER_3_1936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_3073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2054_ _4429_/Q _2054_/B vssd1 vssd1 vccd1 vccd1 _2054_/X sky130_fd_sc_hd__and2b_1
XFILLER_17_3004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_2394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4682__SET_B fanout236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_4085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3012__B1_N _3005_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_2661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2956_ _4921_/Q _4920_/Q vssd1 vssd1 vccd1 vccd1 _2956_/Y sky130_fd_sc_hd__xnor2_2
X_1907_ _4322_/Q _1907_/B vssd1 vssd1 vccd1 vccd1 _4322_/D sky130_fd_sc_hd__xnor2_1
X_2887_ _4889_/Q _4888_/Q vssd1 vssd1 vccd1 vccd1 _2887_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__3556__A _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_2569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4626_ _4626_/CLK _4626_/D fanout236/X vssd1 vssd1 vccd1 vccd1 _4626_/Q sky130_fd_sc_hd__dfrtp_2
X_1838_ _4287_/Q _1838_/B vssd1 vssd1 vccd1 vccd1 _4287_/D sky130_fd_sc_hd__xnor2_1
XFILLER_30_1857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapper_cell_loop\[5\].w1.ro_block_I.ro_pol.tribuf.t_buf _2968_/X _2814_/Y vssd1
+ vssd1 vccd1 vccd1 _5088_/A sky130_fd_sc_hd__ebufn_8
Xwrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
+ _4431_/Q _2096_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XFILLER_28_3133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4557_ input27/X _4557_/D fanout199/X vssd1 vssd1 vccd1 vccd1 _4557_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_2410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1769_ _5027_/Q vssd1 vssd1 vccd1 vccd1 _5027_/D sky130_fd_sc_hd__clkinv_2
XFILLER_11_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_2432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3508_ _4127_/A _4129_/A vssd1 vssd1 vccd1 vccd1 _3508_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_2443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4488_ _5042_/A _4488_/D fanout201/X vssd1 vssd1 vccd1 vccd1 _4488_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3439_ _3445_/A vssd1 vssd1 vccd1 vccd1 _3439_/Y sky130_fd_sc_hd__inv_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2619__B _4742_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_2125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_2086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_3137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_2881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4705__CLK _4718_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_GATE_N _4359_/CLK
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_2745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3466__A _3466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2972__A1 _4003_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4855__CLK _4905_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wrapper_cell_loop\[2\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_A
+ _4619_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput41 _5038_/X vssd1 vssd1 vccd1 vccd1 cclk_I[6] sky130_fd_sc_hd__buf_2
XFILLER_29_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput52 _5049_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_I[1] sky130_fd_sc_hd__buf_2
XFILLER_8_3761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_2014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput63 _5060_/X vssd1 vssd1 vccd1 vccd1 clkdiv2_Q[4] sky130_fd_sc_hd__buf_2
XANTENNA__3913__B _3913_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput74 _5071_/X vssd1 vssd1 vccd1 vccd1 cos_out[7] sky130_fd_sc_hd__buf_2
XFILLER_4_3625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_4129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput85 _5082_/X vssd1 vssd1 vccd1 vccd1 fb1_Q[2] sky130_fd_sc_hd__buf_2
XFILLER_7_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput96 _5093_/X vssd1 vssd1 vccd1 vccd1 sin_out[1] sky130_fd_sc_hd__buf_2
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_4061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_2968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
+ _4489_/Q _2195_/Y vssd1 vssd1 vccd1 vccd1 wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ sky130_fd_sc_hd__ebufn_8
XANTENNA_wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
+ wrapper_cell_loop\[6\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_4058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
+ wrapper_cell_loop\[1\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_2634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2660__B1 _1975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2264__B _4533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_2678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2810_ _3914_/B _2807_/X _2808_/X _2809_/Y vssd1 vssd1 vccd1 vccd1 _2811_/B sky130_fd_sc_hd__a31o_1
XANTENNA__4385__CLK _3845_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_2801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3790_ _4270_/Q vssd1 vssd1 vccd1 vccd1 _4271_/D sky130_fd_sc_hd__inv_2
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2741_ _4803_/Q _4802_/Q _2720_/D _2738_/B vssd1 vssd1 vccd1 vccd1 _2742_/B sky130_fd_sc_hd__a31o_1
XFILLER_31_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3376__A _3393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_2867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn wrapper_cell_loop\[3\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn/D
+ _3659_/A fanout240/X vssd1 vssd1 vccd1 vccd1 _5076_/A sky130_fd_sc_hd__dlrtn_1
XFILLER_16_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2672_ _4767_/Q _2648_/D _2665_/B vssd1 vssd1 vccd1 vccd1 _2673_/B sky130_fd_sc_hd__a21bo_1
XFILLER_25_4007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_4018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4411_ _3932_/A _4411_/D _3221_/Y vssd1 vssd1 vccd1 vccd1 _4411_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_4029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_3317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4342_ _1952_/A1 _4342_/D _3187__71/Y vssd1 vssd1 vccd1 vccd1 _4342_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4273_ _3846_/A _4273_/D _5048_/A vssd1 vssd1 vccd1 vccd1 _4273_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3224_ _3917_/A _3444_/B vssd1 vssd1 vccd1 vccd1 _3224_/Y sky130_fd_sc_hd__xnor2_1
.ends

