** sch_path: /local_disk/fossi_cochlea/xschem/clkgen/comp_clks_1stage.sch
.subckt comp_clks_1stage clk clka clkb vdd vss
*.PININFO clk:I clka:O clkb:O vdd:B vss:B
X1 clk clka vdd vss inv Wpmos=Wpmos Lpmos=Lpmos Wnmos=Wnmos Lnmos=Lnmos
x2 clk clkb vss vdd vdd vss tg Wpmos=0.63 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
.ends

* expanding   symbol:  inv/inv.sym # of pins=4
** sym_path: /local_disk/fossi_cochlea/xschem/inv/inv.sym
** sch_path: /local_disk/fossi_cochlea/xschem/inv/inv.sch
.subckt inv in out vdd vss   Wpmos=Wpmos Lpmos=Lpmos Wnmos=Wnmos Lnmos=Lnmos
*.PININFO in:I out:B vdd:B vss:B
XM1 vss in out vss sky130_fd_pr__nfet_01v8 L=Lnmos W=Wnmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 vdd in out vdd sky130_fd_pr__pfet_01v8 L=Lpmos W=Wpmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  xschem/transmission_gate/tg.sym # of pins=6
** sym_path: /local_disk/fossi_cochlea/xschem/transmission_gate/tg.sym
** sch_path: /local_disk/fossi_cochlea/xschem/transmission_gate/tg.sch
.subckt tg in out ctrl_ ctrl vdd vss   Wpmos=0.63 Lpmos=0.18 Wnmos=0.42 Lnmos=0.18
*.PININFO in:B out:B ctrl_:I ctrl:I vdd:B vss:B
XM1 out ctrl in vss sky130_fd_pr__nfet_01v8 L=Lnmos W=Wnmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out ctrl_ in vdd sky130_fd_pr__pfet_01v8 L=Lpmos W=Wpmos nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
.ends

.end
