magic
tech sky130A
magscale 1 2
timestamp 1654694538
<< obsli1 >>
rect 1104 2159 58880 47345
<< obsm1 >>
rect 14 552 59878 48816
<< metal2 >>
rect 1950 49200 2006 50000
rect 7746 49200 7802 50000
rect 12898 49200 12954 50000
rect 18694 49200 18750 50000
rect 23846 49200 23902 50000
rect 29642 49200 29698 50000
rect 35438 49200 35494 50000
rect 40590 49200 40646 50000
rect 46386 49200 46442 50000
rect 52182 49200 52238 50000
rect 57334 49200 57390 50000
rect 18 0 74 800
rect 5170 0 5226 800
rect 10966 0 11022 800
rect 16118 0 16174 800
rect 21914 0 21970 800
rect 27710 0 27766 800
rect 32862 0 32918 800
rect 38658 0 38714 800
rect 43810 0 43866 800
rect 49606 0 49662 800
rect 55402 0 55458 800
<< obsm2 >>
rect 18 49144 1894 49314
rect 2062 49144 7690 49314
rect 7858 49144 12842 49314
rect 13010 49144 18638 49314
rect 18806 49144 23790 49314
rect 23958 49144 29586 49314
rect 29754 49144 35382 49314
rect 35550 49144 40534 49314
rect 40702 49144 46330 49314
rect 46498 49144 52126 49314
rect 52294 49144 57278 49314
rect 57446 49144 59872 49314
rect 18 856 59872 49144
rect 130 31 5114 856
rect 5282 31 10910 856
rect 11078 31 16062 856
rect 16230 31 21858 856
rect 22026 31 27654 856
rect 27822 31 32806 856
rect 32974 31 38602 856
rect 38770 31 43754 856
rect 43922 31 49550 856
rect 49718 31 55346 856
rect 55514 31 59872 856
<< metal3 >>
rect 59200 46928 60000 47048
rect 0 46248 800 46368
rect 59200 41488 60000 41608
rect 0 40808 800 40928
rect 59200 35368 60000 35488
rect 0 34688 800 34808
rect 0 29248 800 29368
rect 59200 29248 60000 29368
rect 59200 23808 60000 23928
rect 0 23128 800 23248
rect 59200 17688 60000 17808
rect 0 17008 800 17128
rect 59200 12248 60000 12368
rect 0 11568 800 11688
rect 59200 6128 60000 6248
rect 0 5448 800 5568
rect 59200 8 60000 128
<< obsm3 >>
rect 13 47128 59787 49740
rect 13 46848 59120 47128
rect 13 46448 59787 46848
rect 880 46168 59787 46448
rect 13 41688 59787 46168
rect 13 41408 59120 41688
rect 13 41008 59787 41408
rect 880 40728 59787 41008
rect 13 35568 59787 40728
rect 13 35288 59120 35568
rect 13 34888 59787 35288
rect 880 34608 59787 34888
rect 13 29448 59787 34608
rect 880 29168 59120 29448
rect 13 24008 59787 29168
rect 13 23728 59120 24008
rect 13 23328 59787 23728
rect 880 23048 59787 23328
rect 13 17888 59787 23048
rect 13 17608 59120 17888
rect 13 17208 59787 17608
rect 880 16928 59787 17208
rect 13 12448 59787 16928
rect 13 12168 59120 12448
rect 13 11768 59787 12168
rect 880 11488 59787 11768
rect 13 6328 59787 11488
rect 13 6048 59120 6328
rect 13 5648 59787 6048
rect 880 5368 59787 5648
rect 13 208 59787 5368
rect 13 35 59120 208
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
rect 50288 2128 50608 47376
<< obsm4 >>
rect 427 47456 57717 49741
rect 427 2048 4128 47456
rect 4608 2048 19488 47456
rect 19968 2048 34848 47456
rect 35328 2048 50208 47456
rect 50688 2048 57717 47456
rect 427 307 57717 2048
<< labels >>
rlabel metal2 s 38658 0 38714 800 6 cclk_I[0]
port 1 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 cclk_I[1]
port 2 nsew signal output
rlabel metal2 s 40590 49200 40646 50000 6 cclk_Q[0]
port 3 nsew signal output
rlabel metal3 s 59200 23808 60000 23928 6 cclk_Q[1]
port 4 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 clk_master
port 5 nsew signal input
rlabel metal2 s 35438 49200 35494 50000 6 clkdiv2_I[0]
port 6 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 clkdiv2_I[1]
port 7 nsew signal output
rlabel metal2 s 12898 49200 12954 50000 6 clkdiv2_Q[0]
port 8 nsew signal output
rlabel metal3 s 59200 35368 60000 35488 6 clkdiv2_Q[1]
port 9 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 comp_high_I[0]
port 10 nsew signal input
rlabel metal2 s 57334 49200 57390 50000 6 comp_high_I[1]
port 11 nsew signal input
rlabel metal3 s 59200 41488 60000 41608 6 comp_high_Q[0]
port 12 nsew signal input
rlabel metal2 s 18694 49200 18750 50000 6 comp_high_Q[1]
port 13 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 cos_out[0]
port 14 nsew signal output
rlabel metal3 s 59200 6128 60000 6248 6 cos_out[1]
port 15 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 cos_outb[0]
port 16 nsew signal output
rlabel metal3 s 59200 29248 60000 29368 6 cos_outb[1]
port 17 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 fb1_I[0]
port 18 nsew signal output
rlabel metal2 s 18 0 74 800 6 fb1_I[1]
port 19 nsew signal output
rlabel metal2 s 46386 49200 46442 50000 6 fb1_Q[0]
port 20 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 fb1_Q[1]
port 21 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 fb2_I[0]
port 22 nsew signal output
rlabel metal2 s 7746 49200 7802 50000 6 fb2_I[1]
port 23 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 fb2_Q[0]
port 24 nsew signal output
rlabel metal2 s 52182 49200 52238 50000 6 fb2_Q[1]
port 25 nsew signal output
rlabel metal3 s 59200 8 60000 128 6 phi1b_dig_I[0]
port 26 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 phi1b_dig_I[1]
port 27 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 phi1b_dig_Q[0]
port 28 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 phi1b_dig_Q[1]
port 29 nsew signal input
rlabel metal3 s 59200 12248 60000 12368 6 read_out_I[0]
port 30 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 read_out_I[1]
port 31 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 read_out_Q[0]
port 32 nsew signal output
rlabel metal3 s 59200 46928 60000 47048 6 read_out_Q[1]
port 33 nsew signal output
rlabel metal2 s 23846 49200 23902 50000 6 rstb
port 34 nsew signal input
rlabel metal2 s 29642 49200 29698 50000 6 sin_out[0]
port 35 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 sin_out[1]
port 36 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 sin_outb[0]
port 37 nsew signal output
rlabel metal2 s 1950 49200 2006 50000 6 sin_outb[1]
port 38 nsew signal output
rlabel metal3 s 59200 17688 60000 17808 6 ud_en
port 39 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 40 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 40 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 41 nsew ground input
rlabel metal4 s 50288 2128 50608 47376 6 vssd1
port 41 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 60000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6958664
string GDS_FILE /Volumes/export/isn/abhinav/fossi_cochlea/openlane/digital_unison/runs/digital_unison/results/finishing/digital_unison.magic.gds
string GDS_START 442904
<< end >>

