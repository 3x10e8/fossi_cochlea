VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO filter_p_m
  CLASS BLOCK ;
  FOREIGN filter_p_m ;
  ORIGIN 0.130 1.640 ;
  SIZE 253.920 BY 187.340 ;
  PIN vpb
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 111.820 157.200 253.790 157.700 ;
    END
  END vpb
  PIN cclk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.580 165.160 67.860 185.700 ;
    END
  END cclk
  PIN fb1
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.260 175.700 25.540 185.700 ;
    END
  END fb1
  PIN div2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.900 177.350 110.180 185.700 ;
    END
  END div2
  PIN high_buf
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 152.220 177.405 152.500 185.700 ;
    END
  END high_buf
  PIN phi1b_dig
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 194.540 177.285 194.820 185.700 ;
    END
  END phi1b_dig
  PIN lo
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.860 174.915 237.140 185.700 ;
    END
  END lo
  PIN vnb
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 107.615 158.200 253.790 158.700 ;
    END
  END vnb
  PIN th1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 129.955 153.430 253.790 153.930 ;
    END
  END th1
  PIN inm
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 235.010 4.805 253.790 5.800 ;
    END
  END inm
  PIN inp
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT -0.130 1.300 253.790 2.900 ;
    END
  END inp
  PIN vccd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 196.710 154.430 253.790 154.930 ;
    END
  END vccd1
  PIN th2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 131.855 152.430 253.790 152.930 ;
    END
  END th2
  PIN vssd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 234.450 147.745 253.790 148.245 ;
    END
  END vssd1
  PIN vdda1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 237.920 146.790 253.790 147.290 ;
    END
  END vdda1
  OBS
      LAYER li1 ;
        RECT 3.100 125.140 237.280 175.850 ;
      LAYER met1 ;
        RECT 2.435 125.505 237.945 177.380 ;
      LAYER met2 ;
        RECT 2.460 175.420 24.980 177.450 ;
        RECT 25.820 175.420 67.300 177.450 ;
        RECT 2.460 164.880 67.300 175.420 ;
        RECT 68.140 177.070 109.620 177.450 ;
        RECT 110.460 177.125 151.940 177.450 ;
        RECT 152.780 177.125 194.260 177.450 ;
        RECT 110.460 177.070 194.260 177.125 ;
        RECT 68.140 177.005 194.260 177.070 ;
        RECT 195.100 177.005 236.580 177.450 ;
        RECT 68.140 174.635 236.580 177.005 ;
        RECT 237.420 174.635 237.920 177.450 ;
        RECT 68.140 164.880 237.920 174.635 ;
        RECT 2.460 126.325 237.920 164.880 ;
      LAYER met3 ;
        RECT -0.130 159.100 239.820 177.430 ;
        RECT -0.130 158.700 107.215 159.100 ;
        RECT -0.130 158.590 107.615 158.700 ;
        RECT -0.130 158.290 107.315 158.590 ;
        RECT -0.130 158.200 107.615 158.290 ;
        RECT -0.130 157.800 107.215 158.200 ;
        RECT -0.130 157.700 111.420 157.800 ;
        RECT -0.130 157.570 111.820 157.700 ;
        RECT -0.130 157.270 111.520 157.570 ;
        RECT -0.130 157.200 111.820 157.270 ;
        RECT -0.130 156.800 111.420 157.200 ;
        RECT -0.130 155.330 239.820 156.800 ;
        RECT -0.130 154.330 196.310 155.330 ;
        RECT -0.130 153.930 129.555 154.330 ;
        RECT -0.130 153.825 129.955 153.930 ;
        RECT -0.130 153.790 129.675 153.825 ;
        RECT -0.130 153.510 129.555 153.790 ;
        RECT -0.130 153.430 129.955 153.510 ;
        RECT -0.130 153.030 129.555 153.430 ;
        RECT -0.130 152.930 131.455 153.030 ;
        RECT -0.130 152.850 131.855 152.930 ;
        RECT -0.130 152.570 131.455 152.850 ;
        RECT -0.130 152.560 131.575 152.570 ;
        RECT -0.130 152.430 131.855 152.560 ;
        RECT -0.130 152.030 131.455 152.430 ;
        RECT -0.130 148.645 239.820 152.030 ;
        RECT -0.130 148.245 234.050 148.645 ;
        RECT -0.130 148.240 234.450 148.245 ;
        RECT -0.130 147.750 234.050 148.240 ;
        RECT -0.130 147.745 234.450 147.750 ;
        RECT -0.130 147.345 234.050 147.745 ;
        RECT -0.130 147.290 237.520 147.345 ;
        RECT -0.130 147.280 237.920 147.290 ;
        RECT -0.130 146.390 237.520 147.280 ;
        RECT -0.130 0.000 239.820 146.390 ;
      LAYER met4 ;
        RECT -0.130 6.200 253.790 177.430 ;
        RECT -0.130 5.800 234.610 6.200 ;
        RECT -0.130 5.770 235.010 5.800 ;
        RECT -0.130 4.825 234.610 5.770 ;
        RECT -0.130 4.805 235.010 4.825 ;
        RECT -0.130 4.405 234.610 4.805 ;
        RECT -0.130 -1.640 253.790 4.405 ;
      LAYER met5 ;
        RECT -0.130 4.500 253.790 140.315 ;
        RECT -0.130 -1.640 253.790 -0.300 ;
  END
END filter_p_m
END LIBRARY

