magic
tech sky130A
magscale 1 2
timestamp 1654672330
<< metal1 >>
rect 20794 36889 23521 36899
rect 20794 36837 23463 36889
rect 23515 36837 23521 36889
rect 20794 36827 23521 36837
rect 20796 36406 23372 36416
rect 20796 36354 23314 36406
rect 23366 36354 23372 36406
rect 20796 36344 23372 36354
rect 20793 35798 23222 35808
rect 20793 35746 23164 35798
rect 23216 35746 23222 35798
rect 20793 35736 23222 35746
rect 20799 35314 23072 35324
rect 20799 35262 23014 35314
rect 23066 35262 23072 35314
rect 20799 35252 23072 35262
rect 20796 34716 22922 34726
rect 20796 34664 22864 34716
rect 22916 34664 22922 34716
rect 20796 34654 22922 34664
rect 20800 34226 22772 34236
rect 20800 34174 22714 34226
rect 22766 34174 22772 34226
rect 20800 34164 22772 34174
rect 21221 33072 25095 33112
rect 21219 32952 25093 32992
rect 22710 32881 22763 32887
rect 21122 32832 21174 32872
rect 21219 32832 22710 32872
rect 22763 32832 25093 32872
rect 22710 32823 22763 32829
rect 22861 32754 22914 32760
rect 21224 32712 22861 32752
rect 22914 32712 25098 32752
rect 22861 32696 22914 32702
rect 23312 32639 23365 32645
rect 21224 32592 23312 32632
rect 23365 32592 25098 32632
rect 23312 32581 23365 32587
rect 23462 32518 23515 32524
rect 21226 32472 23462 32512
rect 23515 32472 25100 32512
rect 23462 32460 23515 32466
rect 23011 32399 23064 32405
rect 21225 32352 23011 32392
rect 23064 32352 25099 32392
rect 23011 32341 23064 32347
rect 23164 32280 23217 32286
rect 21231 32232 23164 32272
rect 23217 32232 25105 32272
rect 23164 32222 23217 32228
<< via1 >>
rect 23463 36837 23515 36889
rect 23314 36354 23366 36406
rect 23164 35746 23216 35798
rect 23014 35262 23066 35314
rect 22864 34664 22916 34716
rect 22714 34174 22766 34226
rect 22710 32829 22763 32881
rect 22861 32702 22914 32754
rect 23312 32587 23365 32639
rect 23462 32466 23515 32518
rect 23011 32347 23064 32399
rect 23164 32228 23217 32280
<< metal2 >>
rect 23463 36889 23521 36899
rect 23515 36837 23521 36889
rect 23463 36827 23521 36837
rect 23314 36406 23372 36416
rect 23366 36354 23372 36406
rect 23314 36344 23372 36354
rect 23164 35798 23222 35808
rect 23216 35746 23222 35798
rect 23164 35736 23222 35746
rect 23014 35314 23072 35324
rect 23066 35262 23072 35314
rect 23014 35252 23072 35262
rect 22864 34716 22922 34726
rect 22916 34664 22922 34716
rect 22864 34654 22922 34664
rect 22714 34226 22772 34236
rect 22766 34174 22772 34226
rect 22714 34164 22772 34174
rect 22714 32887 22764 34164
rect 22710 32881 22764 32887
rect 22763 32829 22764 32881
rect 22710 32823 22764 32829
rect 22864 32760 22914 34654
rect 22861 32754 22914 32760
rect 22861 32696 22914 32702
rect 23014 32405 23064 35252
rect 23011 32399 23064 32405
rect 23011 32341 23064 32347
rect 23164 32286 23214 35736
rect 23314 32645 23364 36344
rect 23312 32639 23365 32645
rect 23312 32581 23365 32587
rect 23464 32524 23514 36827
rect 23462 32518 23515 32524
rect 23462 32460 23515 32466
rect 23164 32280 23217 32286
rect 23164 32222 23217 32228
rect 45385 28796 46137 28837
rect 45385 28648 45437 28796
rect 162 28529 821 28572
<< metal3 >>
rect 23124 3422 23125 3742
rect 23124 2782 23125 3102
<< metal4 >>
rect 21753 27742 22287 27822
rect 23946 27744 24480 27824
rect 21753 26296 21849 27742
rect 24384 26318 24480 27744
rect 23124 3483 23125 3682
rect 23124 2842 23125 3041
<< metal5 >>
rect 23124 3422 23125 3742
rect 23124 2782 23125 3102
use comparator  comparator_0 ~/Documents/fossi_cochlea/mag/final_designs/comparator
timestamp 1654672330
transform 1 0 22977 0 1 28070
box -1348 -1057 1627 897
use filter  filter_0
timestamp 1654667219
transform 1 0 358 0 1 0
box -1160 2522 22766 33127
use filter  filter_1
timestamp 1654667219
transform -1 0 45891 0 1 0
box -1160 2522 22766 33127
use filter_clkgen  filter_clkgen_0 ~/Documents/fossi_cochlea/mag/final_designs/clkgen
timestamp 1654584312
transform 1 0 17727 0 1 35989
box -1661 -2136 3360 1229
<< end >>
